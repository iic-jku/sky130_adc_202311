magic
tech sky130A
magscale 1 2
timestamp 1698999411
<< error_s >>
rect 2997 276 3984 345
rect 185 -470 261 -461
rect 620 -468 695 -459
rect 185 -526 190 -470
rect 620 -524 634 -468
rect 185 -533 261 -526
rect 620 -531 695 -524
rect 3447 -970 3481 -936
rect 3519 -970 3553 -936
rect 3591 -970 3625 -936
rect 3663 -970 3697 -936
rect 3735 -970 3769 -936
rect 2926 -1202 3145 -984
rect 3180 -1202 3830 -1108
rect 2926 -1238 3866 -1202
rect 3145 -1312 3866 -1238
<< nwell >>
rect 878 186 3984 276
rect 878 177 3024 186
rect 3068 177 3984 186
rect 878 -73 2727 177
rect 3145 -65 3165 177
rect -676 -144 2727 -73
rect -676 -413 2656 -144
rect -676 -480 -190 -413
rect -674 -482 -190 -480
rect -674 -566 -218 -482
rect 2787 -1276 2825 -1238
rect 2863 -1276 2901 -1238
rect 2939 -1276 2977 -1238
rect 3015 -1276 3053 -1238
rect 3180 -1276 3830 -1238
<< pwell >>
rect -678 1896 -504 2072
rect -312 2038 -138 2214
rect 236 2038 410 2214
rect 784 2038 958 2214
rect 1332 2038 1506 2214
rect 1880 2038 2054 2214
rect 2410 2038 2584 2214
rect 2958 2038 3132 2214
rect 3508 2038 3682 2214
rect 4327 1826 4501 2002
rect -678 1422 -504 1598
rect 4327 1350 4501 1526
rect -678 948 -504 1124
rect 4327 876 4501 1052
rect -678 474 -504 650
rect 4325 408 4499 578
rect -142 -547 -56 -543
rect 938 -547 1024 -543
rect -142 -1300 1024 -547
rect 4325 -684 4499 -508
rect 1437 -783 2115 -762
rect 1349 -1300 2203 -783
rect 4325 -1158 4499 -982
rect -142 -1398 2219 -1300
rect -672 -1864 -498 -1688
rect 4325 -1894 4499 -1718
rect -672 -2338 -498 -2162
rect 4325 -2368 4499 -2192
rect -672 -2812 -498 -2636
rect 4325 -2842 4499 -2666
rect -142 -3372 32 -3196
rect 406 -3372 580 -3196
rect 954 -3372 1128 -3196
rect 1502 -3372 1676 -3196
rect 2050 -3372 2224 -3196
rect 2598 -3372 2772 -3196
rect 3148 -3372 3322 -3196
<< nmos >>
rect 30 -1170 60 -1070
rect 118 -1170 148 -1070
rect 206 -1170 236 -1070
rect 294 -1170 324 -1070
rect 382 -1170 412 -1070
rect 470 -1170 500 -1070
rect 558 -1170 588 -1070
rect 646 -1170 676 -1070
rect 734 -1170 764 -1070
rect 822 -1170 852 -1070
rect 1525 -1188 1555 -788
rect 1617 -1188 1647 -788
rect 1713 -1188 1743 -788
rect 1809 -1188 1839 -788
rect 1905 -1188 1935 -788
rect 1997 -1188 2027 -788
<< pmos >>
rect 12 -343 42 -243
rect 104 -343 134 -243
rect 196 -343 226 -243
rect 288 -343 318 -243
rect 380 -343 410 -243
rect 472 -343 502 -243
rect 564 -343 594 -243
rect 656 -343 686 -243
rect 748 -343 778 -243
rect 840 -343 870 -243
rect 1148 -348 1178 52
rect 1236 -348 1266 52
rect 1324 -348 1354 52
rect 1412 -348 1442 52
rect 1500 -348 1530 52
rect 1588 -348 1618 52
rect 1935 -348 1965 52
rect 2023 -348 2053 52
rect 2111 -348 2141 52
rect 2199 -348 2229 52
rect 2287 -348 2317 52
rect 2375 -348 2405 52
<< nmoslvt >>
rect 30 -973 60 -573
rect 118 -973 148 -573
rect 206 -973 236 -573
rect 294 -973 324 -573
rect 382 -973 412 -573
rect 470 -973 500 -573
rect 558 -973 588 -573
rect 646 -973 676 -573
rect 734 -973 764 -573
rect 822 -973 852 -573
<< ndiff >>
rect -28 -586 30 -573
rect -28 -620 -16 -586
rect 18 -620 30 -586
rect -28 -654 30 -620
rect -28 -688 -16 -654
rect 18 -688 30 -654
rect -28 -722 30 -688
rect -28 -756 -16 -722
rect 18 -756 30 -722
rect -28 -790 30 -756
rect -28 -824 -16 -790
rect 18 -824 30 -790
rect -28 -858 30 -824
rect -28 -892 -16 -858
rect 18 -892 30 -858
rect -28 -926 30 -892
rect -28 -960 -16 -926
rect 18 -960 30 -926
rect -28 -973 30 -960
rect 60 -586 118 -573
rect 60 -620 72 -586
rect 106 -620 118 -586
rect 60 -654 118 -620
rect 60 -688 72 -654
rect 106 -688 118 -654
rect 60 -722 118 -688
rect 60 -756 72 -722
rect 106 -756 118 -722
rect 60 -790 118 -756
rect 60 -824 72 -790
rect 106 -824 118 -790
rect 60 -858 118 -824
rect 60 -892 72 -858
rect 106 -892 118 -858
rect 60 -926 118 -892
rect 60 -960 72 -926
rect 106 -960 118 -926
rect 60 -973 118 -960
rect 148 -586 206 -573
rect 148 -620 160 -586
rect 194 -620 206 -586
rect 148 -654 206 -620
rect 148 -688 160 -654
rect 194 -688 206 -654
rect 148 -722 206 -688
rect 148 -756 160 -722
rect 194 -756 206 -722
rect 148 -790 206 -756
rect 148 -824 160 -790
rect 194 -824 206 -790
rect 148 -858 206 -824
rect 148 -892 160 -858
rect 194 -892 206 -858
rect 148 -926 206 -892
rect 148 -960 160 -926
rect 194 -960 206 -926
rect 148 -973 206 -960
rect 236 -586 294 -573
rect 236 -620 248 -586
rect 282 -620 294 -586
rect 236 -654 294 -620
rect 236 -688 248 -654
rect 282 -688 294 -654
rect 236 -722 294 -688
rect 236 -756 248 -722
rect 282 -756 294 -722
rect 236 -790 294 -756
rect 236 -824 248 -790
rect 282 -824 294 -790
rect 236 -858 294 -824
rect 236 -892 248 -858
rect 282 -892 294 -858
rect 236 -926 294 -892
rect 236 -960 248 -926
rect 282 -960 294 -926
rect 236 -973 294 -960
rect 324 -586 382 -573
rect 324 -620 336 -586
rect 370 -620 382 -586
rect 324 -654 382 -620
rect 324 -688 336 -654
rect 370 -688 382 -654
rect 324 -722 382 -688
rect 324 -756 336 -722
rect 370 -756 382 -722
rect 324 -790 382 -756
rect 324 -824 336 -790
rect 370 -824 382 -790
rect 324 -858 382 -824
rect 324 -892 336 -858
rect 370 -892 382 -858
rect 324 -926 382 -892
rect 324 -960 336 -926
rect 370 -960 382 -926
rect 324 -973 382 -960
rect 412 -586 470 -573
rect 412 -620 424 -586
rect 458 -620 470 -586
rect 412 -654 470 -620
rect 412 -688 424 -654
rect 458 -688 470 -654
rect 412 -722 470 -688
rect 412 -756 424 -722
rect 458 -756 470 -722
rect 412 -790 470 -756
rect 412 -824 424 -790
rect 458 -824 470 -790
rect 412 -858 470 -824
rect 412 -892 424 -858
rect 458 -892 470 -858
rect 412 -926 470 -892
rect 412 -960 424 -926
rect 458 -960 470 -926
rect 412 -973 470 -960
rect 500 -586 558 -573
rect 500 -620 512 -586
rect 546 -620 558 -586
rect 500 -654 558 -620
rect 500 -688 512 -654
rect 546 -688 558 -654
rect 500 -722 558 -688
rect 500 -756 512 -722
rect 546 -756 558 -722
rect 500 -790 558 -756
rect 500 -824 512 -790
rect 546 -824 558 -790
rect 500 -858 558 -824
rect 500 -892 512 -858
rect 546 -892 558 -858
rect 500 -926 558 -892
rect 500 -960 512 -926
rect 546 -960 558 -926
rect 500 -973 558 -960
rect 588 -586 646 -573
rect 588 -620 600 -586
rect 634 -620 646 -586
rect 588 -654 646 -620
rect 588 -688 600 -654
rect 634 -688 646 -654
rect 588 -722 646 -688
rect 588 -756 600 -722
rect 634 -756 646 -722
rect 588 -790 646 -756
rect 588 -824 600 -790
rect 634 -824 646 -790
rect 588 -858 646 -824
rect 588 -892 600 -858
rect 634 -892 646 -858
rect 588 -926 646 -892
rect 588 -960 600 -926
rect 634 -960 646 -926
rect 588 -973 646 -960
rect 676 -586 734 -573
rect 676 -620 688 -586
rect 722 -620 734 -586
rect 676 -654 734 -620
rect 676 -688 688 -654
rect 722 -688 734 -654
rect 676 -722 734 -688
rect 676 -756 688 -722
rect 722 -756 734 -722
rect 676 -790 734 -756
rect 676 -824 688 -790
rect 722 -824 734 -790
rect 676 -858 734 -824
rect 676 -892 688 -858
rect 722 -892 734 -858
rect 676 -926 734 -892
rect 676 -960 688 -926
rect 722 -960 734 -926
rect 676 -973 734 -960
rect 764 -586 822 -573
rect 764 -620 776 -586
rect 810 -620 822 -586
rect 764 -654 822 -620
rect 764 -688 776 -654
rect 810 -688 822 -654
rect 764 -722 822 -688
rect 764 -756 776 -722
rect 810 -756 822 -722
rect 764 -790 822 -756
rect 764 -824 776 -790
rect 810 -824 822 -790
rect 764 -858 822 -824
rect 764 -892 776 -858
rect 810 -892 822 -858
rect 764 -926 822 -892
rect 764 -960 776 -926
rect 810 -960 822 -926
rect 764 -973 822 -960
rect 852 -586 910 -573
rect 852 -620 864 -586
rect 898 -620 910 -586
rect 852 -654 910 -620
rect 852 -688 864 -654
rect 898 -688 910 -654
rect 852 -722 910 -688
rect 852 -756 864 -722
rect 898 -756 910 -722
rect 852 -790 910 -756
rect 852 -824 864 -790
rect 898 -824 910 -790
rect 852 -858 910 -824
rect 852 -892 864 -858
rect 898 -892 910 -858
rect 852 -926 910 -892
rect 852 -960 864 -926
rect 898 -960 910 -926
rect 852 -973 910 -960
rect 1463 -801 1525 -788
rect -28 -1103 30 -1070
rect -28 -1137 -16 -1103
rect 18 -1137 30 -1103
rect -28 -1170 30 -1137
rect 60 -1103 118 -1070
rect 60 -1137 72 -1103
rect 106 -1137 118 -1103
rect 60 -1170 118 -1137
rect 148 -1103 206 -1070
rect 148 -1137 160 -1103
rect 194 -1137 206 -1103
rect 148 -1170 206 -1137
rect 236 -1103 294 -1070
rect 236 -1137 248 -1103
rect 282 -1137 294 -1103
rect 236 -1170 294 -1137
rect 324 -1103 382 -1070
rect 324 -1137 336 -1103
rect 370 -1137 382 -1103
rect 324 -1170 382 -1137
rect 412 -1103 470 -1070
rect 412 -1137 424 -1103
rect 458 -1137 470 -1103
rect 412 -1170 470 -1137
rect 500 -1103 558 -1070
rect 500 -1137 512 -1103
rect 546 -1137 558 -1103
rect 500 -1170 558 -1137
rect 588 -1103 646 -1070
rect 588 -1137 600 -1103
rect 634 -1137 646 -1103
rect 588 -1170 646 -1137
rect 676 -1103 734 -1070
rect 676 -1137 688 -1103
rect 722 -1137 734 -1103
rect 676 -1170 734 -1137
rect 764 -1103 822 -1070
rect 764 -1137 776 -1103
rect 810 -1137 822 -1103
rect 764 -1170 822 -1137
rect 852 -1103 910 -1070
rect 852 -1137 864 -1103
rect 898 -1137 910 -1103
rect 852 -1170 910 -1137
rect 1463 -835 1475 -801
rect 1509 -835 1525 -801
rect 1463 -869 1525 -835
rect 1463 -903 1475 -869
rect 1509 -903 1525 -869
rect 1463 -937 1525 -903
rect 1463 -971 1475 -937
rect 1509 -971 1525 -937
rect 1463 -1005 1525 -971
rect 1463 -1039 1475 -1005
rect 1509 -1039 1525 -1005
rect 1463 -1073 1525 -1039
rect 1463 -1107 1475 -1073
rect 1509 -1107 1525 -1073
rect 1463 -1141 1525 -1107
rect 1463 -1175 1475 -1141
rect 1509 -1175 1525 -1141
rect 1463 -1188 1525 -1175
rect 1555 -801 1617 -788
rect 1555 -835 1567 -801
rect 1601 -835 1617 -801
rect 1555 -869 1617 -835
rect 1555 -903 1567 -869
rect 1601 -903 1617 -869
rect 1555 -937 1617 -903
rect 1555 -971 1567 -937
rect 1601 -971 1617 -937
rect 1555 -1005 1617 -971
rect 1555 -1039 1567 -1005
rect 1601 -1039 1617 -1005
rect 1555 -1073 1617 -1039
rect 1555 -1107 1567 -1073
rect 1601 -1107 1617 -1073
rect 1555 -1141 1617 -1107
rect 1555 -1175 1567 -1141
rect 1601 -1175 1617 -1141
rect 1555 -1188 1617 -1175
rect 1647 -801 1713 -788
rect 1647 -835 1663 -801
rect 1697 -835 1713 -801
rect 1647 -869 1713 -835
rect 1647 -903 1663 -869
rect 1697 -903 1713 -869
rect 1647 -937 1713 -903
rect 1647 -971 1663 -937
rect 1697 -971 1713 -937
rect 1647 -1005 1713 -971
rect 1647 -1039 1663 -1005
rect 1697 -1039 1713 -1005
rect 1647 -1073 1713 -1039
rect 1647 -1107 1663 -1073
rect 1697 -1107 1713 -1073
rect 1647 -1141 1713 -1107
rect 1647 -1175 1663 -1141
rect 1697 -1175 1713 -1141
rect 1647 -1188 1713 -1175
rect 1743 -801 1809 -788
rect 1743 -835 1759 -801
rect 1793 -835 1809 -801
rect 1743 -869 1809 -835
rect 1743 -903 1759 -869
rect 1793 -903 1809 -869
rect 1743 -937 1809 -903
rect 1743 -971 1759 -937
rect 1793 -971 1809 -937
rect 1743 -1005 1809 -971
rect 1743 -1039 1759 -1005
rect 1793 -1039 1809 -1005
rect 1743 -1073 1809 -1039
rect 1743 -1107 1759 -1073
rect 1793 -1107 1809 -1073
rect 1743 -1141 1809 -1107
rect 1743 -1175 1759 -1141
rect 1793 -1175 1809 -1141
rect 1743 -1188 1809 -1175
rect 1839 -801 1905 -788
rect 1839 -835 1855 -801
rect 1889 -835 1905 -801
rect 1839 -869 1905 -835
rect 1839 -903 1855 -869
rect 1889 -903 1905 -869
rect 1839 -937 1905 -903
rect 1839 -971 1855 -937
rect 1889 -971 1905 -937
rect 1839 -1005 1905 -971
rect 1839 -1039 1855 -1005
rect 1889 -1039 1905 -1005
rect 1839 -1073 1905 -1039
rect 1839 -1107 1855 -1073
rect 1889 -1107 1905 -1073
rect 1839 -1141 1905 -1107
rect 1839 -1175 1855 -1141
rect 1889 -1175 1905 -1141
rect 1839 -1188 1905 -1175
rect 1935 -801 1997 -788
rect 1935 -835 1951 -801
rect 1985 -835 1997 -801
rect 1935 -869 1997 -835
rect 1935 -903 1951 -869
rect 1985 -903 1997 -869
rect 1935 -937 1997 -903
rect 1935 -971 1951 -937
rect 1985 -971 1997 -937
rect 1935 -1005 1997 -971
rect 1935 -1039 1951 -1005
rect 1985 -1039 1997 -1005
rect 1935 -1073 1997 -1039
rect 1935 -1107 1951 -1073
rect 1985 -1107 1997 -1073
rect 1935 -1141 1997 -1107
rect 1935 -1175 1951 -1141
rect 1985 -1175 1997 -1141
rect 1935 -1188 1997 -1175
rect 2027 -801 2089 -788
rect 2027 -835 2043 -801
rect 2077 -835 2089 -801
rect 2027 -869 2089 -835
rect 2027 -903 2043 -869
rect 2077 -903 2089 -869
rect 2027 -937 2089 -903
rect 2027 -971 2043 -937
rect 2077 -971 2089 -937
rect 2027 -1005 2089 -971
rect 2027 -1039 2043 -1005
rect 2077 -1039 2089 -1005
rect 2027 -1073 2089 -1039
rect 2027 -1107 2043 -1073
rect 2077 -1107 2089 -1073
rect 2027 -1141 2089 -1107
rect 2027 -1175 2043 -1141
rect 2077 -1175 2089 -1141
rect 2027 -1188 2089 -1175
<< pdiff >>
rect 1090 39 1148 52
rect 1090 5 1102 39
rect 1136 5 1148 39
rect 1090 -29 1148 5
rect 1090 -63 1102 -29
rect 1136 -63 1148 -29
rect 1090 -97 1148 -63
rect 1090 -131 1102 -97
rect 1136 -131 1148 -97
rect 1090 -165 1148 -131
rect 1090 -199 1102 -165
rect 1136 -199 1148 -165
rect 1090 -233 1148 -199
rect -50 -276 12 -243
rect -50 -310 -38 -276
rect -4 -310 12 -276
rect -50 -343 12 -310
rect 42 -276 104 -243
rect 42 -310 54 -276
rect 88 -310 104 -276
rect 42 -343 104 -310
rect 134 -276 196 -243
rect 134 -310 148 -276
rect 182 -310 196 -276
rect 134 -343 196 -310
rect 226 -276 288 -243
rect 226 -310 240 -276
rect 274 -310 288 -276
rect 226 -343 288 -310
rect 318 -276 380 -243
rect 318 -310 332 -276
rect 366 -310 380 -276
rect 318 -343 380 -310
rect 410 -276 472 -243
rect 410 -310 424 -276
rect 458 -310 472 -276
rect 410 -343 472 -310
rect 502 -276 564 -243
rect 502 -310 516 -276
rect 550 -310 564 -276
rect 502 -343 564 -310
rect 594 -276 656 -243
rect 594 -310 608 -276
rect 642 -310 656 -276
rect 594 -343 656 -310
rect 686 -276 748 -243
rect 686 -310 700 -276
rect 734 -310 748 -276
rect 686 -343 748 -310
rect 778 -276 840 -243
rect 778 -310 794 -276
rect 828 -310 840 -276
rect 778 -343 840 -310
rect 870 -276 932 -243
rect 870 -310 886 -276
rect 920 -310 932 -276
rect 870 -343 932 -310
rect 1090 -267 1102 -233
rect 1136 -267 1148 -233
rect 1090 -301 1148 -267
rect 1090 -335 1102 -301
rect 1136 -335 1148 -301
rect 1090 -348 1148 -335
rect 1178 39 1236 52
rect 1178 5 1190 39
rect 1224 5 1236 39
rect 1178 -29 1236 5
rect 1178 -63 1190 -29
rect 1224 -63 1236 -29
rect 1178 -97 1236 -63
rect 1178 -131 1190 -97
rect 1224 -131 1236 -97
rect 1178 -165 1236 -131
rect 1178 -199 1190 -165
rect 1224 -199 1236 -165
rect 1178 -233 1236 -199
rect 1178 -267 1190 -233
rect 1224 -267 1236 -233
rect 1178 -301 1236 -267
rect 1178 -335 1190 -301
rect 1224 -335 1236 -301
rect 1178 -348 1236 -335
rect 1266 39 1324 52
rect 1266 5 1278 39
rect 1312 5 1324 39
rect 1266 -29 1324 5
rect 1266 -63 1278 -29
rect 1312 -63 1324 -29
rect 1266 -97 1324 -63
rect 1266 -131 1278 -97
rect 1312 -131 1324 -97
rect 1266 -165 1324 -131
rect 1266 -199 1278 -165
rect 1312 -199 1324 -165
rect 1266 -233 1324 -199
rect 1266 -267 1278 -233
rect 1312 -267 1324 -233
rect 1266 -301 1324 -267
rect 1266 -335 1278 -301
rect 1312 -335 1324 -301
rect 1266 -348 1324 -335
rect 1354 39 1412 52
rect 1354 5 1366 39
rect 1400 5 1412 39
rect 1354 -29 1412 5
rect 1354 -63 1366 -29
rect 1400 -63 1412 -29
rect 1354 -97 1412 -63
rect 1354 -131 1366 -97
rect 1400 -131 1412 -97
rect 1354 -165 1412 -131
rect 1354 -199 1366 -165
rect 1400 -199 1412 -165
rect 1354 -233 1412 -199
rect 1354 -267 1366 -233
rect 1400 -267 1412 -233
rect 1354 -301 1412 -267
rect 1354 -335 1366 -301
rect 1400 -335 1412 -301
rect 1354 -348 1412 -335
rect 1442 39 1500 52
rect 1442 5 1454 39
rect 1488 5 1500 39
rect 1442 -29 1500 5
rect 1442 -63 1454 -29
rect 1488 -63 1500 -29
rect 1442 -97 1500 -63
rect 1442 -131 1454 -97
rect 1488 -131 1500 -97
rect 1442 -165 1500 -131
rect 1442 -199 1454 -165
rect 1488 -199 1500 -165
rect 1442 -233 1500 -199
rect 1442 -267 1454 -233
rect 1488 -267 1500 -233
rect 1442 -301 1500 -267
rect 1442 -335 1454 -301
rect 1488 -335 1500 -301
rect 1442 -348 1500 -335
rect 1530 39 1588 52
rect 1530 5 1542 39
rect 1576 5 1588 39
rect 1530 -29 1588 5
rect 1530 -63 1542 -29
rect 1576 -63 1588 -29
rect 1530 -97 1588 -63
rect 1530 -131 1542 -97
rect 1576 -131 1588 -97
rect 1530 -165 1588 -131
rect 1530 -199 1542 -165
rect 1576 -199 1588 -165
rect 1530 -233 1588 -199
rect 1530 -267 1542 -233
rect 1576 -267 1588 -233
rect 1530 -301 1588 -267
rect 1530 -335 1542 -301
rect 1576 -335 1588 -301
rect 1530 -348 1588 -335
rect 1618 39 1676 52
rect 1618 5 1630 39
rect 1664 5 1676 39
rect 1618 -29 1676 5
rect 1618 -63 1630 -29
rect 1664 -63 1676 -29
rect 1618 -97 1676 -63
rect 1618 -131 1630 -97
rect 1664 -131 1676 -97
rect 1618 -165 1676 -131
rect 1618 -199 1630 -165
rect 1664 -199 1676 -165
rect 1618 -233 1676 -199
rect 1618 -267 1630 -233
rect 1664 -267 1676 -233
rect 1618 -301 1676 -267
rect 1618 -335 1630 -301
rect 1664 -335 1676 -301
rect 1618 -348 1676 -335
rect 1877 39 1935 52
rect 1877 5 1889 39
rect 1923 5 1935 39
rect 1877 -29 1935 5
rect 1877 -63 1889 -29
rect 1923 -63 1935 -29
rect 1877 -97 1935 -63
rect 1877 -131 1889 -97
rect 1923 -131 1935 -97
rect 1877 -165 1935 -131
rect 1877 -199 1889 -165
rect 1923 -199 1935 -165
rect 1877 -233 1935 -199
rect 1877 -267 1889 -233
rect 1923 -267 1935 -233
rect 1877 -301 1935 -267
rect 1877 -335 1889 -301
rect 1923 -335 1935 -301
rect 1877 -348 1935 -335
rect 1965 39 2023 52
rect 1965 5 1977 39
rect 2011 5 2023 39
rect 1965 -29 2023 5
rect 1965 -63 1977 -29
rect 2011 -63 2023 -29
rect 1965 -97 2023 -63
rect 1965 -131 1977 -97
rect 2011 -131 2023 -97
rect 1965 -165 2023 -131
rect 1965 -199 1977 -165
rect 2011 -199 2023 -165
rect 1965 -233 2023 -199
rect 1965 -267 1977 -233
rect 2011 -267 2023 -233
rect 1965 -301 2023 -267
rect 1965 -335 1977 -301
rect 2011 -335 2023 -301
rect 1965 -348 2023 -335
rect 2053 39 2111 52
rect 2053 5 2065 39
rect 2099 5 2111 39
rect 2053 -29 2111 5
rect 2053 -63 2065 -29
rect 2099 -63 2111 -29
rect 2053 -97 2111 -63
rect 2053 -131 2065 -97
rect 2099 -131 2111 -97
rect 2053 -165 2111 -131
rect 2053 -199 2065 -165
rect 2099 -199 2111 -165
rect 2053 -233 2111 -199
rect 2053 -267 2065 -233
rect 2099 -267 2111 -233
rect 2053 -301 2111 -267
rect 2053 -335 2065 -301
rect 2099 -335 2111 -301
rect 2053 -348 2111 -335
rect 2141 39 2199 52
rect 2141 5 2153 39
rect 2187 5 2199 39
rect 2141 -29 2199 5
rect 2141 -63 2153 -29
rect 2187 -63 2199 -29
rect 2141 -97 2199 -63
rect 2141 -131 2153 -97
rect 2187 -131 2199 -97
rect 2141 -165 2199 -131
rect 2141 -199 2153 -165
rect 2187 -199 2199 -165
rect 2141 -233 2199 -199
rect 2141 -267 2153 -233
rect 2187 -267 2199 -233
rect 2141 -301 2199 -267
rect 2141 -335 2153 -301
rect 2187 -335 2199 -301
rect 2141 -348 2199 -335
rect 2229 39 2287 52
rect 2229 5 2241 39
rect 2275 5 2287 39
rect 2229 -29 2287 5
rect 2229 -63 2241 -29
rect 2275 -63 2287 -29
rect 2229 -97 2287 -63
rect 2229 -131 2241 -97
rect 2275 -131 2287 -97
rect 2229 -165 2287 -131
rect 2229 -199 2241 -165
rect 2275 -199 2287 -165
rect 2229 -233 2287 -199
rect 2229 -267 2241 -233
rect 2275 -267 2287 -233
rect 2229 -301 2287 -267
rect 2229 -335 2241 -301
rect 2275 -335 2287 -301
rect 2229 -348 2287 -335
rect 2317 39 2375 52
rect 2317 5 2329 39
rect 2363 5 2375 39
rect 2317 -29 2375 5
rect 2317 -63 2329 -29
rect 2363 -63 2375 -29
rect 2317 -97 2375 -63
rect 2317 -131 2329 -97
rect 2363 -131 2375 -97
rect 2317 -165 2375 -131
rect 2317 -199 2329 -165
rect 2363 -199 2375 -165
rect 2317 -233 2375 -199
rect 2317 -267 2329 -233
rect 2363 -267 2375 -233
rect 2317 -301 2375 -267
rect 2317 -335 2329 -301
rect 2363 -335 2375 -301
rect 2317 -348 2375 -335
rect 2405 39 2463 52
rect 2405 5 2417 39
rect 2451 5 2463 39
rect 2405 -29 2463 5
rect 2405 -63 2417 -29
rect 2451 -63 2463 -29
rect 2405 -97 2463 -63
rect 2405 -131 2417 -97
rect 2451 -131 2463 -97
rect 2405 -165 2463 -131
rect 2405 -199 2417 -165
rect 2451 -199 2463 -165
rect 2405 -233 2463 -199
rect 2405 -267 2417 -233
rect 2451 -267 2463 -233
rect 2405 -301 2463 -267
rect 2405 -335 2417 -301
rect 2451 -335 2463 -301
rect 2405 -348 2463 -335
<< ndiffc >>
rect -16 -620 18 -586
rect -16 -688 18 -654
rect -16 -756 18 -722
rect -16 -824 18 -790
rect -16 -892 18 -858
rect -16 -960 18 -926
rect 72 -620 106 -586
rect 72 -688 106 -654
rect 72 -756 106 -722
rect 72 -824 106 -790
rect 72 -892 106 -858
rect 72 -960 106 -926
rect 160 -620 194 -586
rect 160 -688 194 -654
rect 160 -756 194 -722
rect 160 -824 194 -790
rect 160 -892 194 -858
rect 160 -960 194 -926
rect 248 -620 282 -586
rect 248 -688 282 -654
rect 248 -756 282 -722
rect 248 -824 282 -790
rect 248 -892 282 -858
rect 248 -960 282 -926
rect 336 -620 370 -586
rect 336 -688 370 -654
rect 336 -756 370 -722
rect 336 -824 370 -790
rect 336 -892 370 -858
rect 336 -960 370 -926
rect 424 -620 458 -586
rect 424 -688 458 -654
rect 424 -756 458 -722
rect 424 -824 458 -790
rect 424 -892 458 -858
rect 424 -960 458 -926
rect 512 -620 546 -586
rect 512 -688 546 -654
rect 512 -756 546 -722
rect 512 -824 546 -790
rect 512 -892 546 -858
rect 512 -960 546 -926
rect 600 -620 634 -586
rect 600 -688 634 -654
rect 600 -756 634 -722
rect 600 -824 634 -790
rect 600 -892 634 -858
rect 600 -960 634 -926
rect 688 -620 722 -586
rect 688 -688 722 -654
rect 688 -756 722 -722
rect 688 -824 722 -790
rect 688 -892 722 -858
rect 688 -960 722 -926
rect 776 -620 810 -586
rect 776 -688 810 -654
rect 776 -756 810 -722
rect 776 -824 810 -790
rect 776 -892 810 -858
rect 776 -960 810 -926
rect 864 -620 898 -586
rect 864 -688 898 -654
rect 864 -756 898 -722
rect 864 -824 898 -790
rect 864 -892 898 -858
rect 864 -960 898 -926
rect -16 -1137 18 -1103
rect 72 -1137 106 -1103
rect 160 -1137 194 -1103
rect 248 -1137 282 -1103
rect 336 -1137 370 -1103
rect 424 -1137 458 -1103
rect 512 -1137 546 -1103
rect 600 -1137 634 -1103
rect 688 -1137 722 -1103
rect 776 -1137 810 -1103
rect 864 -1137 898 -1103
rect 1475 -835 1509 -801
rect 1475 -903 1509 -869
rect 1475 -971 1509 -937
rect 1475 -1039 1509 -1005
rect 1475 -1107 1509 -1073
rect 1475 -1175 1509 -1141
rect 1567 -835 1601 -801
rect 1567 -903 1601 -869
rect 1567 -971 1601 -937
rect 1567 -1039 1601 -1005
rect 1567 -1107 1601 -1073
rect 1567 -1175 1601 -1141
rect 1663 -835 1697 -801
rect 1663 -903 1697 -869
rect 1663 -971 1697 -937
rect 1663 -1039 1697 -1005
rect 1663 -1107 1697 -1073
rect 1663 -1175 1697 -1141
rect 1759 -835 1793 -801
rect 1759 -903 1793 -869
rect 1759 -971 1793 -937
rect 1759 -1039 1793 -1005
rect 1759 -1107 1793 -1073
rect 1759 -1175 1793 -1141
rect 1855 -835 1889 -801
rect 1855 -903 1889 -869
rect 1855 -971 1889 -937
rect 1855 -1039 1889 -1005
rect 1855 -1107 1889 -1073
rect 1855 -1175 1889 -1141
rect 1951 -835 1985 -801
rect 1951 -903 1985 -869
rect 1951 -971 1985 -937
rect 1951 -1039 1985 -1005
rect 1951 -1107 1985 -1073
rect 1951 -1175 1985 -1141
rect 2043 -835 2077 -801
rect 2043 -903 2077 -869
rect 2043 -971 2077 -937
rect 2043 -1039 2077 -1005
rect 2043 -1107 2077 -1073
rect 2043 -1175 2077 -1141
<< pdiffc >>
rect 1102 5 1136 39
rect 1102 -63 1136 -29
rect 1102 -131 1136 -97
rect 1102 -199 1136 -165
rect -38 -310 -4 -276
rect 54 -310 88 -276
rect 148 -310 182 -276
rect 240 -310 274 -276
rect 332 -310 366 -276
rect 424 -310 458 -276
rect 516 -310 550 -276
rect 608 -310 642 -276
rect 700 -310 734 -276
rect 794 -310 828 -276
rect 886 -310 920 -276
rect 1102 -267 1136 -233
rect 1102 -335 1136 -301
rect 1190 5 1224 39
rect 1190 -63 1224 -29
rect 1190 -131 1224 -97
rect 1190 -199 1224 -165
rect 1190 -267 1224 -233
rect 1190 -335 1224 -301
rect 1278 5 1312 39
rect 1278 -63 1312 -29
rect 1278 -131 1312 -97
rect 1278 -199 1312 -165
rect 1278 -267 1312 -233
rect 1278 -335 1312 -301
rect 1366 5 1400 39
rect 1366 -63 1400 -29
rect 1366 -131 1400 -97
rect 1366 -199 1400 -165
rect 1366 -267 1400 -233
rect 1366 -335 1400 -301
rect 1454 5 1488 39
rect 1454 -63 1488 -29
rect 1454 -131 1488 -97
rect 1454 -199 1488 -165
rect 1454 -267 1488 -233
rect 1454 -335 1488 -301
rect 1542 5 1576 39
rect 1542 -63 1576 -29
rect 1542 -131 1576 -97
rect 1542 -199 1576 -165
rect 1542 -267 1576 -233
rect 1542 -335 1576 -301
rect 1630 5 1664 39
rect 1630 -63 1664 -29
rect 1630 -131 1664 -97
rect 1630 -199 1664 -165
rect 1630 -267 1664 -233
rect 1630 -335 1664 -301
rect 1889 5 1923 39
rect 1889 -63 1923 -29
rect 1889 -131 1923 -97
rect 1889 -199 1923 -165
rect 1889 -267 1923 -233
rect 1889 -335 1923 -301
rect 1977 5 2011 39
rect 1977 -63 2011 -29
rect 1977 -131 2011 -97
rect 1977 -199 2011 -165
rect 1977 -267 2011 -233
rect 1977 -335 2011 -301
rect 2065 5 2099 39
rect 2065 -63 2099 -29
rect 2065 -131 2099 -97
rect 2065 -199 2099 -165
rect 2065 -267 2099 -233
rect 2065 -335 2099 -301
rect 2153 5 2187 39
rect 2153 -63 2187 -29
rect 2153 -131 2187 -97
rect 2153 -199 2187 -165
rect 2153 -267 2187 -233
rect 2153 -335 2187 -301
rect 2241 5 2275 39
rect 2241 -63 2275 -29
rect 2241 -131 2275 -97
rect 2241 -199 2275 -165
rect 2241 -267 2275 -233
rect 2241 -335 2275 -301
rect 2329 5 2363 39
rect 2329 -63 2363 -29
rect 2329 -131 2363 -97
rect 2329 -199 2363 -165
rect 2329 -267 2363 -233
rect 2329 -335 2363 -301
rect 2417 5 2451 39
rect 2417 -63 2451 -29
rect 2417 -131 2451 -97
rect 2417 -199 2451 -165
rect 2417 -267 2451 -233
rect 2417 -335 2451 -301
<< psubdiff >>
rect -286 2142 -164 2188
rect -286 2108 -242 2142
rect -208 2108 -164 2142
rect -286 2064 -164 2108
rect 262 2142 384 2188
rect 262 2108 306 2142
rect 340 2108 384 2142
rect 262 2064 384 2108
rect 810 2142 932 2188
rect 810 2108 854 2142
rect 888 2108 932 2142
rect 810 2064 932 2108
rect 1358 2142 1480 2188
rect 1358 2108 1402 2142
rect 1436 2108 1480 2142
rect 1358 2064 1480 2108
rect 1906 2142 2028 2188
rect 1906 2108 1950 2142
rect 1984 2108 2028 2142
rect 1906 2064 2028 2108
rect 2436 2142 2558 2188
rect 2436 2108 2480 2142
rect 2514 2108 2558 2142
rect 2436 2064 2558 2108
rect 2984 2142 3106 2188
rect 2984 2108 3028 2142
rect 3062 2108 3106 2142
rect 2984 2064 3106 2108
rect 3534 2142 3656 2188
rect 3534 2108 3578 2142
rect 3612 2108 3656 2142
rect 3534 2064 3656 2108
rect -652 2000 -530 2046
rect -652 1966 -608 2000
rect -574 1966 -530 2000
rect -652 1922 -530 1966
rect 4353 1930 4475 1976
rect 4353 1896 4397 1930
rect 4431 1896 4475 1930
rect 4353 1852 4475 1896
rect -652 1526 -530 1572
rect -652 1492 -608 1526
rect -574 1492 -530 1526
rect -652 1448 -530 1492
rect 4353 1454 4475 1500
rect 4353 1420 4397 1454
rect 4431 1420 4475 1454
rect 4353 1376 4475 1420
rect -652 1052 -530 1098
rect -652 1018 -608 1052
rect -574 1018 -530 1052
rect -652 974 -530 1018
rect 4353 980 4475 1026
rect 4353 946 4397 980
rect 4431 946 4475 980
rect 4353 902 4475 946
rect -652 578 -530 624
rect -652 544 -608 578
rect -574 544 -530 578
rect -652 500 -530 544
rect 4351 506 4473 552
rect 4351 472 4395 506
rect 4429 472 4473 506
rect 4351 434 4473 472
rect -116 -643 -82 -569
rect -116 -712 -82 -677
rect -116 -781 -82 -746
rect -116 -850 -82 -815
rect -116 -919 -82 -884
rect -116 -988 -82 -953
rect 964 -633 998 -569
rect 4351 -580 4473 -534
rect 4351 -614 4395 -580
rect 4429 -614 4473 -580
rect 964 -702 998 -667
rect 964 -771 998 -736
rect 4351 -658 4473 -614
rect 964 -840 998 -805
rect 964 -909 998 -874
rect 964 -978 998 -943
rect -116 -1057 -82 -1022
rect 964 -1047 998 -1012
rect -116 -1126 -82 -1091
rect -116 -1195 -82 -1160
rect 964 -1116 998 -1081
rect -116 -1264 -82 -1229
rect 964 -1185 998 -1150
rect 964 -1254 998 -1219
rect -116 -1326 -82 -1298
rect 964 -1326 998 -1288
rect 1375 -844 1409 -809
rect 1375 -913 1409 -878
rect 1375 -982 1409 -947
rect 1375 -1051 1409 -1016
rect 1375 -1120 1409 -1085
rect 1375 -1189 1409 -1154
rect 2143 -844 2177 -809
rect 2143 -913 2177 -878
rect 2143 -982 2177 -947
rect 2143 -1051 2177 -1016
rect 2143 -1120 2177 -1085
rect 4351 -1054 4473 -1008
rect 4351 -1088 4395 -1054
rect 4429 -1088 4473 -1054
rect 4351 -1132 4473 -1088
rect 1375 -1258 1409 -1223
rect 2143 -1189 2177 -1154
rect 2143 -1258 2177 -1223
rect 1375 -1326 1409 -1292
rect 2143 -1326 2177 -1292
rect -116 -1327 2193 -1326
rect -116 -1333 1122 -1327
rect -116 -1367 101 -1333
rect 135 -1367 219 -1333
rect 253 -1367 337 -1333
rect 371 -1367 455 -1333
rect 489 -1367 573 -1333
rect 607 -1367 691 -1333
rect 725 -1367 809 -1333
rect 843 -1361 1122 -1333
rect 1156 -1361 1214 -1327
rect 1248 -1361 1306 -1327
rect 1340 -1361 1398 -1327
rect 1432 -1361 1490 -1327
rect 1524 -1361 1582 -1327
rect 1616 -1361 1674 -1327
rect 1708 -1361 1770 -1327
rect 1804 -1361 1858 -1327
rect 1892 -1361 1950 -1327
rect 1984 -1361 2042 -1327
rect 2076 -1361 2134 -1327
rect 2168 -1361 2193 -1327
rect 843 -1367 2193 -1361
rect -116 -1372 2193 -1367
rect -646 -1760 -524 -1714
rect -646 -1794 -602 -1760
rect -568 -1794 -524 -1760
rect -646 -1838 -524 -1794
rect 4351 -1790 4473 -1744
rect 4351 -1824 4395 -1790
rect 4429 -1824 4473 -1790
rect 4351 -1868 4473 -1824
rect -646 -2234 -524 -2188
rect -646 -2268 -602 -2234
rect -568 -2268 -524 -2234
rect -646 -2312 -524 -2268
rect 4351 -2264 4473 -2218
rect 4351 -2298 4395 -2264
rect 4429 -2298 4473 -2264
rect 4351 -2342 4473 -2298
rect -646 -2708 -524 -2662
rect -646 -2742 -602 -2708
rect -568 -2742 -524 -2708
rect -646 -2786 -524 -2742
rect 4351 -2738 4473 -2692
rect 4351 -2772 4395 -2738
rect 4429 -2772 4473 -2738
rect 4351 -2816 4473 -2772
rect -116 -3268 6 -3222
rect -116 -3302 -72 -3268
rect -38 -3302 6 -3268
rect -116 -3346 6 -3302
rect 432 -3268 554 -3222
rect 432 -3302 476 -3268
rect 510 -3302 554 -3268
rect 432 -3346 554 -3302
rect 980 -3268 1102 -3222
rect 980 -3302 1024 -3268
rect 1058 -3302 1102 -3268
rect 980 -3346 1102 -3302
rect 1528 -3268 1650 -3222
rect 1528 -3302 1572 -3268
rect 1606 -3302 1650 -3268
rect 1528 -3346 1650 -3302
rect 2076 -3268 2198 -3222
rect 2076 -3302 2120 -3268
rect 2154 -3302 2198 -3268
rect 2076 -3346 2198 -3302
rect 2624 -3268 2746 -3222
rect 2624 -3302 2668 -3268
rect 2702 -3302 2746 -3268
rect 2624 -3346 2746 -3302
rect 3174 -3268 3296 -3222
rect 3174 -3302 3218 -3268
rect 3252 -3302 3296 -3268
rect 3174 -3346 3296 -3302
<< nsubdiff >>
rect 935 226 3068 234
rect 935 210 1084 226
rect 935 176 939 210
rect 973 192 1084 210
rect 1118 192 1168 226
rect 1202 192 1252 226
rect 1286 192 1336 226
rect 1370 192 1420 226
rect 1454 192 1504 226
rect 1538 192 1588 226
rect 1622 192 1672 226
rect 1706 192 1840 226
rect 1874 192 1924 226
rect 1958 192 2008 226
rect 2042 192 2080 226
rect 2114 192 2164 226
rect 2198 192 2248 226
rect 2282 192 2320 226
rect 2354 192 2404 226
rect 2438 192 2476 226
rect 2510 192 2632 226
rect 2666 192 3068 226
rect 973 186 3068 192
rect 973 176 980 186
rect 935 127 980 176
rect 935 93 939 127
rect 973 93 980 127
rect 935 44 980 93
rect 1753 127 1799 186
rect 1753 93 1759 127
rect 1793 93 1799 127
rect 935 10 939 44
rect 973 10 980 44
rect 935 -39 980 10
rect 935 -73 939 -39
rect 973 -73 980 -39
rect 935 -122 980 -73
rect -640 -130 980 -122
rect -640 -164 -600 -130
rect -566 -164 -444 -130
rect -410 -164 -290 -130
rect -256 -164 -146 -130
rect -112 -164 -32 -130
rect 2 -164 82 -130
rect 116 -164 166 -130
rect 200 -164 250 -130
rect 284 -164 334 -130
rect 368 -164 418 -130
rect 452 -164 502 -130
rect 536 -164 586 -130
rect 620 -164 670 -130
rect 704 -164 754 -130
rect 788 -164 838 -130
rect 872 -164 922 -130
rect 956 -164 980 -130
rect -640 -177 980 -164
rect 1753 44 1799 93
rect 2573 127 2619 186
rect 2573 93 2579 127
rect 2613 93 2619 127
rect 1753 10 1759 44
rect 1793 10 1799 44
rect 1753 -39 1799 10
rect 1753 -73 1759 -39
rect 1793 -73 1799 -39
rect 1753 -127 1799 -73
rect 1753 -161 1759 -127
rect 1793 -161 1799 -127
rect 1753 -210 1799 -161
rect 1753 -244 1759 -210
rect 1793 -244 1799 -210
rect 1753 -293 1799 -244
rect 1753 -327 1759 -293
rect 1793 -327 1799 -293
rect 1753 -370 1799 -327
rect 2573 44 2619 93
rect 2573 10 2579 44
rect 2613 10 2619 44
rect 2573 -39 2619 10
rect 2573 -73 2579 -39
rect 2613 -73 2619 -39
rect 2573 -122 2619 -73
rect 2573 -156 2579 -122
rect 2613 -156 2619 -122
rect 2573 -191 2619 -156
rect 2787 -1240 2825 -1238
rect 2787 -1274 2789 -1240
rect 2823 -1274 2825 -1240
rect 2787 -1276 2825 -1274
rect 2863 -1240 2901 -1238
rect 2863 -1274 2865 -1240
rect 2899 -1274 2901 -1240
rect 2863 -1276 2901 -1274
rect 2939 -1240 2977 -1238
rect 2939 -1274 2941 -1240
rect 2975 -1274 2977 -1240
rect 2939 -1276 2977 -1274
rect 3015 -1240 3053 -1238
rect 3015 -1274 3017 -1240
rect 3051 -1274 3053 -1240
rect 3015 -1276 3053 -1274
rect 3180 -1240 3830 -1238
rect 3180 -1274 3206 -1240
rect 3240 -1274 3282 -1240
rect 3316 -1274 3358 -1240
rect 3392 -1274 3434 -1240
rect 3468 -1274 3510 -1240
rect 3544 -1274 3586 -1240
rect 3620 -1274 3662 -1240
rect 3696 -1274 3738 -1240
rect 3772 -1274 3830 -1240
rect 3180 -1276 3830 -1274
<< psubdiffcont >>
rect -242 2108 -208 2142
rect 306 2108 340 2142
rect 854 2108 888 2142
rect 1402 2108 1436 2142
rect 1950 2108 1984 2142
rect 2480 2108 2514 2142
rect 3028 2108 3062 2142
rect 3578 2108 3612 2142
rect -608 1966 -574 2000
rect 4397 1896 4431 1930
rect -608 1492 -574 1526
rect 4397 1420 4431 1454
rect -608 1018 -574 1052
rect 4397 946 4431 980
rect -608 544 -574 578
rect 4395 472 4429 506
rect -116 -677 -82 -643
rect -116 -746 -82 -712
rect -116 -815 -82 -781
rect -116 -884 -82 -850
rect -116 -953 -82 -919
rect 4395 -614 4429 -580
rect 964 -667 998 -633
rect 964 -736 998 -702
rect 964 -805 998 -771
rect 964 -874 998 -840
rect 964 -943 998 -909
rect -116 -1022 -82 -988
rect 964 -1012 998 -978
rect -116 -1091 -82 -1057
rect -116 -1160 -82 -1126
rect 964 -1081 998 -1047
rect 964 -1150 998 -1116
rect -116 -1229 -82 -1195
rect -116 -1298 -82 -1264
rect 964 -1219 998 -1185
rect 964 -1288 998 -1254
rect 1375 -878 1409 -844
rect 1375 -947 1409 -913
rect 1375 -1016 1409 -982
rect 1375 -1085 1409 -1051
rect 1375 -1154 1409 -1120
rect 2143 -878 2177 -844
rect 2143 -947 2177 -913
rect 2143 -1016 2177 -982
rect 2143 -1085 2177 -1051
rect 2143 -1154 2177 -1120
rect 4395 -1088 4429 -1054
rect 1375 -1223 1409 -1189
rect 2143 -1223 2177 -1189
rect 1375 -1292 1409 -1258
rect 2143 -1292 2177 -1258
rect 101 -1367 135 -1333
rect 219 -1367 253 -1333
rect 337 -1367 371 -1333
rect 455 -1367 489 -1333
rect 573 -1367 607 -1333
rect 691 -1367 725 -1333
rect 809 -1367 843 -1333
rect 1122 -1361 1156 -1327
rect 1214 -1361 1248 -1327
rect 1306 -1361 1340 -1327
rect 1398 -1361 1432 -1327
rect 1490 -1361 1524 -1327
rect 1582 -1361 1616 -1327
rect 1674 -1361 1708 -1327
rect 1770 -1361 1804 -1327
rect 1858 -1361 1892 -1327
rect 1950 -1361 1984 -1327
rect 2042 -1361 2076 -1327
rect 2134 -1361 2168 -1327
rect -602 -1794 -568 -1760
rect 4395 -1824 4429 -1790
rect -602 -2268 -568 -2234
rect 4395 -2298 4429 -2264
rect -602 -2742 -568 -2708
rect 4395 -2772 4429 -2738
rect -72 -3302 -38 -3268
rect 476 -3302 510 -3268
rect 1024 -3302 1058 -3268
rect 1572 -3302 1606 -3268
rect 2120 -3302 2154 -3268
rect 2668 -3302 2702 -3268
rect 3218 -3302 3252 -3268
<< nsubdiffcont >>
rect 939 176 973 210
rect 1084 192 1118 226
rect 1168 192 1202 226
rect 1252 192 1286 226
rect 1336 192 1370 226
rect 1420 192 1454 226
rect 1504 192 1538 226
rect 1588 192 1622 226
rect 1672 192 1706 226
rect 1840 192 1874 226
rect 1924 192 1958 226
rect 2008 192 2042 226
rect 2080 192 2114 226
rect 2164 192 2198 226
rect 2248 192 2282 226
rect 2320 192 2354 226
rect 2404 192 2438 226
rect 2476 192 2510 226
rect 2632 192 2666 226
rect 939 93 973 127
rect 1759 93 1793 127
rect 939 10 973 44
rect 939 -73 973 -39
rect -600 -164 -566 -130
rect -444 -164 -410 -130
rect -290 -164 -256 -130
rect -146 -164 -112 -130
rect -32 -164 2 -130
rect 82 -164 116 -130
rect 166 -164 200 -130
rect 250 -164 284 -130
rect 334 -164 368 -130
rect 418 -164 452 -130
rect 502 -164 536 -130
rect 586 -164 620 -130
rect 670 -164 704 -130
rect 754 -164 788 -130
rect 838 -164 872 -130
rect 922 -164 956 -130
rect 2579 93 2613 127
rect 1759 10 1793 44
rect 1759 -73 1793 -39
rect 1759 -161 1793 -127
rect 1759 -244 1793 -210
rect 1759 -327 1793 -293
rect 2579 10 2613 44
rect 2579 -73 2613 -39
rect 2579 -156 2613 -122
rect 2789 -1274 2823 -1240
rect 2865 -1274 2899 -1240
rect 2941 -1274 2975 -1240
rect 3017 -1274 3051 -1240
rect 3206 -1274 3240 -1240
rect 3282 -1274 3316 -1240
rect 3358 -1274 3392 -1240
rect 3434 -1274 3468 -1240
rect 3510 -1274 3544 -1240
rect 3586 -1274 3620 -1240
rect 3662 -1274 3696 -1240
rect 3738 -1274 3772 -1240
<< poly >>
rect 1148 52 1178 78
rect 1236 52 1266 78
rect 1324 52 1354 78
rect 1412 52 1442 78
rect 1500 52 1530 78
rect 1588 52 1618 78
rect 12 -243 42 -217
rect 104 -243 134 -217
rect 196 -243 226 -217
rect 288 -243 318 -217
rect 380 -243 410 -217
rect 472 -243 502 -217
rect 564 -243 594 -217
rect 656 -243 686 -217
rect 748 -243 778 -217
rect 840 -243 870 -217
rect 12 -369 42 -343
rect 104 -369 134 -343
rect 196 -369 226 -343
rect 288 -369 318 -343
rect 380 -369 410 -343
rect 12 -393 410 -369
rect 12 -427 28 -393
rect 62 -399 410 -393
rect 472 -369 502 -343
rect 564 -369 594 -343
rect 656 -369 686 -343
rect 748 -369 778 -343
rect 840 -369 870 -343
rect 1935 52 1965 78
rect 2023 52 2053 78
rect 2111 52 2141 78
rect 2199 52 2229 78
rect 2287 52 2317 78
rect 2375 52 2405 78
rect 472 -393 870 -369
rect 472 -399 813 -393
rect 62 -427 80 -399
rect 12 -446 80 -427
rect 797 -427 813 -399
rect 847 -399 870 -393
rect 1148 -374 1178 -348
rect 1236 -374 1266 -348
rect 1324 -374 1354 -348
rect 847 -427 865 -399
rect 1148 -402 1354 -374
rect 1148 -404 1191 -402
rect 797 -446 865 -427
rect 1174 -436 1191 -404
rect 1225 -404 1354 -402
rect 1412 -374 1442 -348
rect 1500 -374 1530 -348
rect 1588 -374 1618 -348
rect 1412 -404 1618 -374
rect 1225 -436 1244 -404
rect 1174 -446 1244 -436
rect 1530 -413 1618 -404
rect 1530 -447 1558 -413
rect 1592 -447 1618 -413
rect 1530 -463 1618 -447
rect 1935 -374 1965 -348
rect 2023 -374 2053 -348
rect 2111 -374 2141 -348
rect 1935 -404 2141 -374
rect 2199 -374 2229 -348
rect 2287 -370 2317 -348
rect 2375 -370 2405 -348
rect 2287 -374 2405 -370
rect 2199 -402 2405 -374
rect 2199 -404 2329 -402
rect 1935 -413 2023 -404
rect 1935 -447 1963 -413
rect 1997 -447 2023 -413
rect 2313 -436 2329 -404
rect 2363 -404 2405 -402
rect 2363 -436 2379 -404
rect 2313 -446 2379 -436
rect 1935 -463 2023 -447
rect 180 -492 260 -482
rect 180 -516 203 -492
rect 30 -526 203 -516
rect 237 -516 260 -492
rect 622 -490 702 -480
rect 622 -514 645 -490
rect 237 -526 412 -516
rect 30 -547 412 -526
rect 30 -573 60 -547
rect 118 -573 148 -547
rect 206 -573 236 -547
rect 294 -573 324 -547
rect 382 -573 412 -547
rect 470 -524 645 -514
rect 679 -514 702 -490
rect 679 -524 852 -514
rect 470 -545 852 -524
rect 470 -573 500 -545
rect 558 -573 588 -545
rect 646 -573 676 -545
rect 734 -573 764 -545
rect 822 -573 852 -545
rect 1649 -662 1743 -624
rect 1649 -696 1677 -662
rect 1711 -696 1743 -662
rect 1649 -719 1743 -696
rect 1525 -788 1555 -762
rect 1617 -788 1647 -762
rect 1713 -788 1743 -719
rect 1809 -662 1903 -624
rect 1809 -696 1843 -662
rect 1877 -696 1903 -662
rect 1809 -719 1903 -696
rect 1809 -788 1839 -719
rect 1905 -788 1935 -762
rect 1997 -788 2027 -762
rect 30 -1001 60 -973
rect 118 -1001 148 -973
rect 206 -1001 236 -973
rect 294 -1001 324 -973
rect 382 -1001 412 -973
rect 470 -1001 500 -973
rect 558 -1001 588 -973
rect 646 -1001 676 -973
rect 734 -1001 764 -973
rect 822 -1001 852 -973
rect 30 -1070 60 -1044
rect 118 -1070 148 -1044
rect 206 -1070 236 -1044
rect 294 -1070 324 -1044
rect 382 -1070 412 -1044
rect 470 -1070 500 -1044
rect 558 -1070 588 -1044
rect 646 -1070 676 -1044
rect 734 -1070 764 -1044
rect 822 -1070 852 -1044
rect 30 -1196 60 -1170
rect 118 -1196 148 -1170
rect 30 -1238 148 -1196
rect 30 -1272 72 -1238
rect 106 -1272 148 -1238
rect 30 -1298 148 -1272
rect 206 -1196 236 -1170
rect 294 -1196 324 -1170
rect 206 -1238 324 -1196
rect 206 -1272 248 -1238
rect 282 -1272 324 -1238
rect 206 -1298 324 -1272
rect 382 -1196 412 -1170
rect 470 -1196 500 -1170
rect 382 -1238 500 -1196
rect 382 -1272 424 -1238
rect 458 -1272 500 -1238
rect 382 -1298 500 -1272
rect 558 -1196 588 -1170
rect 646 -1196 676 -1170
rect 558 -1238 676 -1196
rect 558 -1272 600 -1238
rect 634 -1272 676 -1238
rect 558 -1298 676 -1272
rect 734 -1196 764 -1170
rect 822 -1196 852 -1170
rect 734 -1238 852 -1196
rect 734 -1272 776 -1238
rect 810 -1272 852 -1238
rect 734 -1298 852 -1272
rect 1525 -1227 1555 -1188
rect 1617 -1226 1647 -1188
rect 1713 -1214 1743 -1188
rect 1809 -1214 1839 -1188
rect 1905 -1226 1935 -1188
rect 1997 -1226 2027 -1188
rect 1462 -1241 1555 -1227
rect 1462 -1275 1491 -1241
rect 1525 -1275 1555 -1241
rect 1462 -1290 1555 -1275
rect 1611 -1242 1671 -1226
rect 1611 -1276 1621 -1242
rect 1655 -1276 1671 -1242
rect 1611 -1292 1671 -1276
rect 1883 -1242 1943 -1226
rect 1883 -1276 1893 -1242
rect 1927 -1276 1943 -1242
rect 1883 -1292 1943 -1276
rect 1997 -1240 2090 -1226
rect 1997 -1274 2026 -1240
rect 2060 -1274 2090 -1240
rect 1997 -1289 2090 -1274
<< polycont >>
rect 28 -427 62 -393
rect 813 -427 847 -393
rect 1191 -436 1225 -402
rect 1558 -447 1592 -413
rect 1963 -447 1997 -413
rect 2329 -436 2363 -402
rect 203 -526 237 -492
rect 645 -524 679 -490
rect 1677 -696 1711 -662
rect 1843 -696 1877 -662
rect 72 -1272 106 -1238
rect 248 -1272 282 -1238
rect 424 -1272 458 -1238
rect 600 -1272 634 -1238
rect 776 -1272 810 -1238
rect 1491 -1275 1525 -1241
rect 1621 -1276 1655 -1242
rect 1893 -1276 1927 -1242
rect 2026 -1274 2060 -1240
<< locali >>
rect -686 2142 4515 2218
rect -686 2108 -242 2142
rect -208 2108 306 2142
rect 340 2108 854 2142
rect 888 2108 1402 2142
rect 1436 2108 1950 2142
rect 1984 2108 2480 2142
rect 2514 2108 3028 2142
rect 3062 2108 3578 2142
rect 3612 2108 4515 2142
rect -686 2020 4515 2108
rect -686 2000 -450 2020
rect 200 2000 660 2020
rect 2780 2000 3240 2020
rect -686 1967 -608 2000
rect -574 1967 -450 2000
rect -686 1573 -638 1967
rect -532 1573 -450 1967
rect -686 1530 -450 1573
rect 4317 1930 4515 2020
rect 4317 1896 4397 1930
rect 4431 1896 4515 1930
rect -686 1526 -488 1530
rect -686 1492 -608 1526
rect -574 1492 -488 1526
rect -686 1407 -488 1492
rect -686 1013 -651 1407
rect -545 1013 -488 1407
rect 4317 1454 4515 1896
rect 4317 1420 4397 1454
rect 4431 1420 4515 1454
rect 4048 1225 4147 1260
rect 4048 1191 4080 1225
rect 4114 1191 4147 1225
rect 4048 1156 4147 1191
rect -686 852 -488 1013
rect -686 458 -641 852
rect -535 458 -488 852
rect -686 420 -488 458
rect 4317 980 4515 1420
rect 4317 946 4397 980
rect 4431 946 4515 980
rect 4317 506 4515 946
rect 4317 472 4395 506
rect 4429 472 4515 506
rect 935 227 4179 234
rect 935 226 3299 227
rect 935 210 1084 226
rect 935 176 939 210
rect 973 192 1084 210
rect 1118 192 1168 226
rect 1202 192 1252 226
rect 1286 192 1336 226
rect 1370 192 1420 226
rect 1454 192 1504 226
rect 1538 192 1588 226
rect 1622 192 1672 226
rect 1706 192 1840 226
rect 1874 192 1924 226
rect 1958 192 2008 226
rect 2042 192 2080 226
rect 2114 192 2164 226
rect 2198 192 2248 226
rect 2282 192 2320 226
rect 2354 192 2404 226
rect 2438 192 2476 226
rect 2510 192 2632 226
rect 2666 192 2716 226
rect 2750 192 2788 226
rect 2822 192 2917 226
rect 2951 192 2989 226
rect 3023 193 3299 226
rect 3333 193 3371 227
rect 3405 193 3443 227
rect 3477 193 3515 227
rect 3549 193 3587 227
rect 3621 193 3659 227
rect 3693 193 3732 227
rect 3766 193 3804 227
rect 3838 193 3876 227
rect 3910 193 3948 227
rect 3982 193 4020 227
rect 4054 193 4092 227
rect 4126 193 4179 227
rect 3023 192 4179 193
rect 973 186 4179 192
rect 973 176 980 186
rect 935 127 980 176
rect 935 93 939 127
rect 973 93 980 127
rect 935 44 980 93
rect 1753 127 1799 186
rect 1753 93 1759 127
rect 1793 93 1799 127
rect 935 10 939 44
rect 973 10 980 44
rect 935 -39 980 10
rect 935 -73 939 -39
rect 973 -73 980 -39
rect 935 -122 980 -73
rect -640 -130 980 -122
rect -640 -164 -600 -130
rect -566 -164 -444 -130
rect -410 -164 -290 -130
rect -256 -164 -146 -130
rect -112 -164 -32 -130
rect 2 -164 82 -130
rect 116 -164 166 -130
rect 200 -164 250 -130
rect 284 -164 334 -130
rect 368 -164 418 -130
rect 452 -164 502 -130
rect 536 -164 586 -130
rect 620 -164 670 -130
rect 704 -164 754 -130
rect 788 -164 838 -130
rect 872 -164 922 -130
rect 956 -164 980 -130
rect -640 -177 980 -164
rect 1102 39 1136 56
rect 1102 -29 1136 5
rect 1102 -97 1136 -70
rect 1102 -165 1136 -131
rect 1102 -233 1136 -199
rect -38 -276 -4 -239
rect -38 -347 -4 -310
rect 54 -276 88 -239
rect 54 -347 88 -310
rect 148 -276 182 -239
rect 148 -347 182 -327
rect 240 -276 274 -239
rect 240 -347 274 -310
rect 332 -276 366 -239
rect 332 -347 366 -327
rect 424 -276 458 -239
rect 424 -347 458 -310
rect 516 -276 550 -239
rect 516 -347 550 -327
rect 608 -276 642 -239
rect 608 -347 642 -310
rect 700 -276 734 -239
rect 700 -347 734 -327
rect 794 -276 828 -239
rect 794 -347 828 -310
rect 886 -276 920 -239
rect 886 -347 920 -310
rect 1102 -301 1136 -267
rect 1102 -352 1136 -335
rect 1190 39 1224 56
rect 1190 -29 1224 5
rect 1190 -97 1224 -70
rect 1190 -165 1224 -131
rect 1190 -233 1224 -199
rect 1190 -301 1224 -267
rect 1190 -352 1224 -335
rect 1278 39 1312 56
rect 1278 -29 1312 5
rect 1278 -97 1312 -63
rect 1278 -165 1312 -131
rect 1278 -233 1312 -199
rect 1278 -268 1312 -267
rect 1278 -352 1312 -335
rect 1366 39 1400 56
rect 1366 -29 1400 5
rect 1366 -97 1400 -70
rect 1366 -165 1400 -131
rect 1366 -233 1400 -199
rect 1366 -301 1400 -267
rect 1366 -352 1400 -335
rect 1454 39 1488 56
rect 1454 -29 1488 3
rect 1454 -97 1488 -63
rect 1454 -165 1488 -131
rect 1454 -233 1488 -199
rect 1454 -301 1488 -267
rect 1454 -352 1488 -335
rect 1542 39 1576 56
rect 1542 -29 1576 5
rect 1542 -97 1576 -70
rect 1542 -165 1576 -131
rect 1542 -233 1576 -199
rect 1542 -301 1576 -267
rect 1542 -352 1576 -335
rect 1630 39 1664 56
rect 1630 -29 1664 5
rect 1630 -97 1664 -70
rect 1630 -165 1664 -131
rect 1630 -233 1664 -199
rect 1630 -301 1664 -267
rect 1630 -352 1664 -335
rect 1753 44 1799 93
rect 2573 127 2619 186
rect 2573 93 2579 127
rect 2613 93 2619 127
rect 1753 10 1759 44
rect 1793 10 1799 44
rect 1753 -39 1799 10
rect 1753 -73 1759 -39
rect 1793 -73 1799 -39
rect 1753 -127 1799 -73
rect 1753 -161 1759 -127
rect 1793 -161 1799 -127
rect 1753 -210 1799 -161
rect 1753 -244 1759 -210
rect 1793 -244 1799 -210
rect 1753 -293 1799 -244
rect 1753 -327 1759 -293
rect 1793 -327 1799 -293
rect 6 -393 85 -389
rect 6 -427 28 -393
rect 62 -427 85 -393
rect 6 -431 85 -427
rect 791 -393 870 -390
rect 791 -427 813 -393
rect 847 -427 870 -393
rect 791 -430 870 -427
rect 1174 -402 1244 -386
rect 1174 -436 1191 -402
rect 1225 -436 1244 -402
rect 1174 -446 1244 -436
rect 1530 -413 1618 -397
rect 1753 -413 1799 -327
rect 1889 39 1923 56
rect 1889 -29 1923 5
rect 1889 -97 1923 -70
rect 1889 -165 1923 -131
rect 1889 -233 1923 -199
rect 1889 -301 1923 -267
rect 1889 -352 1923 -335
rect 1977 39 2011 56
rect 1977 -29 2011 5
rect 1977 -97 2011 -70
rect 1977 -165 2011 -131
rect 1977 -233 2011 -199
rect 1977 -301 2011 -267
rect 1977 -352 2011 -335
rect 2065 39 2099 56
rect 2065 -29 2099 0
rect 2065 -97 2099 -63
rect 2065 -165 2099 -131
rect 2065 -233 2099 -199
rect 2065 -301 2099 -267
rect 2065 -352 2099 -335
rect 2153 39 2187 56
rect 2153 -29 2187 5
rect 2153 -97 2187 -70
rect 2153 -165 2187 -131
rect 2153 -233 2187 -199
rect 2153 -301 2187 -267
rect 2153 -352 2187 -335
rect 2241 39 2275 56
rect 2241 -29 2275 5
rect 2241 -97 2275 -63
rect 2241 -165 2275 -131
rect 2241 -233 2275 -199
rect 2241 -268 2275 -267
rect 2241 -352 2275 -335
rect 2329 39 2363 56
rect 2329 -29 2363 5
rect 2329 -97 2363 -70
rect 2329 -165 2363 -131
rect 2329 -233 2363 -199
rect 2329 -301 2363 -267
rect 2329 -352 2363 -335
rect 2417 39 2451 56
rect 2417 -29 2451 5
rect 2417 -97 2451 -70
rect 2417 -165 2451 -131
rect 2573 44 2619 93
rect 2573 10 2579 44
rect 2613 10 2619 44
rect 2573 -39 2619 10
rect 2573 -73 2579 -39
rect 2613 -73 2619 -39
rect 2573 -122 2619 -73
rect 2573 -156 2579 -122
rect 2613 -156 2619 -122
rect 2573 -191 2619 -156
rect 2417 -233 2451 -199
rect 2417 -301 2451 -267
rect 2417 -352 2451 -335
rect 3429 -358 3803 -314
rect 3429 -359 3633 -358
rect 1935 -413 2023 -397
rect 1182 -448 1226 -446
rect 1530 -447 1558 -413
rect 1592 -447 1618 -413
rect 1530 -463 1618 -447
rect 1935 -447 1963 -413
rect 1997 -447 2023 -413
rect 2313 -402 2379 -386
rect 2313 -436 2329 -402
rect 2363 -436 2379 -402
rect 3429 -393 3463 -359
rect 3497 -393 3549 -359
rect 3583 -392 3633 -359
rect 3667 -359 3803 -358
rect 3667 -392 3717 -359
rect 3583 -393 3717 -392
rect 3751 -393 3803 -359
rect 3429 -436 3803 -393
rect 2313 -446 2379 -436
rect 1935 -463 2023 -447
rect 2325 -448 2367 -446
rect 180 -492 260 -482
rect 180 -526 203 -492
rect 237 -526 260 -492
rect 180 -533 260 -526
rect 622 -490 702 -480
rect 622 -524 645 -490
rect 679 -524 702 -490
rect 622 -531 702 -524
rect 2695 -509 3119 -462
rect 2695 -510 2806 -509
rect 2695 -544 2721 -510
rect 2755 -543 2806 -510
rect 2840 -510 2978 -509
rect 2840 -543 2890 -510
rect 2755 -544 2890 -543
rect 2924 -543 2978 -510
rect 3012 -543 3061 -509
rect 3095 -543 3119 -509
rect 2924 -544 3119 -543
rect -116 -643 -74 -569
rect -82 -677 -74 -643
rect -116 -712 -74 -677
rect -82 -746 -74 -712
rect -116 -781 -74 -746
rect -82 -815 -74 -781
rect -116 -850 -74 -815
rect -82 -884 -74 -850
rect -116 -919 -74 -884
rect -82 -953 -74 -919
rect -116 -988 -74 -953
rect -16 -586 18 -569
rect -16 -654 18 -620
rect -16 -722 18 -688
rect -16 -790 18 -756
rect -16 -858 18 -824
rect -16 -914 18 -892
rect -16 -977 18 -960
rect 72 -586 106 -569
rect 72 -654 106 -620
rect 72 -722 106 -688
rect 72 -790 106 -756
rect 72 -858 106 -824
rect 72 -914 106 -892
rect 72 -977 106 -960
rect 160 -586 194 -568
rect 160 -654 194 -620
rect 160 -722 194 -688
rect 160 -790 194 -756
rect 160 -858 194 -824
rect 160 -926 194 -892
rect 160 -977 194 -960
rect 248 -586 282 -569
rect 248 -654 282 -620
rect 248 -722 282 -688
rect 248 -790 282 -756
rect 248 -858 282 -824
rect 248 -914 282 -892
rect 248 -977 282 -960
rect 336 -585 370 -568
rect 336 -586 376 -585
rect 424 -586 458 -569
rect 512 -585 546 -568
rect 506 -586 546 -585
rect 336 -654 370 -620
rect 336 -722 370 -688
rect 336 -790 370 -756
rect 336 -858 370 -824
rect 336 -926 370 -892
rect 336 -977 370 -960
rect 424 -654 458 -620
rect 424 -722 458 -688
rect 424 -790 458 -756
rect 424 -858 458 -824
rect 424 -914 458 -892
rect 424 -977 458 -960
rect 512 -654 546 -620
rect 512 -722 546 -688
rect 512 -790 546 -756
rect 512 -858 546 -824
rect 512 -926 546 -892
rect 512 -977 546 -960
rect 600 -586 634 -569
rect 600 -654 634 -620
rect 600 -722 634 -688
rect 600 -790 634 -756
rect 600 -858 634 -824
rect 600 -914 634 -892
rect 600 -977 634 -960
rect 688 -586 722 -568
rect 688 -654 722 -620
rect 688 -722 722 -688
rect 688 -790 722 -756
rect 688 -858 722 -824
rect 688 -926 722 -892
rect 688 -977 722 -960
rect 776 -586 810 -569
rect 776 -654 810 -620
rect 776 -722 810 -688
rect 776 -790 810 -756
rect 776 -858 810 -824
rect 776 -914 810 -892
rect 776 -977 810 -960
rect 864 -586 898 -569
rect 864 -654 898 -620
rect 864 -722 898 -688
rect 864 -790 898 -756
rect 864 -858 898 -824
rect 864 -914 898 -892
rect 864 -977 898 -960
rect 956 -633 998 -569
rect 2695 -590 3119 -544
rect 4317 -580 4515 472
rect 956 -667 964 -633
rect 4317 -614 4395 -580
rect 4429 -614 4515 -580
rect 956 -702 998 -667
rect 956 -736 964 -702
rect 1654 -662 1734 -652
rect 1654 -697 1677 -662
rect 1711 -697 1734 -662
rect 1654 -707 1734 -697
rect 1820 -662 1900 -652
rect 1820 -697 1843 -662
rect 1877 -697 1900 -662
rect 1820 -707 1900 -697
rect 956 -771 998 -736
rect 956 -805 964 -771
rect 956 -840 998 -805
rect 1475 -801 1509 -784
rect 956 -874 964 -840
rect 956 -909 998 -874
rect 956 -943 964 -909
rect -82 -1022 -74 -988
rect -116 -1057 -74 -1022
rect -82 -1091 -74 -1057
rect 956 -978 998 -943
rect 956 -1012 964 -978
rect 956 -1047 998 -1012
rect -116 -1126 -74 -1091
rect -82 -1160 -74 -1126
rect -116 -1195 -74 -1160
rect -16 -1103 18 -1064
rect -16 -1174 18 -1137
rect 72 -1103 106 -1064
rect 72 -1174 106 -1137
rect 160 -1103 194 -1064
rect -82 -1229 -74 -1195
rect -116 -1264 -74 -1229
rect -82 -1298 -74 -1264
rect 52 -1238 126 -1226
rect 52 -1272 72 -1238
rect 106 -1272 126 -1238
rect 52 -1282 126 -1272
rect -116 -1316 -74 -1298
rect 160 -1316 194 -1137
rect 248 -1103 282 -1064
rect 248 -1174 282 -1137
rect 336 -1103 370 -1064
rect 228 -1238 302 -1226
rect 228 -1272 248 -1238
rect 282 -1272 302 -1238
rect 228 -1282 302 -1272
rect 336 -1316 370 -1137
rect 424 -1103 458 -1064
rect 424 -1174 458 -1137
rect 512 -1103 546 -1064
rect 404 -1238 478 -1226
rect 404 -1272 424 -1238
rect 458 -1272 478 -1238
rect 404 -1282 478 -1272
rect 512 -1316 546 -1137
rect 600 -1103 634 -1064
rect 600 -1174 634 -1137
rect 688 -1103 722 -1064
rect 580 -1238 654 -1226
rect 580 -1272 600 -1238
rect 634 -1272 654 -1238
rect 580 -1282 654 -1272
rect 688 -1316 722 -1137
rect 776 -1103 810 -1064
rect 776 -1174 810 -1137
rect 864 -1103 898 -1064
rect 864 -1174 898 -1137
rect 956 -1081 964 -1047
rect 956 -1116 998 -1081
rect 956 -1150 964 -1116
rect 956 -1185 998 -1150
rect 956 -1219 964 -1185
rect 756 -1238 830 -1226
rect 756 -1272 776 -1238
rect 810 -1272 830 -1238
rect 756 -1282 830 -1272
rect 956 -1254 998 -1219
rect 956 -1288 964 -1254
rect 956 -1316 998 -1288
rect 1375 -844 1417 -809
rect 1409 -878 1417 -844
rect 1375 -913 1417 -878
rect 1409 -947 1417 -913
rect 1375 -982 1417 -947
rect 1409 -1016 1417 -982
rect 1375 -1051 1417 -1016
rect 1409 -1085 1417 -1051
rect 1375 -1120 1417 -1085
rect 1409 -1154 1417 -1120
rect 1375 -1189 1417 -1154
rect 1409 -1223 1417 -1189
rect 1475 -869 1509 -835
rect 1475 -937 1509 -903
rect 1475 -1005 1509 -971
rect 1475 -1073 1509 -1039
rect 1475 -1137 1509 -1107
rect 1475 -1192 1509 -1175
rect 1567 -801 1601 -784
rect 1567 -869 1601 -835
rect 1567 -937 1601 -903
rect 1567 -1005 1601 -971
rect 1567 -1073 1601 -1039
rect 1567 -1137 1601 -1107
rect 1567 -1192 1601 -1175
rect 1663 -801 1697 -784
rect 1663 -869 1697 -835
rect 1663 -937 1697 -903
rect 1663 -1005 1697 -971
rect 1663 -1073 1697 -1052
rect 1663 -1141 1697 -1107
rect 1663 -1192 1697 -1175
rect 1759 -801 1793 -784
rect 1759 -869 1793 -835
rect 1759 -937 1793 -903
rect 1759 -1005 1793 -971
rect 1759 -1073 1793 -1039
rect 1759 -1137 1793 -1107
rect 1759 -1192 1793 -1175
rect 1855 -801 1889 -784
rect 1855 -869 1889 -835
rect 1855 -933 1889 -903
rect 1855 -1005 1889 -971
rect 1855 -1073 1889 -1039
rect 1855 -1141 1889 -1107
rect 1855 -1192 1889 -1175
rect 1951 -801 1985 -784
rect 1951 -869 1985 -835
rect 1951 -937 1985 -903
rect 1951 -1005 1985 -971
rect 1951 -1073 1985 -1039
rect 1951 -1137 1985 -1107
rect 1951 -1192 1985 -1175
rect 2043 -801 2077 -784
rect 2043 -869 2077 -835
rect 2043 -937 2077 -903
rect 2043 -1005 2077 -971
rect 2043 -1073 2077 -1039
rect 2043 -1137 2077 -1107
rect 2043 -1192 2077 -1175
rect 2135 -844 2177 -809
rect 2135 -878 2143 -844
rect 2135 -913 2177 -878
rect 2135 -947 2143 -913
rect 2135 -982 2177 -947
rect 2135 -1016 2143 -982
rect 2135 -1051 2177 -1016
rect 2135 -1085 2143 -1051
rect 2135 -1120 2177 -1085
rect 2135 -1154 2143 -1120
rect 2135 -1189 2177 -1154
rect 1375 -1258 1417 -1223
rect 2135 -1223 2143 -1189
rect 1409 -1292 1417 -1258
rect 1375 -1316 1417 -1292
rect -116 -1326 1417 -1316
rect 1462 -1241 1555 -1227
rect 1462 -1275 1491 -1241
rect 1525 -1275 1555 -1241
rect 1462 -1326 1555 -1275
rect 1611 -1238 1697 -1226
rect 1611 -1242 1649 -1238
rect 1611 -1276 1621 -1242
rect 1683 -1272 1697 -1238
rect 1655 -1276 1697 -1272
rect 1611 -1292 1697 -1276
rect 1857 -1238 1943 -1226
rect 1857 -1272 1871 -1238
rect 1905 -1242 1943 -1238
rect 1857 -1276 1893 -1272
rect 1927 -1276 1943 -1242
rect 1857 -1292 1943 -1276
rect 1997 -1240 2090 -1226
rect 1997 -1274 2026 -1240
rect 2060 -1274 2090 -1240
rect 1997 -1326 2090 -1274
rect 2135 -1258 2177 -1223
rect 4317 -1054 4515 -614
rect 4317 -1088 4395 -1054
rect 4429 -1088 4515 -1054
rect 4317 -1222 4515 -1088
rect 2135 -1292 2143 -1258
rect 2787 -1240 2825 -1238
rect 2787 -1274 2789 -1240
rect 2823 -1274 2825 -1240
rect 2787 -1276 2825 -1274
rect 2863 -1240 2901 -1238
rect 2863 -1274 2865 -1240
rect 2899 -1274 2901 -1240
rect 2863 -1276 2901 -1274
rect 2939 -1240 2977 -1238
rect 2939 -1274 2941 -1240
rect 2975 -1274 2977 -1240
rect 2939 -1276 2977 -1274
rect 3015 -1240 3053 -1238
rect 3015 -1274 3017 -1240
rect 3051 -1274 3053 -1240
rect 3015 -1276 3053 -1274
rect 3104 -1240 3830 -1238
rect 3104 -1274 3206 -1240
rect 3240 -1274 3282 -1240
rect 3316 -1274 3358 -1240
rect 3392 -1274 3434 -1240
rect 3468 -1274 3510 -1240
rect 3544 -1274 3586 -1240
rect 3620 -1274 3662 -1240
rect 3696 -1274 3738 -1240
rect 3772 -1274 3830 -1240
rect 3104 -1276 3830 -1274
rect 2135 -1311 2177 -1292
rect 2135 -1326 3240 -1311
rect -686 -1366 -488 -1326
rect -686 -1510 -670 -1366
rect -492 -1472 -488 -1366
rect -116 -1327 3240 -1326
rect -116 -1333 1122 -1327
rect -116 -1367 101 -1333
rect 135 -1367 219 -1333
rect 253 -1367 337 -1333
rect 371 -1367 455 -1333
rect 489 -1367 573 -1333
rect 607 -1367 691 -1333
rect 725 -1367 809 -1333
rect 843 -1367 1122 -1333
rect -116 -1375 1122 -1367
rect 1156 -1375 1214 -1327
rect 1248 -1375 1306 -1327
rect 1340 -1375 1398 -1327
rect 1432 -1375 1490 -1327
rect 1524 -1375 1582 -1327
rect 1616 -1375 1674 -1327
rect 1708 -1375 1770 -1327
rect 1804 -1375 1858 -1327
rect 1892 -1375 1950 -1327
rect 1984 -1375 2042 -1327
rect 2076 -1375 2134 -1327
rect 2168 -1345 3240 -1327
rect 2168 -1375 2287 -1345
rect -116 -1379 2287 -1375
rect 2321 -1379 2361 -1345
rect 2395 -1379 2441 -1345
rect 2475 -1379 2521 -1345
rect 2555 -1379 2596 -1345
rect 2630 -1379 2670 -1345
rect 2704 -1379 2750 -1345
rect 2784 -1379 2830 -1345
rect 2864 -1379 2904 -1345
rect 2938 -1379 2984 -1345
rect 3018 -1379 3064 -1345
rect 3098 -1379 3144 -1345
rect 3178 -1379 3240 -1345
rect -116 -1395 3240 -1379
rect -686 -1544 -672 -1510
rect -494 -1544 -488 -1472
rect -686 -1628 -488 -1544
rect 200 -1590 660 -1395
rect 2278 -1396 3240 -1395
rect 2780 -1590 3240 -1396
rect 4317 -1544 4331 -1222
rect 4509 -1544 4515 -1222
rect -686 -2022 -642 -1628
rect -536 -2022 -488 -1628
rect -686 -2183 -488 -2022
rect -686 -2577 -648 -2183
rect -542 -2577 -488 -2183
rect 4317 -1790 4515 -1544
rect 4317 -1824 4395 -1790
rect 4429 -1824 4515 -1790
rect 4317 -2264 4515 -1824
rect 4317 -2298 4395 -2264
rect 4429 -2298 4515 -2264
rect 4048 -2365 4147 -2330
rect 4048 -2399 4080 -2365
rect 4114 -2399 4147 -2365
rect 4048 -2434 4147 -2399
rect -686 -2708 -488 -2577
rect -686 -2738 -602 -2708
rect -568 -2738 -488 -2708
rect -686 -3132 -633 -2738
rect -527 -3132 -488 -2738
rect -686 -3180 -488 -3132
rect 4317 -2738 4515 -2298
rect 4317 -2772 4395 -2738
rect 4429 -2772 4515 -2738
rect 200 -3180 660 -3170
rect 2780 -3180 3240 -3170
rect 4317 -3180 4515 -2772
rect -686 -3268 4515 -3180
rect -686 -3302 -72 -3268
rect -38 -3302 476 -3268
rect 510 -3302 1024 -3268
rect 1058 -3302 1572 -3268
rect 1606 -3302 2120 -3268
rect 2154 -3302 2668 -3268
rect 2702 -3302 3218 -3268
rect 3252 -3302 4515 -3268
rect -686 -3378 4515 -3302
<< viali >>
rect -638 1966 -608 1967
rect -608 1966 -574 1967
rect -574 1966 -532 1967
rect -638 1573 -532 1966
rect -651 1052 -545 1407
rect -651 1018 -608 1052
rect -608 1018 -574 1052
rect -574 1018 -545 1052
rect -651 1013 -545 1018
rect 4080 1191 4114 1225
rect -641 578 -535 852
rect -641 544 -608 578
rect -608 544 -574 578
rect -574 544 -535 578
rect -641 458 -535 544
rect 939 176 973 210
rect 1084 192 1118 226
rect 1168 192 1202 226
rect 1252 192 1286 226
rect 1336 192 1370 226
rect 1420 192 1454 226
rect 1504 192 1538 226
rect 1588 192 1622 226
rect 1672 192 1706 226
rect 1840 192 1874 226
rect 1924 192 1958 226
rect 2008 192 2042 226
rect 2080 192 2114 226
rect 2164 192 2198 226
rect 2248 192 2282 226
rect 2320 192 2354 226
rect 2404 192 2438 226
rect 2476 192 2510 226
rect 2632 192 2666 226
rect 2716 192 2750 226
rect 2788 192 2822 226
rect 2917 192 2951 226
rect 2989 192 3023 226
rect 3299 193 3333 227
rect 3371 193 3405 227
rect 3443 193 3477 227
rect 3515 193 3549 227
rect 3587 193 3621 227
rect 3659 193 3693 227
rect 3732 193 3766 227
rect 3804 193 3838 227
rect 3876 193 3910 227
rect 3948 193 3982 227
rect 4020 193 4054 227
rect 4092 193 4126 227
rect 939 93 973 127
rect 939 10 973 44
rect 939 -73 973 -39
rect -600 -164 -566 -130
rect -444 -164 -410 -130
rect -290 -164 -256 -130
rect -146 -164 -112 -130
rect -32 -164 2 -130
rect 82 -164 116 -130
rect 166 -164 200 -130
rect 250 -164 284 -130
rect 334 -164 368 -130
rect 418 -164 452 -130
rect 502 -164 536 -130
rect 586 -164 620 -130
rect 670 -164 704 -130
rect 754 -164 788 -130
rect 838 -164 872 -130
rect 922 -164 956 -130
rect 1102 -63 1136 -36
rect 1102 -70 1136 -63
rect -38 -310 -4 -276
rect 54 -310 88 -276
rect 148 -310 182 -293
rect 148 -327 182 -310
rect 240 -310 274 -276
rect 332 -310 366 -293
rect 332 -327 366 -310
rect 424 -310 458 -276
rect 516 -310 550 -293
rect 516 -327 550 -310
rect 608 -310 642 -276
rect 700 -310 734 -293
rect 700 -327 734 -310
rect 794 -310 828 -276
rect 886 -310 920 -276
rect 1190 -63 1224 -36
rect 1190 -70 1224 -63
rect 1278 -301 1312 -268
rect 1278 -302 1312 -301
rect 1366 -63 1400 -36
rect 1366 -70 1400 -63
rect 1454 5 1488 37
rect 1454 3 1488 5
rect 1542 -63 1576 -36
rect 1542 -70 1576 -63
rect 1630 -63 1664 -36
rect 1630 -70 1664 -63
rect 2579 93 2613 127
rect 28 -427 62 -393
rect 813 -427 847 -393
rect 1191 -436 1225 -402
rect 1889 -63 1923 -36
rect 1889 -70 1923 -63
rect 1977 -63 2011 -36
rect 1977 -70 2011 -63
rect 2065 5 2099 34
rect 2065 0 2099 5
rect 2153 -63 2187 -36
rect 2153 -70 2187 -63
rect 2241 -301 2275 -268
rect 2241 -302 2275 -301
rect 2329 -63 2363 -36
rect 2329 -70 2363 -63
rect 2417 -63 2451 -36
rect 2417 -70 2451 -63
rect 2579 10 2613 44
rect 2579 -73 2613 -39
rect 2579 -156 2613 -122
rect 1558 -447 1592 -413
rect 1963 -447 1997 -413
rect 2329 -436 2363 -402
rect 3463 -393 3497 -359
rect 3549 -393 3583 -359
rect 3633 -392 3667 -358
rect 3717 -393 3751 -359
rect 203 -526 237 -492
rect 645 -524 679 -490
rect 2721 -544 2755 -510
rect 2806 -543 2840 -509
rect 2890 -544 2924 -510
rect 2978 -543 3012 -509
rect 3061 -543 3095 -509
rect -16 -926 18 -914
rect -16 -948 18 -926
rect 72 -926 106 -914
rect 72 -948 106 -926
rect 160 -620 194 -586
rect 248 -926 282 -914
rect 248 -948 282 -926
rect 342 -620 370 -586
rect 370 -620 376 -586
rect 506 -620 512 -586
rect 512 -620 540 -586
rect 424 -926 458 -914
rect 424 -948 458 -926
rect 600 -926 634 -914
rect 600 -948 634 -926
rect 688 -620 722 -586
rect 776 -926 810 -914
rect 776 -948 810 -926
rect 864 -926 898 -914
rect 864 -948 898 -926
rect 1677 -696 1711 -663
rect 1677 -697 1711 -696
rect 1843 -696 1877 -663
rect 1843 -697 1877 -696
rect -16 -1137 18 -1103
rect 72 -1137 106 -1103
rect 160 -1137 194 -1103
rect 72 -1272 106 -1238
rect 248 -1137 282 -1103
rect 336 -1137 370 -1103
rect 248 -1272 282 -1238
rect 424 -1137 458 -1103
rect 512 -1137 546 -1103
rect 424 -1272 458 -1238
rect 600 -1137 634 -1103
rect 688 -1137 722 -1103
rect 600 -1272 634 -1238
rect 776 -1137 810 -1103
rect 864 -1137 898 -1103
rect 776 -1272 810 -1238
rect 1475 -1141 1509 -1137
rect 1475 -1171 1509 -1141
rect 1567 -1141 1601 -1137
rect 1567 -1171 1601 -1141
rect 1663 -1039 1697 -1018
rect 1663 -1052 1697 -1039
rect 1759 -1141 1793 -1137
rect 1759 -1171 1793 -1141
rect 1855 -937 1889 -933
rect 1855 -967 1889 -937
rect 1951 -1141 1985 -1137
rect 1951 -1171 1985 -1141
rect 2043 -1141 2077 -1137
rect 2043 -1171 2077 -1141
rect 3447 -970 3481 -936
rect 3519 -970 3553 -936
rect 3591 -970 3625 -936
rect 3663 -970 3697 -936
rect 3735 -970 3769 -936
rect 1649 -1242 1683 -1238
rect 1649 -1272 1655 -1242
rect 1655 -1272 1683 -1242
rect 1871 -1242 1905 -1238
rect 1871 -1272 1893 -1242
rect 1893 -1272 1905 -1242
rect 2789 -1274 2823 -1240
rect 2865 -1274 2899 -1240
rect 2941 -1274 2975 -1240
rect 3017 -1274 3051 -1240
rect 3206 -1274 3240 -1240
rect 3282 -1274 3316 -1240
rect 3358 -1274 3392 -1240
rect 3434 -1274 3468 -1240
rect 3510 -1274 3544 -1240
rect 3586 -1274 3620 -1240
rect 3662 -1274 3696 -1240
rect 3738 -1274 3772 -1240
rect -670 -1472 -492 -1366
rect 101 -1367 135 -1333
rect 219 -1367 253 -1333
rect 337 -1367 371 -1333
rect 455 -1367 489 -1333
rect 573 -1367 607 -1333
rect 691 -1367 725 -1333
rect 809 -1367 843 -1333
rect 1122 -1361 1156 -1341
rect 1122 -1375 1156 -1361
rect 1214 -1361 1248 -1341
rect 1214 -1375 1248 -1361
rect 1306 -1361 1340 -1341
rect 1306 -1375 1340 -1361
rect 1398 -1361 1432 -1341
rect 1398 -1375 1432 -1361
rect 1490 -1361 1524 -1341
rect 1490 -1375 1524 -1361
rect 1582 -1361 1616 -1341
rect 1582 -1375 1616 -1361
rect 1674 -1361 1708 -1341
rect 1674 -1375 1708 -1361
rect 1770 -1361 1804 -1341
rect 1770 -1375 1804 -1361
rect 1858 -1361 1892 -1341
rect 1858 -1375 1892 -1361
rect 1950 -1361 1984 -1341
rect 1950 -1375 1984 -1361
rect 2042 -1361 2076 -1341
rect 2042 -1375 2076 -1361
rect 2134 -1361 2168 -1341
rect 2134 -1375 2168 -1361
rect 2287 -1379 2321 -1345
rect 2361 -1379 2395 -1345
rect 2441 -1379 2475 -1345
rect 2521 -1379 2555 -1345
rect 2596 -1379 2630 -1345
rect 2670 -1379 2704 -1345
rect 2750 -1379 2784 -1345
rect 2830 -1379 2864 -1345
rect 2904 -1379 2938 -1345
rect 2984 -1379 3018 -1345
rect 3064 -1379 3098 -1345
rect 3144 -1379 3178 -1345
rect -670 -1510 -494 -1472
rect -672 -1544 -494 -1510
rect 4331 -1544 4509 -1222
rect -642 -1760 -536 -1628
rect -642 -1794 -602 -1760
rect -602 -1794 -568 -1760
rect -568 -1794 -536 -1760
rect -642 -2022 -536 -1794
rect -648 -2234 -542 -2183
rect -648 -2268 -602 -2234
rect -602 -2268 -568 -2234
rect -568 -2268 -542 -2234
rect -648 -2577 -542 -2268
rect 4080 -2399 4114 -2365
rect -633 -2742 -602 -2738
rect -602 -2742 -568 -2738
rect -568 -2742 -527 -2738
rect -633 -3132 -527 -2742
<< metal1 >>
rect -686 1967 -450 2000
rect -686 1956 -638 1967
rect -532 1956 -450 1967
rect -686 1584 -643 1956
rect -527 1584 -450 1956
rect -686 1573 -638 1584
rect -532 1573 -450 1584
rect -686 1530 -450 1573
rect 3890 1520 4154 1651
rect -686 1428 -510 1450
rect -686 992 -656 1428
rect -540 992 -510 1428
rect -686 970 -510 992
rect 4042 1234 4154 1520
rect 4042 1182 4071 1234
rect 4123 1182 4154 1234
rect 4042 900 4154 1182
rect -686 852 -450 890
rect -686 458 -641 852
rect -535 458 -450 852
rect 3890 769 4154 900
rect -686 420 -450 458
rect 809 368 4978 392
rect 809 227 4696 368
rect 809 226 3299 227
rect 809 210 1084 226
rect 809 176 939 210
rect 973 192 1084 210
rect 1118 192 1168 226
rect 1202 192 1252 226
rect 1286 192 1336 226
rect 1370 192 1420 226
rect 1454 192 1504 226
rect 1538 192 1588 226
rect 1622 192 1672 226
rect 1706 192 1840 226
rect 1874 192 1924 226
rect 1958 192 2008 226
rect 2042 192 2080 226
rect 2114 192 2164 226
rect 2198 192 2248 226
rect 2282 192 2320 226
rect 2354 192 2404 226
rect 2438 192 2476 226
rect 2510 192 2632 226
rect 2666 192 2716 226
rect 2750 192 2788 226
rect 2822 192 2917 226
rect 2951 192 2989 226
rect 3023 193 3299 226
rect 3333 193 3371 227
rect 3405 193 3443 227
rect 3477 193 3515 227
rect 3549 193 3587 227
rect 3621 193 3659 227
rect 3693 193 3732 227
rect 3766 193 3804 227
rect 3838 193 3876 227
rect 3910 193 3948 227
rect 3982 193 4020 227
rect 4054 193 4092 227
rect 4126 193 4696 227
rect 3023 192 4696 193
rect 973 188 4696 192
rect 4940 188 4978 368
rect 973 186 4978 188
rect 973 176 980 186
rect 809 127 980 176
rect 809 93 939 127
rect 973 93 980 127
rect 809 44 980 93
rect 809 10 939 44
rect 973 10 980 44
rect 809 -39 980 10
rect 1448 37 1494 186
rect 1448 3 1454 37
rect 1488 3 1494 37
rect 1448 -9 1494 3
rect 2059 34 2105 186
rect 2059 0 2065 34
rect 2099 0 2105 34
rect 2059 -12 2105 0
rect 2573 127 2619 186
rect 2573 93 2579 127
rect 2613 93 2619 127
rect 2573 44 2619 93
rect 2573 10 2579 44
rect 2613 10 2619 44
rect 809 -73 939 -39
rect 973 -73 980 -39
rect -641 -122 80 -101
rect 809 -122 980 -73
rect 1096 -36 1142 -16
rect 1096 -70 1102 -36
rect 1136 -41 1142 -36
rect 1184 -36 1230 -16
rect 1184 -41 1190 -36
rect 1136 -69 1190 -41
rect 1136 -70 1142 -69
rect 1096 -90 1142 -70
rect 1184 -70 1190 -69
rect 1224 -41 1230 -36
rect 1360 -36 1406 -16
rect 1360 -41 1366 -36
rect 1224 -69 1366 -41
rect 1224 -70 1230 -69
rect 1184 -90 1230 -70
rect 1360 -70 1366 -69
rect 1400 -41 1406 -36
rect 1536 -36 1582 -16
rect 1536 -41 1542 -36
rect 1400 -69 1542 -41
rect 1400 -70 1406 -69
rect 1360 -90 1406 -70
rect 1536 -70 1542 -69
rect 1576 -41 1582 -36
rect 1624 -36 1670 -16
rect 1624 -41 1630 -36
rect 1576 -69 1630 -41
rect 1576 -70 1582 -69
rect 1536 -90 1582 -70
rect 1624 -70 1630 -69
rect 1664 -70 1670 -36
rect 1624 -90 1670 -70
rect 1883 -36 1929 -16
rect 1883 -70 1889 -36
rect 1923 -41 1929 -36
rect 1971 -36 2017 -16
rect 1971 -41 1977 -36
rect 1923 -69 1977 -41
rect 1923 -70 1929 -69
rect 1883 -90 1929 -70
rect 1971 -70 1977 -69
rect 2011 -41 2017 -36
rect 2147 -36 2193 -16
rect 2147 -41 2153 -36
rect 2011 -69 2153 -41
rect 2011 -70 2017 -69
rect 1971 -90 2017 -70
rect 2147 -70 2153 -69
rect 2187 -41 2193 -36
rect 2323 -36 2369 -16
rect 2323 -41 2329 -36
rect 2187 -69 2329 -41
rect 2187 -70 2193 -69
rect 2147 -90 2193 -70
rect 2323 -70 2329 -69
rect 2363 -41 2369 -36
rect 2411 -36 2457 -16
rect 2411 -41 2417 -36
rect 2363 -69 2417 -41
rect 2363 -70 2369 -69
rect 2323 -90 2369 -70
rect 2411 -70 2417 -69
rect 2451 -70 2457 -36
rect 2411 -90 2457 -70
rect 2573 -39 2619 10
rect 2573 -73 2579 -39
rect 2613 -73 2619 -39
rect -641 -130 980 -122
rect -641 -164 -600 -130
rect -566 -164 -444 -130
rect -410 -164 -290 -130
rect -256 -164 -146 -130
rect -112 -164 -32 -130
rect 2 -164 82 -130
rect 116 -164 166 -130
rect 200 -164 250 -130
rect 284 -164 334 -130
rect 368 -164 418 -130
rect 452 -164 502 -130
rect 536 -164 586 -130
rect 620 -164 670 -130
rect 704 -164 754 -130
rect 788 -164 838 -130
rect 872 -164 922 -130
rect 956 -164 980 -130
rect -641 -177 980 -164
rect 2573 -122 2619 -73
rect 2573 -156 2579 -122
rect 2613 -156 2619 -122
rect 48 -239 94 -177
rect -44 -276 94 -239
rect 233 -253 280 -177
rect -44 -310 -38 -276
rect -4 -310 54 -276
rect 88 -310 94 -276
rect 234 -276 280 -253
rect -44 -347 94 -310
rect 142 -293 188 -277
rect 142 -327 148 -293
rect 182 -327 188 -293
rect 142 -375 188 -327
rect 234 -310 240 -276
rect 274 -310 280 -276
rect 418 -276 464 -177
rect 234 -347 280 -310
rect 326 -293 372 -277
rect 326 -327 332 -293
rect 366 -327 372 -293
rect 326 -375 372 -327
rect 418 -310 424 -276
rect 458 -310 464 -276
rect 602 -276 648 -177
rect 418 -347 464 -310
rect 510 -293 556 -277
rect 510 -327 516 -293
rect 550 -327 556 -293
rect -99 -384 81 -383
rect -99 -436 -84 -384
rect -32 -393 81 -384
rect -32 -427 28 -393
rect 62 -427 81 -393
rect 142 -407 372 -375
rect -32 -436 81 -427
rect -99 -437 81 -436
rect 327 -450 372 -407
rect 510 -379 556 -327
rect 602 -310 608 -276
rect 642 -310 648 -276
rect 788 -239 834 -177
rect 2573 -191 2619 -156
rect 2651 -212 2721 -184
rect 788 -276 926 -239
rect 602 -347 648 -310
rect 694 -293 740 -277
rect 694 -327 700 -293
rect 734 -327 740 -293
rect 694 -379 740 -327
rect 788 -310 794 -276
rect 828 -310 886 -276
rect 920 -310 926 -276
rect 788 -347 926 -310
rect 1269 -268 1321 -240
rect 1269 -302 1278 -268
rect 1312 -302 1321 -268
rect 1269 -316 1321 -302
rect 2232 -268 2284 -241
rect 2232 -302 2241 -268
rect 2275 -302 2284 -268
rect 2232 -316 2284 -302
rect 510 -407 740 -379
rect 795 -384 984 -383
rect 795 -393 917 -384
rect 510 -450 555 -407
rect 795 -427 813 -393
rect 847 -427 917 -393
rect 795 -436 917 -427
rect 969 -436 984 -384
rect 795 -437 984 -436
rect 1174 -396 1244 -386
rect 327 -456 383 -450
rect 180 -526 193 -474
rect 245 -526 260 -474
rect 180 -533 260 -526
rect 379 -508 383 -456
rect 154 -586 206 -568
rect 154 -620 160 -586
rect 194 -604 206 -586
rect 327 -586 383 -508
rect 327 -604 342 -586
rect 194 -620 342 -604
rect 376 -620 383 -586
rect 154 -632 383 -620
rect 499 -456 555 -450
rect 1174 -448 1181 -396
rect 1233 -448 1244 -396
rect 1174 -453 1244 -448
rect 499 -508 503 -456
rect 499 -586 555 -508
rect 622 -524 636 -472
rect 688 -524 702 -472
rect 622 -531 702 -524
rect 1272 -548 1318 -316
rect 1530 -413 1618 -397
rect 1530 -447 1558 -413
rect 1592 -430 1618 -413
rect 1935 -413 2023 -397
rect 1935 -430 1963 -413
rect 1592 -447 1684 -430
rect 1530 -463 1684 -447
rect 1678 -482 1684 -463
rect 1736 -482 1742 -430
rect 1811 -482 1817 -430
rect 1869 -447 1963 -430
rect 1997 -447 2023 -413
rect 1869 -463 2023 -447
rect 1869 -482 1875 -463
rect 1811 -548 1839 -482
rect 2235 -548 2281 -316
rect 2313 -396 2379 -386
rect 2651 -396 2679 -212
rect 2313 -448 2321 -396
rect 2373 -448 2379 -396
rect 2313 -454 2379 -448
rect 2637 -428 2679 -396
rect 3307 -358 4157 -314
rect 3307 -359 3633 -358
rect 3307 -393 3463 -359
rect 3497 -393 3549 -359
rect 3583 -392 3633 -359
rect 3667 -359 4157 -358
rect 3667 -392 3717 -359
rect 3583 -393 3717 -392
rect 3751 -361 4157 -359
rect 3751 -393 3981 -361
rect 3307 -413 3981 -393
rect 4033 -413 4060 -361
rect 4112 -413 4157 -361
rect 499 -620 506 -586
rect 540 -603 555 -586
rect 676 -586 728 -567
rect 1272 -576 1624 -548
rect 676 -603 688 -586
rect 540 -620 688 -603
rect 722 -620 728 -586
rect 1618 -600 1624 -576
rect 1676 -576 1839 -548
rect 1676 -600 1682 -576
rect 1867 -600 1873 -548
rect 1925 -576 2281 -548
rect 1925 -600 1931 -576
rect 499 -632 728 -620
rect 1654 -663 1734 -646
rect 1654 -697 1677 -663
rect 1711 -697 1734 -663
rect 1654 -708 1734 -697
rect 1654 -760 1670 -708
rect 1722 -760 1734 -708
rect 1654 -766 1734 -760
rect 1820 -663 1900 -646
rect 1820 -697 1843 -663
rect 1877 -697 1900 -663
rect 1820 -708 1900 -697
rect 1820 -760 1833 -708
rect 1885 -760 1900 -708
rect 1820 -766 1900 -760
rect -22 -914 24 -867
rect -22 -948 -16 -914
rect 18 -948 24 -914
rect -486 -964 -398 -953
rect -486 -1016 -468 -964
rect -416 -1016 -398 -964
rect -486 -1027 -398 -1016
rect -22 -1004 24 -948
rect 66 -914 112 -867
rect 66 -948 72 -914
rect 106 -948 112 -914
rect 66 -1004 112 -948
rect 242 -914 288 -867
rect 242 -948 248 -914
rect 282 -948 288 -914
rect 242 -1004 288 -948
rect 418 -914 464 -867
rect 418 -948 424 -914
rect 458 -948 464 -914
rect 418 -1004 464 -948
rect 594 -914 640 -867
rect 594 -948 600 -914
rect 634 -948 640 -914
rect 594 -1004 640 -948
rect 770 -914 816 -867
rect 770 -948 776 -914
rect 810 -948 816 -914
rect 770 -1004 816 -948
rect 858 -914 904 -867
rect 858 -948 864 -914
rect 898 -948 904 -914
rect 858 -1004 904 -948
rect 1648 -923 1712 -921
rect 1648 -950 1654 -923
rect 1353 -975 1654 -950
rect 1706 -950 1712 -923
rect 1839 -933 1903 -921
rect 1839 -950 1855 -933
rect 1706 -967 1855 -950
rect 1889 -950 1903 -933
rect 2637 -950 2665 -428
rect 3307 -436 4157 -413
rect 3307 -462 3367 -436
rect 2695 -509 3367 -462
rect 2695 -510 2806 -509
rect 2695 -544 2721 -510
rect 2755 -543 2806 -510
rect 2840 -510 2978 -509
rect 2840 -543 2890 -510
rect 2755 -544 2890 -543
rect 2924 -543 2978 -510
rect 3012 -543 3061 -509
rect 3095 -525 3367 -509
rect 3095 -543 3119 -525
rect 2924 -544 3119 -543
rect 2695 -590 3119 -544
rect 1889 -967 2665 -950
rect 1706 -975 2665 -967
rect 1353 -978 2665 -975
rect -22 -1036 904 -1004
rect 2693 -1006 2721 -840
rect 3407 -936 3825 -928
rect 3407 -970 3447 -936
rect 3481 -970 3519 -936
rect 3553 -970 3591 -936
rect 3625 -970 3663 -936
rect 3697 -970 3735 -936
rect 3769 -970 3825 -936
rect 3407 -978 3825 -970
rect 1353 -1008 2721 -1006
rect 1353 -1018 1845 -1008
rect 1353 -1034 1663 -1018
rect -22 -1103 24 -1036
rect -22 -1137 -16 -1103
rect 18 -1137 24 -1103
rect -22 -1174 24 -1137
rect 66 -1103 112 -1036
rect 66 -1137 72 -1103
rect 106 -1137 112 -1103
rect 66 -1174 112 -1137
rect 154 -1103 200 -1064
rect 154 -1137 160 -1103
rect 194 -1137 200 -1103
rect 154 -1174 200 -1137
rect 242 -1103 288 -1036
rect 242 -1137 248 -1103
rect 282 -1137 288 -1103
rect 242 -1174 288 -1137
rect 330 -1103 376 -1064
rect 330 -1137 336 -1103
rect 370 -1137 376 -1103
rect 330 -1174 376 -1137
rect 418 -1103 464 -1036
rect 418 -1137 424 -1103
rect 458 -1137 464 -1103
rect 418 -1174 464 -1137
rect 506 -1103 552 -1064
rect 506 -1137 512 -1103
rect 546 -1137 552 -1103
rect 506 -1174 552 -1137
rect 594 -1103 640 -1036
rect 594 -1137 600 -1103
rect 634 -1137 640 -1103
rect 594 -1174 640 -1137
rect 682 -1103 728 -1064
rect 682 -1137 688 -1103
rect 722 -1137 728 -1103
rect 682 -1174 728 -1137
rect 770 -1103 816 -1036
rect 770 -1137 776 -1103
rect 810 -1137 816 -1103
rect 770 -1174 816 -1137
rect 858 -1103 904 -1036
rect 1648 -1052 1663 -1034
rect 1697 -1034 1845 -1018
rect 1697 -1052 1712 -1034
rect 1648 -1063 1712 -1052
rect 1839 -1060 1845 -1034
rect 1897 -1034 2721 -1008
rect 3697 -980 3825 -978
rect 3697 -1032 3703 -980
rect 3755 -1032 3767 -980
rect 3819 -1032 3825 -980
rect 1897 -1060 1903 -1034
rect 1839 -1063 1903 -1060
rect 858 -1137 864 -1103
rect 898 -1137 904 -1103
rect 858 -1174 904 -1137
rect 1463 -1137 1607 -1118
rect 1463 -1171 1475 -1137
rect 1509 -1171 1567 -1137
rect 1601 -1171 1607 -1137
rect 1463 -1182 1607 -1171
rect 30 -1238 852 -1226
rect 30 -1244 72 -1238
rect -99 -1296 -91 -1244
rect -39 -1272 72 -1244
rect 106 -1272 248 -1238
rect 282 -1272 424 -1238
rect 458 -1272 600 -1238
rect 634 -1272 776 -1238
rect 810 -1244 852 -1238
rect 810 -1272 925 -1244
rect -39 -1296 925 -1272
rect 977 -1296 984 -1244
rect -99 -1298 984 -1296
rect 1561 -1326 1607 -1182
rect 1753 -1137 1799 -1118
rect 1753 -1171 1759 -1137
rect 1793 -1171 1799 -1137
rect 1635 -1226 1705 -1218
rect 1635 -1278 1644 -1226
rect 1696 -1278 1705 -1226
rect 1635 -1284 1705 -1278
rect 1753 -1326 1799 -1171
rect 1945 -1137 2089 -1118
rect 1945 -1171 1951 -1137
rect 1985 -1171 2043 -1137
rect 2077 -1171 2089 -1137
rect 1945 -1182 2089 -1171
rect 1847 -1226 1917 -1218
rect 1847 -1278 1855 -1226
rect 1907 -1278 1917 -1226
rect 1847 -1284 1917 -1278
rect 1945 -1326 1991 -1182
rect 3681 -1192 3830 -1156
rect 3681 -1234 3730 -1192
rect 2762 -1240 3730 -1234
rect 2762 -1274 2789 -1240
rect 2823 -1274 2865 -1240
rect 2899 -1274 2941 -1240
rect 2975 -1274 3017 -1240
rect 3051 -1274 3206 -1240
rect 3240 -1274 3282 -1240
rect 3316 -1274 3358 -1240
rect 3392 -1274 3434 -1240
rect 3468 -1274 3510 -1240
rect 3544 -1274 3586 -1240
rect 3620 -1274 3662 -1240
rect 3696 -1244 3730 -1240
rect 3782 -1244 3830 -1192
rect 3696 -1274 3738 -1244
rect 3772 -1274 3830 -1244
rect 2762 -1280 3830 -1274
rect 4317 -1222 4515 -1202
rect 4317 -1326 4331 -1222
rect -686 -1333 4331 -1326
rect -686 -1366 101 -1333
rect -686 -1510 -670 -1366
rect -492 -1367 101 -1366
rect 135 -1367 219 -1333
rect 253 -1367 337 -1333
rect 371 -1367 455 -1333
rect 489 -1367 573 -1333
rect 607 -1367 691 -1333
rect 725 -1367 809 -1333
rect 843 -1340 4331 -1333
rect 843 -1341 1750 -1340
rect 1802 -1341 4331 -1340
rect 843 -1367 1122 -1341
rect -492 -1375 1122 -1367
rect 1156 -1375 1214 -1341
rect 1248 -1375 1306 -1341
rect 1340 -1375 1398 -1341
rect 1432 -1375 1490 -1341
rect 1524 -1375 1582 -1341
rect 1616 -1375 1674 -1341
rect 1708 -1375 1750 -1341
rect 1804 -1375 1858 -1341
rect 1892 -1375 1950 -1341
rect 1984 -1375 2042 -1341
rect 2076 -1375 2134 -1341
rect 2168 -1345 4331 -1341
rect 2168 -1375 2287 -1345
rect -492 -1379 1750 -1375
rect -492 -1472 -398 -1379
rect -494 -1495 -398 -1472
rect 102 -1392 1750 -1379
rect 1802 -1379 2287 -1375
rect 2321 -1379 2361 -1345
rect 2395 -1379 2441 -1345
rect 2475 -1379 2521 -1345
rect 2555 -1379 2596 -1345
rect 2630 -1379 2670 -1345
rect 2704 -1379 2750 -1345
rect 2784 -1379 2830 -1345
rect 2864 -1379 2904 -1345
rect 2938 -1379 2984 -1345
rect 3018 -1379 3064 -1345
rect 3098 -1379 3144 -1345
rect 3178 -1379 4331 -1345
rect 1802 -1392 4331 -1379
rect 102 -1495 4331 -1392
rect -686 -1544 -672 -1510
rect -494 -1544 4331 -1495
rect 4509 -1326 4515 -1222
rect 4509 -1355 4588 -1326
rect 4509 -1407 4526 -1355
rect 4578 -1407 4588 -1355
rect 4509 -1419 4588 -1407
rect 4509 -1471 4526 -1419
rect 4578 -1471 4588 -1419
rect 4509 -1483 4588 -1471
rect 4509 -1535 4526 -1483
rect 4578 -1535 4588 -1483
rect 4509 -1544 4588 -1535
rect -686 -1558 4588 -1544
rect -686 -1628 -450 -1590
rect -686 -2022 -642 -1628
rect -536 -2022 -450 -1628
rect -686 -2060 -450 -2022
rect 3890 -2070 4154 -1939
rect -686 -2162 -510 -2140
rect -686 -2598 -653 -2162
rect -537 -2598 -510 -2162
rect -686 -2620 -510 -2598
rect 4042 -2356 4154 -2070
rect 4042 -2408 4071 -2356
rect 4123 -2408 4154 -2356
rect 4042 -2690 4154 -2408
rect -686 -2738 -450 -2700
rect -686 -2749 -633 -2738
rect -686 -3121 -652 -2749
rect -686 -3132 -633 -3121
rect -527 -3132 -450 -2738
rect 3890 -2821 4154 -2690
rect -686 -3170 -450 -3132
<< via1 >>
rect -643 1584 -638 1956
rect -638 1584 -532 1956
rect -532 1584 -527 1956
rect -656 1407 -540 1428
rect -656 1013 -651 1407
rect -651 1013 -545 1407
rect -545 1013 -540 1407
rect -656 992 -540 1013
rect 4071 1225 4123 1234
rect 4071 1191 4080 1225
rect 4080 1191 4114 1225
rect 4114 1191 4123 1225
rect 4071 1182 4123 1191
rect 4696 188 4940 368
rect -84 -436 -32 -384
rect 917 -436 969 -384
rect 193 -492 245 -474
rect 193 -526 203 -492
rect 203 -526 237 -492
rect 237 -526 245 -492
rect 327 -508 379 -456
rect 1181 -402 1233 -396
rect 1181 -436 1191 -402
rect 1191 -436 1225 -402
rect 1225 -436 1233 -402
rect 1181 -448 1233 -436
rect 503 -508 555 -456
rect 636 -490 688 -472
rect 636 -524 645 -490
rect 645 -524 679 -490
rect 679 -524 688 -490
rect 1684 -482 1736 -430
rect 1817 -482 1869 -430
rect 2321 -402 2373 -396
rect 2321 -436 2329 -402
rect 2329 -436 2363 -402
rect 2363 -436 2373 -402
rect 2321 -448 2373 -436
rect 3981 -413 4033 -361
rect 4060 -413 4112 -361
rect 1624 -600 1676 -548
rect 1873 -600 1925 -548
rect 1670 -760 1722 -708
rect 1833 -760 1885 -708
rect -468 -1016 -416 -964
rect 1654 -975 1706 -923
rect 1845 -1060 1897 -1008
rect 3703 -1032 3755 -980
rect 3767 -1032 3819 -980
rect -91 -1296 -39 -1244
rect 925 -1296 977 -1244
rect 1644 -1238 1696 -1226
rect 1644 -1272 1649 -1238
rect 1649 -1272 1683 -1238
rect 1683 -1272 1696 -1238
rect 1644 -1278 1696 -1272
rect 1855 -1238 1907 -1226
rect 1855 -1272 1871 -1238
rect 1871 -1272 1905 -1238
rect 1905 -1272 1907 -1238
rect 1855 -1278 1907 -1272
rect 3730 -1240 3782 -1192
rect 3730 -1244 3738 -1240
rect 3738 -1244 3772 -1240
rect 3772 -1244 3782 -1240
rect 1750 -1341 1802 -1340
rect 1750 -1375 1770 -1341
rect 1770 -1375 1802 -1341
rect -398 -1495 102 -1379
rect 1750 -1392 1802 -1375
rect 4526 -1407 4578 -1355
rect 4526 -1471 4578 -1419
rect 4526 -1535 4578 -1483
rect -653 -2183 -537 -2162
rect -653 -2577 -648 -2183
rect -648 -2577 -542 -2183
rect -542 -2577 -537 -2183
rect -653 -2598 -537 -2577
rect 4071 -2365 4123 -2356
rect 4071 -2399 4080 -2365
rect 4080 -2399 4114 -2365
rect 4114 -2399 4123 -2365
rect 4071 -2408 4123 -2399
rect -652 -3121 -633 -2749
rect -633 -3121 -536 -2749
<< metal2 >>
rect -686 1958 -450 2000
rect -686 1956 -613 1958
rect -557 1956 -450 1958
rect -686 1584 -643 1956
rect -527 1584 -450 1956
rect -686 1582 -613 1584
rect -557 1582 -450 1584
rect -686 1530 -450 1582
rect -686 1428 -510 1450
rect -686 1398 -656 1428
rect -540 1398 -510 1428
rect -686 1022 -666 1398
rect -530 1022 -510 1398
rect 4042 1234 4154 1265
rect 4042 1182 4071 1234
rect 4123 1182 4154 1234
rect 4042 1149 4154 1182
rect -686 992 -656 1022
rect -540 992 -510 1022
rect -686 970 -510 992
rect 1744 335 1808 420
rect 1744 279 1748 335
rect 1804 279 1808 335
rect 1744 266 1808 279
rect 4658 368 4978 392
rect 4658 188 4696 368
rect 4940 188 4978 368
rect 4658 162 4978 188
rect 3967 -362 3981 -361
rect -99 -384 -17 -383
rect -99 -436 -84 -384
rect -32 -436 -17 -384
rect -99 -437 -17 -436
rect 902 -384 984 -383
rect 902 -436 917 -384
rect 969 -436 984 -384
rect 902 -437 984 -436
rect -486 -962 -398 -953
rect -486 -1018 -470 -962
rect -414 -1018 -398 -962
rect -486 -1027 -398 -1018
rect -99 -1244 -71 -437
rect 327 -456 383 -450
rect 179 -470 261 -460
rect 179 -526 190 -470
rect 246 -526 261 -470
rect 179 -533 261 -526
rect 379 -477 383 -456
rect 327 -542 383 -533
rect 499 -456 555 -450
rect 499 -477 503 -456
rect 620 -468 702 -458
rect 620 -524 634 -468
rect 690 -524 702 -468
rect 620 -531 702 -524
rect 499 -542 555 -533
rect 956 -1244 984 -437
rect 1174 -396 1244 -386
rect 1174 -448 1181 -396
rect 1233 -413 1244 -396
rect 2313 -396 2379 -386
rect 2313 -413 2321 -396
rect 1233 -422 1354 -413
rect 1233 -448 1298 -422
rect 1174 -453 1298 -448
rect 2198 -422 2321 -413
rect 1678 -454 1684 -430
rect 1298 -487 1354 -478
rect 1561 -482 1684 -454
rect 1736 -482 1742 -430
rect 1561 -708 1589 -482
rect 1710 -548 1742 -482
rect 1811 -482 1817 -430
rect 1869 -454 1875 -430
rect 1869 -482 1988 -454
rect 1811 -519 1839 -482
rect 1618 -600 1624 -548
rect 1676 -600 1682 -548
rect 1710 -576 1873 -548
rect 1867 -600 1873 -576
rect 1925 -600 1931 -548
rect 1960 -708 1988 -482
rect 2254 -448 2321 -422
rect 2373 -448 2379 -396
rect 3967 -418 3976 -362
rect 4033 -413 4060 -361
rect 4112 -362 4126 -361
rect 4032 -418 4060 -413
rect 4116 -418 4126 -362
rect 3967 -419 4126 -418
rect 2254 -454 2379 -448
rect 2198 -487 2254 -478
rect 1561 -736 1670 -708
rect 1664 -760 1670 -736
rect 1722 -760 1728 -708
rect 1827 -760 1833 -708
rect 1885 -736 1988 -708
rect 1885 -760 1891 -736
rect 1678 -897 1706 -760
rect 1654 -923 1706 -897
rect 1654 -1066 1706 -975
rect 1845 -897 1873 -760
rect 1845 -1008 1897 -897
rect 1845 -1066 1897 -1060
rect 3681 -980 3830 -978
rect 3681 -1032 3703 -980
rect 3755 -1032 3767 -980
rect 3819 -1032 3830 -980
rect 1746 -1079 1806 -1070
rect 1746 -1135 1748 -1079
rect 1804 -1135 1806 -1079
rect -99 -1296 -91 -1244
rect -39 -1296 -31 -1244
rect -99 -1298 -31 -1296
rect 916 -1296 925 -1244
rect 977 -1296 984 -1244
rect 1633 -1222 1707 -1218
rect 1633 -1278 1642 -1222
rect 1698 -1278 1707 -1222
rect 1633 -1284 1707 -1278
rect 916 -1298 984 -1296
rect -450 -1369 190 -1326
rect -450 -1505 -416 -1369
rect 120 -1505 190 -1369
rect 1746 -1340 1806 -1135
rect 3681 -1107 3830 -1032
rect 3681 -1163 3727 -1107
rect 3783 -1163 3830 -1107
rect 3681 -1192 3830 -1163
rect 3681 -1210 3730 -1192
rect 3782 -1210 3830 -1192
rect 1844 -1222 1918 -1215
rect 1844 -1278 1853 -1222
rect 1909 -1278 1918 -1222
rect 1844 -1287 1918 -1278
rect 3681 -1266 3728 -1210
rect 3784 -1266 3830 -1210
rect 3681 -1280 3830 -1266
rect 1746 -1392 1750 -1340
rect 1802 -1392 1806 -1340
rect 1746 -1400 1806 -1392
rect 4268 -1355 4588 -1326
rect 4268 -1377 4526 -1355
rect -450 -1590 190 -1505
rect 1744 -1447 1808 -1434
rect 1744 -1503 1748 -1447
rect 1804 -1503 1808 -1447
rect 1744 -1590 1808 -1503
rect 4268 -1513 4325 -1377
rect 4578 -1407 4588 -1355
rect 4541 -1419 4588 -1407
rect 4578 -1471 4588 -1419
rect 4541 -1483 4588 -1471
rect 4268 -1535 4526 -1513
rect 4578 -1535 4588 -1483
rect 4268 -1558 4588 -1535
rect -686 -2162 -510 -2140
rect -686 -2598 -653 -2162
rect -537 -2598 -510 -2162
rect 4042 -2356 4154 -2325
rect 4042 -2408 4071 -2356
rect 4123 -2408 4154 -2356
rect 4042 -2441 4154 -2408
rect -686 -2620 -510 -2598
rect -686 -2747 -450 -2700
rect -686 -2749 -622 -2747
rect -566 -2749 -450 -2747
rect -686 -3121 -652 -2749
rect -536 -3121 -450 -2749
rect -686 -3123 -622 -3121
rect -566 -3123 -450 -3121
rect -686 -3170 -450 -3123
<< via2 >>
rect -613 1956 -557 1958
rect -613 1902 -557 1956
rect -613 1822 -557 1878
rect -613 1742 -557 1798
rect -613 1662 -557 1718
rect -613 1584 -557 1638
rect -613 1582 -557 1584
rect -666 1022 -656 1398
rect -656 1022 -540 1398
rect -540 1022 -530 1398
rect 1748 279 1804 335
rect 4710 207 4926 343
rect -470 -964 -414 -962
rect -470 -1016 -468 -964
rect -468 -1016 -416 -964
rect -416 -1016 -414 -964
rect -470 -1018 -414 -1016
rect 190 -474 246 -470
rect 190 -526 193 -474
rect 193 -526 245 -474
rect 245 -526 246 -474
rect 327 -508 379 -477
rect 379 -508 383 -477
rect 327 -533 383 -508
rect 499 -508 503 -477
rect 503 -508 555 -477
rect 499 -533 555 -508
rect 634 -472 690 -468
rect 634 -524 636 -472
rect 636 -524 688 -472
rect 688 -524 690 -472
rect 1298 -478 1354 -422
rect 2198 -478 2254 -422
rect 3976 -413 3981 -362
rect 3981 -413 4032 -362
rect 4060 -413 4112 -362
rect 4112 -413 4116 -362
rect 3976 -418 4032 -413
rect 4060 -418 4116 -413
rect 1748 -1135 1804 -1079
rect 1642 -1226 1698 -1222
rect 1642 -1278 1644 -1226
rect 1644 -1278 1696 -1226
rect 1696 -1278 1698 -1226
rect -416 -1379 120 -1369
rect -416 -1495 -398 -1379
rect -398 -1495 102 -1379
rect 102 -1495 120 -1379
rect -416 -1505 120 -1495
rect 3727 -1163 3783 -1107
rect 1853 -1226 1909 -1222
rect 1853 -1278 1855 -1226
rect 1855 -1278 1907 -1226
rect 1907 -1278 1909 -1226
rect 3728 -1244 3730 -1210
rect 3730 -1244 3782 -1210
rect 3782 -1244 3784 -1210
rect 3728 -1266 3784 -1244
rect 1748 -1503 1804 -1447
rect 4325 -1407 4526 -1377
rect 4526 -1407 4541 -1377
rect 4325 -1419 4541 -1407
rect 4325 -1471 4526 -1419
rect 4526 -1471 4541 -1419
rect 4325 -1483 4541 -1471
rect 4325 -1513 4526 -1483
rect 4526 -1513 4541 -1483
rect -623 -2248 -567 -2192
rect -623 -2328 -567 -2272
rect -623 -2408 -567 -2352
rect -623 -2488 -567 -2432
rect -623 -2568 -567 -2512
rect -622 -2749 -566 -2747
rect -622 -2803 -566 -2749
rect -622 -2883 -566 -2827
rect -622 -2963 -566 -2907
rect -622 -3043 -566 -2987
rect -622 -3121 -566 -3067
rect -622 -3123 -566 -3121
<< metal3 >>
rect -686 1962 -512 2000
rect -686 1898 -617 1962
rect -553 1898 -512 1962
rect -686 1882 -512 1898
rect -686 1818 -617 1882
rect -553 1818 -512 1882
rect -686 1802 -512 1818
rect -686 1738 -617 1802
rect -553 1738 -512 1802
rect -686 1722 -512 1738
rect -686 1658 -617 1722
rect -553 1658 -512 1722
rect -686 1642 -512 1658
rect -686 1578 -617 1642
rect -553 1578 -512 1642
rect -686 1530 -512 1578
rect -686 1402 -510 1450
rect -686 1398 -630 1402
rect -566 1398 -510 1402
rect -686 1022 -666 1398
rect -530 1022 -510 1398
rect 3890 1240 4588 1265
rect 3890 1176 4321 1240
rect 4385 1176 4401 1240
rect 4465 1176 4481 1240
rect 4545 1176 4588 1240
rect 3890 1149 4588 1176
rect -686 1018 -630 1022
rect -566 1018 -510 1022
rect -686 970 -510 1018
rect 1724 339 1824 357
rect 1724 275 1744 339
rect 1808 275 1824 339
rect 1724 261 1824 275
rect 4658 347 4978 392
rect 4658 203 4706 347
rect 4930 203 4978 347
rect 1291 -422 1361 -415
rect 185 -470 261 -461
rect 185 -526 190 -470
rect 246 -526 261 -470
rect 185 -533 261 -526
rect 322 -477 390 -459
rect 322 -533 327 -477
rect 383 -533 390 -477
rect 322 -560 390 -533
rect 320 -855 390 -560
rect 384 -919 390 -855
rect 320 -925 390 -919
rect 492 -477 560 -459
rect 492 -533 499 -477
rect 555 -533 560 -477
rect 620 -468 695 -459
rect 620 -524 634 -468
rect 690 -524 695 -468
rect 620 -531 695 -524
rect 1043 -483 1107 -470
rect 492 -560 560 -533
rect 492 -729 562 -560
rect 492 -793 498 -729
rect 492 -925 562 -793
rect 1043 -729 1107 -547
rect 1043 -925 1107 -793
rect 1167 -609 1231 -473
rect 1167 -855 1231 -673
rect 1291 -478 1298 -422
rect 1354 -478 1361 -422
rect 1746 -423 1806 201
rect 4658 162 4978 203
rect 3963 -358 4130 -356
rect 2191 -422 2261 -415
rect 1291 -483 1361 -478
rect 1291 -547 1294 -483
rect 1358 -547 1361 -483
rect 1291 -679 1361 -547
rect 1556 -733 1996 -423
rect 2191 -478 2198 -422
rect 2254 -478 2261 -422
rect 3963 -422 3969 -358
rect 4033 -422 4060 -358
rect 4124 -422 4130 -358
rect 3963 -424 4130 -422
rect 2191 -609 2261 -478
rect 2191 -673 2194 -609
rect 2258 -673 2261 -609
rect 2191 -679 2261 -673
rect 2322 -483 2386 -470
rect 2322 -729 2386 -547
rect 1167 -925 1231 -919
rect -486 -960 -398 -953
rect -486 -962 -165 -960
rect -486 -1018 -470 -962
rect -414 -1018 -165 -962
rect -486 -1020 -165 -1018
rect -486 -1027 -398 -1020
rect -230 -1204 -165 -1020
rect 1743 -1079 1809 -733
rect 2322 -925 2386 -793
rect 2448 -609 2512 -473
rect 2448 -855 2512 -673
rect 2448 -925 2512 -919
rect 1743 -1135 1748 -1079
rect 1804 -1135 1809 -1079
rect 4658 -1057 4978 -1022
rect 4658 -1087 4709 -1057
rect 1743 -1144 1809 -1135
rect 3681 -1107 4709 -1087
rect 3681 -1163 3727 -1107
rect 3783 -1121 4709 -1107
rect 4773 -1121 4789 -1057
rect 4853 -1121 4869 -1057
rect 4933 -1121 4978 -1057
rect 3783 -1156 4978 -1121
rect 3783 -1163 3830 -1156
rect -230 -1222 1918 -1204
rect -230 -1264 1642 -1222
rect 1630 -1278 1642 -1264
rect 1698 -1278 1853 -1222
rect 1909 -1278 1918 -1222
rect 1630 -1288 1918 -1278
rect 3681 -1210 3830 -1163
rect 3681 -1266 3728 -1210
rect 3784 -1266 3830 -1210
rect 3681 -1280 3830 -1266
rect -450 -1369 180 -1326
rect -450 -1505 -416 -1369
rect 120 -1505 180 -1369
rect 4268 -1373 4588 -1326
rect -450 -1526 180 -1505
rect 1724 -1443 1825 -1432
rect 1724 -1507 1744 -1443
rect 1808 -1507 1825 -1443
rect 1724 -1528 1825 -1507
rect 4268 -1517 4321 -1373
rect 4545 -1517 4588 -1373
rect 4268 -1558 4588 -1517
rect -686 -2188 -510 -2140
rect -686 -2252 -627 -2188
rect -563 -2252 -510 -2188
rect -686 -2268 -510 -2252
rect -686 -2332 -627 -2268
rect -563 -2332 -510 -2268
rect -686 -2348 -510 -2332
rect -686 -2412 -627 -2348
rect -563 -2412 -510 -2348
rect -686 -2428 -510 -2412
rect -686 -2492 -627 -2428
rect -563 -2492 -510 -2428
rect 3889 -2353 4588 -2325
rect 3889 -2417 4321 -2353
rect 4385 -2417 4401 -2353
rect 4465 -2417 4481 -2353
rect 4545 -2417 4588 -2353
rect 3889 -2442 4588 -2417
rect -686 -2508 -510 -2492
rect -686 -2572 -627 -2508
rect -563 -2572 -510 -2508
rect -686 -2620 -510 -2572
rect -686 -2743 -514 -2700
rect -686 -2807 -626 -2743
rect -562 -2807 -514 -2743
rect -686 -2823 -514 -2807
rect -686 -2887 -626 -2823
rect -562 -2887 -514 -2823
rect -686 -2903 -514 -2887
rect -686 -2967 -626 -2903
rect -562 -2967 -514 -2903
rect -686 -2983 -514 -2967
rect -686 -3047 -626 -2983
rect -562 -3047 -514 -2983
rect -686 -3063 -514 -3047
rect -686 -3127 -626 -3063
rect -562 -3127 -514 -3063
rect -686 -3170 -514 -3127
<< via3 >>
rect -617 1958 -553 1962
rect -617 1902 -613 1958
rect -613 1902 -557 1958
rect -557 1902 -553 1958
rect -617 1898 -553 1902
rect -617 1878 -553 1882
rect -617 1822 -613 1878
rect -613 1822 -557 1878
rect -557 1822 -553 1878
rect -617 1818 -553 1822
rect -617 1798 -553 1802
rect -617 1742 -613 1798
rect -613 1742 -557 1798
rect -557 1742 -553 1798
rect -617 1738 -553 1742
rect -617 1718 -553 1722
rect -617 1662 -613 1718
rect -613 1662 -557 1718
rect -557 1662 -553 1718
rect -617 1658 -553 1662
rect -617 1638 -553 1642
rect -617 1582 -613 1638
rect -613 1582 -557 1638
rect -557 1582 -553 1638
rect -617 1578 -553 1582
rect -630 1398 -566 1402
rect -630 1338 -566 1398
rect -630 1258 -566 1322
rect -630 1178 -566 1242
rect -630 1098 -566 1162
rect -630 1022 -566 1082
rect 4321 1176 4385 1240
rect 4401 1176 4465 1240
rect 4481 1176 4545 1240
rect -630 1018 -566 1022
rect 1744 335 1808 339
rect 1744 279 1748 335
rect 1748 279 1804 335
rect 1804 279 1808 335
rect 1744 275 1808 279
rect 4706 343 4930 347
rect 4706 207 4710 343
rect 4710 207 4926 343
rect 4926 207 4930 343
rect 4706 203 4930 207
rect 320 -919 384 -855
rect 1043 -547 1107 -483
rect 498 -793 562 -729
rect 1043 -793 1107 -729
rect 1167 -673 1231 -609
rect 1294 -547 1358 -483
rect 3969 -362 4033 -358
rect 3969 -418 3976 -362
rect 3976 -418 4032 -362
rect 4032 -418 4033 -362
rect 3969 -422 4033 -418
rect 4060 -362 4124 -358
rect 4060 -418 4116 -362
rect 4116 -418 4124 -362
rect 4060 -422 4124 -418
rect 2194 -673 2258 -609
rect 2322 -547 2386 -483
rect 1167 -919 1231 -855
rect 2322 -793 2386 -729
rect 2448 -673 2512 -609
rect 2448 -919 2512 -855
rect 4709 -1121 4773 -1057
rect 4789 -1121 4853 -1057
rect 4869 -1121 4933 -1057
rect 1744 -1447 1808 -1443
rect 1744 -1503 1748 -1447
rect 1748 -1503 1804 -1447
rect 1804 -1503 1808 -1447
rect 1744 -1507 1808 -1503
rect 4321 -1377 4545 -1373
rect 4321 -1513 4325 -1377
rect 4325 -1513 4541 -1377
rect 4541 -1513 4545 -1377
rect 4321 -1517 4545 -1513
rect -627 -2192 -563 -2188
rect -627 -2248 -623 -2192
rect -623 -2248 -567 -2192
rect -567 -2248 -563 -2192
rect -627 -2252 -563 -2248
rect -627 -2272 -563 -2268
rect -627 -2328 -623 -2272
rect -623 -2328 -567 -2272
rect -567 -2328 -563 -2272
rect -627 -2332 -563 -2328
rect -627 -2352 -563 -2348
rect -627 -2408 -623 -2352
rect -623 -2408 -567 -2352
rect -567 -2408 -563 -2352
rect -627 -2412 -563 -2408
rect -627 -2432 -563 -2428
rect -627 -2488 -623 -2432
rect -623 -2488 -567 -2432
rect -567 -2488 -563 -2432
rect -627 -2492 -563 -2488
rect 4321 -2417 4385 -2353
rect 4401 -2417 4465 -2353
rect 4481 -2417 4545 -2353
rect -627 -2512 -563 -2508
rect -627 -2568 -623 -2512
rect -623 -2568 -567 -2512
rect -567 -2568 -563 -2512
rect -627 -2572 -563 -2568
rect -626 -2747 -562 -2743
rect -626 -2803 -622 -2747
rect -622 -2803 -566 -2747
rect -566 -2803 -562 -2747
rect -626 -2807 -562 -2803
rect -626 -2827 -562 -2823
rect -626 -2883 -622 -2827
rect -622 -2883 -566 -2827
rect -566 -2883 -562 -2827
rect -626 -2887 -562 -2883
rect -626 -2907 -562 -2903
rect -626 -2963 -622 -2907
rect -622 -2963 -566 -2907
rect -566 -2963 -562 -2907
rect -626 -2967 -562 -2963
rect -626 -2987 -562 -2983
rect -626 -3043 -622 -2987
rect -622 -3043 -566 -2987
rect -566 -3043 -562 -2987
rect -626 -3047 -562 -3043
rect -626 -3067 -562 -3063
rect -626 -3123 -622 -3067
rect -622 -3123 -566 -3067
rect -566 -3123 -562 -3067
rect -626 -3127 -562 -3123
<< metal4 >>
rect -686 1962 -450 2000
rect -686 1898 -617 1962
rect -553 1898 -450 1962
rect -686 1882 -450 1898
rect -686 1818 -617 1882
rect -553 1818 -450 1882
rect -686 1802 -450 1818
rect -686 1738 -617 1802
rect -553 1738 -450 1802
rect -686 1722 -450 1738
rect -686 1658 -617 1722
rect -553 1658 -450 1722
rect -686 1642 -450 1658
rect 4268 1651 4588 2218
rect -686 1578 -617 1642
rect -553 1578 -450 1642
rect -686 1530 -450 1578
rect 3890 1530 4588 1651
rect -686 1402 -450 1450
rect -686 1338 -630 1402
rect -566 1338 -450 1402
rect -686 1322 -450 1338
rect -686 1258 -630 1322
rect -566 1258 -450 1322
rect -686 1242 -450 1258
rect -686 1178 -630 1242
rect -566 1178 -450 1242
rect -686 1162 -450 1178
rect -686 1098 -630 1162
rect -566 1098 -450 1162
rect -686 1082 -450 1098
rect -686 1018 -630 1082
rect -566 1018 -450 1082
rect -686 970 -450 1018
rect 4268 1240 4588 1530
rect 4268 1176 4321 1240
rect 4385 1176 4401 1240
rect 4465 1176 4481 1240
rect 4545 1176 4588 1240
rect 4268 890 4588 1176
rect 3890 769 4588 890
rect 1743 339 1809 340
rect 1743 275 1744 339
rect 1808 275 1809 339
rect 1743 274 1809 275
rect 1042 -483 1108 -482
rect 1042 -547 1043 -483
rect 1107 -488 1108 -483
rect 1293 -483 1359 -482
rect 1293 -488 1294 -483
rect 1107 -547 1294 -488
rect 1358 -488 1359 -483
rect 1746 -488 1806 274
rect 4268 -356 4588 769
rect 3963 -358 4588 -356
rect 3963 -422 3969 -358
rect 4033 -422 4060 -358
rect 4124 -422 4588 -358
rect 3963 -424 4588 -422
rect 2195 -488 2261 -482
rect 2321 -483 2387 -482
rect 2321 -488 2322 -483
rect 1358 -547 2322 -488
rect 2386 -488 2387 -483
rect 2386 -547 2513 -488
rect 1042 -548 2513 -547
rect 1042 -609 2513 -608
rect 1042 -668 1167 -609
rect 1166 -673 1167 -668
rect 1231 -668 2194 -609
rect 1231 -673 1232 -668
rect 1166 -674 1232 -673
rect 319 -729 563 -728
rect 319 -734 498 -729
rect -156 -793 498 -734
rect 562 -734 563 -729
rect 1042 -729 1108 -728
rect 1042 -734 1043 -729
rect 562 -793 1043 -734
rect 1107 -734 1108 -729
rect 1107 -793 1232 -734
rect -156 -794 1232 -793
rect -156 -855 1232 -854
rect -156 -914 320 -855
rect 319 -919 320 -914
rect 384 -914 1167 -855
rect 384 -919 563 -914
rect 319 -920 563 -919
rect 1166 -919 1167 -914
rect 1231 -919 1232 -855
rect 1166 -920 1232 -919
rect 1746 -1437 1806 -668
rect 2193 -673 2194 -668
rect 2258 -668 2448 -609
rect 2258 -673 2259 -668
rect 2193 -674 2259 -673
rect 2447 -673 2448 -668
rect 2512 -673 2513 -609
rect 2447 -674 2513 -673
rect 2321 -729 2387 -728
rect 2321 -793 2322 -729
rect 2386 -734 2387 -729
rect 2386 -793 2513 -734
rect 2321 -794 2513 -793
rect 2321 -855 2513 -854
rect 2321 -914 2448 -855
rect 2447 -919 2448 -914
rect 2512 -919 2513 -855
rect 2447 -920 2513 -919
rect 4268 -1373 4588 -424
rect 1743 -1443 1809 -1437
rect 1743 -1507 1744 -1443
rect 1808 -1507 1809 -1443
rect 1743 -1509 1809 -1507
rect 4268 -1517 4321 -1373
rect 4545 -1517 4588 -1373
rect 4268 -1939 4588 -1517
rect 3890 -2060 4588 -1939
rect -686 -2188 -450 -2140
rect -686 -2252 -627 -2188
rect -563 -2252 -450 -2188
rect -686 -2268 -450 -2252
rect -686 -2332 -627 -2268
rect -563 -2332 -450 -2268
rect -686 -2348 -450 -2332
rect -686 -2412 -627 -2348
rect -563 -2412 -450 -2348
rect -686 -2428 -450 -2412
rect -686 -2492 -627 -2428
rect -563 -2492 -450 -2428
rect -686 -2508 -450 -2492
rect -686 -2572 -627 -2508
rect -563 -2572 -450 -2508
rect -686 -2620 -450 -2572
rect 4268 -2353 4588 -2060
rect 4268 -2417 4321 -2353
rect 4385 -2417 4401 -2353
rect 4465 -2417 4481 -2353
rect 4545 -2417 4588 -2353
rect 4268 -2700 4588 -2417
rect -686 -2743 -450 -2700
rect -686 -2807 -626 -2743
rect -562 -2807 -450 -2743
rect -686 -2823 -450 -2807
rect 3890 -2821 4588 -2700
rect -686 -2887 -626 -2823
rect -562 -2887 -450 -2823
rect -686 -2903 -450 -2887
rect -686 -2967 -626 -2903
rect -562 -2967 -450 -2903
rect -686 -2983 -450 -2967
rect -686 -3047 -626 -2983
rect -562 -3047 -450 -2983
rect -686 -3063 -450 -3047
rect -686 -3127 -626 -3063
rect -562 -3127 -450 -3063
rect -686 -3170 -450 -3127
rect 4268 -3378 4588 -2821
rect 4658 347 4978 2218
rect 4658 203 4706 347
rect 4930 203 4978 347
rect 4658 -1057 4978 203
rect 4658 -1121 4709 -1057
rect 4773 -1121 4789 -1057
rect 4853 -1121 4869 -1057
rect 4933 -1121 4978 -1057
rect 4658 -3378 4978 -1121
use adc_comp_buffer  adc_comp_buffer_0
timestamp 1698999411
transform 1 0 2737 0 1 -192
box -68 -332 408 452
use adc_comp_buffer  adc_comp_buffer_1
timestamp 1698999411
transform 1 0 2737 0 -1 -860
box -68 -332 408 452
use adc_noise_decoup_cell2  adc_noise_decoup_cell2_0
timestamp 1698999411
transform 1 0 -450 0 1 -3170
box 0 0 4340 1580
use adc_noise_decoup_cell2  adc_noise_decoup_cell2_1
timestamp 1698999411
transform 1 0 -450 0 1 420
box 0 0 4340 1580
<< labels >>
flabel metal1 s 1272 -469 1318 -427 0 FreeSans 200 180 0 0 bp
port 1 nsew
flabel metal1 s 2235 -477 2281 -435 0 FreeSans 200 180 0 0 bn
port 2 nsew
flabel metal4 s 1427 -548 1487 -488 0 FreeSans 200 0 0 0 on
port 3 nsew
flabel metal4 s 1425 -668 1485 -608 0 FreeSans 200 0 0 0 op
port 4 nsew
flabel metal4 s 4658 -3378 4978 2218 0 FreeSans 1000 90 0 0 VPWR
port 5 nsew
flabel metal4 s 4268 -3378 4588 2218 0 FreeSans 1000 90 0 0 VGND
port 6 nsew
<< end >>
