magic
tech sky130A
magscale 1 2
timestamp 1695643842
<< error_p >>
rect -701 -538 -643 -532
rect -509 -538 -451 -532
rect -317 -538 -259 -532
rect -125 -538 -67 -532
rect 67 -538 125 -532
rect 259 -538 317 -532
rect 451 -538 509 -532
rect 643 -538 701 -532
rect -701 -572 -689 -538
rect -509 -572 -497 -538
rect -317 -572 -305 -538
rect -125 -572 -113 -538
rect 67 -572 79 -538
rect 259 -572 271 -538
rect 451 -572 463 -538
rect 643 -572 655 -538
rect -701 -578 -643 -572
rect -509 -578 -451 -572
rect -317 -578 -259 -572
rect -125 -578 -67 -572
rect 67 -578 125 -572
rect 259 -578 317 -572
rect 451 -578 509 -572
rect 643 -578 701 -572
<< pwell >>
rect -983 -710 983 710
<< nmos >>
rect -783 -500 -753 500
rect -687 -500 -657 500
rect -591 -500 -561 500
rect -495 -500 -465 500
rect -399 -500 -369 500
rect -303 -500 -273 500
rect -207 -500 -177 500
rect -111 -500 -81 500
rect -15 -500 15 500
rect 81 -500 111 500
rect 177 -500 207 500
rect 273 -500 303 500
rect 369 -500 399 500
rect 465 -500 495 500
rect 561 -500 591 500
rect 657 -500 687 500
rect 753 -500 783 500
<< ndiff >>
rect -845 488 -783 500
rect -845 -488 -833 488
rect -799 -488 -783 488
rect -845 -500 -783 -488
rect -753 488 -687 500
rect -753 -488 -737 488
rect -703 -488 -687 488
rect -753 -500 -687 -488
rect -657 488 -591 500
rect -657 -488 -641 488
rect -607 -488 -591 488
rect -657 -500 -591 -488
rect -561 488 -495 500
rect -561 -488 -545 488
rect -511 -488 -495 488
rect -561 -500 -495 -488
rect -465 488 -399 500
rect -465 -488 -449 488
rect -415 -488 -399 488
rect -465 -500 -399 -488
rect -369 488 -303 500
rect -369 -488 -353 488
rect -319 -488 -303 488
rect -369 -500 -303 -488
rect -273 488 -207 500
rect -273 -488 -257 488
rect -223 -488 -207 488
rect -273 -500 -207 -488
rect -177 488 -111 500
rect -177 -488 -161 488
rect -127 -488 -111 488
rect -177 -500 -111 -488
rect -81 488 -15 500
rect -81 -488 -65 488
rect -31 -488 -15 488
rect -81 -500 -15 -488
rect 15 488 81 500
rect 15 -488 31 488
rect 65 -488 81 488
rect 15 -500 81 -488
rect 111 488 177 500
rect 111 -488 127 488
rect 161 -488 177 488
rect 111 -500 177 -488
rect 207 488 273 500
rect 207 -488 223 488
rect 257 -488 273 488
rect 207 -500 273 -488
rect 303 488 369 500
rect 303 -488 319 488
rect 353 -488 369 488
rect 303 -500 369 -488
rect 399 488 465 500
rect 399 -488 415 488
rect 449 -488 465 488
rect 399 -500 465 -488
rect 495 488 561 500
rect 495 -488 511 488
rect 545 -488 561 488
rect 495 -500 561 -488
rect 591 488 657 500
rect 591 -488 607 488
rect 641 -488 657 488
rect 591 -500 657 -488
rect 687 488 753 500
rect 687 -488 703 488
rect 737 -488 753 488
rect 687 -500 753 -488
rect 783 488 845 500
rect 783 -488 799 488
rect 833 -488 845 488
rect 783 -500 845 -488
<< ndiffc >>
rect -833 -488 -799 488
rect -737 -488 -703 488
rect -641 -488 -607 488
rect -545 -488 -511 488
rect -449 -488 -415 488
rect -353 -488 -319 488
rect -257 -488 -223 488
rect -161 -488 -127 488
rect -65 -488 -31 488
rect 31 -488 65 488
rect 127 -488 161 488
rect 223 -488 257 488
rect 319 -488 353 488
rect 415 -488 449 488
rect 511 -488 545 488
rect 607 -488 641 488
rect 703 -488 737 488
rect 799 -488 833 488
<< psubdiff >>
rect -947 640 -851 674
rect 851 640 947 674
rect -947 578 -913 640
rect 913 578 947 640
rect -947 -640 -913 -578
rect 913 -640 947 -578
rect -947 -674 -851 -640
rect 851 -674 947 -640
<< psubdiffcont >>
rect -851 640 851 674
rect -947 -578 -913 578
rect 913 -578 947 578
rect -851 -674 851 -640
<< poly >>
rect -783 500 -753 526
rect -687 500 -657 526
rect -591 500 -561 526
rect -495 500 -465 526
rect -399 500 -369 526
rect -303 500 -273 526
rect -207 500 -177 526
rect -111 500 -81 526
rect -15 500 15 526
rect 81 500 111 526
rect 177 500 207 526
rect 273 500 303 526
rect 369 500 399 526
rect 465 500 495 526
rect 561 500 591 526
rect 657 500 687 526
rect 753 500 783 526
rect -783 -522 -753 -500
rect -687 -522 -657 -500
rect -591 -522 -561 -500
rect -495 -522 -465 -500
rect -399 -522 -369 -500
rect -303 -522 -273 -500
rect -207 -522 -177 -500
rect -111 -522 -81 -500
rect -15 -522 15 -500
rect 81 -522 111 -500
rect 177 -522 207 -500
rect 273 -522 303 -500
rect 369 -522 399 -500
rect 465 -522 495 -500
rect 561 -522 591 -500
rect 657 -522 687 -500
rect 753 -522 783 -500
rect -819 -538 -753 -522
rect -819 -572 -803 -538
rect -769 -572 -753 -538
rect -819 -588 -753 -572
rect -705 -538 705 -522
rect -705 -572 -689 -538
rect -655 -572 -497 -538
rect -463 -572 -305 -538
rect -271 -572 -113 -538
rect -79 -572 79 -538
rect 113 -572 271 -538
rect 305 -572 463 -538
rect 497 -572 655 -538
rect 689 -572 705 -538
rect -705 -588 705 -572
rect 753 -538 819 -522
rect 753 -572 769 -538
rect 803 -572 819 -538
rect 753 -588 819 -572
<< polycont >>
rect -803 -572 -769 -538
rect -689 -572 -655 -538
rect -497 -572 -463 -538
rect -305 -572 -271 -538
rect -113 -572 -79 -538
rect 79 -572 113 -538
rect 271 -572 305 -538
rect 463 -572 497 -538
rect 655 -572 689 -538
rect 769 -572 803 -538
<< locali >>
rect -947 640 -851 674
rect 851 640 947 674
rect -947 578 -913 640
rect 913 578 947 640
rect -833 488 -799 504
rect -833 -504 -799 -488
rect -737 488 -703 504
rect -737 -504 -703 -488
rect -641 488 -607 504
rect -641 -504 -607 -488
rect -545 488 -511 504
rect -545 -504 -511 -488
rect -449 488 -415 504
rect -449 -504 -415 -488
rect -353 488 -319 504
rect -353 -504 -319 -488
rect -257 488 -223 504
rect -257 -504 -223 -488
rect -161 488 -127 504
rect -161 -504 -127 -488
rect -65 488 -31 504
rect -65 -504 -31 -488
rect 31 488 65 504
rect 31 -504 65 -488
rect 127 488 161 504
rect 127 -504 161 -488
rect 223 488 257 504
rect 223 -504 257 -488
rect 319 488 353 504
rect 319 -504 353 -488
rect 415 488 449 504
rect 415 -504 449 -488
rect 511 488 545 504
rect 511 -504 545 -488
rect 607 488 641 504
rect 607 -504 641 -488
rect 703 488 737 504
rect 703 -504 737 -488
rect 799 488 833 504
rect 799 -504 833 -488
rect -819 -572 -803 -538
rect -769 -572 -753 -538
rect -705 -572 -689 -538
rect -655 -572 -639 -538
rect -513 -572 -497 -538
rect -463 -572 -447 -538
rect -321 -572 -305 -538
rect -271 -572 -255 -538
rect -129 -572 -113 -538
rect -79 -572 -63 -538
rect 63 -572 79 -538
rect 113 -572 129 -538
rect 255 -572 271 -538
rect 305 -572 321 -538
rect 447 -572 463 -538
rect 497 -572 513 -538
rect 639 -572 655 -538
rect 689 -572 705 -538
rect 753 -572 769 -538
rect 803 -572 819 -538
rect -947 -640 -913 -578
rect 913 -640 947 -578
rect -947 -674 -851 -640
rect 851 -674 947 -640
<< viali >>
rect -833 -488 -799 488
rect -737 -488 -703 488
rect -641 -488 -607 488
rect -545 -488 -511 488
rect -449 -488 -415 488
rect -353 -488 -319 488
rect -257 -488 -223 488
rect -161 -488 -127 488
rect -65 -488 -31 488
rect 31 -488 65 488
rect 127 -488 161 488
rect 223 -488 257 488
rect 319 -488 353 488
rect 415 -488 449 488
rect 511 -488 545 488
rect 607 -488 641 488
rect 703 -488 737 488
rect 799 -488 833 488
rect -689 -572 -655 -538
rect -497 -572 -463 -538
rect -305 -572 -271 -538
rect -113 -572 -79 -538
rect 79 -572 113 -538
rect 271 -572 305 -538
rect 463 -572 497 -538
rect 655 -572 689 -538
<< metal1 >>
rect -839 488 -793 500
rect -839 -488 -833 488
rect -799 -488 -793 488
rect -839 -500 -793 -488
rect -743 488 -697 500
rect -743 -488 -737 488
rect -703 -488 -697 488
rect -743 -500 -697 -488
rect -647 488 -601 500
rect -647 -488 -641 488
rect -607 -488 -601 488
rect -647 -500 -601 -488
rect -551 488 -505 500
rect -551 -488 -545 488
rect -511 -488 -505 488
rect -551 -500 -505 -488
rect -455 488 -409 500
rect -455 -488 -449 488
rect -415 -488 -409 488
rect -455 -500 -409 -488
rect -359 488 -313 500
rect -359 -488 -353 488
rect -319 -488 -313 488
rect -359 -500 -313 -488
rect -263 488 -217 500
rect -263 -488 -257 488
rect -223 -488 -217 488
rect -263 -500 -217 -488
rect -167 488 -121 500
rect -167 -488 -161 488
rect -127 -488 -121 488
rect -167 -500 -121 -488
rect -71 488 -25 500
rect -71 -488 -65 488
rect -31 -488 -25 488
rect -71 -500 -25 -488
rect 25 488 71 500
rect 25 -488 31 488
rect 65 -488 71 488
rect 25 -500 71 -488
rect 121 488 167 500
rect 121 -488 127 488
rect 161 -488 167 488
rect 121 -500 167 -488
rect 217 488 263 500
rect 217 -488 223 488
rect 257 -488 263 488
rect 217 -500 263 -488
rect 313 488 359 500
rect 313 -488 319 488
rect 353 -488 359 488
rect 313 -500 359 -488
rect 409 488 455 500
rect 409 -488 415 488
rect 449 -488 455 488
rect 409 -500 455 -488
rect 505 488 551 500
rect 505 -488 511 488
rect 545 -488 551 488
rect 505 -500 551 -488
rect 601 488 647 500
rect 601 -488 607 488
rect 641 -488 647 488
rect 601 -500 647 -488
rect 697 488 743 500
rect 697 -488 703 488
rect 737 -488 743 488
rect 697 -500 743 -488
rect 793 488 839 500
rect 793 -488 799 488
rect 833 -488 839 488
rect 793 -500 839 -488
rect -701 -538 -643 -532
rect -701 -572 -689 -538
rect -655 -572 -643 -538
rect -701 -578 -643 -572
rect -509 -538 -451 -532
rect -509 -572 -497 -538
rect -463 -572 -451 -538
rect -509 -578 -451 -572
rect -317 -538 -259 -532
rect -317 -572 -305 -538
rect -271 -572 -259 -538
rect -317 -578 -259 -572
rect -125 -538 -67 -532
rect -125 -572 -113 -538
rect -79 -572 -67 -538
rect -125 -578 -67 -572
rect 67 -538 125 -532
rect 67 -572 79 -538
rect 113 -572 125 -538
rect 67 -578 125 -572
rect 259 -538 317 -532
rect 259 -572 271 -538
rect 305 -572 317 -538
rect 259 -578 317 -572
rect 451 -538 509 -532
rect 451 -572 463 -538
rect 497 -572 509 -538
rect 451 -578 509 -572
rect 643 -538 701 -532
rect 643 -572 655 -538
rect 689 -572 701 -538
rect 643 -578 701 -572
<< properties >>
string FIXED_BBOX -930 -657 930 657
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 5 l 0.150 m 1 nf 17 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
