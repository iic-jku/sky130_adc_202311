magic
tech sky130A
magscale 1 2
timestamp 1515178157
<< checkpaint >>
rect -1212 8512 2818 22558
<< pwell >>
rect 624 15490 1094 15704
rect 690 15234 1022 15490
<< nmos >>
rect 788 15260 930 15398
<< ndiff >>
rect 716 15380 788 15398
rect 716 15346 736 15380
rect 770 15346 788 15380
rect 716 15312 788 15346
rect 716 15278 736 15312
rect 770 15278 788 15312
rect 716 15260 788 15278
rect 930 15379 996 15398
rect 930 15345 946 15379
rect 980 15345 996 15379
rect 930 15311 996 15345
rect 930 15277 946 15311
rect 980 15277 996 15311
rect 930 15260 996 15277
<< ndiffc >>
rect 736 15346 770 15380
rect 736 15278 770 15312
rect 946 15345 980 15379
rect 946 15277 980 15311
<< psubdiff >>
rect 650 15610 1068 15678
rect 650 15576 741 15610
rect 775 15576 809 15610
rect 843 15576 877 15610
rect 911 15576 945 15610
rect 979 15576 1068 15610
rect 650 15516 1068 15576
<< psubdiffcont >>
rect 741 15576 775 15610
rect 809 15576 843 15610
rect 877 15576 911 15610
rect 945 15576 979 15610
<< poly >>
rect 788 15398 930 15448
rect 788 15199 930 15260
rect 788 15165 808 15199
rect 842 15165 876 15199
rect 910 15165 930 15199
rect 788 15140 930 15165
<< polycont >>
rect 808 15165 842 15199
rect 876 15165 910 15199
<< locali >>
rect 658 15648 1068 15674
rect 658 15542 738 15648
rect 988 15542 1068 15648
rect 658 15514 1068 15542
rect 728 15380 782 15514
rect 940 15414 988 15514
rect 728 15346 736 15380
rect 770 15346 782 15380
rect 728 15312 782 15346
rect 728 15278 736 15312
rect 770 15278 782 15312
rect 728 15252 782 15278
rect 934 15379 988 15414
rect 934 15345 946 15379
rect 980 15345 988 15379
rect 934 15311 988 15345
rect 934 15277 946 15311
rect 980 15277 988 15311
rect 934 15252 988 15277
rect 788 15199 930 15218
rect 788 15197 808 15199
rect 788 15163 806 15197
rect 842 15165 876 15199
rect 910 15197 930 15199
rect 840 15163 878 15165
rect 912 15163 930 15197
rect 788 15140 930 15163
<< viali >>
rect 738 15610 988 15648
rect 738 15576 741 15610
rect 741 15576 775 15610
rect 775 15576 809 15610
rect 809 15576 843 15610
rect 843 15576 877 15610
rect 877 15576 911 15610
rect 911 15576 945 15610
rect 945 15576 979 15610
rect 979 15576 988 15610
rect 738 15542 988 15576
rect 806 15165 808 15197
rect 808 15165 840 15197
rect 878 15165 910 15197
rect 910 15165 912 15197
rect 806 15163 840 15165
rect 878 15163 912 15165
<< metal1 >>
rect 658 15648 1068 15674
rect 658 15621 738 15648
rect 988 15621 1068 15648
rect 658 15569 709 15621
rect 1017 15569 1068 15621
rect 658 15542 738 15569
rect 988 15542 1068 15569
rect 658 15514 1068 15542
rect 788 15206 930 15218
rect 788 15197 833 15206
rect 885 15197 930 15206
rect 788 15163 806 15197
rect 912 15163 930 15197
rect 788 15154 833 15163
rect 885 15154 930 15163
rect 788 15140 930 15154
<< via1 >>
rect 709 15569 738 15621
rect 738 15569 761 15621
rect 773 15569 825 15621
rect 837 15569 889 15621
rect 901 15569 953 15621
rect 965 15569 988 15621
rect 988 15569 1017 15621
rect 833 15197 885 15206
rect 833 15163 840 15197
rect 840 15163 878 15197
rect 878 15163 885 15197
rect 833 15154 885 15163
<< metal2 >>
rect 658 15623 1068 15674
rect 658 15621 715 15623
rect 771 15621 795 15623
rect 851 15621 875 15623
rect 931 15621 955 15623
rect 1011 15621 1068 15623
rect 658 15569 709 15621
rect 771 15569 773 15621
rect 953 15569 955 15621
rect 1017 15569 1068 15621
rect 658 15567 715 15569
rect 771 15567 795 15569
rect 851 15567 875 15569
rect 931 15567 955 15569
rect 1011 15567 1068 15569
rect 658 15514 1068 15567
rect 788 15208 930 15218
rect 788 15152 831 15208
rect 887 15152 930 15208
rect 788 15140 930 15152
<< via2 >>
rect 715 15621 771 15623
rect 795 15621 851 15623
rect 875 15621 931 15623
rect 955 15621 1011 15623
rect 715 15569 761 15621
rect 761 15569 771 15621
rect 795 15569 825 15621
rect 825 15569 837 15621
rect 837 15569 851 15621
rect 875 15569 889 15621
rect 889 15569 901 15621
rect 901 15569 931 15621
rect 955 15569 965 15621
rect 965 15569 1011 15621
rect 715 15567 771 15569
rect 795 15567 851 15569
rect 875 15567 931 15569
rect 955 15567 1011 15569
rect 831 15206 887 15208
rect 831 15154 833 15206
rect 833 15154 885 15206
rect 885 15154 887 15206
rect 831 15152 887 15154
<< metal3 >>
rect 50 15630 1558 15676
rect 50 15566 171 15630
rect 235 15566 251 15630
rect 315 15566 331 15630
rect 395 15566 411 15630
rect 475 15623 1558 15630
rect 475 15567 715 15623
rect 771 15567 795 15623
rect 851 15567 875 15623
rect 931 15567 955 15623
rect 1011 15567 1558 15623
rect 475 15566 1558 15567
rect 50 15514 1558 15566
rect 48 15362 1556 15412
rect 48 15298 1095 15362
rect 1159 15298 1175 15362
rect 1239 15298 1255 15362
rect 1319 15298 1335 15362
rect 1399 15298 1556 15362
rect 48 15250 1556 15298
rect 788 15208 930 15250
rect 788 15152 831 15208
rect 887 15152 930 15208
rect 788 15140 930 15152
<< via3 >>
rect 171 15566 235 15630
rect 251 15566 315 15630
rect 331 15566 395 15630
rect 411 15566 475 15630
rect 1095 15298 1159 15362
rect 1175 15298 1239 15362
rect 1255 15298 1319 15362
rect 1335 15298 1399 15362
<< metal4 >>
rect 144 15630 502 21290
rect 144 15566 171 15630
rect 235 15566 251 15630
rect 315 15566 331 15630
rect 395 15566 411 15630
rect 475 15566 502 15630
rect 144 9772 502 15566
rect 1068 15362 1426 21298
rect 1068 15298 1095 15362
rect 1159 15298 1175 15362
rect 1239 15298 1255 15362
rect 1319 15298 1335 15362
rect 1399 15298 1426 15362
rect 1068 9780 1426 15298
<< labels >>
flabel metal4 s 144 9772 502 21290 0 FreeSans 2000 0 0 0 VSS
port 1 nsew
flabel metal4 s 1068 9780 1424 21298 0 FreeSans 2000 0 0 0 VDD
port 2 nsew
<< properties >>
string FIXED_BBOX 0 0 1600 32000
string GDS_END 734862
string GDS_FILE adc_top.gds.gz
string GDS_START 730762
<< end >>
