magic
tech sky130A
magscale 1 2
timestamp 1697705955
<< pwell >>
rect -134 188 -24 938
rect 1050 188 1160 938
rect 30 14 96 150
rect 930 14 996 150
<< locali >>
rect -134 188 16 938
rect 1010 188 1160 938
rect 30 14 96 150
rect 930 14 996 150
<< metal1 >>
rect 9 1300 57 1588
rect 103 1582 155 1588
rect 103 1476 155 1482
rect 7 1294 59 1300
rect 7 1188 59 1194
rect 9 926 57 1188
rect 105 926 153 1476
rect 201 1444 249 1588
rect 199 1438 251 1444
rect 199 1332 251 1338
rect 201 926 249 1332
rect 297 1300 345 1588
rect 393 1444 441 1588
rect 487 1582 539 1588
rect 487 1476 539 1482
rect 391 1438 443 1444
rect 391 1332 443 1338
rect 295 1294 347 1300
rect 295 1188 347 1194
rect 297 926 345 1188
rect 393 926 441 1332
rect 489 926 537 1476
rect 585 1444 633 1588
rect 583 1438 635 1444
rect 583 1332 635 1338
rect 585 926 633 1332
rect 681 1300 729 1588
rect 777 1444 825 1588
rect 871 1582 923 1588
rect 871 1476 923 1482
rect 775 1438 827 1444
rect 775 1332 827 1338
rect 679 1294 731 1300
rect 679 1188 731 1194
rect 681 926 729 1188
rect 777 926 825 1332
rect 873 926 921 1476
rect 969 1300 1017 1588
rect 967 1294 1019 1300
rect 967 1188 1019 1194
rect 969 926 1017 1188
rect 153 -206 201 156
rect 258 110 384 156
rect 450 110 576 156
rect 642 110 768 156
rect 321 -62 369 110
rect 319 -68 371 -62
rect 319 -174 371 -168
rect 151 -212 203 -206
rect 151 -318 203 -312
rect 321 -318 369 -174
rect 489 -206 537 110
rect 657 -62 705 110
rect 655 -68 707 -62
rect 655 -174 707 -168
rect 487 -212 539 -206
rect 487 -318 539 -312
rect 657 -318 705 -174
rect 825 -206 873 156
rect 823 -212 875 -206
rect 823 -318 875 -312
<< via1 >>
rect 103 1482 155 1582
rect 7 1194 59 1294
rect 199 1338 251 1438
rect 487 1482 539 1582
rect 391 1338 443 1438
rect 295 1194 347 1294
rect 583 1338 635 1438
rect 871 1482 923 1582
rect 775 1338 827 1438
rect 679 1194 731 1294
rect 967 1194 1019 1294
rect 319 -168 371 -68
rect 151 -312 203 -212
rect 655 -168 707 -68
rect 487 -312 539 -212
rect 823 -312 875 -212
<< metal2 >>
rect 103 1582 155 1588
rect -134 1484 103 1580
rect 487 1582 539 1588
rect 155 1484 487 1580
rect 103 1476 155 1482
rect 871 1582 923 1588
rect 539 1484 871 1580
rect 487 1476 539 1482
rect 923 1484 1160 1580
rect 871 1476 923 1482
rect 199 1438 251 1444
rect -134 1340 199 1436
rect 391 1438 443 1444
rect 251 1340 391 1436
rect 199 1332 251 1338
rect 583 1438 635 1444
rect 443 1340 583 1436
rect 391 1332 443 1338
rect 775 1438 827 1444
rect 635 1340 775 1436
rect 583 1332 635 1338
rect 827 1340 1160 1436
rect 775 1332 827 1338
rect 7 1294 59 1300
rect -134 1196 7 1292
rect 295 1294 347 1300
rect 59 1196 295 1292
rect 7 1188 59 1194
rect 679 1294 731 1300
rect 347 1196 679 1292
rect 295 1188 347 1194
rect 967 1294 1019 1300
rect 731 1196 967 1292
rect 679 1188 731 1194
rect 1019 1196 1160 1292
rect 967 1188 1019 1194
rect 319 -68 371 -62
rect -134 -166 319 -70
rect 655 -68 707 -62
rect 371 -166 655 -70
rect 319 -174 371 -168
rect 707 -166 1160 -70
rect 655 -174 707 -168
rect 151 -212 203 -206
rect -134 -310 151 -214
rect 487 -212 539 -206
rect 203 -310 487 -214
rect 151 -318 203 -312
rect 823 -212 875 -206
rect 539 -310 823 -214
rect 487 -318 539 -312
rect 875 -310 1160 -214
rect 823 -318 875 -312
use sky130_fd_pr__nfet_01v8_QMBXET  sky130_fd_pr__nfet_01v8_QMBXET_0
timestamp 1697705955
transform 1 0 513 0 1 563
box -647 -585 647 585
<< labels >>
flabel locali -134 188 16 938 0 FreeSans 320 0 0 0 VSUB
port 0 nsew
flabel locali 1010 188 1160 938 0 FreeSans 320 0 0 0 VSUB
port 0 nsew
flabel metal2 -134 1484 1160 1580 0 FreeSans 400 0 0 0 M1D
port 3 nsew
flabel metal2 -134 -310 1160 -214 0 FreeSans 400 0 0 0 M1G
port 1 nsew
flabel metal2 -134 -166 1160 -70 0 FreeSans 400 0 0 0 M2G
port 2 nsew
<< end >>
