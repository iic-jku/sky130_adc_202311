magic
tech sky130A
magscale 1 2
timestamp 1699097993
<< error_s >>
rect 582340 640944 582394 640978
rect 584806 640944 584860 641038
rect 582340 630826 582394 630918
rect 584806 630826 584860 630978
rect 582340 182510 582394 182644
rect 584806 182510 584860 182704
<< metal3 >>
rect 582334 640944 582340 643404
rect 584800 640944 584806 643404
rect 582334 630826 582340 633286
rect 584800 630826 584806 633286
rect 582186 589482 582830 589542
rect 583014 589482 583520 589542
rect 582388 500138 583028 500140
rect 582388 500114 583034 500138
rect 582418 500080 583034 500114
rect 583200 500080 583520 500140
rect 582454 455652 583018 455712
rect 583200 455652 583520 455712
rect 582540 411272 583046 411274
rect 581312 411248 583046 411272
rect 581358 411238 583046 411248
rect 581358 411212 583036 411238
rect 583220 411212 583520 411272
rect 580752 364796 582996 364858
rect 583186 364796 583520 364858
rect 582554 319578 583032 319638
rect 583210 319578 583520 319638
rect 582406 275156 583038 275216
rect 583224 275156 583520 275216
rect 582334 182510 582340 184970
rect 584800 182510 584806 184970
rect 583104 95152 583238 95212
rect 583416 95152 583520 95212
rect 583024 50484 583276 50544
rect 583448 50484 583520 50544
use adc_wrapper  adc_wrapper_0
timestamp 1699054381
transform 1 0 483822 0 1 345788
box -21565 -296491 100978 298237
use sky130_fd_pr__res_generic_m3_R56YQM  sky130_fd_pr__res_generic_m3_R56YQM_0
timestamp 1699054381
transform 0 1 582923 -1 0 589512
box -30 -117 30 117
use sky130_fd_pr__res_generic_m3_R56YQM  sky130_fd_pr__res_generic_m3_R56YQM_1
timestamp 1699054381
transform 0 1 583361 -1 0 50514
box -30 -117 30 117
use sky130_fd_pr__res_generic_m3_R56YQM  sky130_fd_pr__res_generic_m3_R56YQM_2
timestamp 1699054381
transform 0 1 583333 -1 0 95182
box -30 -117 30 117
use sky130_fd_pr__res_generic_m3_R56YQM  sky130_fd_pr__res_generic_m3_R56YQM_3
timestamp 1699054381
transform 0 1 583133 -1 0 275186
box -30 -117 30 117
use sky130_fd_pr__res_generic_m3_R56YQM  sky130_fd_pr__res_generic_m3_R56YQM_4
timestamp 1699054381
transform 0 1 583121 -1 0 319608
box -30 -117 30 117
use sky130_fd_pr__res_generic_m3_R56YQM  sky130_fd_pr__res_generic_m3_R56YQM_5
timestamp 1699054381
transform 0 1 583095 -1 0 364828
box -30 -117 30 117
use sky130_fd_pr__res_generic_m3_R56YQM  sky130_fd_pr__res_generic_m3_R56YQM_6
timestamp 1699054381
transform 0 1 583129 -1 0 411242
box -30 -117 30 117
use sky130_fd_pr__res_generic_m3_R56YQM  sky130_fd_pr__res_generic_m3_R56YQM_7
timestamp 1699054381
transform 0 1 583107 -1 0 455682
box -30 -117 30 117
use sky130_fd_pr__res_generic_m3_R56YQM  sky130_fd_pr__res_generic_m3_R56YQM_8
timestamp 1699054381
transform 0 1 583111 -1 0 500110
box -30 -117 30 117
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
