magic
tech sky130A
magscale 1 2
timestamp 1699972208
<< nwell >>
rect 1021 22396 2579 22717
rect -177 2754 3825 3075
rect -179 1239 26 1341
rect 3610 1239 3825 1341
rect -179 1152 55 1239
rect 3578 1152 3825 1239
rect -179 1020 26 1152
rect 3610 1020 3825 1152
<< pwell >>
rect 1021 22775 2579 23018
rect -175 3159 3825 3376
rect -175 3133 3344 3159
rect 3524 3133 3825 3159
rect -175 1618 95 1642
rect 3572 1618 3825 1642
rect -175 1399 3825 1618
<< psubdiff >>
rect 1140 22944 1184 22968
rect 1140 22802 1184 22826
rect 2416 22944 2460 22968
rect 2416 22802 2460 22826
rect -96 3302 -52 3326
rect -96 3160 -52 3184
rect 3662 3302 3706 3326
rect 3662 3160 3706 3184
rect -96 1568 -52 1592
rect -96 1426 -52 1450
rect 3662 1568 3706 1592
rect 3662 1426 3706 1450
<< nsubdiff >>
rect 1091 22531 1115 22618
rect 1265 22531 1289 22618
rect 2344 22531 2368 22618
rect 2518 22531 2542 22618
rect -141 2911 -117 2998
rect 33 2911 57 2998
rect 3578 2911 3602 2998
rect 3752 2911 3776 2998
rect -143 1152 -119 1239
rect 31 1152 55 1239
rect 3578 1152 3602 1239
rect 3752 1152 3776 1239
<< psubdiffcont >>
rect 1140 22826 1184 22944
rect 2416 22826 2460 22944
rect -96 3184 -52 3302
rect 3662 3184 3706 3302
rect -96 1450 -52 1568
rect 3662 1450 3706 1568
<< nsubdiffcont >>
rect 1115 22531 1265 22618
rect 2368 22531 2518 22618
rect -117 2911 33 2998
rect 3602 2911 3752 2998
rect -119 1152 31 1239
rect 3602 1152 3752 1239
<< locali >>
rect 1135 22962 1401 22970
rect 2262 22962 2465 22976
rect 1135 22944 1494 22962
rect 1135 22826 1140 22944
rect 1184 22826 1494 22944
rect 1135 22770 1494 22826
rect 1348 22762 1494 22770
rect 2116 22944 2465 22962
rect 2116 22826 2416 22944
rect 2460 22826 2465 22944
rect 2116 22770 2465 22826
rect 2116 22762 2262 22770
rect 1700 22716 1860 22760
rect 2245 22618 2380 22654
rect 1091 22531 1115 22618
rect 1265 22531 1289 22618
rect 1236 22426 1289 22531
rect 2245 22531 2368 22618
rect 2518 22531 2542 22618
rect 2245 22500 2380 22531
rect 2216 22435 2380 22500
rect 1236 22417 1282 22426
rect 1088 21829 1418 21932
rect 2190 21829 2520 21932
rect 962 21482 1042 21782
rect 1464 21482 1544 21782
rect 1950 21482 2030 21782
rect 2064 21482 2144 21782
rect 2566 21482 2646 21782
rect 962 20750 1042 20850
rect 1164 20750 1244 20850
rect 1278 20750 1358 20850
rect 2364 20750 2444 20850
rect 2566 20750 2646 20850
rect 1070 20610 1136 20712
rect 2472 20610 2538 20712
rect 1223 20440 1563 20576
rect 763 20420 1563 20440
rect 763 6974 783 20420
rect 1223 20230 1563 20420
rect 2045 20440 2385 20576
rect 1657 20268 1723 20370
rect 1885 20268 1951 20370
rect 2045 20230 2845 20440
rect 1223 20030 1739 20230
rect 1965 20030 2845 20230
rect 1223 19208 1563 20030
rect 1643 20029 1739 20030
rect 1657 19246 1723 19348
rect 1885 19246 1951 19348
rect 2045 19208 2845 20030
rect 1223 19008 1739 19208
rect 1965 19008 2845 19208
rect 1223 18186 1563 19008
rect 1643 19007 1739 19008
rect 1657 18224 1723 18326
rect 1885 18224 1951 18326
rect 2045 18186 2845 19008
rect 1223 17986 1739 18186
rect 1965 17986 2845 18186
rect 1223 17034 1563 17986
rect 1643 17985 1739 17986
rect 1657 17072 1723 17174
rect 1885 17072 1951 17174
rect 2045 17034 2845 17986
rect 1223 16834 1739 17034
rect 1965 16834 2845 17034
rect 1223 16012 1563 16834
rect 1643 16833 1739 16834
rect 1657 16050 1723 16152
rect 1885 16050 1951 16152
rect 2045 16012 2845 16834
rect 1223 15812 1739 16012
rect 1965 15812 2845 16012
rect 1223 14860 1563 15812
rect 1643 15811 1739 15812
rect 1657 14898 1723 15000
rect 1885 14898 1951 15000
rect 2045 14860 2845 15812
rect 1223 14660 1739 14860
rect 1965 14660 2845 14860
rect 1223 12816 1563 14660
rect 1643 14659 1739 14660
rect 1657 12854 1723 12956
rect 1885 12854 1951 12956
rect 2045 12816 2845 14660
rect 1223 12616 1739 12816
rect 1965 12616 2845 12816
rect 1223 10642 1563 12616
rect 1643 12615 1739 12616
rect 1657 10680 1723 10782
rect 1885 10680 1951 10782
rect 2045 10642 2845 12616
rect 1223 10442 1739 10642
rect 1965 10442 2845 10642
rect 1223 8598 1563 10442
rect 1643 10441 1739 10442
rect 1657 8636 1723 8738
rect 1885 8636 1951 8738
rect 2045 8598 2845 10442
rect 1223 8398 1739 8598
rect 1965 8398 2845 8598
rect 1223 6974 1563 8398
rect 1643 8397 1739 8398
rect 763 6954 1563 6974
rect 2045 6954 2845 8398
rect 763 6238 1243 6954
rect 1349 5697 1499 5897
rect 2013 5697 2259 5897
rect 1522 5548 1570 5650
rect 2038 5548 2086 5650
rect 1349 4374 1499 4388
rect 1349 4298 1364 4374
rect 1424 4298 1499 4374
rect 1349 4288 1499 4298
rect 2013 4288 2259 4388
rect 1522 4148 1570 4250
rect 2038 4148 2086 4250
rect -96 3322 82 3326
rect -96 3320 198 3322
rect -96 3302 250 3320
rect -52 3184 250 3302
rect -96 3166 250 3184
rect 104 3104 250 3166
rect 360 3104 506 3320
rect 3136 3288 3250 3334
rect 710 3072 918 3120
rect 1222 3072 1430 3120
rect 2190 3072 2388 3120
rect 2692 3072 2900 3120
rect 3104 3118 3250 3288
rect 3360 3302 3711 3334
rect 3360 3184 3662 3302
rect 3706 3184 3711 3302
rect 3360 3159 3711 3184
rect 3360 3118 3506 3159
rect -141 2911 -117 2998
rect 33 2911 57 2998
rect 3578 2911 3602 2998
rect 3752 2911 3776 2998
rect 3602 2809 3646 2911
rect -16 2775 38 2809
rect 3572 2775 3646 2809
rect -96 1586 108 1592
rect 3477 1586 3711 1600
rect -96 1568 248 1586
rect -52 1450 248 1568
rect -96 1432 248 1450
rect 102 1370 248 1432
rect 3360 1568 3711 1586
rect 3360 1450 3662 1568
rect 3706 1450 3711 1568
rect 438 1350 615 1386
rect 1934 1376 2002 1378
rect 1934 1340 1950 1376
rect 1984 1340 2002 1376
rect 1934 1322 2002 1340
rect 2750 1331 2804 1405
rect 3360 1394 3711 1450
rect 3016 1350 3156 1386
rect 3360 1370 3506 1394
rect -143 1152 -119 1239
rect 31 1152 55 1239
rect 3578 1152 3602 1239
rect 3752 1152 3776 1239
rect -16 1075 31 1152
rect 3602 1075 3650 1152
rect -16 1041 36 1075
rect 3572 1041 3650 1075
<< viali >>
rect 1588 22718 1622 22752
rect 1958 22726 1992 22760
rect 783 6974 1223 20420
rect 1364 4298 1424 4374
rect 597 3079 631 3123
rect 981 3075 1015 3119
rect 1102 3078 1136 3122
rect 1486 3080 1520 3120
rect 1612 3082 1646 3116
rect 1725 3080 1759 3114
rect 1948 3078 1982 3122
rect 2088 3080 2122 3120
rect 2460 3078 2494 3122
rect 2596 3076 2630 3120
rect 2972 3078 3006 3122
rect 346 1338 380 1374
rect 738 1336 772 1372
rect 860 1338 894 1374
rect 988 1338 1022 1374
rect 1798 1340 1832 1376
rect 1950 1340 1984 1376
rect 2070 1334 2104 1370
rect 2836 1336 2870 1372
rect 3228 1336 3262 1372
rect 1500 1210 1534 1246
<< metal1 >>
rect -38 22996 3646 23026
rect -38 22756 -8 22996
rect 412 22930 3646 22996
rect 412 22756 442 22930
rect -38 22726 442 22756
rect 1566 22772 1638 22780
rect 1566 22716 1574 22772
rect 1630 22716 1638 22772
rect 1566 22708 1638 22716
rect 1950 22772 2022 22780
rect 1950 22716 1958 22772
rect 2014 22716 2022 22772
rect 1950 22708 2022 22716
rect -38 22452 3646 22482
rect -38 22386 3196 22452
rect 3166 22212 3196 22386
rect 3616 22212 3646 22452
rect 3166 22182 3646 22212
rect 1714 21882 1894 21888
rect 1714 21869 1720 21882
rect 1704 21830 1720 21869
rect 1888 21869 1894 21882
rect 1888 21830 1904 21869
rect 1704 21823 1904 21830
rect -38 21482 1042 21782
rect 1351 20850 1399 21334
rect 1651 21150 1699 21482
rect 1780 21294 1828 21823
rect 2572 21752 3646 21782
rect 2572 21512 3196 21752
rect 3616 21512 3646 21752
rect 2572 21482 3646 21512
rect 1778 21288 1830 21294
rect 1778 21182 1830 21188
rect 1649 21144 1701 21150
rect 1649 21038 1701 21044
rect 1651 20998 1699 21038
rect 1780 20718 1828 21182
rect 1909 20998 1957 21482
rect 2209 21150 2257 21334
rect 2207 21144 2259 21150
rect 2207 21038 2259 21044
rect 2209 20850 2257 21038
rect 1404 20672 2204 20718
rect -38 20420 1243 20440
rect -38 20410 783 20420
rect -38 20170 -8 20410
rect 412 20170 783 20410
rect -38 20140 783 20170
rect 763 6974 783 20140
rect 1223 6974 1243 20420
rect 1813 20218 1891 20224
rect 1813 20042 1819 20218
rect 1885 20042 1891 20218
rect 2210 20140 2365 20440
rect 2845 20140 3646 20440
rect 1813 20036 1891 20042
rect 1293 19952 1837 19998
rect 1813 19196 1891 19202
rect 1813 19020 1819 19196
rect 1885 19020 1891 19196
rect 1813 19014 1891 19020
rect 1293 18930 1837 18976
rect 1813 18174 1891 18180
rect 1813 17998 1819 18174
rect 1885 17998 1891 18174
rect 1813 17992 1891 17998
rect 1293 17908 1837 17954
rect 1813 17022 1891 17028
rect 1813 16846 1819 17022
rect 1885 16846 1891 17022
rect 1813 16840 1891 16846
rect 1293 16756 1837 16802
rect 1393 15780 1439 16756
rect 1813 16000 1891 16006
rect 1813 15824 1819 16000
rect 1885 15824 1891 16000
rect 1813 15818 1891 15824
rect 1393 15734 1837 15780
rect 1813 14848 1891 14854
rect 1813 14672 1819 14848
rect 1885 14672 1891 14848
rect 1813 14666 1891 14672
rect 1293 14582 1837 14628
rect 1393 12584 1439 14582
rect 1813 12804 1891 12810
rect 1813 12628 1819 12804
rect 1885 12628 1891 12804
rect 1813 12622 1891 12628
rect 1393 12538 1837 12584
rect 1813 10630 1891 10636
rect 1813 10454 1819 10630
rect 1885 10454 1891 10630
rect 1813 10448 1891 10454
rect 1293 10364 1837 10410
rect 1393 8366 1439 10364
rect 1813 8586 1891 8592
rect 1813 8410 1819 8586
rect 1885 8410 1891 8586
rect 1813 8404 1891 8410
rect 1393 8320 1837 8366
rect 763 3384 1243 6974
rect 1396 6410 1444 6554
rect 1394 6404 1446 6410
rect 1394 6302 1446 6308
rect 1396 5292 1444 6302
rect 1492 5888 1540 6554
rect 1588 6410 1636 6554
rect 1682 6548 1734 6554
rect 1682 6446 1734 6452
rect 1586 6404 1638 6410
rect 1586 6302 1638 6308
rect 1588 5888 1636 6302
rect 1684 5888 1732 6446
rect 1780 6266 1828 6554
rect 1874 6548 1926 6554
rect 1874 6446 1926 6452
rect 1778 6260 1830 6266
rect 1778 6158 1830 6164
rect 1780 5888 1828 6158
rect 1876 5888 1924 6446
rect 1972 5888 2020 6554
rect 2068 5897 2116 6554
rect 2164 5897 2212 6554
rect 2068 5888 2259 5897
rect 2083 5844 2259 5888
rect 2083 5835 2260 5844
rect 2083 5759 2126 5835
rect 2250 5759 2260 5835
rect 2083 5750 2260 5759
rect 2083 5697 2259 5750
rect 1588 5436 1636 5656
rect 1586 5430 1638 5436
rect 1586 5328 1638 5334
rect 1394 5286 1446 5292
rect 1394 5184 1446 5190
rect 1588 5184 1636 5328
rect 1780 5292 1828 5656
rect 1972 5436 2020 5656
rect 1970 5430 2022 5436
rect 1970 5328 2022 5334
rect 1778 5286 1830 5292
rect 1778 5184 1830 5190
rect 1972 5184 2020 5328
rect 2164 5184 2212 5697
rect 1396 4388 1444 5036
rect 1492 4388 1540 5036
rect 1588 4892 1636 5036
rect 1682 5030 1734 5036
rect 1682 4928 1734 4934
rect 1586 4886 1638 4892
rect 1586 4784 1638 4790
rect 1588 4388 1636 4784
rect 1684 4388 1732 4928
rect 1780 4748 1828 5036
rect 1874 5030 1926 5036
rect 1874 4928 1926 4934
rect 1778 4742 1830 4748
rect 1778 4640 1830 4646
rect 1780 4388 1828 4640
rect 1876 4388 1924 4928
rect 1972 4388 2020 5036
rect 2068 4388 2116 5036
rect 2164 4892 2212 5036
rect 2162 4886 2214 4892
rect 2162 4784 2214 4790
rect 1349 4374 1494 4388
rect 1349 4298 1359 4374
rect 1482 4298 1494 4374
rect 1349 4288 1494 4298
rect 1396 3784 1444 4288
rect 1588 4036 1636 4256
rect 1586 4030 1638 4036
rect 1586 3928 1638 3934
rect 1588 3784 1636 3928
rect 1780 3892 1828 4256
rect 1972 4036 2020 4256
rect 1970 4030 2022 4036
rect 1970 3928 2022 3934
rect 1778 3886 1830 3892
rect 1778 3784 1830 3790
rect 1972 3784 2020 3928
rect 2164 3892 2212 4784
rect 2162 3886 2214 3892
rect 2162 3784 2214 3790
rect 2365 3384 2845 4422
rect -175 3374 38 3384
rect -175 3298 -104 3374
rect 0 3298 38 3374
rect -175 3288 38 3298
rect 3543 3288 3825 3384
rect 578 3128 650 3134
rect 578 3072 586 3128
rect 642 3072 650 3128
rect 578 3066 650 3072
rect 962 3128 1034 3136
rect 962 3072 970 3128
rect 1026 3072 1034 3128
rect 962 3064 1034 3072
rect 1090 3128 1162 3136
rect 1090 3072 1098 3128
rect 1154 3072 1162 3128
rect 1090 3064 1162 3072
rect 1474 3128 1546 3136
rect 1474 3072 1482 3128
rect 1538 3072 1546 3128
rect 1474 3064 1546 3072
rect 1602 3128 1674 3136
rect 1602 3072 1610 3128
rect 1666 3072 1674 3128
rect 1602 3064 1674 3072
rect 1713 3128 1841 3136
rect 1713 3114 1777 3128
rect 1713 3080 1725 3114
rect 1759 3080 1777 3114
rect 1713 3072 1777 3080
rect 1833 3072 1841 3128
rect 1713 3064 1841 3072
rect 1936 3128 2008 3136
rect 1936 3072 1944 3128
rect 2000 3072 2008 3128
rect 1936 3064 2008 3072
rect 2064 3128 2136 3136
rect 2064 3072 2072 3128
rect 2128 3072 2136 3128
rect 2064 3064 2136 3072
rect 2448 3128 2520 3136
rect 2448 3072 2456 3128
rect 2512 3072 2520 3128
rect 2448 3064 2520 3072
rect 2576 3126 2648 3132
rect 2576 3070 2585 3126
rect 2641 3070 2648 3126
rect 2576 3064 2648 3070
rect 2960 3128 3032 3136
rect 2960 3072 2968 3128
rect 3024 3072 3032 3128
rect 2960 3064 3032 3072
rect 3571 2830 3825 2840
rect 3571 2754 3612 2830
rect 3716 2754 3825 2830
rect 3571 2744 3825 2754
rect -110 1640 36 1650
rect -110 1564 -102 1640
rect 2 1564 36 1640
rect -110 1554 36 1564
rect 322 1378 394 1384
rect 322 1322 330 1378
rect 386 1322 394 1378
rect 322 1316 394 1322
rect 706 1378 778 1384
rect 706 1322 714 1378
rect 770 1372 778 1378
rect 772 1336 778 1372
rect 770 1322 778 1336
rect 706 1316 778 1322
rect 834 1378 906 1384
rect 834 1322 842 1378
rect 898 1322 906 1378
rect 834 1316 906 1322
rect 962 1378 1034 1384
rect 962 1322 970 1378
rect 1026 1322 1034 1378
rect 962 1316 1034 1322
rect 1772 1378 1844 1384
rect 1772 1322 1780 1378
rect 1836 1322 1844 1378
rect 1474 1312 1546 1319
rect 1772 1316 1844 1322
rect 1938 1378 2010 1384
rect 1938 1322 1946 1378
rect 2002 1322 2010 1378
rect 1938 1316 2010 1322
rect 2056 1378 2124 1384
rect 2056 1322 2062 1378
rect 2118 1322 2124 1378
rect 2056 1316 2124 1322
rect 2830 1378 2906 1384
rect 2830 1372 2842 1378
rect 2830 1336 2836 1372
rect 2830 1322 2842 1336
rect 2898 1322 2906 1378
rect 2830 1316 2906 1322
rect 3218 1378 3290 1384
rect 3218 1322 3226 1378
rect 3282 1322 3290 1378
rect 3218 1316 3290 1322
rect 1474 1256 1482 1312
rect 1538 1256 1546 1312
rect 1474 1246 1546 1256
rect 1474 1210 1500 1246
rect 1534 1210 1546 1246
rect 1474 1199 1546 1210
rect -111 1010 36 1106
rect 3572 1096 3722 1106
rect 3572 1020 3610 1096
rect 3714 1020 3722 1096
rect 3572 1010 3722 1020
<< via1 >>
rect -8 22756 412 22996
rect 1574 22752 1630 22772
rect 1574 22718 1588 22752
rect 1588 22718 1622 22752
rect 1622 22718 1630 22752
rect 1574 22716 1630 22718
rect 1958 22760 2014 22772
rect 1958 22726 1992 22760
rect 1992 22726 2014 22760
rect 1958 22716 2014 22726
rect 3196 22212 3616 22452
rect 1720 21830 1888 21882
rect 3196 21512 3616 21752
rect 1778 21188 1830 21288
rect 1649 21044 1701 21144
rect 2207 21044 2259 21144
rect -8 20170 412 20410
rect 783 6974 1223 20420
rect 1819 20042 1885 20218
rect 1819 19020 1885 19196
rect 1819 17998 1885 18174
rect 1819 16846 1885 17022
rect 1819 15824 1885 16000
rect 1819 14672 1885 14848
rect 1819 12628 1885 12804
rect 1819 10454 1885 10630
rect 1819 8410 1885 8586
rect 1394 6308 1446 6404
rect 1682 6452 1734 6548
rect 1586 6308 1638 6404
rect 1874 6452 1926 6548
rect 1778 6164 1830 6260
rect 2126 5759 2250 5835
rect 1586 5334 1638 5430
rect 1394 5190 1446 5286
rect 1970 5334 2022 5430
rect 1778 5190 1830 5286
rect 1682 4934 1734 5030
rect 1586 4790 1638 4886
rect 1874 4934 1926 5030
rect 1778 4646 1830 4742
rect 2162 4790 2214 4886
rect 1359 4298 1364 4374
rect 1364 4298 1424 4374
rect 1424 4298 1482 4374
rect 1586 3934 1638 4030
rect 1970 3934 2022 4030
rect 1778 3790 1830 3886
rect 2162 3790 2214 3886
rect -104 3298 0 3374
rect 586 3123 642 3128
rect 586 3079 597 3123
rect 597 3079 631 3123
rect 631 3079 642 3123
rect 586 3072 642 3079
rect 970 3119 1026 3128
rect 970 3075 981 3119
rect 981 3075 1015 3119
rect 1015 3075 1026 3119
rect 970 3072 1026 3075
rect 1098 3122 1154 3128
rect 1098 3078 1102 3122
rect 1102 3078 1136 3122
rect 1136 3078 1154 3122
rect 1098 3072 1154 3078
rect 1482 3120 1538 3128
rect 1482 3080 1486 3120
rect 1486 3080 1520 3120
rect 1520 3080 1538 3120
rect 1482 3072 1538 3080
rect 1610 3116 1666 3128
rect 1610 3082 1612 3116
rect 1612 3082 1646 3116
rect 1646 3082 1666 3116
rect 1610 3072 1666 3082
rect 1777 3072 1833 3128
rect 1944 3122 2000 3128
rect 1944 3078 1948 3122
rect 1948 3078 1982 3122
rect 1982 3078 2000 3122
rect 1944 3072 2000 3078
rect 2072 3120 2128 3128
rect 2072 3080 2088 3120
rect 2088 3080 2122 3120
rect 2122 3080 2128 3120
rect 2072 3072 2128 3080
rect 2456 3122 2512 3128
rect 2456 3078 2460 3122
rect 2460 3078 2494 3122
rect 2494 3078 2512 3122
rect 2456 3072 2512 3078
rect 2585 3120 2641 3126
rect 2585 3076 2596 3120
rect 2596 3076 2630 3120
rect 2630 3076 2641 3120
rect 2585 3070 2641 3076
rect 2968 3122 3024 3128
rect 2968 3078 2972 3122
rect 2972 3078 3006 3122
rect 3006 3078 3024 3122
rect 2968 3072 3024 3078
rect 3612 2754 3716 2830
rect -102 1564 2 1640
rect 330 1374 386 1378
rect 330 1338 346 1374
rect 346 1338 380 1374
rect 380 1338 386 1374
rect 330 1322 386 1338
rect 714 1372 770 1378
rect 714 1336 738 1372
rect 738 1336 770 1372
rect 714 1322 770 1336
rect 842 1374 898 1378
rect 842 1338 860 1374
rect 860 1338 894 1374
rect 894 1338 898 1374
rect 842 1322 898 1338
rect 970 1374 1026 1378
rect 970 1338 988 1374
rect 988 1338 1022 1374
rect 1022 1338 1026 1374
rect 970 1322 1026 1338
rect 1780 1376 1836 1378
rect 1780 1340 1798 1376
rect 1798 1340 1832 1376
rect 1832 1340 1836 1376
rect 1780 1322 1836 1340
rect 1946 1376 2002 1378
rect 1946 1340 1950 1376
rect 1950 1340 1984 1376
rect 1984 1340 2002 1376
rect 1946 1322 2002 1340
rect 2062 1370 2118 1378
rect 2062 1334 2070 1370
rect 2070 1334 2104 1370
rect 2104 1334 2118 1370
rect 2062 1322 2118 1334
rect 2842 1372 2898 1378
rect 2842 1336 2870 1372
rect 2870 1336 2898 1372
rect 2842 1322 2898 1336
rect 3226 1372 3282 1378
rect 3226 1336 3228 1372
rect 3228 1336 3262 1372
rect 3262 1336 3282 1372
rect 3226 1322 3282 1336
rect 1482 1256 1538 1312
rect 3610 1020 3714 1096
<< metal2 >>
rect -38 22996 442 23026
rect -38 22756 -8 22996
rect 412 22756 442 22996
rect -38 22726 442 22756
rect 1566 22772 1638 22780
rect 1566 22716 1574 22772
rect 1630 22716 1638 22772
rect 1566 22140 1638 22716
rect 1950 22772 2022 22780
rect 1950 22716 1958 22772
rect 2014 22716 2022 22772
rect 1950 22332 2022 22716
rect 1950 22248 1954 22332
rect 2018 22248 2022 22332
rect 1566 22056 1570 22140
rect 1634 22056 1638 22140
rect 1566 22002 1638 22056
rect 1714 22136 1894 22146
rect 1714 22060 1724 22136
rect 1884 22060 1894 22136
rect 1714 21882 1894 22060
rect 1950 22002 2022 22248
rect 3166 22452 3646 22482
rect 3166 22212 3196 22452
rect 3616 22212 3646 22452
rect 3166 22182 3646 22212
rect 1714 21830 1720 21882
rect 1888 21830 1894 21882
rect 1714 21824 1894 21830
rect 3166 21752 3646 21782
rect 3166 21512 3196 21752
rect 3616 21512 3646 21752
rect 3166 21482 3646 21512
rect 1778 21288 1830 21294
rect 763 21190 793 21286
rect 1213 21190 1778 21286
rect 1830 21190 2716 21286
rect 1778 21182 1830 21188
rect 1649 21144 1701 21150
rect 892 21046 1649 21142
rect 2207 21144 2259 21150
rect 1701 21046 2207 21142
rect 1649 21038 1701 21044
rect 2259 21046 2395 21142
rect 2815 21046 2845 21142
rect 2207 21038 2259 21044
rect -38 20420 1243 20440
rect -38 20410 783 20420
rect -38 20170 -8 20410
rect 412 20170 783 20410
rect -38 20140 783 20170
rect 763 6974 783 20140
rect 1223 6974 1243 20420
rect 1493 20218 2115 20230
rect 1493 20210 1819 20218
rect 1885 20210 2115 20218
rect 1493 20050 1513 20210
rect 2095 20050 2115 20210
rect 1493 20042 1819 20050
rect 1885 20042 2115 20050
rect 1493 20030 2115 20042
rect 2365 20140 3646 20440
rect 1493 19196 2115 19208
rect 1493 19188 1819 19196
rect 1885 19188 2115 19196
rect 1493 19028 1513 19188
rect 2095 19028 2115 19188
rect 1493 19020 1819 19028
rect 1885 19020 2115 19028
rect 1493 19008 2115 19020
rect 1493 18174 2115 18186
rect 1493 18166 1819 18174
rect 1885 18166 2115 18174
rect 1493 18006 1513 18166
rect 2095 18006 2115 18166
rect 1493 17998 1819 18006
rect 1885 17998 2115 18006
rect 1493 17986 2115 17998
rect 1493 17022 2115 17034
rect 1493 17014 1819 17022
rect 1885 17014 2115 17022
rect 1493 16854 1513 17014
rect 2095 16854 2115 17014
rect 1493 16846 1819 16854
rect 1885 16846 2115 16854
rect 1493 16834 2115 16846
rect 1493 16000 2115 16012
rect 1493 15992 1819 16000
rect 1885 15992 2115 16000
rect 1493 15832 1513 15992
rect 2095 15832 2115 15992
rect 1493 15824 1819 15832
rect 1885 15824 2115 15832
rect 1493 15812 2115 15824
rect 1493 14848 2115 14860
rect 1493 14840 1819 14848
rect 1885 14840 2115 14848
rect 1493 14680 1513 14840
rect 2095 14680 2115 14840
rect 1493 14672 1819 14680
rect 1885 14672 2115 14680
rect 1493 14660 2115 14672
rect 1493 12804 2115 12816
rect 1493 12796 1819 12804
rect 1885 12796 2115 12804
rect 1493 12636 1513 12796
rect 2095 12636 2115 12796
rect 1493 12628 1819 12636
rect 1885 12628 2115 12636
rect 1493 12616 2115 12628
rect 1493 10630 2115 10642
rect 1493 10622 1819 10630
rect 1885 10622 2115 10630
rect 1493 10462 1513 10622
rect 2095 10462 2115 10622
rect 1493 10454 1819 10462
rect 1885 10454 2115 10462
rect 1493 10442 2115 10454
rect 1493 8586 2115 8598
rect 1493 8578 1819 8586
rect 1885 8578 2115 8586
rect 1493 8418 1513 8578
rect 2095 8418 2115 8578
rect 1493 8410 1819 8418
rect 1885 8410 2115 8418
rect 1493 8398 2115 8410
rect -110 3854 442 3884
rect -110 3514 -8 3854
rect 412 3514 442 3854
rect -110 3484 442 3514
rect -110 3374 10 3484
rect 763 3384 1243 6974
rect 1682 6548 1734 6554
rect 1874 6548 1926 6554
rect 1349 6452 1682 6548
rect 1734 6452 1874 6548
rect 1926 6452 2259 6548
rect 1682 6446 1734 6452
rect 1874 6446 1926 6452
rect 1394 6404 1446 6410
rect 1586 6404 1638 6410
rect 1349 6308 1394 6404
rect 1446 6308 1586 6404
rect 1638 6308 2259 6404
rect 1586 6302 1638 6308
rect 1778 6260 1830 6266
rect 1348 6250 1778 6260
rect 1348 6174 1358 6250
rect 1482 6174 1778 6250
rect 1348 6164 1778 6174
rect 1830 6164 2260 6260
rect 1778 6158 1830 6164
rect 2116 5835 2260 5844
rect 2116 5759 2126 5835
rect 2250 5759 2260 5835
rect 2116 5750 2260 5759
rect 1586 5430 1638 5436
rect 1970 5430 2022 5436
rect 1349 5334 1586 5430
rect 1638 5420 1970 5430
rect 1738 5344 1970 5420
rect 1638 5334 1970 5344
rect 2022 5334 2259 5430
rect 1586 5328 1638 5334
rect 1970 5328 2022 5334
rect 1394 5286 1446 5292
rect 1778 5286 1830 5292
rect 1349 5190 1394 5286
rect 1446 5190 1778 5286
rect 1830 5276 2259 5286
rect 1830 5200 1870 5276
rect 1994 5200 2259 5276
rect 1830 5190 2259 5200
rect 1394 5184 1446 5190
rect 1778 5184 1830 5190
rect 1682 5030 1734 5036
rect 1874 5030 1926 5036
rect 1349 4934 1682 5030
rect 1734 4934 1874 5030
rect 1926 4934 2259 5030
rect 2365 4950 2845 20140
rect 1682 4928 1734 4934
rect 1874 4928 1926 4934
rect 1586 4886 1638 4892
rect 2162 4886 2214 4892
rect 1349 4790 1586 4886
rect 1638 4790 2162 4886
rect 2214 4790 2259 4886
rect 1586 4784 1638 4790
rect 2162 4784 2214 4790
rect 1778 4742 1830 4748
rect 1349 4646 1778 4742
rect 1830 4732 2259 4742
rect 1830 4656 2126 4732
rect 2250 4656 2259 4732
rect 1830 4646 2259 4656
rect 1778 4640 1830 4646
rect 1349 4374 1492 4388
rect 1349 4298 1358 4374
rect 1482 4298 1492 4374
rect 1349 4288 1492 4298
rect 1586 4030 1638 4036
rect 1970 4030 2022 4036
rect 1349 3934 1586 4030
rect 1638 4020 1970 4030
rect 1738 3944 1970 4020
rect 1638 3934 1970 3944
rect 2022 3934 2259 4030
rect 1586 3928 1638 3934
rect 1970 3928 2022 3934
rect 1778 3886 1830 3892
rect 2162 3886 2214 3892
rect 1349 3790 1778 3886
rect 1830 3876 2162 3886
rect 1830 3800 1870 3876
rect 1994 3800 2162 3876
rect 1830 3790 2162 3800
rect 2214 3790 2259 3886
rect 1778 3784 1830 3790
rect 2162 3784 2214 3790
rect 2365 3384 2845 4422
rect 3166 3854 3722 3884
rect 3166 3514 3196 3854
rect 3616 3514 3722 3854
rect 3166 3484 3722 3514
rect -110 3298 -104 3374
rect 0 3298 10 3374
rect -110 1640 10 3298
rect 66 1744 138 3328
rect 194 1744 266 3328
rect 322 1744 394 3328
rect 450 1744 522 3328
rect 578 3128 650 3328
rect 578 3072 586 3128
rect 642 3072 650 3128
rect 578 1874 650 3072
rect 578 1790 582 1874
rect 646 1790 650 1874
rect 578 1744 650 1790
rect 706 1744 778 3328
rect 834 1744 906 3328
rect 962 3128 1034 3328
rect 962 3072 970 3128
rect 1026 3072 1034 3128
rect 962 2066 1034 3072
rect 962 1982 966 2066
rect 1030 1982 1034 2066
rect 962 1744 1034 1982
rect 1090 3128 1162 3328
rect 1090 3072 1098 3128
rect 1154 3072 1162 3128
rect 1090 2258 1162 3072
rect 1090 2174 1094 2258
rect 1158 2174 1162 2258
rect 1090 1744 1162 2174
rect 1218 1744 1290 3328
rect 1346 1744 1418 3328
rect 1474 3128 1546 3328
rect 1474 3072 1482 3128
rect 1538 3072 1546 3128
rect 1474 2450 1546 3072
rect 1474 2366 1478 2450
rect 1542 2366 1546 2450
rect 1474 1744 1546 2366
rect 1602 3308 1674 3328
rect 1602 3146 1609 3308
rect 1665 3146 1674 3308
rect 1602 3128 1674 3146
rect 1602 3072 1610 3128
rect 1666 3072 1674 3128
rect 1602 1744 1674 3072
rect 1769 3128 1841 3328
rect 1769 3072 1777 3128
rect 1833 3072 1841 3128
rect 1769 3020 1841 3072
rect 1769 2858 1778 3020
rect 1834 2858 1841 3020
rect 1769 1744 1841 2858
rect 1936 3128 2008 3328
rect 1936 3072 1944 3128
rect 2000 3072 2008 3128
rect 1936 2642 2008 3072
rect 1936 2558 1940 2642
rect 2004 2558 2008 2642
rect 1936 1744 2008 2558
rect 2064 3128 2136 3328
rect 2064 3072 2072 3128
rect 2128 3072 2136 3128
rect 2064 2642 2136 3072
rect 2064 2558 2068 2642
rect 2132 2558 2136 2642
rect 2064 1744 2136 2558
rect 2192 1744 2264 3328
rect 2320 1744 2392 3328
rect 2448 3128 2520 3328
rect 2448 3072 2456 3128
rect 2512 3072 2520 3128
rect 2448 2450 2520 3072
rect 2448 2366 2452 2450
rect 2516 2366 2520 2450
rect 2448 1744 2520 2366
rect 2576 3126 2648 3328
rect 2576 3070 2585 3126
rect 2641 3070 2648 3126
rect 2576 2258 2648 3070
rect 2576 2174 2580 2258
rect 2644 2174 2648 2258
rect 2576 1744 2648 2174
rect 2704 1744 2776 3328
rect 2832 1744 2904 3328
rect 2960 3128 3032 3328
rect 2960 3072 2968 3128
rect 3024 3072 3032 3128
rect 2960 2066 3032 3072
rect 2960 1982 2964 2066
rect 3028 1982 3032 2066
rect 2960 1744 3032 1982
rect 3088 1744 3160 3328
rect 3216 1744 3288 3328
rect 3344 1744 3416 3328
rect 3472 1744 3544 3328
rect 3602 2830 3722 3484
rect 3602 2754 3612 2830
rect 3716 2754 3722 2830
rect -110 1564 -102 1640
rect 2 1564 10 1640
rect -110 1010 10 1564
rect 66 2 138 1402
rect 194 2 266 1402
rect 322 1378 394 1402
rect 322 1322 330 1378
rect 386 1322 394 1378
rect 322 2 394 1322
rect 450 2 522 1402
rect 578 2 650 1402
rect 706 1378 778 1402
rect 706 1322 714 1378
rect 770 1322 778 1378
rect 706 140 778 1322
rect 706 56 710 140
rect 774 56 778 140
rect 706 2 778 56
rect 834 1378 906 1402
rect 834 1322 842 1378
rect 898 1322 906 1378
rect 834 716 906 1322
rect 834 632 838 716
rect 902 632 906 716
rect 834 2 906 632
rect 962 1378 1034 1402
rect 962 1322 970 1378
rect 1026 1322 1034 1378
rect 962 908 1034 1322
rect 962 824 966 908
rect 1030 824 1034 908
rect 962 2 1034 824
rect 1090 2 1162 1402
rect 1218 2 1290 1402
rect 1346 2 1418 1402
rect 1474 1312 1546 1402
rect 1474 1256 1482 1312
rect 1538 1256 1546 1312
rect 1474 2 1546 1256
rect 1602 2 1674 1402
rect 1772 1378 1844 1402
rect 1772 1322 1780 1378
rect 1836 1322 1844 1378
rect 1772 332 1844 1322
rect 1772 248 1776 332
rect 1840 248 1844 332
rect 1772 2 1844 248
rect 1938 1378 2010 1402
rect 1938 1322 1946 1378
rect 2002 1322 2010 1378
rect 1938 524 2010 1322
rect 2056 1378 2138 1402
rect 2056 1322 2062 1378
rect 2118 1322 2138 1378
rect 2056 1316 2138 1322
rect 1938 440 1942 524
rect 2006 440 2010 524
rect 1938 2 2010 440
rect 2066 2 2138 1316
rect 2194 2 2266 1402
rect 2322 2 2394 1402
rect 2450 2 2522 1402
rect 2578 2 2650 1402
rect 2706 2 2778 1402
rect 2834 1378 2906 1402
rect 2834 1322 2842 1378
rect 2898 1322 2906 1378
rect 2834 2 2906 1322
rect 2962 2 3034 1402
rect 3090 2 3162 1402
rect 3218 1378 3290 1402
rect 3218 1322 3226 1378
rect 3282 1322 3290 1378
rect 3218 2 3290 1322
rect 3346 2 3418 1402
rect 3474 2 3546 1402
rect 3602 1096 3722 2754
rect 3602 1020 3610 1096
rect 3714 1020 3722 1096
rect 3602 1010 3722 1020
<< via2 >>
rect -8 22756 412 22996
rect 1954 22248 2018 22332
rect 1570 22056 1634 22140
rect 1724 22060 1884 22136
rect 3196 22212 3616 22452
rect 3196 21512 3616 21752
rect 793 21190 1213 21286
rect 2395 21046 2815 21142
rect -8 20170 412 20410
rect 1513 20050 1819 20210
rect 1819 20050 1885 20210
rect 1885 20050 2095 20210
rect 1513 19028 1819 19188
rect 1819 19028 1885 19188
rect 1885 19028 2095 19188
rect 1513 18006 1819 18166
rect 1819 18006 1885 18166
rect 1885 18006 2095 18166
rect 1513 16854 1819 17014
rect 1819 16854 1885 17014
rect 1885 16854 2095 17014
rect 1513 15832 1819 15992
rect 1819 15832 1885 15992
rect 1885 15832 2095 15992
rect 1513 14680 1819 14840
rect 1819 14680 1885 14840
rect 1885 14680 2095 14840
rect 1513 12636 1819 12796
rect 1819 12636 1885 12796
rect 1885 12636 2095 12796
rect 1513 10462 1819 10622
rect 1819 10462 1885 10622
rect 1885 10462 2095 10622
rect 1513 8418 1819 8578
rect 1819 8418 1885 8578
rect 1885 8418 2095 8578
rect -8 3514 412 3854
rect 1358 6174 1482 6250
rect 2126 5759 2250 5835
rect 1614 5344 1638 5420
rect 1638 5344 1738 5420
rect 1870 5200 1994 5276
rect 2126 4656 2250 4732
rect 1358 4298 1359 4374
rect 1359 4298 1482 4374
rect 1614 3944 1638 4020
rect 1638 3944 1738 4020
rect 1870 3800 1994 3876
rect 3196 3514 3616 3854
rect 582 1790 646 1874
rect 966 1982 1030 2066
rect 1094 2174 1158 2258
rect 1478 2366 1542 2450
rect 1609 3146 1665 3308
rect 1778 2858 1834 3020
rect 1940 2558 2004 2642
rect 2068 2558 2132 2642
rect 2452 2366 2516 2450
rect 2580 2174 2644 2258
rect 2964 1982 3028 2066
rect 330 1322 386 1378
rect 710 56 774 140
rect 838 632 902 716
rect 966 824 1030 908
rect 1776 248 1840 332
rect 1942 440 2006 524
rect 3226 1322 3282 1378
<< metal3 >>
rect -38 22996 442 23026
rect -38 22756 -8 22996
rect 412 22756 442 22996
rect -38 22726 442 22756
rect 3166 22452 3646 22482
rect 892 22332 2716 22338
rect 892 22248 1954 22332
rect 2018 22248 2716 22332
rect 892 22242 2716 22248
rect 3166 22212 3196 22452
rect 3616 22212 3646 22452
rect 3166 22182 3646 22212
rect 892 22140 2716 22146
rect 892 22056 1570 22140
rect 1634 22136 2716 22140
rect 1634 22060 1724 22136
rect 1884 22060 2716 22136
rect 1634 22056 2716 22060
rect 892 22050 2716 22056
rect 3166 21752 3646 21782
rect 3166 21512 3196 21752
rect 3616 21512 3646 21752
rect 3166 21482 3646 21512
rect 763 21286 1243 21334
rect 763 21046 793 21286
rect 1213 21046 1243 21286
rect 763 20998 1243 21046
rect 2365 21286 2845 21334
rect 2365 21046 2395 21286
rect 2815 21046 2845 21286
rect 2365 20998 2845 21046
rect -38 20410 442 20440
rect -38 20170 -8 20410
rect 412 20170 442 20410
rect -38 20140 442 20170
rect 1493 20210 2115 20230
rect 1493 20050 1513 20210
rect 2095 20050 2115 20210
rect 1493 20030 2115 20050
rect 1493 19188 2115 19208
rect 1493 19028 1513 19188
rect 2095 19028 2115 19188
rect 1493 19008 2115 19028
rect 1493 18166 2115 18186
rect 1493 18006 1513 18166
rect 2095 18006 2115 18166
rect 1493 17986 2115 18006
rect 1493 17014 2115 17034
rect 1493 16854 1513 17014
rect 2095 16854 2115 17014
rect 1493 16834 2115 16854
rect 1493 15992 2115 16012
rect 1493 15832 1513 15992
rect 2095 15832 2115 15992
rect 1493 15812 2115 15832
rect 1493 14840 2115 14860
rect 1493 14680 1513 14840
rect 2095 14680 2115 14840
rect 1493 14660 2115 14680
rect 1493 12796 2115 12816
rect 1493 12636 1513 12796
rect 2095 12636 2115 12796
rect 1493 12616 2115 12636
rect 1493 10622 2115 10642
rect 1493 10462 1513 10622
rect 2095 10462 2115 10622
rect 1493 10442 2115 10462
rect 1493 8578 2115 8598
rect 1493 8418 1513 8578
rect 2095 8418 2115 8578
rect 1493 8398 2115 8418
rect 1348 6250 1492 6548
rect 1348 6174 1358 6250
rect 1482 6174 1492 6250
rect 1348 4412 1492 6174
rect 1348 4080 1358 4412
rect 1482 4080 1492 4412
rect -38 3854 442 3884
rect -38 3514 -8 3854
rect 412 3514 442 3854
rect 1348 3790 1492 4080
rect 1604 5468 1748 6548
rect 1604 5136 1614 5468
rect 1738 5136 1748 5468
rect 1604 4020 1748 5136
rect 1604 3944 1614 4020
rect 1738 3944 1748 4020
rect 1604 3790 1748 3944
rect 1860 5276 2004 6548
rect 1860 5200 1870 5276
rect 1994 5200 2004 5276
rect 1860 4940 2004 5200
rect 1860 4608 1870 4940
rect 1994 4608 2004 4940
rect 1860 3876 2004 4608
rect 1860 3800 1870 3876
rect 1994 3800 2004 3876
rect 1860 3790 2004 3800
rect 2116 5996 2260 6548
rect 2116 5664 2126 5996
rect 2250 5664 2260 5996
rect 2116 4732 2260 5664
rect 2116 4656 2126 4732
rect 2250 4656 2260 4732
rect 2116 3790 2260 4656
rect 3166 3854 3646 3884
rect -38 3484 442 3514
rect 3166 3514 3196 3854
rect 3616 3514 3646 3854
rect 3166 3484 3646 3514
rect -176 3318 3825 3328
rect -176 3166 1594 3318
rect 2014 3166 3825 3318
rect -176 3146 1609 3166
rect 1665 3146 3825 3166
rect -176 3136 3825 3146
rect -176 2888 793 3040
rect 1213 3020 3825 3040
rect 1213 2888 1778 3020
rect -176 2858 1778 2888
rect 1834 2858 3825 3020
rect -176 2848 3825 2858
rect -175 2642 3825 2648
rect -175 2638 1940 2642
rect -175 2562 1716 2638
rect 1894 2562 1940 2638
rect -175 2558 1940 2562
rect 2004 2558 2068 2642
rect 2132 2558 3825 2642
rect -175 2552 3825 2558
rect -175 2450 3825 2456
rect -175 2366 1478 2450
rect 1542 2446 2452 2450
rect 1542 2370 2330 2446
rect 1542 2366 2452 2370
rect 2516 2366 3825 2450
rect -175 2360 3825 2366
rect -175 2258 3825 2264
rect -175 2174 1094 2258
rect 1158 2254 2580 2258
rect 1278 2178 2580 2254
rect 1158 2174 2580 2178
rect 2644 2174 3825 2258
rect -175 2168 3825 2174
rect -175 2066 3825 2072
rect -175 1982 966 2066
rect 1030 2062 2964 2066
rect 1030 1986 2842 2062
rect 1030 1982 2964 1986
rect 3028 1982 3825 2066
rect -175 1976 3825 1982
rect -175 1874 3825 1880
rect -175 1790 582 1874
rect 646 1870 3825 1874
rect 766 1794 3825 1870
rect 646 1790 3825 1794
rect -175 1784 3825 1790
rect 266 1392 394 1402
rect 266 1284 276 1392
rect 384 1378 394 1392
rect 386 1322 394 1378
rect 384 1284 394 1322
rect 266 1274 394 1284
rect 3218 1392 3346 1402
rect 3218 1378 3228 1392
rect 3218 1322 3226 1378
rect 3218 1284 3228 1322
rect 3336 1284 3346 1392
rect 3218 1274 3346 1284
rect -143 1152 55 1239
rect 3578 1152 3776 1239
rect -175 908 3825 914
rect -175 824 966 908
rect 1030 904 3825 908
rect 1030 828 2330 904
rect 2508 828 3825 904
rect 1030 824 3825 828
rect -175 818 3825 824
rect -175 716 3825 722
rect -175 632 838 716
rect 902 712 3825 716
rect 902 636 1100 712
rect 1278 636 3825 712
rect 902 632 3825 636
rect -175 626 3825 632
rect -175 524 3825 530
rect -175 440 1942 524
rect 2006 520 3825 524
rect 2006 444 2842 520
rect 3020 444 3825 520
rect 2006 440 3825 444
rect -175 434 3825 440
rect -175 332 3825 338
rect -175 328 1776 332
rect -175 252 588 328
rect 766 252 1776 328
rect -175 248 1776 252
rect 1840 248 3825 332
rect -175 242 3825 248
rect -175 140 3825 146
rect -175 56 710 140
rect 774 136 3825 140
rect 774 60 1716 136
rect 1894 60 3825 136
rect 774 56 3825 60
rect -175 50 3825 56
<< via3 >>
rect -8 22756 412 22996
rect 3196 22212 3616 22452
rect 3196 21512 3616 21752
rect 793 21190 1213 21286
rect 793 21046 1213 21190
rect 2395 21142 2815 21286
rect 2395 21046 2815 21142
rect -8 20170 412 20410
rect 1513 20050 2095 20190
rect 1513 19028 2095 19168
rect 1513 18006 2095 18166
rect 1513 16854 2095 17014
rect 1513 15832 2095 15992
rect 1513 14680 2095 14840
rect 1513 12636 2095 12796
rect 1513 10462 2095 10622
rect 1513 8418 2095 8578
rect 1358 4374 1482 4412
rect 1358 4298 1482 4374
rect 1358 4080 1482 4298
rect -8 3514 412 3854
rect 1614 5420 1738 5468
rect 1614 5344 1738 5420
rect 1614 5136 1738 5344
rect 1870 4608 1994 4940
rect 2126 5835 2250 5996
rect 2126 5759 2250 5835
rect 2126 5664 2250 5759
rect 3196 3514 3616 3854
rect 1594 3308 2014 3318
rect 1594 3166 1609 3308
rect 1609 3166 1665 3308
rect 1665 3166 2014 3308
rect 793 2888 1213 3040
rect 1716 2562 1894 2638
rect 2330 2370 2452 2446
rect 2452 2370 2508 2446
rect 1100 2178 1158 2254
rect 1158 2178 1278 2254
rect 2842 1986 2964 2062
rect 2964 1986 3020 2062
rect 588 1794 646 1870
rect 646 1794 766 1870
rect 276 1378 384 1392
rect 276 1322 330 1378
rect 330 1322 384 1378
rect 276 1284 384 1322
rect 3228 1378 3336 1392
rect 3228 1322 3282 1378
rect 3282 1322 3336 1378
rect 3228 1284 3336 1322
rect 2330 828 2508 904
rect 1100 636 1278 712
rect 2842 444 3020 520
rect 588 252 766 328
rect 1716 60 1894 136
<< metal4 >>
rect -38 22996 442 23026
rect -38 22756 -8 22996
rect 412 22756 442 22996
rect -38 22726 442 22756
rect 3166 22452 3646 22482
rect 3166 22212 3196 22452
rect 3616 22212 3646 22452
rect 3166 22182 3646 22212
rect 3166 21752 3646 21782
rect 3166 21512 3196 21752
rect 3616 21512 3646 21752
rect 3166 21482 3646 21512
rect 763 21286 1243 21334
rect 763 21046 793 21286
rect 1213 21046 1243 21286
rect 763 20998 1243 21046
rect 2365 21286 2845 21334
rect 2365 21046 2395 21286
rect 2815 21046 2845 21286
rect 2365 20998 2845 21046
rect -38 20410 442 20440
rect -38 20170 -8 20410
rect 412 20170 442 20410
rect -38 20140 442 20170
rect 763 20190 2845 20440
rect 763 20140 1513 20190
rect 1493 20050 1513 20140
rect 2095 20140 2845 20190
rect 2095 20050 2115 20140
rect 1493 20030 2115 20050
rect 763 19878 2845 19908
rect 763 19638 2395 19878
rect 2815 19638 2845 19878
rect 763 19608 2845 19638
rect 763 19241 2845 19418
rect 763 19168 2842 19241
rect 763 19118 1513 19168
rect 1493 19028 1513 19118
rect 2095 19118 2842 19168
rect 2095 19028 2115 19118
rect 1493 19008 2115 19028
rect 763 18856 2845 18886
rect 763 18616 2395 18856
rect 2815 18616 2845 18856
rect 763 18586 2845 18616
rect 33 18166 3575 18396
rect 33 18096 1513 18166
rect 1493 18006 1513 18096
rect 2095 18096 3575 18166
rect 2095 18006 2115 18096
rect 1493 17986 2115 18006
rect 33 17834 3575 17864
rect 33 17594 2395 17834
rect 2815 17594 3575 17834
rect 33 17564 3575 17594
rect 33 17214 3575 17244
rect 33 17014 1594 17214
rect 2014 17014 3575 17214
rect 33 16944 1513 17014
rect 1493 16854 1513 16944
rect 2095 16944 3575 17014
rect 2095 16854 2115 16944
rect 1493 16834 2115 16854
rect 33 16442 2395 16662
rect 2815 16442 3575 16662
rect 33 16412 3575 16442
rect 33 16192 3575 16222
rect 33 15992 1594 16192
rect 2014 15992 3575 16192
rect 33 15922 1513 15992
rect 1493 15832 1513 15922
rect 2095 15922 3575 15992
rect 2095 15832 2115 15922
rect 1493 15812 2115 15832
rect 33 15660 3575 15690
rect 33 15420 2395 15660
rect 2815 15420 3575 15660
rect 33 15390 3575 15420
rect 33 15040 3575 15070
rect 33 14840 1594 15040
rect 2014 14840 3575 15040
rect 33 14770 1513 14840
rect 1493 14680 1513 14770
rect 2095 14770 3575 14840
rect 2095 14680 2115 14770
rect 1493 14660 2115 14680
rect 33 14508 3575 14538
rect 33 14268 2395 14508
rect 2815 14268 3575 14508
rect 33 14238 3575 14268
rect 33 14018 3575 14048
rect 33 13778 1594 14018
rect 2014 13778 3575 14018
rect 33 13748 3575 13778
rect 33 13486 3575 13516
rect 33 13246 2395 13486
rect 2815 13246 3575 13486
rect 33 13216 3575 13246
rect 33 12996 3575 13026
rect 33 12796 1594 12996
rect 2014 12796 3575 12996
rect 33 12726 1513 12796
rect 1493 12636 1513 12726
rect 2095 12726 3575 12796
rect 2095 12636 2115 12726
rect 1493 12616 2115 12636
rect 33 12464 3575 12494
rect 33 12224 2395 12464
rect 2815 12224 3575 12464
rect 33 12194 3575 12224
rect 33 11974 3575 12004
rect 33 11734 1594 11974
rect 2014 11734 3575 11974
rect 33 11704 3575 11734
rect 33 11442 3575 11472
rect 33 11202 2395 11442
rect 2815 11202 3575 11442
rect 33 11172 3575 11202
rect 33 10822 3575 10852
rect 33 10622 1594 10822
rect 2014 10622 3575 10822
rect 33 10552 1513 10622
rect 1493 10462 1513 10552
rect 2095 10552 3575 10622
rect 2095 10462 2115 10552
rect 1493 10442 2115 10462
rect 33 10290 3575 10320
rect 33 10050 2395 10290
rect 2815 10050 3575 10290
rect 33 10020 3575 10050
rect 33 9800 3575 9830
rect 33 9560 1594 9800
rect 2014 9560 3575 9800
rect 33 9530 3575 9560
rect 33 9268 3575 9298
rect 33 9028 2395 9268
rect 2815 9028 3575 9268
rect 33 8998 3575 9028
rect 33 8778 3575 8808
rect 33 8578 1594 8778
rect 2014 8578 3575 8778
rect 33 8508 1513 8578
rect 1493 8418 1513 8508
rect 2095 8508 3575 8578
rect 2095 8418 2115 8508
rect 1493 8398 2115 8418
rect 33 8246 3575 8276
rect 33 8006 2395 8246
rect 2815 8006 3575 8246
rect 33 7976 3575 8006
rect 33 7756 3575 7786
rect 33 7516 1594 7756
rect 2014 7516 3575 7756
rect 33 7486 3575 7516
rect 33 7224 3575 7254
rect 33 6984 2395 7224
rect 2815 6984 3575 7224
rect 33 6954 3575 6984
rect -38 5996 3646 6006
rect -38 5664 2126 5996
rect 2250 5976 3646 5996
rect 2250 5684 3196 5976
rect 3616 5684 3646 5976
rect 2250 5664 3646 5684
rect -38 5654 3646 5664
rect -38 5468 3646 5478
rect -38 5136 1614 5468
rect 1738 5448 3646 5468
rect 1738 5156 2395 5448
rect 2815 5156 3646 5448
rect 1738 5136 3646 5156
rect -38 5126 3646 5136
rect -38 4940 3646 4950
rect -38 4920 1870 4940
rect 1994 4920 3646 4940
rect -38 4628 1594 4920
rect 2014 4628 3646 4920
rect -38 4608 1870 4628
rect 1994 4608 3646 4628
rect -38 4598 3646 4608
rect -38 4412 3646 4422
rect -38 4392 1358 4412
rect -38 4100 -8 4392
rect 412 4100 1358 4392
rect -38 4080 1358 4100
rect 1482 4080 3646 4412
rect -38 4070 3646 4080
rect -38 3854 442 3884
rect -38 3514 -8 3854
rect 412 3514 442 3854
rect -38 3484 442 3514
rect 2366 3854 3646 3884
rect 2366 3514 2396 3854
rect 2816 3514 3196 3854
rect 3616 3514 3646 3854
rect 2366 3484 3646 3514
rect 763 3354 1243 3384
rect 763 2878 793 3354
rect 1213 2878 1243 3354
rect 763 2848 1243 2878
rect 1564 3354 2044 3384
rect 1564 2878 1594 3354
rect 2014 2878 2044 3354
rect 1564 2848 2044 2878
rect 66 1402 266 2648
rect 578 1870 778 2648
rect 578 1794 588 1870
rect 766 1794 778 1870
rect 66 1392 394 1402
rect 66 1284 276 1392
rect 384 1284 394 1392
rect 66 1274 394 1284
rect 66 2 266 1274
rect 578 328 778 1794
rect 578 252 588 328
rect 766 252 778 328
rect 578 2 778 252
rect 1090 2254 1290 2648
rect 1090 2178 1100 2254
rect 1278 2178 1290 2254
rect 1090 712 1290 2178
rect 1090 636 1100 712
rect 1278 636 1290 712
rect 1090 2 1290 636
rect 1705 2638 1905 2648
rect 1705 2562 1716 2638
rect 1894 2562 1905 2638
rect 1705 136 1905 2562
rect 1705 60 1716 136
rect 1894 60 1905 136
rect 1705 2 1905 60
rect 2320 2446 2520 2648
rect 2320 2370 2330 2446
rect 2508 2370 2520 2446
rect 2320 904 2520 2370
rect 2320 828 2330 904
rect 2508 828 2520 904
rect 2320 2 2520 828
rect 2832 2062 3032 2648
rect 2832 1986 2842 2062
rect 3020 1986 3032 2062
rect 2832 520 3032 1986
rect 3344 1402 3544 2648
rect 3218 1392 3544 1402
rect 3218 1284 3228 1392
rect 3336 1284 3544 1392
rect 3218 1274 3544 1284
rect 2832 444 2842 520
rect 3020 444 3032 520
rect 2832 2 3032 444
rect 3344 2 3544 1274
<< via4 >>
rect -8 22756 412 22996
rect 3196 22212 3616 22452
rect 3196 21512 3616 21752
rect 793 21046 1213 21286
rect 2395 21046 2815 21286
rect -8 20170 412 20410
rect 2395 19638 2815 19878
rect 2395 18616 2815 18856
rect 2395 17594 2815 17834
rect 1594 17014 2014 17214
rect 1594 16974 2014 17014
rect 2395 16442 2815 16682
rect 1594 15992 2014 16192
rect 1594 15952 2014 15992
rect 2395 15420 2815 15660
rect 1594 14840 2014 15040
rect 1594 14800 2014 14840
rect 2395 14268 2815 14508
rect 1594 13778 2014 14018
rect 2395 13246 2815 13486
rect 1594 12796 2014 12996
rect 1594 12756 2014 12796
rect 2395 12224 2815 12464
rect 1594 11734 2014 11974
rect 2395 11202 2815 11442
rect 1594 10622 2014 10822
rect 1594 10582 2014 10622
rect 2395 10050 2815 10290
rect 1594 9560 2014 9800
rect 2395 9028 2815 9268
rect 1594 8578 2014 8778
rect 1594 8538 2014 8578
rect 2395 8006 2815 8246
rect 1594 7516 2014 7756
rect 2395 6984 2815 7224
rect 3196 5684 3616 5976
rect 2395 5156 2815 5448
rect 1594 4628 1870 4920
rect 1870 4628 1994 4920
rect 1994 4628 2014 4920
rect -8 4100 412 4392
rect -8 3514 412 3854
rect 2396 3514 2816 3854
rect 3196 3514 3616 3854
rect 793 3040 1213 3354
rect 793 2888 1213 3040
rect 793 2878 1213 2888
rect 1594 3318 2014 3354
rect 1594 3166 2014 3318
rect 1594 2878 2014 3166
<< metal5 >>
rect -38 22996 442 23026
rect -38 22756 -8 22996
rect 412 22756 442 22996
rect -38 20410 442 22756
rect 3166 22452 3646 23026
rect 3166 22212 3196 22452
rect 3616 22212 3646 22452
rect 3166 21752 3646 22212
rect 3166 21512 3196 21752
rect 3616 21512 3646 21752
rect -38 20170 -8 20410
rect 412 20170 442 20410
rect -38 4392 442 20170
rect -38 4100 -8 4392
rect 412 4100 442 4392
rect -38 3854 442 4100
rect -38 3514 -8 3854
rect 412 3514 442 3854
rect -38 2848 442 3514
rect 763 21286 1243 21334
rect 763 21046 793 21286
rect 1213 21046 1243 21286
rect 763 3354 1243 21046
rect 2365 21286 2845 21334
rect 2365 21046 2395 21286
rect 2815 21046 2845 21286
rect 1564 17564 2044 20440
rect 2365 19878 2845 21046
rect 2365 19638 2395 19878
rect 2815 19638 2845 19878
rect 2365 18856 2845 19638
rect 2365 18616 2395 18856
rect 2815 18616 2845 18856
rect 2365 17834 2845 18616
rect 2365 17594 2395 17834
rect 2815 17594 2845 17834
rect 1564 17214 2044 17244
rect 1564 16974 1594 17214
rect 2014 16974 2044 17214
rect 1564 16192 2044 16974
rect 1564 15952 1594 16192
rect 2014 15952 2044 16192
rect 1564 15390 2044 15952
rect 2365 16682 2845 17594
rect 2365 16442 2395 16682
rect 2815 16442 2845 16682
rect 2365 15660 2845 16442
rect 2365 15420 2395 15660
rect 2815 15420 2845 15660
rect 1564 15040 2044 15070
rect 1564 14800 1594 15040
rect 2014 14800 2044 15040
rect 1564 14018 2044 14800
rect 1564 13778 1594 14018
rect 2014 13778 2044 14018
rect 1564 12996 2044 13778
rect 1564 12756 1594 12996
rect 2014 12756 2044 12996
rect 1564 11974 2044 12756
rect 1564 11734 1594 11974
rect 2014 11734 2044 11974
rect 1564 11172 2044 11734
rect 2365 14508 2845 15420
rect 2365 14268 2395 14508
rect 2815 14268 2845 14508
rect 2365 13486 2845 14268
rect 2365 13246 2395 13486
rect 2815 13246 2845 13486
rect 2365 12464 2845 13246
rect 2365 12224 2395 12464
rect 2815 12224 2845 12464
rect 2365 11442 2845 12224
rect 2365 11202 2395 11442
rect 2815 11202 2845 11442
rect 1564 10822 2044 10852
rect 1564 10582 1594 10822
rect 2014 10582 2044 10822
rect 1564 9800 2044 10582
rect 1564 9560 1594 9800
rect 2014 9560 2044 9800
rect 1564 8778 2044 9560
rect 1564 8538 1594 8778
rect 2014 8538 2044 8778
rect 1564 7756 2044 8538
rect 1564 7516 1594 7756
rect 2014 7516 2044 7756
rect 1564 6954 2044 7516
rect 2365 10290 2845 11202
rect 2365 10050 2395 10290
rect 2815 10050 2845 10290
rect 2365 9268 2845 10050
rect 2365 9028 2395 9268
rect 2815 9028 2845 9268
rect 2365 8246 2845 9028
rect 2365 8006 2395 8246
rect 2815 8006 2845 8246
rect 2365 7224 2845 8006
rect 2365 6984 2395 7224
rect 2815 6984 2845 7224
rect 2365 5448 2845 6984
rect 2365 5156 2395 5448
rect 2815 5156 2845 5448
rect 2365 4950 2845 5156
rect 3166 5976 3646 21512
rect 3166 5684 3196 5976
rect 3616 5684 3646 5976
rect 763 2878 793 3354
rect 1213 2878 1243 3354
rect 763 2848 1243 2878
rect 1564 4920 2044 4950
rect 1564 4628 1594 4920
rect 2014 4628 2044 4920
rect 1564 3354 2044 4628
rect 1564 2878 1594 3354
rect 2014 2878 2044 3354
rect 1564 2848 2044 2878
rect 2365 3854 2845 4422
rect 2365 3514 2396 3854
rect 2816 3514 2845 3854
rect 2365 -352 2845 3514
rect 3166 3854 3646 5684
rect 3166 3514 3196 3854
rect 3616 3514 3646 3854
rect 3166 2848 3646 3514
use sky130_fd_pr__cap_mim_m3_1_FJFAMD  sky130_fd_pr__cap_mim_m3_1_FJFAMD_0
timestamp 1696948209
transform 0 -1 2605 -1 0 11618
box -386 -240 386 240
use sky130_fd_pr__cap_mim_m3_1_FJFAMD  sky130_fd_pr__cap_mim_m3_1_FJFAMD_1
timestamp 1696948209
transform 0 1 1003 -1 0 19032
box -386 -240 386 240
use sky130_fd_pr__cap_mim_m3_1_FJFAMD  sky130_fd_pr__cap_mim_m3_1_FJFAMD_2
timestamp 1696948209
transform 0 -1 3335 1 0 15836
box -386 -240 386 240
use sky130_fd_pr__cap_mim_m3_1_FJFAMD  sky130_fd_pr__cap_mim_m3_1_FJFAMD_3
timestamp 1696948209
transform 0 1 1003 -1 0 20054
box -386 -240 386 240
use sky130_fd_pr__cap_mim_m3_1_FJFAMD  sky130_fd_pr__cap_mim_m3_1_FJFAMD_4
timestamp 1696948209
transform 0 -1 2605 -1 0 20054
box -386 -240 386 240
use sky130_fd_pr__cap_mim_m3_1_FJFAMD  sky130_fd_pr__cap_mim_m3_1_FJFAMD_5
timestamp 1696948209
transform 0 -1 2605 -1 0 15836
box -386 -240 386 240
use sky130_fd_pr__cap_mim_m3_1_FJFAMD  sky130_fd_pr__cap_mim_m3_1_FJFAMD_6
timestamp 1696948209
transform 0 1 1003 -1 0 15836
box -386 -240 386 240
use sky130_fd_pr__cap_mim_m3_1_FJFAMD  sky130_fd_pr__cap_mim_m3_1_FJFAMD_7
timestamp 1696948209
transform 0 -1 2605 -1 0 19032
box -386 -240 386 240
use sky130_fd_pr__cap_mim_m3_1_FJFAMD  sky130_fd_pr__cap_mim_m3_1_FJFAMD_8
timestamp 1696948209
transform 0 1 273 1 0 18010
box -386 -240 386 240
use sky130_fd_pr__cap_mim_m3_1_FJFAMD  sky130_fd_pr__cap_mim_m3_1_FJFAMD_9
timestamp 1696948209
transform 0 1 1003 -1 0 18010
box -386 -240 386 240
use sky130_fd_pr__cap_mim_m3_1_FJFAMD  sky130_fd_pr__cap_mim_m3_1_FJFAMD_10
timestamp 1696948209
transform 0 -1 2605 -1 0 18010
box -386 -240 386 240
use sky130_fd_pr__cap_mim_m3_1_FJFAMD  sky130_fd_pr__cap_mim_m3_1_FJFAMD_11
timestamp 1696948209
transform 0 -1 3335 1 0 18010
box -386 -240 386 240
use sky130_fd_pr__cap_mim_m3_1_FJFAMD  sky130_fd_pr__cap_mim_m3_1_FJFAMD_12
timestamp 1696948209
transform 0 1 273 1 0 15836
box -386 -240 386 240
use sky130_fd_pr__cap_mim_m3_1_FJFAMD  sky130_fd_pr__cap_mim_m3_1_FJFAMD_13
timestamp 1696948209
transform 0 1 1003 -1 0 11618
box -386 -240 386 240
use sky130_fd_pr__cap_mim_m3_1_FJFAMD  sky130_fd_pr__cap_mim_m3_1_FJFAMD_14
timestamp 1696948209
transform 0 1 273 1 0 11618
box -386 -240 386 240
use sky130_fd_pr__cap_mim_m3_1_FJFAMD  sky130_fd_pr__cap_mim_m3_1_FJFAMD_15
timestamp 1696948209
transform 0 -1 2605 -1 0 12640
box -386 -240 386 240
use sky130_fd_pr__cap_mim_m3_1_FJFAMD  sky130_fd_pr__cap_mim_m3_1_FJFAMD_16
timestamp 1696948209
transform 0 1 273 1 0 16858
box -386 -240 386 240
use sky130_fd_pr__cap_mim_m3_1_FJFAMD  sky130_fd_pr__cap_mim_m3_1_FJFAMD_17
timestamp 1696948209
transform 0 1 1003 -1 0 16858
box -386 -240 386 240
use sky130_fd_pr__cap_mim_m3_1_FJFAMD  sky130_fd_pr__cap_mim_m3_1_FJFAMD_18
timestamp 1696948209
transform 0 -1 2605 -1 0 16858
box -386 -240 386 240
use sky130_fd_pr__cap_mim_m3_1_FJFAMD  sky130_fd_pr__cap_mim_m3_1_FJFAMD_19
timestamp 1696948209
transform 0 -1 3335 1 0 16858
box -386 -240 386 240
use sky130_fd_pr__cap_mim_m3_1_FJFAMD  sky130_fd_pr__cap_mim_m3_1_FJFAMD_20
timestamp 1696948209
transform 0 1 1003 -1 0 12640
box -386 -240 386 240
use sky130_fd_pr__cap_mim_m3_1_FJFAMD  sky130_fd_pr__cap_mim_m3_1_FJFAMD_21
timestamp 1696948209
transform 0 1 273 1 0 12640
box -386 -240 386 240
use sky130_fd_pr__cap_mim_m3_1_FJFAMD  sky130_fd_pr__cap_mim_m3_1_FJFAMD_22
timestamp 1696948209
transform 0 -1 3335 1 0 11618
box -386 -240 386 240
use sky130_fd_pr__cap_mim_m3_1_FJFAMD  sky130_fd_pr__cap_mim_m3_1_FJFAMD_23
timestamp 1696948209
transform 0 -1 3335 1 0 12640
box -386 -240 386 240
use sky130_fd_pr__cap_mim_m3_1_FJFAMD  sky130_fd_pr__cap_mim_m3_1_FJFAMD_24
timestamp 1696948209
transform 0 -1 3335 1 0 9444
box -386 -240 386 240
use sky130_fd_pr__cap_mim_m3_1_FJFAMD  sky130_fd_pr__cap_mim_m3_1_FJFAMD_25
timestamp 1696948209
transform 0 1 273 1 0 9444
box -386 -240 386 240
use sky130_fd_pr__cap_mim_m3_1_FJFAMD  sky130_fd_pr__cap_mim_m3_1_FJFAMD_26
timestamp 1696948209
transform 0 1 1003 -1 0 9444
box -386 -240 386 240
use sky130_fd_pr__cap_mim_m3_1_FJFAMD  sky130_fd_pr__cap_mim_m3_1_FJFAMD_27
timestamp 1696948209
transform 0 -1 2605 -1 0 9444
box -386 -240 386 240
use sky130_fd_pr__cap_mim_m3_1_FJFAMD  sky130_fd_pr__cap_mim_m3_1_FJFAMD_28
timestamp 1696948209
transform 0 -1 2605 -1 0 8422
box -386 -240 386 240
use sky130_fd_pr__cap_mim_m3_1_FJFAMD  sky130_fd_pr__cap_mim_m3_1_FJFAMD_29
timestamp 1696948209
transform 0 1 1003 -1 0 8422
box -386 -240 386 240
use sky130_fd_pr__cap_mim_m3_1_FJFAMD  sky130_fd_pr__cap_mim_m3_1_FJFAMD_30
timestamp 1696948209
transform 0 1 273 1 0 8422
box -386 -240 386 240
use sky130_fd_pr__cap_mim_m3_1_FJFAMD  sky130_fd_pr__cap_mim_m3_1_FJFAMD_31
timestamp 1696948209
transform 0 -1 3335 1 0 8422
box -386 -240 386 240
use sky130_fd_pr__cap_mim_m3_1_FJFAMD  sky130_fd_pr__cap_mim_m3_1_FJFAMD_32
timestamp 1696948209
transform 0 -1 2605 -1 0 7400
box -386 -240 386 240
use sky130_fd_pr__cap_mim_m3_1_FJFAMD  sky130_fd_pr__cap_mim_m3_1_FJFAMD_33
timestamp 1696948209
transform 0 1 1003 -1 0 7400
box -386 -240 386 240
use sky130_fd_pr__cap_mim_m3_1_FJFAMD  sky130_fd_pr__cap_mim_m3_1_FJFAMD_34
timestamp 1696948209
transform 0 1 273 1 0 7400
box -386 -240 386 240
use sky130_fd_pr__cap_mim_m3_1_FJFAMD  sky130_fd_pr__cap_mim_m3_1_FJFAMD_35
timestamp 1696948209
transform 0 -1 3335 1 0 7400
box -386 -240 386 240
use sky130_fd_pr__cap_mim_m3_1_FJFAMD  sky130_fd_pr__cap_mim_m3_1_FJFAMD_36
timestamp 1696948209
transform 0 1 273 1 0 10466
box -386 -240 386 240
use sky130_fd_pr__cap_mim_m3_1_FJFAMD  sky130_fd_pr__cap_mim_m3_1_FJFAMD_37
timestamp 1696948209
transform 0 1 1003 -1 0 10466
box -386 -240 386 240
use sky130_fd_pr__cap_mim_m3_1_FJFAMD  sky130_fd_pr__cap_mim_m3_1_FJFAMD_38
timestamp 1696948209
transform 0 -1 2605 -1 0 10466
box -386 -240 386 240
use sky130_fd_pr__cap_mim_m3_1_FJFAMD  sky130_fd_pr__cap_mim_m3_1_FJFAMD_39
timestamp 1696948209
transform 0 -1 3335 1 0 10466
box -386 -240 386 240
use sky130_fd_pr__cap_mim_m3_1_FJFAMD  sky130_fd_pr__cap_mim_m3_1_FJFAMD_40
timestamp 1696948209
transform 0 1 1003 -1 0 13662
box -386 -240 386 240
use sky130_fd_pr__cap_mim_m3_1_FJFAMD  sky130_fd_pr__cap_mim_m3_1_FJFAMD_41
timestamp 1696948209
transform 0 1 273 1 0 13662
box -386 -240 386 240
use sky130_fd_pr__cap_mim_m3_1_FJFAMD  sky130_fd_pr__cap_mim_m3_1_FJFAMD_42
timestamp 1696948209
transform 0 -1 2605 -1 0 13662
box -386 -240 386 240
use sky130_fd_pr__cap_mim_m3_1_FJFAMD  sky130_fd_pr__cap_mim_m3_1_FJFAMD_43
timestamp 1696948209
transform 0 1 273 1 0 14684
box -386 -240 386 240
use sky130_fd_pr__cap_mim_m3_1_FJFAMD  sky130_fd_pr__cap_mim_m3_1_FJFAMD_44
timestamp 1696948209
transform 0 1 1003 -1 0 14684
box -386 -240 386 240
use sky130_fd_pr__cap_mim_m3_1_FJFAMD  sky130_fd_pr__cap_mim_m3_1_FJFAMD_45
timestamp 1696948209
transform 0 -1 2605 -1 0 14684
box -386 -240 386 240
use sky130_fd_pr__cap_mim_m3_1_FJFAMD  sky130_fd_pr__cap_mim_m3_1_FJFAMD_46
timestamp 1696948209
transform 0 -1 3335 1 0 14684
box -386 -240 386 240
use sky130_fd_pr__cap_mim_m3_1_FJFAMD  sky130_fd_pr__cap_mim_m3_1_FJFAMD_47
timestamp 1696948209
transform 0 -1 3335 1 0 13662
box -386 -240 386 240
use sky130_fd_pr__nfet_01v8_722GYZ  sky130_fd_pr__nfet_01v8_722GYZ_0
timestamp 1696948209
transform 1 0 1804 0 -1 12716
box -311 -310 311 310
use sky130_fd_pr__nfet_01v8_722GYZ  sky130_fd_pr__nfet_01v8_722GYZ_1
timestamp 1696948209
transform 1 0 1804 0 -1 19108
box -311 -310 311 310
use sky130_fd_pr__nfet_01v8_722GYZ  sky130_fd_pr__nfet_01v8_722GYZ_2
timestamp 1696948209
transform 1 0 1804 0 -1 20130
box -311 -310 311 310
use sky130_fd_pr__nfet_01v8_722GYZ  sky130_fd_pr__nfet_01v8_722GYZ_3
timestamp 1696948209
transform 1 0 1804 0 -1 18086
box -311 -310 311 310
use sky130_fd_pr__nfet_01v8_722GYZ  sky130_fd_pr__nfet_01v8_722GYZ_4
timestamp 1696948209
transform 1 0 1804 0 -1 15912
box -311 -310 311 310
use sky130_fd_pr__nfet_01v8_722GYZ  sky130_fd_pr__nfet_01v8_722GYZ_5
timestamp 1696948209
transform 1 0 1804 0 -1 8498
box -311 -310 311 310
use sky130_fd_pr__nfet_01v8_722GYZ  sky130_fd_pr__nfet_01v8_722GYZ_6
timestamp 1696948209
transform 1 0 1804 0 -1 16934
box -311 -310 311 310
use sky130_fd_pr__nfet_01v8_722GYZ  sky130_fd_pr__nfet_01v8_722GYZ_7
timestamp 1696948209
transform 1 0 1804 0 -1 14760
box -311 -310 311 310
use sky130_fd_pr__nfet_01v8_722GYZ  sky130_fd_pr__nfet_01v8_722GYZ_8
timestamp 1696948209
transform 1 0 1804 0 -1 10542
box -311 -310 311 310
use sky130_fd_pr__nfet_01v8_DGP55P  sky130_fd_pr__nfet_01v8_DGP55P_0
timestamp 1696943242
transform 1 0 1804 0 1 20769
box -596 -229 596 229
use sky130_fd_pr__nfet_01v8_L9WNCD  sky130_fd_pr__nfet_01v8_L9WNCD_0
timestamp 1696943731
transform 1 0 2505 0 1 20769
box -211 -229 211 229
use sky130_fd_pr__nfet_01v8_L9WNCD  sky130_fd_pr__nfet_01v8_L9WNCD_1
timestamp 1696943731
transform 1 0 1103 0 1 20769
box -211 -229 211 229
use sky130_fd_pr__nfet_01v8_QWA63T  sky130_fd_pr__nfet_01v8_QWA63T_1
timestamp 1696930192
transform -1 0 1804 0 1 4338
box -455 -260 455 260
use sky130_fd_pr__pfet_01v8_4N94TK  sky130_fd_pr__pfet_01v8_4N94TK_0
timestamp 1696943242
transform 1 0 2355 0 1 21668
box -361 -334 361 334
use sky130_fd_pr__pfet_01v8_4N94TK  sky130_fd_pr__pfet_01v8_4N94TK_1
timestamp 1696943242
transform 1 0 1253 0 1 21668
box -361 -334 361 334
use sky130_fd_pr__pfet_01v8_ADYTEV  sky130_fd_pr__pfet_01v8_ADYTEV_0
timestamp 1696943242
transform 1 0 1804 0 1 21668
box -296 -334 296 334
use sky130_fd_pr__pfet_01v8_UAU7GH  sky130_fd_pr__pfet_01v8_UAU7GH_0
timestamp 1696931086
transform -1 0 1804 0 1 5797
box -455 -319 455 319
use sky130_fd_sc_hd__buf_1  sky130_fd_sc_hd__buf_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform -1 0 838 0 -1 1602
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform -1 0 568 0 -1 1602
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_1
timestamp 1694700623
transform 1 0 2016 0 -1 3336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_2
timestamp 1694700623
transform 1 0 2784 0 -1 3336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_3
timestamp 1694700623
transform -1 0 570 0 -1 3336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_4
timestamp 1694700623
transform -1 0 1594 0 -1 3336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_5
timestamp 1694700623
transform -1 0 1338 0 -1 3336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_6
timestamp 1694700623
transform -1 0 1082 0 -1 3336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_7
timestamp 1694700623
transform -1 0 826 0 -1 3336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_8
timestamp 1694700623
transform 1 0 3296 0 -1 3336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_9
timestamp 1694700623
transform -1 0 314 0 -1 3336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_10
timestamp 1694700623
transform 1 0 3296 0 -1 1602
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_11
timestamp 1694700623
transform -1 0 312 0 -1 1602
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_12
timestamp 1694700623
transform -1 0 1558 0 -1 22978
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_13
timestamp 1694700623
transform -1 0 2326 0 -1 22978
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_14
timestamp 1694700623
transform -1 0 2070 0 -1 22978
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_15
timestamp 1694700623
transform -1 0 1814 0 -1 22978
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  x2
timestamp 1694700623
transform 1 0 3040 0 -1 3336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  x3
timestamp 1694700623
transform 1 0 3040 0 -1 1602
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_1  x7 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 838 0 -1 1602
box -38 -48 1970 592
use sky130_fd_sc_hd__inv_1  x8
timestamp 1694700623
transform 1 0 2528 0 -1 3336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  x9
timestamp 1694700623
transform 1 0 2272 0 -1 3336
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  x11
timestamp 1694700623
transform 1 0 2770 0 -1 1602
box -38 -48 314 592
use sky130_fd_sc_hd__nand2b_1  x18 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 1574 0 -1 3336
box -38 -48 498 592
<< labels >>
flabel metal1 2579 22930 3166 23026 0 FreeSans 320 0 0 0 vss_startup
port 0 nsew
flabel metal1 2579 22386 3166 22482 0 FreeSans 320 0 0 0 vdd_startup
port 1 nsew
flabel metal3 892 22242 2716 22338 0 FreeSans 320 0 0 0 uwb_trigger
port 2 nsew
flabel metal1 1293 14582 1837 14628 0 FreeSans 240 0 0 0 delay_line[4]
port 4 nsew
flabel metal1 1293 16756 1837 16802 0 FreeSans 240 0 0 0 delay_line[3]
port 5 nsew
flabel metal1 1293 17908 1837 17954 0 FreeSans 240 0 0 0 delay_line[2]
port 6 nsew
flabel metal1 1293 18930 1837 18976 0 FreeSans 240 0 0 0 delay_line[1]
port 7 nsew
flabel metal1 1293 19952 1837 19998 0 FreeSans 240 0 0 0 delay_line[0]
port 8 nsew
flabel metal2 2066 2 2138 1322 0 FreeSans 240 90 0 0 trigger_line[1]
port 9 nsew
flabel metal2 1474 2 1546 1256 0 FreeSans 240 90 0 0 trigger_line[0]
port 10 nsew
flabel metal4 3344 2 3544 2648 0 FreeSans 1600 90 0 0 osc_trigger2
port 12 nsew
flabel metal4 66 2 266 2648 0 FreeSans 1600 90 0 0 osc_trigger1
port 11 nsew
flabel metal1 1293 10364 1837 10410 0 FreeSans 240 0 0 0 delay_line[5]
port 3 nsew
<< end >>
