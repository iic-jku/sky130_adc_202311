magic
tech sky130A
magscale 1 2
timestamp 1697705955
<< pwell >>
rect -134 188 -24 938
rect 1050 188 1160 938
rect 30 14 96 150
rect 921 109 927 161
rect 930 14 996 150
<< locali >>
rect -134 188 16 938
rect 1010 188 1160 938
rect 30 14 96 150
rect 930 14 996 150
<< metal1 >>
rect -87 1588 -39 1732
rect -89 1582 -37 1588
rect -89 1476 -37 1482
rect -87 -62 -39 1476
rect 9 1300 57 1732
rect 103 1726 155 1732
rect 103 1620 155 1626
rect 7 1294 59 1300
rect 7 1188 59 1194
rect 9 926 57 1188
rect 105 926 153 1620
rect 201 1444 249 1732
rect 199 1438 251 1444
rect 199 1332 251 1338
rect 201 926 249 1332
rect 297 1300 345 1732
rect 393 1444 441 1732
rect 487 1726 539 1732
rect 487 1620 539 1626
rect 489 1588 537 1620
rect 487 1582 539 1588
rect 487 1476 539 1482
rect 391 1438 443 1444
rect 391 1332 443 1338
rect 295 1294 347 1300
rect 295 1188 347 1194
rect 297 926 345 1188
rect 393 926 441 1332
rect 489 926 537 1476
rect 585 1444 633 1732
rect 583 1438 635 1444
rect 583 1332 635 1338
rect 585 926 633 1332
rect 681 1300 729 1732
rect 777 1444 825 1732
rect 873 1588 921 1732
rect 871 1582 923 1588
rect 871 1476 923 1482
rect 775 1438 827 1444
rect 775 1332 827 1338
rect 679 1294 731 1300
rect 679 1188 731 1194
rect 681 926 729 1188
rect 777 926 825 1332
rect 873 926 921 1476
rect 969 1300 1017 1732
rect 1063 1726 1115 1732
rect 1063 1620 1115 1626
rect 967 1294 1019 1300
rect 967 1188 1019 1194
rect 969 926 1017 1188
rect 105 110 206 156
rect 258 110 345 156
rect 369 110 384 156
rect 450 110 576 156
rect 642 110 768 156
rect 820 110 921 156
rect 105 -62 153 110
rect -89 -68 -37 -62
rect -89 -174 -37 -168
rect 103 -68 155 -62
rect 103 -174 155 -168
rect -87 -465 -39 -174
rect 105 -465 153 -174
rect 297 -465 345 110
rect 489 -62 537 110
rect 487 -68 539 -62
rect 487 -174 539 -168
rect 489 -465 537 -174
rect 681 -465 729 110
rect 873 -62 921 110
rect 1065 -62 1113 1620
rect 871 -68 923 -62
rect 871 -174 923 -168
rect 1063 -68 1115 -62
rect 1063 -174 1115 -168
rect 873 -465 921 -174
rect 1065 -465 1113 -174
<< via1 >>
rect -89 1482 -37 1582
rect 103 1626 155 1726
rect 7 1194 59 1294
rect 199 1338 251 1438
rect 487 1626 539 1726
rect 487 1482 539 1582
rect 391 1338 443 1438
rect 295 1194 347 1294
rect 583 1338 635 1438
rect 871 1482 923 1582
rect 775 1338 827 1438
rect 679 1194 731 1294
rect 1063 1626 1115 1726
rect 967 1194 1019 1294
rect -89 -168 -37 -68
rect 103 -168 155 -68
rect 487 -168 539 -68
rect 871 -168 923 -68
rect 1063 -168 1115 -68
<< metal2 >>
rect 103 1726 155 1732
rect -134 1628 103 1724
rect 487 1726 539 1732
rect 155 1628 487 1724
rect 103 1620 155 1626
rect 487 1620 539 1626
rect 1063 1726 1115 1732
rect 1115 1628 1160 1724
rect 1063 1620 1115 1626
rect -89 1582 -37 1588
rect -134 1484 -89 1580
rect -89 1476 -37 1482
rect 487 1582 539 1588
rect 871 1582 923 1588
rect 539 1484 871 1580
rect 487 1476 539 1482
rect 923 1484 1160 1580
rect 871 1476 923 1482
rect 199 1438 251 1444
rect -94 1340 199 1436
rect 391 1438 443 1444
rect 251 1340 391 1436
rect 199 1332 251 1338
rect 583 1438 635 1444
rect 443 1340 583 1436
rect 391 1332 443 1338
rect 775 1438 827 1444
rect 635 1340 775 1436
rect 583 1332 635 1338
rect 827 1340 1118 1436
rect 775 1332 827 1338
rect 7 1294 59 1300
rect -134 1196 7 1292
rect 295 1294 347 1300
rect 59 1196 295 1292
rect 7 1188 59 1194
rect 679 1294 731 1300
rect 347 1196 679 1292
rect 295 1188 347 1194
rect 967 1294 1019 1300
rect 731 1196 967 1292
rect 679 1188 731 1194
rect 1019 1196 1160 1292
rect 967 1188 1019 1194
rect -89 -68 -37 -62
rect -94 -166 -89 -70
rect 103 -68 155 -62
rect -37 -166 103 -70
rect -89 -174 -37 -168
rect 487 -68 539 -62
rect 155 -166 487 -70
rect 103 -174 155 -168
rect 871 -68 923 -62
rect 539 -166 871 -70
rect 487 -174 539 -168
rect 1063 -68 1115 -62
rect 923 -166 1063 -70
rect 871 -174 923 -168
rect 1115 -166 1120 -70
rect 1063 -174 1115 -168
rect -134 -310 1160 -214
rect -134 -454 1160 -358
use sky130_fd_pr__nfet_01v8_QMBXET  sky130_fd_pr__nfet_01v8_QMBXET_0
timestamp 1697705955
transform 1 0 513 0 1 563
box -647 -585 647 585
<< labels >>
flabel locali -134 188 16 938 0 FreeSans 320 0 0 0 VSUB
port 0 nsew
flabel locali 1010 188 1160 938 0 FreeSans 320 0 0 0 VSUB
port 0 nsew
flabel metal2 -134 1628 -89 1724 0 FreeSans 128 0 0 0 drain
port 2 nsew
flabel metal2 -134 1484 -89 1580 0 FreeSans 128 0 0 0 gate
port 1 nsew
flabel metal2 -134 -310 -89 -214 0 FreeSans 176 0 0 0 en1
port 3 nsew
flabel metal2 -134 -454 -89 -358 0 FreeSans 176 0 0 0 en2
port 4 nsew
<< end >>
