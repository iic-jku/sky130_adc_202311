magic
tech sky130A
magscale 1 2
timestamp 1697439515
<< nwell >>
rect 7361 -28333 7562 -28012
rect 11146 -28333 11361 -28012
rect 7361 -30067 11361 -29746
<< pwell >>
rect 7361 -28610 11361 -28391
rect 7361 -28634 7631 -28610
rect 11108 -28634 11361 -28610
rect 7361 -30368 11361 -30125
<< psubdiff >>
rect 7440 -28442 7484 -28418
rect 7440 -28584 7484 -28560
rect 11198 -28442 11242 -28418
rect 11198 -28584 11242 -28560
rect 7440 -30176 7484 -30152
rect 7440 -30318 7484 -30294
rect 11198 -30176 11242 -30152
rect 11198 -30318 11242 -30294
<< nsubdiff >>
rect 7398 -28076 7520 -28051
rect 7398 -28297 7520 -28270
rect 11162 -28076 11284 -28051
rect 11162 -28297 11284 -28270
rect 7398 -29810 7520 -29785
rect 7398 -30031 7520 -30004
rect 11162 -29810 11284 -29785
rect 11162 -30031 11284 -30004
<< psubdiffcont >>
rect 7440 -28560 7484 -28442
rect 11198 -28560 11242 -28442
rect 7440 -30294 7484 -30176
rect 11198 -30294 11242 -30176
<< nsubdiffcont >>
rect 7398 -28270 7520 -28076
rect 11162 -28270 11284 -28076
rect 7398 -30004 7520 -29810
rect 11162 -30004 11284 -29810
<< locali >>
rect 7379 -28076 7659 -28042
rect 7379 -28270 7398 -28076
rect 7520 -28270 7659 -28076
rect 7379 -28301 7659 -28270
rect 11009 -28076 11284 -28051
rect 11009 -28270 11162 -28076
rect 11009 -28297 11284 -28270
rect 7638 -28424 7784 -28362
rect 7974 -28378 8151 -28342
rect 9470 -28332 9538 -28314
rect 9470 -28368 9486 -28332
rect 9520 -28368 9538 -28332
rect 9470 -28370 9538 -28368
rect 10286 -28397 10340 -28323
rect 10552 -28378 10692 -28342
rect 10896 -28386 11042 -28362
rect 7440 -28442 7784 -28424
rect 7484 -28560 7784 -28442
rect 7440 -28578 7784 -28560
rect 10896 -28442 11247 -28386
rect 10896 -28560 11198 -28442
rect 11242 -28560 11247 -28442
rect 10896 -28578 11247 -28560
rect 7440 -28584 7644 -28578
rect 11013 -28592 11247 -28578
rect 7379 -29810 7678 -29776
rect 7379 -30004 7398 -29810
rect 7520 -30004 7678 -29810
rect 7379 -30035 7678 -30004
rect 11026 -29810 11284 -29785
rect 11026 -30004 11162 -29810
rect 11026 -30031 11284 -30004
rect 7640 -30158 7786 -30096
rect 7440 -30176 7786 -30158
rect 7484 -30294 7786 -30176
rect 7440 -30312 7786 -30294
rect 7896 -30312 8042 -30096
rect 8246 -30112 8454 -30064
rect 8758 -30112 8966 -30064
rect 9726 -30112 9924 -30064
rect 10228 -30112 10436 -30064
rect 10640 -30280 10786 -30110
rect 7440 -30314 7734 -30312
rect 7440 -30318 7618 -30314
rect 10672 -30326 10786 -30280
rect 10896 -30120 11042 -30110
rect 10896 -30176 11247 -30120
rect 10896 -30294 11198 -30176
rect 11242 -30294 11247 -30176
rect 10896 -30326 11247 -30294
<< viali >>
rect 7882 -28366 7916 -28330
rect 8274 -28364 8308 -28328
rect 8396 -28366 8430 -28330
rect 8524 -28366 8558 -28330
rect 9022 -28368 9056 -28332
rect 9334 -28368 9368 -28332
rect 9486 -28368 9520 -28332
rect 9606 -28362 9640 -28326
rect 10372 -28364 10406 -28328
rect 10764 -28364 10798 -28328
rect 8638 -30114 8672 -30070
rect 9022 -30112 9056 -30072
rect 9148 -30108 9182 -30074
rect 9261 -30106 9295 -30072
rect 9484 -30114 9518 -30070
rect 9624 -30112 9658 -30072
rect 9996 -30114 10030 -30070
rect 10508 -30114 10542 -30070
<< metal1 >>
rect 7858 -28314 7930 -28308
rect 7858 -28370 7866 -28314
rect 7922 -28370 7930 -28314
rect 7858 -28376 7930 -28370
rect 8242 -28314 8314 -28308
rect 8242 -28370 8250 -28314
rect 8306 -28328 8314 -28314
rect 8308 -28364 8314 -28328
rect 8306 -28370 8314 -28364
rect 8242 -28376 8314 -28370
rect 8370 -28314 8442 -28308
rect 8370 -28370 8378 -28314
rect 8434 -28370 8442 -28314
rect 8370 -28376 8442 -28370
rect 8498 -28314 8570 -28308
rect 8498 -28370 8506 -28314
rect 8562 -28370 8570 -28314
rect 8498 -28376 8570 -28370
rect 9010 -28314 9082 -28306
rect 9010 -28370 9018 -28314
rect 9074 -28370 9082 -28314
rect 9010 -28378 9082 -28370
rect 9308 -28314 9380 -28308
rect 9308 -28370 9316 -28314
rect 9372 -28370 9380 -28314
rect 9308 -28376 9380 -28370
rect 9474 -28314 9546 -28308
rect 9474 -28370 9482 -28314
rect 9538 -28370 9546 -28314
rect 9474 -28376 9546 -28370
rect 9592 -28314 9660 -28308
rect 9592 -28370 9598 -28314
rect 9654 -28370 9660 -28314
rect 9592 -28376 9660 -28370
rect 10366 -28314 10442 -28308
rect 10366 -28328 10378 -28314
rect 10366 -28364 10372 -28328
rect 10366 -28370 10378 -28364
rect 10434 -28370 10442 -28314
rect 10366 -28376 10442 -28370
rect 10754 -28314 10826 -28308
rect 10754 -28370 10762 -28314
rect 10818 -28370 10826 -28314
rect 10754 -28376 10826 -28370
rect 8498 -30064 8570 -30056
rect 8498 -30120 8506 -30064
rect 8562 -30120 8570 -30064
rect 8498 -30128 8570 -30120
rect 8626 -30064 8698 -30056
rect 8626 -30120 8634 -30064
rect 8690 -30120 8698 -30064
rect 8626 -30128 8698 -30120
rect 9010 -30064 9082 -30056
rect 9010 -30120 9018 -30064
rect 9074 -30120 9082 -30064
rect 9010 -30128 9082 -30120
rect 9138 -30064 9210 -30056
rect 9138 -30120 9146 -30064
rect 9202 -30120 9210 -30064
rect 9138 -30128 9210 -30120
rect 9249 -30064 9377 -30056
rect 9249 -30072 9313 -30064
rect 9249 -30106 9261 -30072
rect 9295 -30106 9313 -30072
rect 9249 -30120 9313 -30106
rect 9369 -30120 9377 -30064
rect 9249 -30128 9377 -30120
rect 9472 -30064 9544 -30056
rect 9472 -30120 9480 -30064
rect 9536 -30120 9544 -30064
rect 9472 -30128 9544 -30120
rect 9600 -30064 9672 -30056
rect 9600 -30120 9608 -30064
rect 9664 -30120 9672 -30064
rect 9600 -30128 9672 -30120
rect 9984 -30064 10056 -30056
rect 9984 -30120 9992 -30064
rect 10048 -30120 10056 -30064
rect 9984 -30128 10056 -30120
rect 10496 -30064 10568 -30056
rect 10496 -30120 10504 -30064
rect 10560 -30120 10568 -30064
rect 10496 -30128 10568 -30120
<< via1 >>
rect 7866 -28330 7922 -28314
rect 7866 -28366 7882 -28330
rect 7882 -28366 7916 -28330
rect 7916 -28366 7922 -28330
rect 7866 -28370 7922 -28366
rect 8250 -28328 8306 -28314
rect 8250 -28364 8274 -28328
rect 8274 -28364 8306 -28328
rect 8250 -28370 8306 -28364
rect 8378 -28330 8434 -28314
rect 8378 -28366 8396 -28330
rect 8396 -28366 8430 -28330
rect 8430 -28366 8434 -28330
rect 8378 -28370 8434 -28366
rect 8506 -28330 8562 -28314
rect 8506 -28366 8524 -28330
rect 8524 -28366 8558 -28330
rect 8558 -28366 8562 -28330
rect 8506 -28370 8562 -28366
rect 9018 -28332 9074 -28314
rect 9018 -28368 9022 -28332
rect 9022 -28368 9056 -28332
rect 9056 -28368 9074 -28332
rect 9018 -28370 9074 -28368
rect 9316 -28332 9372 -28314
rect 9316 -28368 9334 -28332
rect 9334 -28368 9368 -28332
rect 9368 -28368 9372 -28332
rect 9316 -28370 9372 -28368
rect 9482 -28332 9538 -28314
rect 9482 -28368 9486 -28332
rect 9486 -28368 9520 -28332
rect 9520 -28368 9538 -28332
rect 9482 -28370 9538 -28368
rect 9598 -28326 9654 -28314
rect 9598 -28362 9606 -28326
rect 9606 -28362 9640 -28326
rect 9640 -28362 9654 -28326
rect 9598 -28370 9654 -28362
rect 10378 -28328 10434 -28314
rect 10378 -28364 10406 -28328
rect 10406 -28364 10434 -28328
rect 10378 -28370 10434 -28364
rect 10762 -28328 10818 -28314
rect 10762 -28364 10764 -28328
rect 10764 -28364 10798 -28328
rect 10798 -28364 10818 -28328
rect 10762 -28370 10818 -28364
rect 8506 -30120 8562 -30064
rect 8634 -30070 8690 -30064
rect 8634 -30114 8638 -30070
rect 8638 -30114 8672 -30070
rect 8672 -30114 8690 -30070
rect 8634 -30120 8690 -30114
rect 9018 -30072 9074 -30064
rect 9018 -30112 9022 -30072
rect 9022 -30112 9056 -30072
rect 9056 -30112 9074 -30072
rect 9018 -30120 9074 -30112
rect 9146 -30074 9202 -30064
rect 9146 -30108 9148 -30074
rect 9148 -30108 9182 -30074
rect 9182 -30108 9202 -30074
rect 9146 -30120 9202 -30108
rect 9313 -30120 9369 -30064
rect 9480 -30070 9536 -30064
rect 9480 -30114 9484 -30070
rect 9484 -30114 9518 -30070
rect 9518 -30114 9536 -30070
rect 9480 -30120 9536 -30114
rect 9608 -30072 9664 -30064
rect 9608 -30112 9624 -30072
rect 9624 -30112 9658 -30072
rect 9658 -30112 9664 -30072
rect 9608 -30120 9664 -30112
rect 9992 -30070 10048 -30064
rect 9992 -30114 9996 -30070
rect 9996 -30114 10030 -30070
rect 10030 -30114 10048 -30070
rect 9992 -30120 10048 -30114
rect 10504 -30070 10560 -30064
rect 10504 -30114 10508 -30070
rect 10508 -30114 10542 -30070
rect 10542 -30114 10560 -30070
rect 10504 -30120 10560 -30114
<< metal2 >>
rect 7602 -28394 7674 -26994
rect 7730 -28394 7802 -26994
rect 7858 -28314 7930 -26994
rect 7858 -28370 7866 -28314
rect 7922 -28370 7930 -28314
rect 7858 -28394 7930 -28370
rect 7986 -28394 8058 -26994
rect 8114 -28394 8186 -26994
rect 8242 -27048 8314 -26994
rect 8242 -27132 8246 -27048
rect 8310 -27132 8314 -27048
rect 8242 -28314 8314 -27132
rect 8242 -28370 8250 -28314
rect 8306 -28370 8314 -28314
rect 8242 -28394 8314 -28370
rect 8370 -27624 8442 -26994
rect 8370 -27708 8374 -27624
rect 8438 -27708 8442 -27624
rect 8370 -28314 8442 -27708
rect 8370 -28370 8378 -28314
rect 8434 -28370 8442 -28314
rect 8370 -28394 8442 -28370
rect 8498 -27816 8570 -26994
rect 8498 -27900 8502 -27816
rect 8566 -27900 8570 -27816
rect 8498 -28314 8570 -27900
rect 8498 -28370 8506 -28314
rect 8562 -28370 8570 -28314
rect 8498 -28394 8570 -28370
rect 8626 -28394 8698 -26994
rect 8754 -28394 8826 -26994
rect 8882 -28394 8954 -26994
rect 9010 -28314 9082 -26994
rect 9010 -28370 9018 -28314
rect 9074 -28370 9082 -28314
rect 9010 -28394 9082 -28370
rect 9138 -28394 9210 -26994
rect 9308 -27240 9380 -26994
rect 9308 -27324 9312 -27240
rect 9376 -27324 9380 -27240
rect 9308 -28314 9380 -27324
rect 9308 -28370 9316 -28314
rect 9372 -28370 9380 -28314
rect 9308 -28394 9380 -28370
rect 9474 -27432 9546 -26994
rect 9474 -27516 9478 -27432
rect 9542 -27516 9546 -27432
rect 9474 -28314 9546 -27516
rect 9602 -28308 9674 -26994
rect 9474 -28370 9482 -28314
rect 9538 -28370 9546 -28314
rect 9474 -28394 9546 -28370
rect 9592 -28314 9674 -28308
rect 9592 -28370 9598 -28314
rect 9654 -28370 9674 -28314
rect 9592 -28394 9674 -28370
rect 9730 -28394 9802 -26994
rect 9858 -28394 9930 -26994
rect 9986 -28394 10058 -26994
rect 10114 -28394 10186 -26994
rect 10242 -28394 10314 -26994
rect 10370 -28314 10442 -26994
rect 10370 -28370 10378 -28314
rect 10434 -28370 10442 -28314
rect 10370 -28394 10442 -28370
rect 10498 -28394 10570 -26994
rect 10626 -28394 10698 -26994
rect 10754 -28314 10826 -26994
rect 10754 -28370 10762 -28314
rect 10818 -28370 10826 -28314
rect 10754 -28394 10826 -28370
rect 10882 -28394 10954 -26994
rect 11010 -28394 11082 -26994
rect 7602 -30320 7674 -28736
rect 7730 -30320 7802 -28736
rect 7858 -30320 7930 -28736
rect 7986 -30320 8058 -28736
rect 8114 -28782 8186 -28736
rect 8114 -28866 8118 -28782
rect 8182 -28866 8186 -28782
rect 8114 -30320 8186 -28866
rect 8242 -28782 8314 -28736
rect 8242 -28866 8246 -28782
rect 8310 -28866 8314 -28782
rect 8242 -30320 8314 -28866
rect 8370 -28782 8442 -28736
rect 8370 -28866 8374 -28782
rect 8438 -28866 8442 -28782
rect 8370 -30320 8442 -28866
rect 8498 -28782 8570 -28736
rect 8498 -28866 8502 -28782
rect 8566 -28866 8570 -28782
rect 8498 -28974 8570 -28866
rect 8498 -29058 8502 -28974
rect 8566 -29058 8570 -28974
rect 8498 -30064 8570 -29058
rect 8498 -30120 8506 -30064
rect 8562 -30120 8570 -30064
rect 8498 -30320 8570 -30120
rect 8626 -29166 8698 -28736
rect 8626 -29250 8630 -29166
rect 8694 -29250 8698 -29166
rect 8626 -30064 8698 -29250
rect 8626 -30120 8634 -30064
rect 8690 -30120 8698 -30064
rect 8626 -30320 8698 -30120
rect 8754 -30320 8826 -28736
rect 8882 -30320 8954 -28736
rect 9010 -29358 9082 -28736
rect 9010 -29442 9014 -29358
rect 9078 -29442 9082 -29358
rect 9010 -30064 9082 -29442
rect 9010 -30120 9018 -30064
rect 9074 -30120 9082 -30064
rect 9010 -30320 9082 -30120
rect 9138 -30064 9210 -28736
rect 9138 -30120 9146 -30064
rect 9202 -30120 9210 -30064
rect 9138 -30320 9210 -30120
rect 9305 -30064 9377 -28736
rect 9305 -30120 9313 -30064
rect 9369 -30120 9377 -30064
rect 9305 -30320 9377 -30120
rect 9472 -29550 9544 -28736
rect 9472 -29634 9476 -29550
rect 9540 -29634 9544 -29550
rect 9472 -30064 9544 -29634
rect 9472 -30120 9480 -30064
rect 9536 -30120 9544 -30064
rect 9472 -30320 9544 -30120
rect 9600 -29550 9672 -28736
rect 9600 -29634 9604 -29550
rect 9668 -29634 9672 -29550
rect 9600 -30064 9672 -29634
rect 9600 -30120 9608 -30064
rect 9664 -30120 9672 -30064
rect 9600 -30320 9672 -30120
rect 9728 -30320 9800 -28736
rect 9856 -30320 9928 -28736
rect 9984 -29358 10056 -28736
rect 9984 -29442 9988 -29358
rect 10052 -29442 10056 -29358
rect 9984 -30064 10056 -29442
rect 9984 -30120 9992 -30064
rect 10048 -30120 10056 -30064
rect 9984 -30320 10056 -30120
rect 10112 -29166 10184 -28736
rect 10112 -29250 10116 -29166
rect 10180 -29250 10184 -29166
rect 10112 -30320 10184 -29250
rect 10240 -30320 10312 -28736
rect 10368 -30320 10440 -28736
rect 10496 -28974 10568 -28736
rect 10496 -29058 10500 -28974
rect 10564 -29058 10568 -28974
rect 10496 -30064 10568 -29058
rect 10496 -30120 10504 -30064
rect 10560 -30120 10568 -30064
rect 10496 -30320 10568 -30120
rect 10624 -30320 10696 -28736
rect 10752 -30320 10824 -28736
rect 10880 -30320 10952 -28736
rect 11008 -30320 11080 -28736
<< via2 >>
rect 7866 -28370 7922 -28314
rect 8246 -27132 8310 -27048
rect 8374 -27708 8438 -27624
rect 8502 -27900 8566 -27816
rect 9312 -27324 9376 -27240
rect 9478 -27516 9542 -27432
rect 10762 -28370 10818 -28314
rect 8118 -28866 8182 -28782
rect 8246 -28866 8310 -28782
rect 8374 -28866 8438 -28782
rect 8502 -28866 8566 -28782
rect 8502 -29058 8566 -28974
rect 8630 -29250 8694 -29166
rect 9014 -29442 9078 -29358
rect 9476 -29634 9540 -29550
rect 9604 -29634 9668 -29550
rect 9988 -29442 10052 -29358
rect 10116 -29250 10180 -29166
rect 10500 -29058 10564 -28974
<< metal3 >>
rect 7361 -27048 11361 -27042
rect 7361 -27132 8246 -27048
rect 8310 -27052 11361 -27048
rect 8310 -27128 9252 -27052
rect 9430 -27128 11361 -27052
rect 8310 -27132 11361 -27128
rect 7361 -27138 11361 -27132
rect 7361 -27240 11361 -27234
rect 7361 -27244 9312 -27240
rect 7361 -27320 8124 -27244
rect 8302 -27320 9312 -27244
rect 7361 -27324 9312 -27320
rect 9376 -27324 11361 -27240
rect 7361 -27330 11361 -27324
rect 7361 -27432 11361 -27426
rect 7361 -27516 9478 -27432
rect 9542 -27436 11361 -27432
rect 9542 -27512 10378 -27436
rect 10556 -27512 11361 -27436
rect 9542 -27516 11361 -27512
rect 7361 -27522 11361 -27516
rect 7361 -27624 11361 -27618
rect 7361 -27708 8374 -27624
rect 8438 -27628 11361 -27624
rect 8438 -27704 8636 -27628
rect 8814 -27704 11361 -27628
rect 8438 -27708 11361 -27704
rect 7361 -27714 11361 -27708
rect 7361 -27816 11361 -27810
rect 7361 -27900 8502 -27816
rect 8566 -27820 11361 -27816
rect 8566 -27896 9866 -27820
rect 10044 -27896 11361 -27820
rect 8566 -27900 11361 -27896
rect 7361 -27906 11361 -27900
rect 7802 -28276 7930 -28266
rect 7802 -28384 7812 -28276
rect 7920 -28314 7930 -28276
rect 7922 -28370 7930 -28314
rect 7920 -28384 7930 -28370
rect 7802 -28394 7930 -28384
rect 10754 -28276 10882 -28266
rect 10754 -28314 10764 -28276
rect 10754 -28370 10762 -28314
rect 10754 -28384 10764 -28370
rect 10872 -28384 10882 -28276
rect 10754 -28394 10882 -28384
rect 7361 -28782 11361 -28776
rect 7361 -28866 8118 -28782
rect 8182 -28786 8246 -28782
rect 8182 -28866 8246 -28862
rect 8310 -28866 8374 -28782
rect 8438 -28866 8502 -28782
rect 8566 -28866 11361 -28782
rect 7361 -28872 11361 -28866
rect 7361 -28974 11361 -28968
rect 7361 -29058 8502 -28974
rect 8566 -28978 10500 -28974
rect 8566 -29054 10378 -28978
rect 8566 -29058 10500 -29054
rect 10564 -29058 11361 -28974
rect 7361 -29064 11361 -29058
rect 7361 -29166 11361 -29160
rect 7361 -29250 8630 -29166
rect 8694 -29170 10116 -29166
rect 8814 -29246 10116 -29170
rect 8694 -29250 10116 -29246
rect 10180 -29250 11361 -29166
rect 7361 -29256 11361 -29250
rect 7361 -29358 11361 -29352
rect 7361 -29442 9014 -29358
rect 9078 -29362 9988 -29358
rect 9078 -29438 9866 -29362
rect 9078 -29442 9988 -29438
rect 10052 -29442 11361 -29358
rect 7361 -29448 11361 -29442
rect 7361 -29550 11361 -29544
rect 7361 -29554 9476 -29550
rect 7361 -29630 9252 -29554
rect 9430 -29630 9476 -29554
rect 7361 -29634 9476 -29630
rect 9540 -29634 9604 -29550
rect 9668 -29634 11361 -29550
rect 7361 -29640 11361 -29634
rect 7360 -30032 11361 -29840
rect 7360 -30320 11361 -30128
<< via3 >>
rect 9252 -27128 9430 -27052
rect 8124 -27320 8302 -27244
rect 10378 -27512 10556 -27436
rect 8636 -27704 8814 -27628
rect 9866 -27896 10044 -27820
rect 7812 -28314 7920 -28276
rect 7812 -28370 7866 -28314
rect 7866 -28370 7920 -28314
rect 7812 -28384 7920 -28370
rect 10764 -28314 10872 -28276
rect 10764 -28370 10818 -28314
rect 10818 -28370 10872 -28314
rect 10764 -28384 10872 -28370
rect 8124 -28862 8182 -28786
rect 8182 -28862 8246 -28786
rect 8246 -28862 8302 -28786
rect 10378 -29054 10500 -28978
rect 10500 -29054 10556 -28978
rect 8636 -29246 8694 -29170
rect 8694 -29246 8814 -29170
rect 9866 -29438 9988 -29362
rect 9988 -29438 10044 -29362
rect 9252 -29630 9430 -29554
<< metal4 >>
rect 7602 -28266 7802 -26994
rect 8114 -27244 8314 -26994
rect 8114 -27320 8124 -27244
rect 8302 -27320 8314 -27244
rect 7602 -28276 7930 -28266
rect 7602 -28384 7812 -28276
rect 7920 -28384 7930 -28276
rect 7602 -28394 7930 -28384
rect 7602 -29640 7802 -28394
rect 8114 -28786 8314 -27320
rect 8114 -28862 8124 -28786
rect 8302 -28862 8314 -28786
rect 8114 -29640 8314 -28862
rect 8626 -27628 8826 -26994
rect 8626 -27704 8636 -27628
rect 8814 -27704 8826 -27628
rect 8626 -29170 8826 -27704
rect 8626 -29246 8636 -29170
rect 8814 -29246 8826 -29170
rect 8626 -29640 8826 -29246
rect 9241 -27052 9441 -26994
rect 9241 -27128 9252 -27052
rect 9430 -27128 9441 -27052
rect 9241 -29554 9441 -27128
rect 9241 -29630 9252 -29554
rect 9430 -29630 9441 -29554
rect 9241 -29640 9441 -29630
rect 9856 -27820 10056 -26994
rect 9856 -27896 9866 -27820
rect 10044 -27896 10056 -27820
rect 9856 -29362 10056 -27896
rect 9856 -29438 9866 -29362
rect 10044 -29438 10056 -29362
rect 9856 -29640 10056 -29438
rect 10368 -27436 10568 -26994
rect 10368 -27512 10378 -27436
rect 10556 -27512 10568 -27436
rect 10368 -28978 10568 -27512
rect 10880 -28266 11080 -26994
rect 10754 -28276 11080 -28266
rect 10754 -28384 10764 -28276
rect 10872 -28384 11080 -28276
rect 10754 -28394 11080 -28384
rect 10368 -29054 10378 -28978
rect 10556 -29054 10568 -28978
rect 10368 -29640 10568 -29054
rect 10880 -29640 11080 -28394
use sky130_fd_sc_hd__buf_1  sky130_fd_sc_hd__buf_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 8374 0 1 -28594
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_0
timestamp 1696857842
transform -1 0 8104 0 1 -28594
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_1
timestamp 1696857842
transform 1 0 9808 0 1 -30328
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_2
timestamp 1696857842
transform 1 0 10320 0 1 -30328
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_3
timestamp 1696857842
transform -1 0 8106 0 1 -30328
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_4
timestamp 1696857842
transform -1 0 9130 0 1 -30328
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_5
timestamp 1696857842
transform -1 0 8874 0 1 -30328
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_6
timestamp 1696857842
transform -1 0 8618 0 1 -30328
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_7
timestamp 1696857842
transform -1 0 8362 0 1 -30328
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_8
timestamp 1696857842
transform 1 0 10832 0 1 -30328
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_9
timestamp 1696857842
transform -1 0 7850 0 1 -30328
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_10
timestamp 1696857842
transform 1 0 10832 0 1 -28594
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_11
timestamp 1696857842
transform -1 0 7848 0 1 -28594
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  x2
timestamp 1696857842
transform 1 0 10576 0 1 -30328
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  x3
timestamp 1696857842
transform 1 0 10576 0 1 -28594
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_1  x7 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 8374 0 1 -28594
box -38 -48 1970 592
use sky130_fd_sc_hd__inv_1  x8
timestamp 1696857842
transform 1 0 10064 0 1 -30328
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  x9
timestamp 1696857842
transform 1 0 9552 0 1 -30328
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  x11
timestamp 1676037725
transform 1 0 10306 0 1 -28594
box -38 -48 314 592
use sky130_fd_sc_hd__nand2b_1  x18 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 9110 0 1 -30328
box -38 -48 498 592
<< end >>
