magic
tech sky130A
magscale 1 2
timestamp 1696579262
<< pwell >>
rect -359 -585 359 585
<< nmos >>
rect -159 -375 -129 375
rect -63 -375 -33 375
rect 33 -375 63 375
rect 129 -375 159 375
<< ndiff >>
rect -221 363 -159 375
rect -221 -363 -209 363
rect -175 -363 -159 363
rect -221 -375 -159 -363
rect -129 363 -63 375
rect -129 -363 -113 363
rect -79 -363 -63 363
rect -129 -375 -63 -363
rect -33 363 33 375
rect -33 -363 -17 363
rect 17 -363 33 363
rect -33 -375 33 -363
rect 63 363 129 375
rect 63 -363 79 363
rect 113 -363 129 363
rect 63 -375 129 -363
rect 159 363 221 375
rect 159 -363 175 363
rect 209 -363 221 363
rect 159 -375 221 -363
<< ndiffc >>
rect -209 -363 -175 363
rect -113 -363 -79 363
rect -17 -363 17 363
rect 79 -363 113 363
rect 175 -363 209 363
<< psubdiff >>
rect -323 515 -227 549
rect 227 515 323 549
rect -323 453 -289 515
rect 289 453 323 515
rect -323 -515 -289 -453
rect 289 -515 323 -453
rect -323 -549 -227 -515
rect 227 -549 323 -515
<< psubdiffcont >>
rect -227 515 227 549
rect -323 -453 -289 453
rect 289 -453 323 453
rect -227 -549 227 -515
<< poly >>
rect -159 375 -129 401
rect -63 375 -33 401
rect 33 375 63 401
rect 129 375 159 401
rect -159 -397 -129 -375
rect -63 -397 -33 -375
rect 33 -397 63 -375
rect 129 -397 159 -375
rect -159 -413 159 -397
rect -159 -447 -143 -413
rect 143 -447 159 -413
rect -159 -463 159 -447
<< polycont >>
rect -143 -447 143 -413
<< locali >>
rect -323 515 -227 549
rect 227 515 323 549
rect -323 453 -289 515
rect 289 453 323 515
rect -209 363 -175 379
rect -209 -379 -175 -363
rect -113 363 -79 379
rect -113 -379 -79 -363
rect -17 363 17 379
rect -17 -379 17 -363
rect 79 363 113 379
rect 79 -379 113 -363
rect 175 363 209 379
rect 175 -379 209 -363
rect -159 -447 -143 -413
rect 143 -447 159 -413
rect -323 -515 -289 -453
rect 289 -515 323 -453
rect -323 -549 -227 -515
rect 227 -549 323 -515
<< viali >>
rect -209 -363 -175 363
rect -113 -363 -79 363
rect -17 -363 17 363
rect 79 -363 113 363
rect 175 -363 209 363
<< metal1 >>
rect -215 363 -169 375
rect -215 -363 -209 363
rect -175 -363 -169 363
rect -215 -375 -169 -363
rect -119 363 -73 375
rect -119 -363 -113 363
rect -79 -363 -73 363
rect -119 -375 -73 -363
rect -23 363 23 375
rect -23 -363 -17 363
rect 17 -363 23 363
rect -23 -375 23 -363
rect 73 363 119 375
rect 73 -363 79 363
rect 113 -363 119 363
rect 73 -375 119 -363
rect 169 363 215 375
rect 169 -363 175 363
rect 209 -363 215 363
rect 169 -375 215 -363
<< properties >>
string FIXED_BBOX -306 -532 306 532
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 3.75 l 0.150 m 1 nf 4 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
