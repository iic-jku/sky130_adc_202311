magic
tech sky130A
magscale 1 2
timestamp 1698999411
<< nwell >>
rect -38 261 866 582
<< pwell >>
rect 12 21 827 203
rect 24 -17 58 21
<< scnmos >>
rect 111 47 141 177
rect 195 47 225 177
rect 279 47 309 177
rect 467 47 497 177
rect 551 47 581 177
rect 635 47 665 177
rect 719 47 749 177
<< scpmoshvt >>
rect 111 297 141 497
rect 207 297 237 497
rect 282 297 312 497
rect 467 297 497 497
rect 539 297 569 497
rect 635 297 665 497
rect 719 297 749 497
<< ndiff >>
rect 38 157 111 177
rect 38 123 50 157
rect 84 123 111 157
rect 38 89 111 123
rect 38 55 50 89
rect 84 55 111 89
rect 38 47 111 55
rect 141 93 195 177
rect 141 59 151 93
rect 185 59 195 93
rect 141 47 195 59
rect 225 163 279 177
rect 225 129 235 163
rect 269 129 279 163
rect 225 47 279 129
rect 309 93 361 177
rect 309 59 319 93
rect 353 59 361 93
rect 309 47 361 59
rect 415 95 467 177
rect 415 61 423 95
rect 457 61 467 95
rect 415 47 467 61
rect 497 163 551 177
rect 497 129 507 163
rect 541 129 551 163
rect 497 95 551 129
rect 497 61 507 95
rect 541 61 551 95
rect 497 47 551 61
rect 581 163 635 177
rect 581 129 591 163
rect 625 129 635 163
rect 581 95 635 129
rect 581 61 591 95
rect 625 61 635 95
rect 581 47 635 61
rect 665 163 719 177
rect 665 129 675 163
rect 709 129 719 163
rect 665 95 719 129
rect 665 61 675 95
rect 709 61 719 95
rect 665 47 719 61
rect 749 95 801 177
rect 749 61 759 95
rect 793 61 801 95
rect 749 47 801 61
<< pdiff >>
rect 46 477 111 497
rect 46 443 66 477
rect 100 443 111 477
rect 46 409 111 443
rect 46 375 66 409
rect 100 375 111 409
rect 46 341 111 375
rect 46 307 66 341
rect 100 307 111 341
rect 46 297 111 307
rect 141 488 207 497
rect 141 454 158 488
rect 192 454 207 488
rect 141 420 207 454
rect 141 386 158 420
rect 192 386 207 420
rect 141 297 207 386
rect 237 297 282 497
rect 312 477 467 497
rect 312 443 322 477
rect 356 443 423 477
rect 457 443 467 477
rect 312 409 467 443
rect 312 375 322 409
rect 356 375 423 409
rect 457 375 467 409
rect 312 297 467 375
rect 497 297 539 497
rect 569 477 635 497
rect 569 443 579 477
rect 613 443 635 477
rect 569 409 635 443
rect 569 375 579 409
rect 613 375 635 409
rect 569 297 635 375
rect 665 477 719 497
rect 665 443 675 477
rect 709 443 719 477
rect 665 409 719 443
rect 665 375 675 409
rect 709 375 719 409
rect 665 297 719 375
rect 749 477 801 497
rect 749 443 759 477
rect 793 443 801 477
rect 749 297 801 443
<< ndiffc >>
rect 50 123 84 157
rect 50 55 84 89
rect 151 59 185 93
rect 235 129 269 163
rect 319 59 353 93
rect 423 61 457 95
rect 507 129 541 163
rect 507 61 541 95
rect 591 129 625 163
rect 591 61 625 95
rect 675 129 709 163
rect 675 61 709 95
rect 759 61 793 95
<< pdiffc >>
rect 66 443 100 477
rect 66 375 100 409
rect 66 307 100 341
rect 158 454 192 488
rect 158 386 192 420
rect 322 443 356 477
rect 423 443 457 477
rect 322 375 356 409
rect 423 375 457 409
rect 579 443 613 477
rect 579 375 613 409
rect 675 443 709 477
rect 675 375 709 409
rect 759 443 793 477
<< poly >>
rect 111 497 141 523
rect 207 497 237 523
rect 282 497 312 523
rect 467 497 497 523
rect 539 497 569 523
rect 635 497 665 523
rect 719 497 749 523
rect 111 265 141 297
rect 207 265 237 297
rect 282 265 312 297
rect 467 265 497 297
rect 25 249 141 265
rect 25 215 35 249
rect 69 215 141 249
rect 25 195 141 215
rect 183 249 237 265
rect 183 215 193 249
rect 227 215 237 249
rect 183 199 237 215
rect 279 249 352 265
rect 279 215 308 249
rect 342 215 352 249
rect 279 199 352 215
rect 423 249 497 265
rect 423 215 433 249
rect 467 215 497 249
rect 423 199 497 215
rect 539 265 569 297
rect 635 265 665 297
rect 719 265 749 297
rect 539 249 593 265
rect 539 215 549 249
rect 583 215 593 249
rect 539 199 593 215
rect 635 249 749 265
rect 635 215 665 249
rect 699 215 749 249
rect 635 199 749 215
rect 111 177 141 195
rect 195 177 225 199
rect 279 177 309 199
rect 467 177 497 199
rect 551 177 581 199
rect 635 177 665 199
rect 719 177 749 199
rect 111 21 141 47
rect 195 21 225 47
rect 279 21 309 47
rect 467 21 497 47
rect 551 21 581 47
rect 635 21 665 47
rect 719 21 749 47
<< polycont >>
rect 35 215 69 249
rect 193 215 227 249
rect 308 215 342 249
rect 433 215 467 249
rect 549 215 583 249
rect 665 215 699 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 828 561
rect 50 477 116 493
rect 50 443 66 477
rect 100 443 116 477
rect 50 409 116 443
rect 50 375 66 409
rect 100 375 116 409
rect 50 341 116 375
rect 150 488 198 527
rect 150 454 158 488
rect 192 454 198 488
rect 150 420 198 454
rect 150 386 158 420
rect 192 386 198 420
rect 310 477 461 493
rect 310 443 322 477
rect 356 443 423 477
rect 457 443 461 477
rect 310 409 461 443
rect 559 477 625 527
rect 559 443 579 477
rect 613 443 625 477
rect 559 409 625 443
rect 150 370 198 386
rect 232 375 322 409
rect 356 375 423 409
rect 457 375 525 409
rect 50 307 66 341
rect 100 334 116 341
rect 232 334 266 375
rect 100 307 266 334
rect 50 299 266 307
rect 109 289 266 299
rect 17 249 69 265
rect 17 215 35 249
rect 17 195 69 215
rect 109 161 143 289
rect 300 255 358 341
rect 177 249 246 255
rect 177 215 193 249
rect 227 215 246 249
rect 280 249 358 255
rect 280 215 308 249
rect 342 215 358 249
rect 396 257 457 341
rect 491 325 525 375
rect 559 375 579 409
rect 613 375 625 409
rect 659 477 709 493
rect 659 443 675 477
rect 743 477 811 527
rect 743 443 759 477
rect 793 443 811 477
rect 659 409 709 443
rect 659 375 675 409
rect 709 375 811 409
rect 559 359 625 375
rect 491 291 683 325
rect 649 257 683 291
rect 396 249 493 257
rect 396 215 433 249
rect 467 215 493 249
rect 527 249 615 257
rect 527 215 549 249
rect 583 215 615 249
rect 649 249 715 257
rect 649 215 665 249
rect 699 215 715 249
rect 749 181 811 375
rect 34 157 143 161
rect 34 123 50 157
rect 84 127 143 157
rect 217 163 557 181
rect 217 129 235 163
rect 269 147 507 163
rect 269 129 294 147
rect 491 129 507 147
rect 541 129 557 163
rect 84 123 100 127
rect 34 89 100 123
rect 423 95 457 111
rect 34 55 50 89
rect 84 55 100 89
rect 134 59 151 93
rect 185 59 319 93
rect 353 59 371 93
rect 34 51 100 55
rect 423 17 457 61
rect 491 95 557 129
rect 491 61 507 95
rect 541 61 557 95
rect 491 54 557 61
rect 591 163 625 181
rect 591 95 625 129
rect 591 17 625 61
rect 659 163 811 181
rect 659 129 675 163
rect 709 147 811 163
rect 709 129 725 147
rect 659 95 725 129
rect 659 61 675 95
rect 709 61 725 95
rect 659 53 725 61
rect 759 95 793 113
rect 759 17 793 61
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 828 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
<< metal1 >>
rect 0 561 828 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 828 561
rect 0 496 828 527
rect 0 17 828 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 828 17
rect 0 -48 828 -17
<< labels >>
flabel metal1 s 24 -17 58 17 0 FreeSans 200 0 0 0 VGND
port 1 nsew
flabel metal1 s 28 527 62 561 0 FreeSans 200 0 0 0 VPWR
port 2 nsew
flabel locali s 300 289 334 323 0 FreeSans 400 0 0 0 B2
port 4 nsew
flabel locali s 396 289 430 323 0 FreeSans 400 0 0 0 A2
port 5 nsew
flabel locali s 396 221 430 255 0 FreeSans 400 0 0 0 A2
port 5 nsew
flabel locali s 764 357 798 391 0 FreeSans 400 0 0 0 X
port 7 nsew
flabel locali s 208 221 242 255 0 FreeSans 400 0 0 0 B1
port 3 nsew
flabel locali s 24 221 58 255 0 FreeSans 400 0 0 0 C1
port 8 nsew
flabel locali s 580 221 614 255 0 FreeSans 400 0 0 0 A1
port 6 nsew
flabel locali s 300 221 334 255 0 FreeSans 400 0 0 0 B2
port 4 nsew
rlabel comment s 0 0 0 0 4 o221a_2
flabel nwell s 28 527 62 561 0 FreeSans 200 0 0 0 VPB
port 10 nsew
flabel pwell s 24 -17 58 17 0 FreeSans 200 0 0 0 VNB
port 11 nsew
<< properties >>
string FIXED_BBOX 0 0 828 544
string path 3.350 1.900 9.275 1.900 
<< end >>
