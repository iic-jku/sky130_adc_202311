magic
tech sky130A
magscale 1 2
timestamp 1698999411
<< nwell >>
rect -38 261 314 582
<< pwell >>
rect 1 21 271 203
rect 30 -17 64 21
<< scnmos >>
rect 79 47 109 177
rect 163 47 193 177
<< scpmoshvt >>
rect 79 297 109 497
rect 151 297 181 497
<< ndiff >>
rect 27 163 79 177
rect 27 129 35 163
rect 69 129 79 163
rect 27 95 79 129
rect 27 61 35 95
rect 69 61 79 95
rect 27 47 79 61
rect 109 163 163 177
rect 109 129 119 163
rect 153 129 163 163
rect 109 95 163 129
rect 109 61 119 95
rect 153 61 163 95
rect 109 47 163 61
rect 193 163 245 177
rect 193 129 203 163
rect 237 129 245 163
rect 193 95 245 129
rect 193 61 203 95
rect 237 61 245 95
rect 193 47 245 61
<< pdiff >>
rect 27 485 79 497
rect 27 451 35 485
rect 69 451 79 485
rect 27 417 79 451
rect 27 383 35 417
rect 69 383 79 417
rect 27 349 79 383
rect 27 315 35 349
rect 69 315 79 349
rect 27 297 79 315
rect 109 297 151 497
rect 181 485 233 497
rect 181 451 191 485
rect 225 451 233 485
rect 181 417 233 451
rect 181 383 191 417
rect 225 383 233 417
rect 181 349 233 383
rect 181 315 191 349
rect 225 315 233 349
rect 181 297 233 315
<< ndiffc >>
rect 35 129 69 163
rect 35 61 69 95
rect 119 129 153 163
rect 119 61 153 95
rect 203 129 237 163
rect 203 61 237 95
<< pdiffc >>
rect 35 451 69 485
rect 35 383 69 417
rect 35 315 69 349
rect 191 451 225 485
rect 191 383 225 417
rect 191 315 225 349
<< poly >>
rect 79 497 109 523
rect 151 497 181 523
rect 79 265 109 297
rect 22 249 109 265
rect 22 215 37 249
rect 71 215 109 249
rect 151 265 181 297
rect 151 249 255 265
rect 151 235 205 249
rect 22 199 109 215
rect 79 177 109 199
rect 163 215 205 235
rect 239 215 255 249
rect 163 199 255 215
rect 163 177 193 199
rect 79 21 109 47
rect 163 21 193 47
<< polycont >>
rect 37 215 71 249
rect 205 215 239 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 276 561
rect 19 485 85 490
rect 19 451 35 485
rect 69 451 85 485
rect 19 417 85 451
rect 19 383 35 417
rect 69 383 85 417
rect 19 349 85 383
rect 19 315 35 349
rect 69 333 85 349
rect 191 485 257 527
rect 225 451 257 485
rect 191 417 257 451
rect 225 383 257 417
rect 191 349 257 383
rect 69 315 155 333
rect 19 299 155 315
rect 225 315 257 349
rect 191 299 257 315
rect 17 249 87 265
rect 17 215 37 249
rect 71 215 87 249
rect 121 179 155 299
rect 189 249 259 265
rect 189 215 205 249
rect 239 215 259 249
rect 21 163 69 179
rect 21 129 35 163
rect 21 95 69 129
rect 21 61 35 95
rect 21 17 69 61
rect 103 163 169 179
rect 103 129 119 163
rect 153 129 169 163
rect 103 95 169 129
rect 103 61 119 95
rect 153 61 169 95
rect 103 51 169 61
rect 203 163 257 179
rect 237 129 257 163
rect 203 95 257 129
rect 237 61 257 95
rect 203 17 257 61
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 276 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
<< metal1 >>
rect 0 561 276 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 276 561
rect 0 496 276 527
rect 0 17 276 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 276 17
rect 0 -48 276 -17
<< labels >>
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 1 nsew
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 2 nsew
flabel locali s 29 221 63 255 0 FreeSans 200 0 0 0 B
port 4 nsew
flabel locali s 30 425 64 459 0 FreeSans 200 0 0 0 Y
port 5 nsew
flabel locali s 213 221 247 255 0 FreeSans 200 0 0 0 A
port 3 nsew
rlabel comment s 0 0 0 0 4 nor2_1
flabel nwell s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 7 nsew
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 8 nsew
<< properties >>
string FIXED_BBOX 0 0 276 544
string path 0.000 0.000 6.900 0.000 
<< end >>
