magic
tech sky130A
magscale 1 2
timestamp 1515178157
<< checkpaint >>
rect -1298 -1308 3506 1852
<< nwell >>
rect -38 414 2246 582
rect -38 247 822 414
rect 1556 247 2246 414
<< pwell >>
rect 937 190 1514 372
rect 29 181 1514 190
rect 29 54 2121 181
rect 121 -17 155 54
rect 673 -17 707 54
rect 937 45 2121 54
rect 949 -17 983 45
rect 1225 -17 1351 45
rect 1777 -17 1811 45
<< scnmos >>
rect 113 80 851 164
rect 1021 71 1430 346
rect 1602 71 1632 155
rect 1698 71 1728 155
rect 1907 71 1937 155
rect 2003 71 2033 155
<< scpmoshvt >>
rect 285 283 569 443
rect 1661 329 1691 489
rect 1757 329 1787 489
rect 1995 329 2025 489
rect 2091 329 2121 489
<< ndiff >>
rect 963 325 1021 346
rect 963 291 975 325
rect 1009 291 1021 325
rect 963 257 1021 291
rect 963 223 975 257
rect 1009 223 1021 257
rect 963 189 1021 223
rect 55 126 113 164
rect 55 92 67 126
rect 101 92 113 126
rect 55 80 113 92
rect 851 135 909 164
rect 851 101 863 135
rect 897 101 909 135
rect 851 80 909 101
rect 963 155 975 189
rect 1009 155 1021 189
rect 963 121 1021 155
rect 963 87 975 121
rect 1009 87 1021 121
rect 963 71 1021 87
rect 1430 325 1488 346
rect 1430 291 1442 325
rect 1476 291 1488 325
rect 1430 257 1488 291
rect 1430 223 1442 257
rect 1476 223 1488 257
rect 1430 189 1488 223
rect 1430 155 1442 189
rect 1476 155 1488 189
rect 1430 121 1488 155
rect 1430 87 1442 121
rect 1476 87 1488 121
rect 1430 71 1488 87
rect 1542 130 1602 155
rect 1542 96 1552 130
rect 1586 96 1602 130
rect 1542 71 1602 96
rect 1632 131 1698 155
rect 1632 97 1648 131
rect 1682 97 1698 131
rect 1632 71 1698 97
rect 1728 131 1786 155
rect 1728 97 1744 131
rect 1778 97 1786 131
rect 1728 71 1786 97
rect 1845 121 1907 155
rect 1845 87 1857 121
rect 1891 87 1907 121
rect 1845 71 1907 87
rect 1937 131 2003 155
rect 1937 97 1953 131
rect 1987 97 2003 131
rect 1937 71 2003 97
rect 2033 131 2095 155
rect 2033 97 2049 131
rect 2083 97 2095 131
rect 2033 71 2095 97
<< pdiff >>
rect 1601 460 1661 489
rect 227 422 285 443
rect 227 388 239 422
rect 273 388 285 422
rect 227 283 285 388
rect 569 419 627 443
rect 569 385 581 419
rect 615 385 627 419
rect 569 351 627 385
rect 569 317 581 351
rect 615 317 627 351
rect 569 283 627 317
rect 1601 426 1611 460
rect 1645 426 1661 460
rect 1601 392 1661 426
rect 1601 358 1611 392
rect 1645 358 1661 392
rect 1601 329 1661 358
rect 1691 465 1757 489
rect 1691 431 1707 465
rect 1741 431 1757 465
rect 1691 397 1757 431
rect 1691 363 1707 397
rect 1741 363 1757 397
rect 1691 329 1757 363
rect 1787 459 1847 489
rect 1787 425 1803 459
rect 1837 425 1847 459
rect 1787 391 1847 425
rect 1787 357 1803 391
rect 1837 357 1847 391
rect 1787 329 1847 357
rect 1933 454 1995 489
rect 1933 420 1945 454
rect 1979 420 1995 454
rect 1933 329 1995 420
rect 2025 459 2091 489
rect 2025 425 2041 459
rect 2075 425 2091 459
rect 2025 391 2091 425
rect 2025 357 2041 391
rect 2075 357 2091 391
rect 2025 329 2091 357
rect 2121 459 2181 489
rect 2121 425 2137 459
rect 2171 425 2181 459
rect 2121 391 2181 425
rect 2121 357 2137 391
rect 2171 357 2181 391
rect 2121 329 2181 357
<< ndiffc >>
rect 975 291 1009 325
rect 975 223 1009 257
rect 67 92 101 126
rect 863 101 897 135
rect 975 155 1009 189
rect 975 87 1009 121
rect 1442 291 1476 325
rect 1442 223 1476 257
rect 1442 155 1476 189
rect 1442 87 1476 121
rect 1552 96 1586 130
rect 1648 97 1682 131
rect 1744 97 1778 131
rect 1857 87 1891 121
rect 1953 97 1987 131
rect 2049 97 2083 131
<< pdiffc >>
rect 239 388 273 422
rect 581 385 615 419
rect 581 317 615 351
rect 1611 426 1645 460
rect 1611 358 1645 392
rect 1707 431 1741 465
rect 1707 363 1741 397
rect 1803 425 1837 459
rect 1803 357 1837 391
rect 1945 420 1979 454
rect 2041 425 2075 459
rect 2041 357 2075 391
rect 2137 425 2171 459
rect 2137 357 2171 391
<< poly >>
rect 1661 489 1691 515
rect 1757 489 1787 515
rect 1995 489 2025 515
rect 2091 489 2121 515
rect 285 443 569 479
rect 650 428 1430 438
rect 649 418 1430 428
rect 649 384 1116 418
rect 1150 384 1184 418
rect 1218 384 1252 418
rect 1286 384 1430 418
rect 649 361 1430 384
rect 113 261 181 281
rect 113 227 129 261
rect 163 228 181 261
rect 285 228 569 283
rect 649 235 943 361
rect 1021 346 1430 361
rect 163 227 569 228
rect 113 190 569 227
rect 113 164 851 190
rect 113 54 851 80
rect 1661 314 1691 329
rect 1757 314 1787 329
rect 1661 284 1787 314
rect 1995 305 2025 329
rect 2091 305 2121 329
rect 1661 248 1691 284
rect 1602 236 1691 248
rect 1995 275 2121 305
rect 1995 265 2088 275
rect 1602 202 1641 236
rect 1675 214 1691 236
rect 1824 227 1890 238
rect 1675 202 1728 214
rect 1602 184 1728 202
rect 1602 155 1632 184
rect 1698 155 1728 184
rect 1824 193 1840 227
rect 1874 219 1890 227
rect 1995 231 2038 265
rect 2072 231 2088 265
rect 1995 219 2088 231
rect 1874 193 2033 219
rect 1824 189 2033 193
rect 1824 182 1937 189
rect 1907 155 1937 182
rect 2003 155 2033 189
rect 1021 32 1430 71
rect 1602 44 1632 71
rect 1698 44 1728 71
rect 1907 44 1937 71
rect 2003 44 2033 71
<< polycont >>
rect 1116 384 1150 418
rect 1184 384 1218 418
rect 1252 384 1286 418
rect 129 227 163 261
rect 1641 202 1675 236
rect 1840 193 1874 227
rect 2038 231 2072 265
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2145 561
rect 2179 527 2208 561
rect 1611 460 1645 527
rect 239 422 273 447
rect 238 388 239 400
rect 238 361 273 388
rect 581 419 615 447
rect 581 351 615 380
rect 581 289 615 308
rect 650 336 1016 460
rect 1095 418 1407 425
rect 1095 384 1116 418
rect 1171 384 1184 418
rect 1218 384 1235 418
rect 1286 384 1407 418
rect 1095 374 1407 384
rect 1611 392 1645 426
rect 1442 336 1476 351
rect 650 325 1476 336
rect 1611 325 1645 358
rect 1707 465 1741 491
rect 1707 416 1741 431
rect 1707 325 1741 363
rect 1803 459 1837 491
rect 1803 391 1837 425
rect 650 291 975 325
rect 1009 291 1442 325
rect 113 264 181 281
rect 21 261 181 264
rect 21 227 129 261
rect 163 227 181 261
rect 21 209 181 227
rect 21 198 75 209
rect 113 195 181 209
rect 650 257 1476 291
rect 650 223 975 257
rect 1009 223 1442 257
rect 1542 268 1576 279
rect 1542 235 1586 268
rect 650 196 1476 223
rect 973 189 1476 196
rect 67 126 101 143
rect 67 76 101 92
rect 863 135 897 160
rect 863 58 897 93
rect 973 155 975 189
rect 1009 155 1442 189
rect 973 121 1476 155
rect 973 87 975 121
rect 1009 87 1442 121
rect 973 17 1476 87
rect 1552 130 1586 235
rect 1620 202 1636 236
rect 1675 202 1691 236
rect 1803 228 1837 357
rect 1871 296 1905 527
rect 1939 454 1979 491
rect 1939 414 1945 454
rect 1939 383 1979 414
rect 2041 459 2075 491
rect 2041 391 2075 425
rect 2041 309 2075 348
rect 2137 459 2177 491
rect 2171 425 2177 459
rect 2137 419 2177 425
rect 2171 357 2177 419
rect 2137 325 2177 357
rect 1871 262 1987 296
rect 1803 227 1890 228
rect 1803 210 1840 227
rect 1744 193 1840 210
rect 1874 193 1890 227
rect 1744 176 1837 193
rect 1552 17 1586 96
rect 1648 141 1682 159
rect 1648 69 1682 97
rect 1744 131 1778 176
rect 1744 69 1778 97
rect 1857 133 1891 143
rect 1857 69 1891 87
rect 1953 131 1987 262
rect 2022 231 2038 265
rect 2072 231 2089 265
rect 2043 193 2089 231
rect 1953 69 1987 97
rect 2049 139 2083 159
rect 2049 69 2083 97
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2145 17
rect 2179 -17 2208 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 1685 527 1719 561
rect 1777 527 1811 561
rect 1869 527 1903 561
rect 1961 527 1995 561
rect 2053 527 2087 561
rect 2145 527 2179 561
rect 239 388 273 422
rect 581 385 615 414
rect 581 380 615 385
rect 581 317 615 342
rect 581 308 615 317
rect 1137 384 1150 418
rect 1150 384 1171 418
rect 1235 384 1252 418
rect 1252 384 1269 418
rect 1707 397 1741 416
rect 1707 382 1741 397
rect 1542 279 1576 313
rect 67 92 101 126
rect 863 101 897 127
rect 863 93 897 101
rect 1636 202 1641 236
rect 1641 202 1670 236
rect 1945 420 1979 448
rect 1945 414 1979 420
rect 2041 357 2075 382
rect 2041 348 2075 357
rect 2137 391 2171 419
rect 2137 385 2171 391
rect 1648 131 1682 141
rect 1648 107 1682 131
rect 1857 121 1891 133
rect 1857 99 1891 121
rect 2049 131 2083 139
rect 2049 105 2083 131
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
rect 1685 -17 1719 17
rect 1777 -17 1811 17
rect 1869 -17 1903 17
rect 1961 -17 1995 17
rect 2053 -17 2087 17
rect 2145 -17 2179 17
<< metal1 >>
rect 0 561 2208 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2145 561
rect 2179 527 2208 561
rect 0 496 2208 527
rect 233 422 279 496
rect 233 388 239 422
rect 273 388 279 422
rect 233 362 279 388
rect 573 414 1016 460
rect 1701 448 2177 458
rect 1701 430 1945 448
rect 573 380 581 414
rect 615 380 1016 414
rect 238 361 273 362
rect 573 342 1016 380
rect 1124 418 1282 424
rect 1124 384 1137 418
rect 1171 384 1235 418
rect 1269 384 1282 418
rect 1124 378 1282 384
rect 1701 416 1747 430
rect 1701 382 1707 416
rect 1741 382 1747 416
rect 1939 414 1945 430
rect 1979 430 2177 448
rect 1979 414 1985 430
rect 1939 400 1985 414
rect 2131 419 2177 430
rect 573 308 581 342
rect 615 336 1016 342
rect 1181 336 1226 378
rect 1701 342 1747 382
rect 2035 382 2081 402
rect 2035 348 2041 382
rect 2075 348 2081 382
rect 2131 385 2137 419
rect 2171 385 2177 419
rect 2131 349 2177 385
rect 615 308 1496 336
rect 573 223 1496 308
rect 1530 314 1582 320
rect 2035 314 2081 348
rect 1530 313 2081 314
rect 1530 279 1542 313
rect 1576 279 2081 313
rect 1530 275 2081 279
rect 1530 273 1582 275
rect 1601 236 1691 242
rect 1601 223 1636 236
rect 573 202 1636 223
rect 1670 202 1691 236
rect 573 196 1691 202
rect 955 184 1691 196
rect 955 142 1496 184
rect 61 126 107 140
rect 61 92 67 126
rect 101 92 107 126
rect 61 48 107 92
rect 856 127 1496 142
rect 856 93 863 127
rect 897 93 1496 127
rect 1642 141 1688 155
rect 1642 107 1648 141
rect 1682 121 1688 141
rect 2037 139 2095 147
rect 1845 133 1903 139
rect 1845 121 1857 133
rect 1682 107 1857 121
rect 1642 99 1857 107
rect 1891 121 1903 133
rect 2037 121 2049 139
rect 1891 105 2049 121
rect 2083 113 2095 139
rect 2083 105 2089 113
rect 1891 99 2089 105
rect 1642 93 2089 99
rect 856 78 940 93
rect 0 17 2208 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2145 17
rect 2179 -17 2208 17
rect 0 -48 2208 -17
<< labels >>
flabel metal1 s 0 496 2208 592 0 FreeSans 200 0 0 0 VPWR
port 1 nsew
flabel metal1 s 673 527 707 561 0 FreeSans 200 0 0 0 VPWR
port 1 nsew
flabel metal1 s 121 527 155 561 0 FreeSans 200 0 0 0 VPWR
port 1 nsew
flabel metal1 s 1409 527 1443 561 0 FreeSans 200 0 0 0 VPWR
port 1 nsew
flabel metal1 s 1869 527 1903 561 0 FreeSans 200 0 0 0 VPWR
port 1 nsew
flabel metal1 s 2053 527 2087 561 0 FreeSans 200 0 0 0 VPWR
port 1 nsew
flabel metal1 s 0 -48 2208 48 0 FreeSans 200 0 0 0 VGND
port 2 nsew
flabel metal1 s 673 -17 707 17 0 FreeSans 200 0 0 0 VGND
port 2 nsew
flabel metal1 s 121 -17 155 17 0 FreeSans 200 0 0 0 VGND
port 2 nsew
flabel metal1 s 1225 -17 1259 17 0 FreeSans 200 0 0 0 VGND
port 2 nsew
flabel metal1 s 1777 -17 1811 17 0 FreeSans 200 0 0 0 VGND
port 2 nsew
flabel metal1 s 1317 -17 1351 17 0 FreeSans 200 0 0 0 VGND
port 2 nsew
flabel metal1 s 949 -17 983 17 0 FreeSans 200 0 0 0 VGND
port 2 nsew
flabel locali s 40 221 74 255 7 FreeSans 200 0 0 0 in
port 3 nsew
flabel locali s 2049 207 2083 241 0 FreeSans 200 0 0 0 out
port 4 nsew
rlabel metal1 s 982 285 982 285 4 mid
port 5 nsew
flabel nwell s 673 527 707 561 0 FreeSans 200 0 0 0 VPB
port 6 nsew
flabel nwell s 121 527 155 561 0 FreeSans 200 0 0 0 VPB
port 6 nsew
flabel nwell s 1409 527 1443 561 0 FreeSans 200 0 0 0 VPB
port 6 nsew
flabel nwell s 1869 527 1903 561 0 FreeSans 200 0 0 0 VPB
port 6 nsew
flabel nwell s 2053 527 2087 561 0 FreeSans 200 0 0 0 VPB
port 6 nsew
flabel pwell s 673 -17 707 17 0 FreeSans 200 0 0 0 VNB
port 7 nsew
flabel pwell s 121 -17 155 17 0 FreeSans 200 0 0 0 VNB
port 7 nsew
flabel pwell s 1225 -17 1259 17 0 FreeSans 200 0 0 0 VNB
port 7 nsew
flabel pwell s 1777 -17 1811 17 0 FreeSans 200 0 0 0 VNB
port 7 nsew
flabel pwell s 1317 -17 1351 17 0 FreeSans 200 0 0 0 VNB
port 7 nsew
flabel pwell s 949 -17 983 17 0 FreeSans 200 0 0 0 VNB
port 7 nsew
<< properties >>
string FIXED_BBOX 0 0 2208 544
string GDS_END 179266
string GDS_FILE adc_top.gds.gz
string GDS_START 161944
<< end >>
