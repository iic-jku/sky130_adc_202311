magic
tech sky130A
magscale 1 2
timestamp 1695643842
<< error_s >>
rect -131 1381 -37 1441
rect 151 133 209 139
rect 343 133 401 139
rect 535 133 593 139
rect 727 133 785 139
rect 919 133 977 139
rect 1111 133 1169 139
rect 1303 133 1361 139
rect 1495 133 1553 139
rect 151 99 163 133
rect 343 99 355 133
rect 535 99 547 133
rect 727 99 739 133
rect 919 99 931 133
rect 1111 99 1123 133
rect 1303 99 1315 133
rect 1495 99 1507 133
rect 151 93 209 99
rect 343 93 401 99
rect 535 93 593 99
rect 727 93 785 99
rect 919 93 977 99
rect 1111 93 1169 99
rect 1303 93 1361 99
rect 1495 93 1553 99
<< locali >>
rect -61 171 115 1171
rect 1589 171 1765 1171
rect -61 99 99 133
rect 1605 99 1765 133
<< metal1 >>
rect 1453 1171 1499 1623
<< metal3 >>
rect -131 1381 -37 1427
use sky130_fd_pr__nfet_01v8_YN9FL4  sky130_fd_pr__nfet_01v8_UDPJLN_0
timestamp 1695643842
transform 1 0 852 0 1 671
box -983 -710 983 710
<< end >>
