magic
tech sky130A
magscale 1 2
timestamp 1698999411
<< nwell >>
rect 160 493 1192 814
<< pwell >>
rect 266 270 568 408
rect 784 270 1086 408
rect 204 184 1148 270
<< nmos >>
rect 354 298 384 382
rect 450 298 480 382
rect 872 298 902 382
rect 968 298 998 382
<< pmos >>
rect 258 530 288 690
rect 354 530 384 690
rect 450 530 480 690
rect 546 530 576 690
rect 776 530 806 690
rect 872 530 902 690
rect 968 530 998 690
rect 1064 530 1094 690
<< ndiff >>
rect 292 357 354 382
rect 292 323 304 357
rect 338 323 354 357
rect 292 298 354 323
rect 384 357 450 382
rect 384 323 400 357
rect 434 323 450 357
rect 384 298 450 323
rect 480 357 542 382
rect 480 323 496 357
rect 530 323 542 357
rect 480 298 542 323
rect 810 357 872 382
rect 810 323 822 357
rect 856 323 872 357
rect 810 298 872 323
rect 902 357 968 382
rect 902 323 918 357
rect 952 323 968 357
rect 902 298 968 323
rect 998 357 1060 382
rect 998 323 1014 357
rect 1048 323 1060 357
rect 998 298 1060 323
<< pdiff >>
rect 196 661 258 690
rect 196 627 208 661
rect 242 627 258 661
rect 196 593 258 627
rect 196 559 208 593
rect 242 559 258 593
rect 196 530 258 559
rect 288 661 354 690
rect 288 627 304 661
rect 338 627 354 661
rect 288 593 354 627
rect 288 559 304 593
rect 338 559 354 593
rect 288 530 354 559
rect 384 661 450 690
rect 384 627 400 661
rect 434 627 450 661
rect 384 593 450 627
rect 384 559 400 593
rect 434 559 450 593
rect 384 530 450 559
rect 480 661 546 690
rect 480 627 496 661
rect 530 627 546 661
rect 480 593 546 627
rect 480 559 496 593
rect 530 559 546 593
rect 480 530 546 559
rect 576 661 638 690
rect 576 627 592 661
rect 626 627 638 661
rect 576 593 638 627
rect 576 559 592 593
rect 626 559 638 593
rect 576 530 638 559
rect 714 661 776 690
rect 714 627 726 661
rect 760 627 776 661
rect 714 593 776 627
rect 714 559 726 593
rect 760 559 776 593
rect 714 530 776 559
rect 806 661 872 690
rect 806 627 822 661
rect 856 627 872 661
rect 806 593 872 627
rect 806 559 822 593
rect 856 559 872 593
rect 806 530 872 559
rect 902 661 968 690
rect 902 627 918 661
rect 952 627 968 661
rect 902 593 968 627
rect 902 559 918 593
rect 952 559 968 593
rect 902 530 968 559
rect 998 661 1064 690
rect 998 627 1014 661
rect 1048 627 1064 661
rect 998 593 1064 627
rect 998 559 1014 593
rect 1048 559 1064 593
rect 998 530 1064 559
rect 1094 661 1156 690
rect 1094 627 1110 661
rect 1144 627 1156 661
rect 1094 593 1156 627
rect 1094 559 1110 593
rect 1144 559 1156 593
rect 1094 530 1156 559
<< ndiffc >>
rect 304 323 338 357
rect 400 323 434 357
rect 496 323 530 357
rect 822 323 856 357
rect 918 323 952 357
rect 1014 323 1048 357
<< pdiffc >>
rect 208 627 242 661
rect 208 559 242 593
rect 304 627 338 661
rect 304 559 338 593
rect 400 627 434 661
rect 400 559 434 593
rect 496 627 530 661
rect 496 559 530 593
rect 592 627 626 661
rect 592 559 626 593
rect 726 627 760 661
rect 726 559 760 593
rect 822 627 856 661
rect 822 559 856 593
rect 918 627 952 661
rect 918 559 952 593
rect 1014 627 1048 661
rect 1014 559 1048 593
rect 1110 627 1144 661
rect 1110 559 1144 593
<< psubdiff >>
rect 230 210 264 244
rect 298 210 332 244
rect 366 210 400 244
rect 434 210 468 244
rect 502 210 536 244
rect 570 210 782 244
rect 816 210 850 244
rect 884 210 918 244
rect 952 210 986 244
rect 1020 210 1054 244
rect 1088 210 1122 244
<< nsubdiff >>
rect 208 744 264 778
rect 298 744 332 778
rect 366 744 400 778
rect 434 744 468 778
rect 502 744 536 778
rect 570 744 782 778
rect 816 744 850 778
rect 884 744 918 778
rect 952 744 986 778
rect 1020 744 1054 778
rect 1088 744 1144 778
<< psubdiffcont >>
rect 264 210 298 244
rect 332 210 366 244
rect 400 210 434 244
rect 468 210 502 244
rect 536 210 570 244
rect 782 210 816 244
rect 850 210 884 244
rect 918 210 952 244
rect 986 210 1020 244
rect 1054 210 1088 244
<< nsubdiffcont >>
rect 264 744 298 778
rect 332 744 366 778
rect 400 744 434 778
rect 468 744 502 778
rect 536 744 570 778
rect 782 744 816 778
rect 850 744 884 778
rect 918 744 952 778
rect 986 744 1020 778
rect 1054 744 1088 778
<< poly >>
rect 258 690 288 717
rect 354 690 384 716
rect 450 690 480 717
rect 546 690 576 716
rect 776 690 806 717
rect 872 690 902 716
rect 968 690 998 717
rect 1064 690 1094 716
rect 258 484 288 530
rect 354 490 384 530
rect 220 468 288 484
rect 220 434 238 468
rect 272 434 288 468
rect 220 424 288 434
rect 330 480 390 490
rect 450 484 480 530
rect 546 490 576 530
rect 330 446 346 480
rect 380 446 390 480
rect 330 430 390 446
rect 444 469 504 484
rect 444 435 454 469
rect 488 435 504 469
rect 354 382 384 430
rect 444 425 504 435
rect 546 480 614 490
rect 776 484 806 530
rect 872 490 902 530
rect 546 446 564 480
rect 598 446 614 480
rect 546 430 614 446
rect 738 468 806 484
rect 738 434 756 468
rect 790 434 806 468
rect 450 382 480 425
rect 738 424 806 434
rect 848 480 908 490
rect 968 484 998 530
rect 1064 490 1094 530
rect 848 446 864 480
rect 898 446 908 480
rect 848 430 908 446
rect 962 469 1022 484
rect 962 435 972 469
rect 1006 435 1022 469
rect 872 382 902 430
rect 962 425 1022 435
rect 1064 480 1132 490
rect 1064 446 1082 480
rect 1116 446 1132 480
rect 1064 430 1132 446
rect 968 382 998 425
rect 354 272 384 298
rect 450 272 480 298
rect 872 272 902 298
rect 968 272 998 298
<< polycont >>
rect 238 434 272 468
rect 346 446 380 480
rect 454 435 488 469
rect 564 446 598 480
rect 756 434 790 468
rect 864 446 898 480
rect 972 435 1006 469
rect 1082 446 1116 480
<< locali >>
rect 208 744 264 778
rect 298 744 332 778
rect 366 744 400 778
rect 434 744 468 778
rect 502 744 536 778
rect 570 744 782 778
rect 816 744 850 778
rect 884 744 918 778
rect 952 744 986 778
rect 1020 744 1054 778
rect 1088 744 1144 778
rect 208 661 242 744
rect 208 593 242 627
rect 208 526 242 559
rect 304 661 338 694
rect 304 593 338 627
rect 304 526 338 559
rect 400 661 434 694
rect 400 593 434 594
rect 400 526 434 559
rect 496 661 530 694
rect 496 593 530 627
rect 496 526 530 559
rect 592 661 626 744
rect 592 593 626 627
rect 592 526 626 559
rect 726 661 760 744
rect 726 593 760 627
rect 726 526 760 559
rect 822 661 856 694
rect 822 593 856 627
rect 822 526 856 559
rect 918 661 952 694
rect 918 593 952 594
rect 918 526 952 559
rect 1014 661 1048 694
rect 1014 593 1048 627
rect 1014 526 1048 559
rect 1110 661 1144 744
rect 1110 593 1144 627
rect 1110 526 1144 559
rect 220 468 288 484
rect 220 434 238 468
rect 272 434 288 468
rect 220 424 288 434
rect 330 480 398 490
rect 330 446 346 480
rect 380 446 398 480
rect 330 430 398 446
rect 436 469 504 484
rect 436 434 454 469
rect 488 434 504 469
rect 436 425 504 434
rect 546 480 614 490
rect 546 446 564 480
rect 598 446 614 480
rect 546 430 614 446
rect 738 468 806 484
rect 738 434 756 468
rect 790 434 806 468
rect 738 424 806 434
rect 848 480 916 490
rect 848 446 864 480
rect 898 446 916 480
rect 848 430 916 446
rect 954 469 1022 484
rect 954 434 972 469
rect 1006 434 1022 469
rect 954 425 1022 434
rect 1064 480 1132 490
rect 1064 446 1082 480
rect 1116 446 1132 480
rect 1064 430 1132 446
rect 304 357 338 386
rect 304 244 338 323
rect 400 357 434 386
rect 400 294 434 302
rect 496 357 530 386
rect 496 244 530 323
rect 822 357 856 386
rect 822 244 856 323
rect 918 357 952 386
rect 918 294 952 302
rect 1014 357 1048 386
rect 1014 244 1048 323
rect 230 210 264 244
rect 298 210 332 244
rect 366 210 400 244
rect 434 210 468 244
rect 502 210 536 244
rect 570 210 782 244
rect 816 210 850 244
rect 884 210 918 244
rect 952 210 986 244
rect 1020 210 1054 244
rect 1088 210 1122 244
<< viali >>
rect 400 627 434 628
rect 400 594 434 627
rect 918 627 952 628
rect 918 594 952 627
rect 238 434 272 468
rect 346 446 380 480
rect 454 435 488 468
rect 454 434 488 435
rect 564 446 598 480
rect 756 434 790 468
rect 864 446 898 480
rect 972 435 1006 468
rect 972 434 1006 435
rect 1082 446 1116 480
rect 400 323 434 336
rect 400 302 434 323
rect 918 323 952 336
rect 918 302 952 323
<< metal1 >>
rect 391 637 443 643
rect 391 579 443 585
rect 909 637 961 643
rect 909 579 961 585
rect 190 508 644 536
rect 708 508 1162 536
rect 336 480 388 508
rect 554 486 618 508
rect 229 468 281 480
rect 229 434 238 468
rect 272 434 281 468
rect 336 446 346 480
rect 380 446 388 480
rect 336 434 388 446
rect 444 468 504 480
rect 444 434 454 468
rect 488 434 504 468
rect 554 434 560 486
rect 612 434 618 486
rect 854 480 906 508
rect 1072 486 1136 508
rect 747 468 799 480
rect 747 434 756 468
rect 790 434 799 468
rect 854 446 864 480
rect 898 446 906 480
rect 854 434 906 446
rect 962 468 1022 480
rect 962 434 972 468
rect 1006 434 1022 468
rect 1072 434 1078 486
rect 1130 434 1136 486
rect 229 405 281 434
rect 444 405 504 434
rect 747 406 799 434
rect 190 377 627 405
rect 391 338 443 348
rect 391 277 443 286
rect 596 305 627 377
rect 655 354 661 406
rect 713 405 799 406
rect 962 405 1022 434
rect 713 377 1162 405
rect 713 354 719 377
rect 909 338 961 348
rect 655 305 661 324
rect 596 277 661 305
rect 655 272 661 277
rect 713 305 719 324
rect 713 277 795 305
rect 909 277 961 286
rect 713 272 719 277
<< via1 >>
rect 391 628 443 637
rect 391 594 400 628
rect 400 594 434 628
rect 434 594 443 628
rect 391 585 443 594
rect 909 628 961 637
rect 909 594 918 628
rect 918 594 952 628
rect 952 594 961 628
rect 909 585 961 594
rect 560 480 612 486
rect 560 446 564 480
rect 564 446 598 480
rect 598 446 612 480
rect 560 434 612 446
rect 1078 480 1130 486
rect 1078 446 1082 480
rect 1082 446 1116 480
rect 1116 446 1130 480
rect 1078 434 1130 446
rect 391 336 443 338
rect 391 302 400 336
rect 400 302 434 336
rect 434 302 443 336
rect 391 286 443 302
rect 661 354 713 406
rect 909 336 961 338
rect 661 272 713 324
rect 909 302 918 336
rect 918 302 952 336
rect 952 302 961 336
rect 909 286 961 302
<< metal2 >>
rect 389 637 445 648
rect 389 585 391 637
rect 443 585 445 637
rect 389 574 445 585
rect 391 338 443 574
rect 618 499 682 638
rect 907 637 963 648
rect 907 585 909 637
rect 961 585 963 637
rect 907 574 963 585
rect 1136 630 1200 639
rect 1136 574 1140 630
rect 1196 574 1200 630
rect 618 486 622 499
rect 554 434 560 486
rect 612 443 622 486
rect 678 443 682 499
rect 612 434 682 443
rect 655 405 661 406
rect 190 286 391 305
rect 596 377 661 405
rect 596 305 627 377
rect 655 354 661 377
rect 713 354 719 406
rect 909 338 961 574
rect 1136 486 1200 574
rect 1072 434 1078 486
rect 1130 434 1200 486
rect 443 286 627 305
rect 190 277 627 286
rect 655 272 661 324
rect 713 305 719 324
rect 713 286 909 305
rect 961 286 1162 305
rect 713 277 1162 286
rect 713 272 719 277
<< via2 >>
rect 1140 574 1196 630
rect 622 443 678 499
<< metal3 >>
rect 618 629 684 642
rect 1134 630 1202 642
rect 1134 629 1140 630
rect 190 574 1140 629
rect 1196 574 1202 630
rect 190 569 1202 574
rect 616 499 684 507
rect 616 494 622 499
rect 190 443 622 494
rect 678 494 684 499
rect 1132 494 1202 507
rect 678 443 1202 494
rect 190 434 1202 443
<< labels >>
flabel metal1 s 1086 377 1162 405 0 FreeSans 200 0 0 0 qn
port 1 nsew
flabel metal1 s 190 377 229 405 0 FreeSans 200 0 0 0 q
port 2 nsew
flabel locali s 208 744 1144 778 0 FreeSans 200 0 0 0 VDD
port 3 nsew
flabel locali s 230 210 1122 244 0 FreeSans 200 0 0 0 VSS
port 4 nsew
flabel metal3 s 190 434 1200 494 0 FreeSans 200 0 0 0 s
port 5 nsew
flabel metal3 s 190 569 1200 629 0 FreeSans 200 0 0 0 r
port 6 nsew
flabel metal2 s 1086 277 1162 305 0 FreeSans 200 0 0 0 q
port 2 nsew
flabel metal2 s 190 277 229 305 0 FreeSans 200 0 0 0 qn
port 1 nsew
<< end >>
