magic
tech sky130A
magscale 1 2
timestamp 1697443344
<< pwell >>
rect 2811 7100 3433 7720
<< nmos >>
rect 3011 7310 3041 7510
rect 3107 7310 3137 7510
rect 3203 7310 3233 7510
<< ndiff >>
rect 2949 7498 3011 7510
rect 2949 7322 2961 7498
rect 2995 7322 3011 7498
rect 2949 7310 3011 7322
rect 3041 7498 3107 7510
rect 3041 7322 3057 7498
rect 3091 7322 3107 7498
rect 3041 7310 3107 7322
rect 3137 7498 3203 7510
rect 3137 7322 3153 7498
rect 3187 7322 3203 7498
rect 3137 7310 3203 7322
rect 3233 7498 3295 7510
rect 3233 7322 3249 7498
rect 3283 7322 3295 7498
rect 3233 7310 3295 7322
<< ndiffc >>
rect 2961 7322 2995 7498
rect 3057 7322 3091 7498
rect 3153 7322 3187 7498
rect 3249 7322 3283 7498
<< psubdiff >>
rect 2847 7650 2943 7684
rect 3301 7650 3397 7684
rect 2847 7588 2881 7650
rect 3363 7588 3397 7650
rect 2847 7170 2881 7232
rect 3363 7170 3397 7232
rect 2847 7136 2943 7170
rect 3301 7136 3397 7170
<< psubdiffcont >>
rect 2943 7650 3301 7684
rect 2847 7232 2881 7588
rect 3363 7232 3397 7588
rect 2943 7136 3301 7170
<< poly >>
rect 2975 7582 3041 7598
rect 2975 7548 2991 7582
rect 3025 7548 3041 7582
rect 2975 7532 3041 7548
rect 3203 7582 3269 7598
rect 3203 7548 3219 7582
rect 3253 7548 3269 7582
rect 3011 7510 3041 7532
rect 3107 7510 3137 7536
rect 3203 7532 3269 7548
rect 3203 7510 3233 7532
rect 3011 7284 3041 7310
rect 3107 7288 3137 7310
rect 3089 7272 3155 7288
rect 3203 7284 3233 7310
rect 3089 7238 3105 7272
rect 3139 7238 3155 7272
rect 3089 7222 3155 7238
<< polycont >>
rect 2991 7548 3025 7582
rect 3219 7548 3253 7582
rect 3105 7238 3139 7272
<< locali >>
rect 2081 11918 2881 11938
rect 2081 -1528 2101 11918
rect 2541 11728 2881 11918
rect 3363 11918 4163 11938
rect 2975 11766 3041 11868
rect 3203 11766 3269 11868
rect 3363 11728 3703 11918
rect 2541 11528 3057 11728
rect 3283 11528 3703 11728
rect 2541 10706 2881 11528
rect 2961 11527 3057 11528
rect 2975 10744 3041 10846
rect 3203 10744 3269 10846
rect 3363 10706 3703 11528
rect 2541 10506 3057 10706
rect 3283 10506 3703 10706
rect 2541 9684 2881 10506
rect 2961 10505 3057 10506
rect 2975 9722 3041 9824
rect 3203 9722 3269 9824
rect 3363 9684 3703 10506
rect 2541 9484 3057 9684
rect 3283 9484 3703 9684
rect 2541 8532 2881 9484
rect 2961 9483 3057 9484
rect 2975 8570 3041 8672
rect 3203 8570 3269 8672
rect 3363 8532 3703 9484
rect 2541 8332 3057 8532
rect 3283 8332 3703 8532
rect 2541 7684 2881 8332
rect 2961 8331 3057 8332
rect 3363 7684 3703 8332
rect 2541 7650 2943 7684
rect 3301 7650 3703 7684
rect 2541 7588 2881 7650
rect 2541 7232 2847 7588
rect 2975 7582 3041 7650
rect 2975 7548 2991 7582
rect 3025 7548 3041 7582
rect 3203 7582 3269 7650
rect 3203 7548 3219 7582
rect 3253 7548 3269 7582
rect 3363 7588 3703 7650
rect 2961 7510 2995 7514
rect 3057 7510 3091 7514
rect 2881 7498 3091 7510
rect 2881 7322 2961 7498
rect 2995 7322 3057 7498
rect 2881 7310 3091 7322
rect 2961 7309 3091 7310
rect 2961 7306 2995 7309
rect 3057 7306 3091 7309
rect 3153 7498 3187 7514
rect 3153 7306 3187 7322
rect 3249 7510 3283 7514
rect 3249 7498 3363 7510
rect 3283 7322 3363 7498
rect 3249 7310 3363 7322
rect 3249 7306 3283 7310
rect 3089 7238 3105 7272
rect 3139 7238 3155 7272
rect 2541 7170 2881 7232
rect 3397 7232 3703 7588
rect 3363 7170 3703 7232
rect 2541 7136 2943 7170
rect 3301 7136 3703 7170
rect 2541 6358 2881 7136
rect 2975 6396 3041 6498
rect 3203 6396 3269 6498
rect 3363 6358 3703 7136
rect 2541 6158 3057 6358
rect 3283 6158 3703 6358
rect 2541 4314 2881 6158
rect 2961 6157 3057 6158
rect 2975 4352 3041 4454
rect 3203 4352 3269 4454
rect 3363 4314 3703 6158
rect 2541 4114 3057 4314
rect 3283 4114 3703 4314
rect 2541 2140 2881 4114
rect 2961 4113 3057 4114
rect 2975 2178 3041 2280
rect 3203 2178 3269 2280
rect 3363 2140 3703 4114
rect 2541 1940 3057 2140
rect 3283 1940 3703 2140
rect 2541 96 2881 1940
rect 2961 1939 3057 1940
rect 2975 134 3041 236
rect 3203 134 3269 236
rect 3363 96 3703 1940
rect 2541 -104 3057 96
rect 3283 -104 3703 96
rect 2541 -1528 2881 -104
rect 2961 -105 3057 -104
rect 2081 -1548 2881 -1528
rect 3363 -1528 3703 -104
rect 4143 -1528 4163 11918
rect 3363 -1548 4163 -1528
<< viali >>
rect 2101 -1528 2541 11918
rect 2961 7322 2995 7498
rect 3057 7322 3091 7498
rect 3153 7322 3187 7498
rect 3249 7322 3283 7498
rect 3105 7238 3139 7272
rect 3703 -1528 4143 11918
<< metal1 >>
rect 2081 11918 2561 11938
rect 2081 -1528 2101 11918
rect 2541 -1528 2561 11918
rect 3683 11918 4163 11938
rect 3131 11716 3209 11722
rect 3131 11540 3137 11716
rect 3203 11540 3209 11716
rect 3131 11534 3209 11540
rect 2811 11450 3155 11496
rect 3131 10694 3209 10700
rect 3131 10518 3137 10694
rect 3203 10518 3209 10694
rect 3131 10512 3209 10518
rect 2811 10428 3155 10474
rect 3131 9672 3209 9678
rect 3131 9496 3137 9672
rect 3203 9496 3209 9672
rect 3131 9490 3209 9496
rect 2811 9406 3155 9452
rect 3131 8520 3209 8526
rect 3131 8344 3137 8520
rect 3203 8344 3209 8520
rect 3131 8338 3209 8344
rect 2811 8254 3155 8300
rect 2955 7498 3001 7510
rect 2955 7322 2961 7498
rect 2995 7322 3001 7498
rect 2955 7310 3001 7322
rect 3051 7498 3097 7510
rect 3147 7504 3193 7510
rect 3051 7322 3057 7498
rect 3091 7322 3097 7498
rect 3051 7310 3097 7322
rect 3131 7498 3209 7504
rect 3131 7322 3137 7498
rect 3203 7322 3209 7498
rect 3131 7316 3209 7322
rect 3243 7498 3289 7510
rect 3243 7322 3249 7498
rect 3283 7322 3289 7498
rect 3147 7310 3193 7316
rect 3243 7310 3289 7322
rect 2811 7272 3155 7278
rect 2811 7238 3105 7272
rect 3139 7238 3155 7272
rect 2811 7232 3155 7238
rect 3131 6346 3209 6352
rect 3131 6170 3137 6346
rect 3203 6170 3209 6346
rect 3131 6164 3209 6170
rect 2811 6080 3155 6126
rect 3131 4302 3209 4308
rect 3131 4126 3137 4302
rect 3203 4126 3209 4302
rect 3131 4120 3209 4126
rect 2811 4036 3155 4082
rect 3131 2128 3209 2134
rect 3131 1952 3137 2128
rect 3203 1952 3209 2128
rect 3131 1946 3209 1952
rect 2811 1862 3155 1908
rect 3131 84 3209 90
rect 3131 -92 3137 84
rect 3203 -92 3209 84
rect 3131 -98 3209 -92
rect 2811 -182 3155 -136
rect 2081 -1548 2561 -1528
rect 3683 -1528 3703 11918
rect 4143 -1528 4163 11918
rect 3683 -1548 4163 -1528
<< via1 >>
rect 2101 -1528 2541 11918
rect 3137 11540 3203 11716
rect 3137 10518 3203 10694
rect 3137 9496 3203 9672
rect 3137 8344 3203 8520
rect 3137 7322 3153 7498
rect 3153 7322 3187 7498
rect 3187 7322 3203 7498
rect 3137 6170 3203 6346
rect 3137 4126 3203 4302
rect 3137 1952 3203 2128
rect 3137 -92 3203 84
rect 3703 -1528 4143 11918
<< metal2 >>
rect 2081 11918 2561 11938
rect 2081 -1528 2101 11918
rect 2541 -1528 2561 11918
rect 3683 11918 4163 11938
rect 2811 11716 3433 11728
rect 2811 11708 3137 11716
rect 3203 11708 3433 11716
rect 2811 11548 2831 11708
rect 3413 11548 3433 11708
rect 2811 11540 3137 11548
rect 3203 11540 3433 11548
rect 2811 11528 3433 11540
rect 2811 10694 3433 10706
rect 2811 10686 3137 10694
rect 3203 10686 3433 10694
rect 2811 10526 2831 10686
rect 3413 10526 3433 10686
rect 2811 10518 3137 10526
rect 3203 10518 3433 10526
rect 2811 10506 3433 10518
rect 2811 9672 3433 9684
rect 2811 9664 3137 9672
rect 3203 9664 3433 9672
rect 2811 9504 2831 9664
rect 3413 9504 3433 9664
rect 2811 9496 3137 9504
rect 3203 9496 3433 9504
rect 2811 9484 3433 9496
rect 2811 8520 3433 8532
rect 2811 8512 3137 8520
rect 3203 8512 3433 8520
rect 2811 8352 2831 8512
rect 3413 8352 3433 8512
rect 2811 8344 3137 8352
rect 3203 8344 3433 8352
rect 2811 8332 3433 8344
rect 2811 7498 3433 7510
rect 2811 7490 3137 7498
rect 3203 7490 3433 7498
rect 2811 7330 2831 7490
rect 3413 7330 3433 7490
rect 2811 7322 3137 7330
rect 3203 7322 3433 7330
rect 2811 7310 3433 7322
rect 2811 6346 3433 6358
rect 2811 6338 3137 6346
rect 3203 6338 3433 6346
rect 2811 6178 2831 6338
rect 3413 6178 3433 6338
rect 2811 6170 3137 6178
rect 3203 6170 3433 6178
rect 2811 6158 3433 6170
rect 2811 4302 3433 4314
rect 2811 4294 3137 4302
rect 3203 4294 3433 4302
rect 2811 4134 2831 4294
rect 3413 4134 3433 4294
rect 2811 4126 3137 4134
rect 3203 4126 3433 4134
rect 2811 4114 3433 4126
rect 2811 2128 3433 2140
rect 2811 2120 3137 2128
rect 3203 2120 3433 2128
rect 2811 1960 2831 2120
rect 3413 1960 3433 2120
rect 2811 1952 3137 1960
rect 3203 1952 3433 1960
rect 2811 1940 3433 1952
rect 2811 84 3433 96
rect 2811 76 3137 84
rect 3203 76 3433 84
rect 2811 -84 2831 76
rect 3413 -84 3433 76
rect 2811 -92 3137 -84
rect 3203 -92 3433 -84
rect 2811 -104 3433 -92
rect 2081 -1548 2561 -1528
rect 3683 -1528 3703 11918
rect 4143 -1528 4163 11918
rect 3683 -1548 4163 -1528
<< via2 >>
rect 2831 11548 3137 11708
rect 3137 11548 3203 11708
rect 3203 11548 3413 11708
rect 2831 10526 3137 10686
rect 3137 10526 3203 10686
rect 3203 10526 3413 10686
rect 2831 9504 3137 9664
rect 3137 9504 3203 9664
rect 3203 9504 3413 9664
rect 2831 8352 3137 8512
rect 3137 8352 3203 8512
rect 3203 8352 3413 8512
rect 2831 7330 3137 7490
rect 3137 7330 3203 7490
rect 3203 7330 3413 7490
rect 2831 6178 3137 6338
rect 3137 6178 3203 6338
rect 3203 6178 3413 6338
rect 2831 4134 3137 4294
rect 3137 4134 3203 4294
rect 3203 4134 3413 4294
rect 2831 1960 3137 2120
rect 3137 1960 3203 2120
rect 3203 1960 3413 2120
rect 2831 -84 3137 76
rect 3137 -84 3203 76
rect 3203 -84 3413 76
<< metal3 >>
rect 2811 11708 3433 11728
rect 2811 11548 2831 11708
rect 3413 11548 3433 11708
rect 2811 11528 3433 11548
rect 2811 10686 3433 10706
rect 2811 10526 2831 10686
rect 3413 10526 3433 10686
rect 2811 10506 3433 10526
rect 2811 9664 3433 9684
rect 2811 9504 2831 9664
rect 3413 9504 3433 9664
rect 2811 9484 3433 9504
rect 2811 8512 3433 8532
rect 2811 8352 2831 8512
rect 3413 8352 3433 8512
rect 2811 8332 3433 8352
rect 2811 7490 3433 7510
rect 2811 7330 2831 7490
rect 3413 7330 3433 7490
rect 2811 7310 3433 7330
rect 2811 6338 3433 6358
rect 2811 6178 2831 6338
rect 3413 6178 3433 6338
rect 2811 6158 3433 6178
rect 2811 4294 3433 4314
rect 2811 4134 2831 4294
rect 3413 4134 3433 4294
rect 2811 4114 3433 4134
rect 2811 2120 3433 2140
rect 2811 1960 2831 2120
rect 3413 1960 3433 2120
rect 2811 1940 3433 1960
rect 2811 76 3433 96
rect 2811 -84 2831 76
rect 3413 -84 3433 76
rect 2811 -104 3433 -84
<< via3 >>
rect 2831 11548 3413 11688
rect 2831 10526 3413 10666
rect 2831 9504 3413 9664
rect 2831 8352 3413 8512
rect 2831 7330 3413 7490
rect 2831 6178 3413 6338
rect 2831 4134 3413 4294
rect 2831 1960 3413 2120
rect 2831 -84 3413 76
<< metal4 >>
rect 2081 11688 4163 11938
rect 2081 11638 2831 11688
rect 2811 11548 2831 11638
rect 3413 11638 4163 11688
rect 3413 11548 3433 11638
rect 2811 11528 3433 11548
rect 2081 11376 4163 11406
rect 2081 11136 3713 11376
rect 4133 11136 4163 11376
rect 2081 11106 4163 11136
rect 2081 10739 4163 10916
rect 2081 10666 4160 10739
rect 2081 10616 2831 10666
rect 2811 10526 2831 10616
rect 3413 10616 4160 10666
rect 3413 10526 3433 10616
rect 2811 10506 3433 10526
rect 2081 10354 4163 10384
rect 2081 10114 3713 10354
rect 4133 10114 4163 10354
rect 2081 10084 4163 10114
rect 1351 9664 4893 9894
rect 1351 9594 2831 9664
rect 2811 9504 2831 9594
rect 3413 9594 4893 9664
rect 3413 9504 3433 9594
rect 2811 9484 3433 9504
rect 1351 9332 4893 9362
rect 1351 9092 3713 9332
rect 4133 9092 4893 9332
rect 1351 9062 4893 9092
rect 1351 8712 4893 8742
rect 1351 8512 2912 8712
rect 3332 8512 4893 8712
rect 1351 8442 2831 8512
rect 2811 8352 2831 8442
rect 3413 8442 4893 8512
rect 3413 8352 3433 8442
rect 2811 8332 3433 8352
rect 1351 7940 3713 8160
rect 4133 7940 4893 8160
rect 1351 7910 4893 7940
rect 1351 7690 4893 7720
rect 1351 7490 2912 7690
rect 3332 7490 4893 7690
rect 1351 7420 2831 7490
rect 2811 7330 2831 7420
rect 3413 7420 4893 7490
rect 3413 7330 3433 7420
rect 2811 7310 3433 7330
rect 1351 7158 4893 7188
rect 1351 6918 3713 7158
rect 4133 6918 4893 7158
rect 1351 6888 4893 6918
rect 1351 6538 4893 6568
rect 1351 6338 2912 6538
rect 3332 6338 4893 6538
rect 1351 6268 2831 6338
rect 2811 6178 2831 6268
rect 3413 6268 4893 6338
rect 3413 6178 3433 6268
rect 2811 6158 3433 6178
rect 1351 6006 4893 6036
rect 1351 5766 3713 6006
rect 4133 5766 4893 6006
rect 1351 5736 4893 5766
rect 1351 5516 4893 5546
rect 1351 5276 2912 5516
rect 3332 5276 4893 5516
rect 1351 5246 4893 5276
rect 1351 4984 4893 5014
rect 1351 4744 3713 4984
rect 4133 4744 4893 4984
rect 1351 4714 4893 4744
rect 1351 4494 4893 4524
rect 1351 4294 2912 4494
rect 3332 4294 4893 4494
rect 1351 4224 2831 4294
rect 2811 4134 2831 4224
rect 3413 4224 4893 4294
rect 3413 4134 3433 4224
rect 2811 4114 3433 4134
rect 1351 3962 4893 3992
rect 1351 3722 3713 3962
rect 4133 3722 4893 3962
rect 1351 3692 4893 3722
rect 1351 3472 4893 3502
rect 1351 3232 2912 3472
rect 3332 3232 4893 3472
rect 1351 3202 4893 3232
rect 1351 2940 4893 2970
rect 1351 2700 3713 2940
rect 4133 2700 4893 2940
rect 1351 2670 4893 2700
rect 1351 2320 4893 2350
rect 1351 2120 2912 2320
rect 3332 2120 4893 2320
rect 1351 2050 2831 2120
rect 2811 1960 2831 2050
rect 3413 2050 4893 2120
rect 3413 1960 3433 2050
rect 2811 1940 3433 1960
rect 1351 1788 4893 1818
rect 1351 1548 3713 1788
rect 4133 1548 4893 1788
rect 1351 1518 4893 1548
rect 1351 1298 4893 1328
rect 1351 1058 2912 1298
rect 3332 1058 4893 1298
rect 1351 1028 4893 1058
rect 1351 766 4893 796
rect 1351 526 3713 766
rect 4133 526 4893 766
rect 1351 496 4893 526
rect 1351 276 4893 306
rect 1351 76 2912 276
rect 3332 76 4893 276
rect 1351 6 2831 76
rect 2811 -84 2831 6
rect 3413 6 4893 76
rect 3413 -84 3433 6
rect 2811 -104 3433 -84
rect 1351 -256 4893 -226
rect 1351 -496 3713 -256
rect 4133 -496 4893 -256
rect 1351 -526 4893 -496
rect 1351 -746 4893 -716
rect 1351 -986 2912 -746
rect 3332 -986 4893 -746
rect 1351 -1016 4893 -986
rect 1351 -1278 4893 -1248
rect 1351 -1518 3713 -1278
rect 4133 -1518 4893 -1278
rect 1351 -1548 4893 -1518
<< via4 >>
rect 3713 11136 4133 11376
rect 3713 10114 4133 10354
rect 3713 9092 4133 9332
rect 2912 8512 3332 8712
rect 2912 8472 3332 8512
rect 3713 7940 4133 8180
rect 2912 7490 3332 7690
rect 2912 7450 3332 7490
rect 3713 6918 4133 7158
rect 2912 6338 3332 6538
rect 2912 6298 3332 6338
rect 3713 5766 4133 6006
rect 2912 5276 3332 5516
rect 3713 4744 4133 4984
rect 2912 4294 3332 4494
rect 2912 4254 3332 4294
rect 3713 3722 4133 3962
rect 2912 3232 3332 3472
rect 3713 2700 4133 2940
rect 2912 2120 3332 2320
rect 2912 2080 3332 2120
rect 3713 1548 4133 1788
rect 2912 1058 3332 1298
rect 3713 526 4133 766
rect 2912 76 3332 276
rect 2912 36 3332 76
rect 3713 -496 4133 -256
rect 2912 -986 3332 -746
rect 3713 -1518 4133 -1278
<< metal5 >>
rect 2081 -1548 2561 11938
rect 2882 9062 3362 11938
rect 3683 11376 4163 11938
rect 3683 11136 3713 11376
rect 4133 11136 4163 11376
rect 3683 10354 4163 11136
rect 3683 10114 3713 10354
rect 4133 10114 4163 10354
rect 3683 9332 4163 10114
rect 3683 9092 3713 9332
rect 4133 9092 4163 9332
rect 2882 8712 3362 8742
rect 2882 8472 2912 8712
rect 3332 8472 3362 8712
rect 2882 7690 3362 8472
rect 2882 7450 2912 7690
rect 3332 7450 3362 7690
rect 2882 6888 3362 7450
rect 3683 8180 4163 9092
rect 3683 7940 3713 8180
rect 4133 7940 4163 8180
rect 3683 7158 4163 7940
rect 3683 6918 3713 7158
rect 4133 6918 4163 7158
rect 2882 6538 3362 6568
rect 2882 6298 2912 6538
rect 3332 6298 3362 6538
rect 2882 5516 3362 6298
rect 2882 5276 2912 5516
rect 3332 5276 3362 5516
rect 2882 4494 3362 5276
rect 2882 4254 2912 4494
rect 3332 4254 3362 4494
rect 2882 3472 3362 4254
rect 2882 3232 2912 3472
rect 3332 3232 3362 3472
rect 2882 2670 3362 3232
rect 3683 6006 4163 6918
rect 3683 5766 3713 6006
rect 4133 5766 4163 6006
rect 3683 4984 4163 5766
rect 3683 4744 3713 4984
rect 4133 4744 4163 4984
rect 3683 3962 4163 4744
rect 3683 3722 3713 3962
rect 4133 3722 4163 3962
rect 3683 2940 4163 3722
rect 3683 2700 3713 2940
rect 4133 2700 4163 2940
rect 2882 2320 3362 2350
rect 2882 2080 2912 2320
rect 3332 2080 3362 2320
rect 2882 1298 3362 2080
rect 2882 1058 2912 1298
rect 3332 1058 3362 1298
rect 2882 276 3362 1058
rect 2882 36 2912 276
rect 3332 36 3362 276
rect 2882 -746 3362 36
rect 2882 -986 2912 -746
rect 3332 -986 3362 -746
rect 2882 -1548 3362 -986
rect 3683 1788 4163 2700
rect 3683 1548 3713 1788
rect 4133 1548 4163 1788
rect 3683 766 4163 1548
rect 3683 526 3713 766
rect 4133 526 4163 766
rect 3683 -256 4163 526
rect 3683 -496 3713 -256
rect 4133 -496 4163 -256
rect 3683 -1278 4163 -496
rect 3683 -1518 3713 -1278
rect 4133 -1518 4163 -1278
rect 3683 -1548 4163 -1518
use sky130_fd_pr__cap_mim_m3_1_FJFAMD  sky130_fd_pr__cap_mim_m3_1_FJFAMD_0
timestamp 1696948209
transform 0 -1 3923 -1 0 3116
box -386 -240 386 240
use sky130_fd_pr__cap_mim_m3_1_FJFAMD  sky130_fd_pr__cap_mim_m3_1_FJFAMD_1
timestamp 1696948209
transform 0 1 2321 1 0 10530
box -386 -240 386 240
use sky130_fd_pr__cap_mim_m3_1_FJFAMD  sky130_fd_pr__cap_mim_m3_1_FJFAMD_2
timestamp 1696948209
transform 0 -1 4653 -1 0 7334
box -386 -240 386 240
use sky130_fd_pr__cap_mim_m3_1_FJFAMD  sky130_fd_pr__cap_mim_m3_1_FJFAMD_3
timestamp 1696948209
transform 0 1 2321 1 0 11552
box -386 -240 386 240
use sky130_fd_pr__cap_mim_m3_1_FJFAMD  sky130_fd_pr__cap_mim_m3_1_FJFAMD_4
timestamp 1696948209
transform 0 -1 3923 -1 0 11552
box -386 -240 386 240
use sky130_fd_pr__cap_mim_m3_1_FJFAMD  sky130_fd_pr__cap_mim_m3_1_FJFAMD_5
timestamp 1696948209
transform 0 -1 3923 -1 0 7334
box -386 -240 386 240
use sky130_fd_pr__cap_mim_m3_1_FJFAMD  sky130_fd_pr__cap_mim_m3_1_FJFAMD_6
timestamp 1696948209
transform 0 1 2321 1 0 7334
box -386 -240 386 240
use sky130_fd_pr__cap_mim_m3_1_FJFAMD  sky130_fd_pr__cap_mim_m3_1_FJFAMD_7
timestamp 1696948209
transform 0 -1 3923 -1 0 10530
box -386 -240 386 240
use sky130_fd_pr__cap_mim_m3_1_FJFAMD  sky130_fd_pr__cap_mim_m3_1_FJFAMD_8
timestamp 1696948209
transform 0 1 1591 -1 0 9508
box -386 -240 386 240
use sky130_fd_pr__cap_mim_m3_1_FJFAMD  sky130_fd_pr__cap_mim_m3_1_FJFAMD_9
timestamp 1696948209
transform 0 1 2321 1 0 9508
box -386 -240 386 240
use sky130_fd_pr__cap_mim_m3_1_FJFAMD  sky130_fd_pr__cap_mim_m3_1_FJFAMD_10
timestamp 1696948209
transform 0 -1 3923 -1 0 9508
box -386 -240 386 240
use sky130_fd_pr__cap_mim_m3_1_FJFAMD  sky130_fd_pr__cap_mim_m3_1_FJFAMD_11
timestamp 1696948209
transform 0 -1 4653 -1 0 9508
box -386 -240 386 240
use sky130_fd_pr__cap_mim_m3_1_FJFAMD  sky130_fd_pr__cap_mim_m3_1_FJFAMD_12
timestamp 1696948209
transform 0 1 1591 -1 0 7334
box -386 -240 386 240
use sky130_fd_pr__cap_mim_m3_1_FJFAMD  sky130_fd_pr__cap_mim_m3_1_FJFAMD_13
timestamp 1696948209
transform 0 1 2321 -1 0 3116
box -386 -240 386 240
use sky130_fd_pr__cap_mim_m3_1_FJFAMD  sky130_fd_pr__cap_mim_m3_1_FJFAMD_14
timestamp 1696948209
transform 0 1 1591 1 0 3116
box -386 -240 386 240
use sky130_fd_pr__cap_mim_m3_1_FJFAMD  sky130_fd_pr__cap_mim_m3_1_FJFAMD_15
timestamp 1696948209
transform 0 -1 3923 -1 0 4138
box -386 -240 386 240
use sky130_fd_pr__cap_mim_m3_1_FJFAMD  sky130_fd_pr__cap_mim_m3_1_FJFAMD_16
timestamp 1696948209
transform 0 1 1591 -1 0 8356
box -386 -240 386 240
use sky130_fd_pr__cap_mim_m3_1_FJFAMD  sky130_fd_pr__cap_mim_m3_1_FJFAMD_17
timestamp 1696948209
transform 0 1 2321 1 0 8356
box -386 -240 386 240
use sky130_fd_pr__cap_mim_m3_1_FJFAMD  sky130_fd_pr__cap_mim_m3_1_FJFAMD_18
timestamp 1696948209
transform 0 -1 3923 -1 0 8356
box -386 -240 386 240
use sky130_fd_pr__cap_mim_m3_1_FJFAMD  sky130_fd_pr__cap_mim_m3_1_FJFAMD_19
timestamp 1696948209
transform 0 -1 4653 -1 0 8356
box -386 -240 386 240
use sky130_fd_pr__cap_mim_m3_1_FJFAMD  sky130_fd_pr__cap_mim_m3_1_FJFAMD_20
timestamp 1696948209
transform 0 1 2321 1 0 4138
box -386 -240 386 240
use sky130_fd_pr__cap_mim_m3_1_FJFAMD  sky130_fd_pr__cap_mim_m3_1_FJFAMD_21
timestamp 1696948209
transform 0 1 1591 1 0 4138
box -386 -240 386 240
use sky130_fd_pr__cap_mim_m3_1_FJFAMD  sky130_fd_pr__cap_mim_m3_1_FJFAMD_22
timestamp 1696948209
transform 0 -1 4653 1 0 3116
box -386 -240 386 240
use sky130_fd_pr__cap_mim_m3_1_FJFAMD  sky130_fd_pr__cap_mim_m3_1_FJFAMD_23
timestamp 1696948209
transform 0 -1 4653 1 0 4138
box -386 -240 386 240
use sky130_fd_pr__cap_mim_m3_1_FJFAMD  sky130_fd_pr__cap_mim_m3_1_FJFAMD_24
timestamp 1696948209
transform 0 -1 4653 1 0 942
box -386 -240 386 240
use sky130_fd_pr__cap_mim_m3_1_FJFAMD  sky130_fd_pr__cap_mim_m3_1_FJFAMD_25
timestamp 1696948209
transform 0 1 1591 1 0 942
box -386 -240 386 240
use sky130_fd_pr__cap_mim_m3_1_FJFAMD  sky130_fd_pr__cap_mim_m3_1_FJFAMD_26
timestamp 1696948209
transform 0 1 2321 -1 0 942
box -386 -240 386 240
use sky130_fd_pr__cap_mim_m3_1_FJFAMD  sky130_fd_pr__cap_mim_m3_1_FJFAMD_27
timestamp 1696948209
transform 0 -1 3923 -1 0 942
box -386 -240 386 240
use sky130_fd_pr__cap_mim_m3_1_FJFAMD  sky130_fd_pr__cap_mim_m3_1_FJFAMD_28
timestamp 1696948209
transform 0 -1 3923 -1 0 -80
box -386 -240 386 240
use sky130_fd_pr__cap_mim_m3_1_FJFAMD  sky130_fd_pr__cap_mim_m3_1_FJFAMD_29
timestamp 1696948209
transform 0 1 2321 -1 0 -80
box -386 -240 386 240
use sky130_fd_pr__cap_mim_m3_1_FJFAMD  sky130_fd_pr__cap_mim_m3_1_FJFAMD_30
timestamp 1696948209
transform 0 1 1591 1 0 -80
box -386 -240 386 240
use sky130_fd_pr__cap_mim_m3_1_FJFAMD  sky130_fd_pr__cap_mim_m3_1_FJFAMD_31
timestamp 1696948209
transform 0 -1 4653 1 0 -80
box -386 -240 386 240
use sky130_fd_pr__cap_mim_m3_1_FJFAMD  sky130_fd_pr__cap_mim_m3_1_FJFAMD_32
timestamp 1696948209
transform 0 -1 3923 -1 0 -1102
box -386 -240 386 240
use sky130_fd_pr__cap_mim_m3_1_FJFAMD  sky130_fd_pr__cap_mim_m3_1_FJFAMD_33
timestamp 1696948209
transform 0 1 2321 -1 0 -1102
box -386 -240 386 240
use sky130_fd_pr__cap_mim_m3_1_FJFAMD  sky130_fd_pr__cap_mim_m3_1_FJFAMD_34
timestamp 1696948209
transform 0 1 1591 1 0 -1102
box -386 -240 386 240
use sky130_fd_pr__cap_mim_m3_1_FJFAMD  sky130_fd_pr__cap_mim_m3_1_FJFAMD_35
timestamp 1696948209
transform 0 -1 4653 1 0 -1102
box -386 -240 386 240
use sky130_fd_pr__cap_mim_m3_1_FJFAMD  sky130_fd_pr__cap_mim_m3_1_FJFAMD_36
timestamp 1696948209
transform 0 1 1591 -1 0 1964
box -386 -240 386 240
use sky130_fd_pr__cap_mim_m3_1_FJFAMD  sky130_fd_pr__cap_mim_m3_1_FJFAMD_37
timestamp 1696948209
transform 0 1 2321 -1 0 1964
box -386 -240 386 240
use sky130_fd_pr__cap_mim_m3_1_FJFAMD  sky130_fd_pr__cap_mim_m3_1_FJFAMD_38
timestamp 1696948209
transform 0 -1 3923 -1 0 1964
box -386 -240 386 240
use sky130_fd_pr__cap_mim_m3_1_FJFAMD  sky130_fd_pr__cap_mim_m3_1_FJFAMD_39
timestamp 1696948209
transform 0 -1 4653 1 0 1964
box -386 -240 386 240
use sky130_fd_pr__cap_mim_m3_1_FJFAMD  sky130_fd_pr__cap_mim_m3_1_FJFAMD_40
timestamp 1696948209
transform 0 1 2321 1 0 5160
box -386 -240 386 240
use sky130_fd_pr__cap_mim_m3_1_FJFAMD  sky130_fd_pr__cap_mim_m3_1_FJFAMD_41
timestamp 1696948209
transform 0 1 1591 1 0 5160
box -386 -240 386 240
use sky130_fd_pr__cap_mim_m3_1_FJFAMD  sky130_fd_pr__cap_mim_m3_1_FJFAMD_42
timestamp 1696948209
transform 0 -1 3923 -1 0 5160
box -386 -240 386 240
use sky130_fd_pr__cap_mim_m3_1_FJFAMD  sky130_fd_pr__cap_mim_m3_1_FJFAMD_43
timestamp 1696948209
transform 0 1 1591 1 0 6182
box -386 -240 386 240
use sky130_fd_pr__cap_mim_m3_1_FJFAMD  sky130_fd_pr__cap_mim_m3_1_FJFAMD_44
timestamp 1696948209
transform 0 1 2321 1 0 6182
box -386 -240 386 240
use sky130_fd_pr__cap_mim_m3_1_FJFAMD  sky130_fd_pr__cap_mim_m3_1_FJFAMD_45
timestamp 1696948209
transform 0 -1 3923 -1 0 6182
box -386 -240 386 240
use sky130_fd_pr__cap_mim_m3_1_FJFAMD  sky130_fd_pr__cap_mim_m3_1_FJFAMD_46
timestamp 1696948209
transform 0 -1 4653 1 0 6182
box -386 -240 386 240
use sky130_fd_pr__cap_mim_m3_1_FJFAMD  sky130_fd_pr__cap_mim_m3_1_FJFAMD_47
timestamp 1696948209
transform 0 -1 4653 1 0 5160
box -386 -240 386 240
use sky130_fd_pr__nfet_01v8_722GYZ  sky130_fd_pr__nfet_01v8_722GYZ_0
timestamp 1696948209
transform 1 0 3122 0 -1 4214
box -311 -310 311 310
use sky130_fd_pr__nfet_01v8_722GYZ  sky130_fd_pr__nfet_01v8_722GYZ_1
timestamp 1696948209
transform 1 0 3122 0 -1 10606
box -311 -310 311 310
use sky130_fd_pr__nfet_01v8_722GYZ  sky130_fd_pr__nfet_01v8_722GYZ_2
timestamp 1696948209
transform 1 0 3122 0 -1 11628
box -311 -310 311 310
use sky130_fd_pr__nfet_01v8_722GYZ  sky130_fd_pr__nfet_01v8_722GYZ_3
timestamp 1696948209
transform 1 0 3122 0 -1 9584
box -311 -310 311 310
use sky130_fd_pr__nfet_01v8_722GYZ  sky130_fd_pr__nfet_01v8_722GYZ_4
timestamp 1696948209
transform 1 0 3122 0 -1 8432
box -311 -310 311 310
use sky130_fd_pr__nfet_01v8_722GYZ  sky130_fd_pr__nfet_01v8_722GYZ_5
timestamp 1696948209
transform 1 0 3122 0 -1 -4
box -311 -310 311 310
use sky130_fd_pr__nfet_01v8_722GYZ  sky130_fd_pr__nfet_01v8_722GYZ_6
timestamp 1696948209
transform 1 0 3122 0 -1 2040
box -311 -310 311 310
use sky130_fd_pr__nfet_01v8_722GYZ  sky130_fd_pr__nfet_01v8_722GYZ_7
timestamp 1696948209
transform 1 0 3122 0 -1 6258
box -311 -310 311 310
<< end >>
