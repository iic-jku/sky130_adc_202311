magic
tech sky130A
magscale 1 2
timestamp 1696596751
<< locali >>
rect 3761 25870 4079 26006
rect 6749 25870 7067 26006
rect 3667 25082 4173 25832
rect 6655 25082 7161 25832
rect 11947 22090 17512 25910
rect 22428 25870 22746 26006
rect 25416 25870 25734 26006
rect 22334 25082 22840 25832
rect 25322 25082 25828 25832
rect 14559 21329 14763 22090
<< metal1 >>
rect 2828 27610 2876 27622
rect 26283 27610 26331 27631
rect 2826 27604 2878 27610
rect 2826 27498 2878 27504
rect 26281 27604 26333 27610
rect 26281 27498 26333 27504
rect 2828 26188 2876 27498
rect 5816 27410 5864 27413
rect 23631 27410 23679 27413
rect 5814 27404 5866 27410
rect 5814 27298 5866 27304
rect 23630 27404 23682 27410
rect 23630 27298 23682 27304
rect 5816 26233 5864 27298
rect 23631 26233 23679 27298
rect 26283 26188 26331 27498
<< via1 >>
rect 2826 27504 2878 27604
rect 26281 27504 26333 27604
rect 5814 27304 5866 27404
rect 23630 27304 23682 27404
<< metal2 >>
rect 2826 27604 2878 27610
rect 2799 27506 2826 27602
rect 26281 27604 26333 27610
rect 2878 27506 26281 27602
rect 2826 27498 2878 27504
rect 26333 27506 26430 27602
rect 26281 27498 26333 27504
rect 5814 27404 5866 27410
rect 5804 27306 5814 27402
rect 23630 27404 23682 27410
rect 5866 27306 23630 27402
rect 5814 27298 5866 27304
rect 23682 27306 23700 27402
rect 23630 27298 23682 27304
rect 2373 26744 12019 26804
rect 2373 26294 2433 26744
rect 7159 26294 12019 26744
rect 2373 26234 12019 26294
rect 17476 26745 27122 26804
rect 17476 26294 22335 26745
rect 27062 26294 27122 26745
rect 17476 26234 27122 26294
rect 12019 26090 18454 26186
rect 22334 26090 22412 26186
rect 25322 26090 25407 26186
rect 27122 26090 27207 26186
rect 2373 24476 12019 24536
rect 2373 24026 2433 24476
rect 10903 24026 12019 24476
rect 2373 23966 12019 24026
rect 17476 24476 27122 24536
rect 17476 24026 18592 24476
rect 26989 24026 27122 24476
rect 17476 23966 27122 24026
rect 2373 23752 11983 23812
rect 2373 23302 2433 23752
rect 7159 23302 11983 23752
rect 2373 23242 11983 23302
rect 17512 23752 27122 23812
rect 17512 23302 22335 23752
rect 27062 23302 27122 23752
rect 17512 23242 27122 23302
rect 2297 23098 2373 23194
rect 11530 23098 17512 23194
rect 27122 23098 27198 23194
rect 2373 21484 11288 21544
rect 2373 21034 2433 21484
rect 10867 21456 11288 21484
rect 17512 21484 27122 21544
rect 10867 21034 11983 21456
rect 2373 20974 11983 21034
rect 17512 21034 18628 21484
rect 27062 21034 27122 21484
rect 17512 20974 27122 21034
<< via2 >>
rect 2433 26294 7159 26744
rect 22335 26294 27062 26745
rect 2433 24026 10903 24476
rect 18592 24026 26989 24476
rect 2433 23302 7159 23752
rect 22335 23302 27062 23752
rect 2433 21034 10867 21484
rect 18628 21034 27062 21484
<< metal3 >>
rect 2373 26744 7219 26804
rect 2373 26294 2433 26744
rect 7159 26294 7219 26744
rect 2373 26234 7219 26294
rect 22275 26745 27122 26804
rect 22275 26294 22335 26745
rect 27062 26294 27122 26745
rect 22275 26234 27122 26294
rect 2373 24476 12019 24536
rect 2373 24026 2433 24476
rect 10903 24026 12019 24476
rect 2373 23966 12019 24026
rect 17476 24476 27122 24536
rect 17476 24026 18592 24476
rect 27062 24026 27122 24476
rect 17476 23966 27122 24026
rect 2373 23752 7219 23812
rect 2373 23302 2433 23752
rect 7159 23302 7219 23752
rect 2373 23242 7219 23302
rect 22275 23752 27122 23812
rect 22275 23302 22335 23752
rect 27062 23302 27122 23752
rect 22275 23242 27122 23302
rect 2373 21484 11288 21544
rect 2373 21034 2433 21484
rect 10867 21456 11288 21484
rect 17476 21484 27122 21544
rect 10867 21034 11983 21456
rect 2373 20974 11983 21034
rect 17476 21034 18628 21484
rect 27062 21034 27122 21484
rect 17476 20974 27122 21034
<< via3 >>
rect 2433 26294 7159 26744
rect 22335 26294 27062 26745
rect 2433 24026 10903 24476
rect 18592 24026 26989 24476
rect 26989 24026 27062 24476
rect 2433 23302 7159 23752
rect 22335 23302 27062 23752
rect 2433 21034 10867 21484
rect 18628 21034 27062 21484
<< metal4 >>
rect 1185 32446 28311 32506
rect 1185 31996 17535 32446
rect 18416 31996 22335 32446
rect 23215 31996 28311 32446
rect 1185 31936 28311 31996
rect 1185 31748 28311 31808
rect 1185 31298 6279 31748
rect 7159 31298 11079 31748
rect 11960 31298 28311 31748
rect 1185 31238 28311 31298
rect 8044 27468 21450 27528
rect 8044 27018 17534 27468
rect 18415 27018 21450 27468
rect 8044 26958 21450 27018
rect 2373 26744 7219 26804
rect 2373 26294 2433 26744
rect 7159 26294 7219 26744
rect 2373 26234 7219 26294
rect 22275 26745 27122 26804
rect 22275 26294 22335 26745
rect 27062 26294 27122 26745
rect 22275 26234 27122 26294
rect 8044 25846 21450 25906
rect 8044 25396 11079 25846
rect 11960 25396 21450 25846
rect 8044 25336 21450 25396
rect 2373 24476 12019 24536
rect 2373 24026 2433 24476
rect 10903 24026 12019 24476
rect 2373 23966 12019 24026
rect 17476 24476 27122 24536
rect 17476 24026 18592 24476
rect 27062 24026 27122 24476
rect 17476 23966 27122 24026
rect 2373 23752 7219 23812
rect 2373 23302 2433 23752
rect 7159 23302 7219 23752
rect 2373 23242 7219 23302
rect 22275 23752 27122 23812
rect 22275 23302 22335 23752
rect 27062 23302 27122 23752
rect 22275 23242 27122 23302
rect 2373 21484 12019 21544
rect 2373 21034 2433 21484
rect 10867 21034 12019 21484
rect 2373 20974 12019 21034
rect 17476 21484 27122 21544
rect 17476 21034 18628 21484
rect 27062 21034 27122 21484
rect 17476 20974 27122 21034
<< via4 >>
rect 17535 31996 18416 32446
rect 22335 31996 23215 32446
rect 6279 31298 7159 31748
rect 11079 31298 11960 31748
rect 17534 27018 18415 27468
rect 6279 26294 7159 26744
rect 22335 26294 23215 26744
rect 11079 25396 11960 25846
rect 6279 23302 7159 23752
rect 22335 23302 23215 23752
<< metal5 >>
rect 6219 31748 7219 32506
rect 6219 31298 6279 31748
rect 7159 31298 7219 31748
rect 6219 26744 7219 31298
rect 11019 31748 12019 35036
rect 11019 31298 11079 31748
rect 11960 31298 12019 31748
rect 11019 31238 12019 31298
rect 17475 32446 18475 35036
rect 17475 31996 17535 32446
rect 18416 31996 18475 32446
rect 17475 31238 18475 31996
rect 22275 32446 23275 32506
rect 22275 31996 22335 32446
rect 23215 31996 23275 32446
rect 6219 26294 6279 26744
rect 7159 26294 7219 26744
rect 6219 23752 7219 26294
rect 6219 23302 6279 23752
rect 7159 23302 7219 23752
rect 6219 23242 7219 23302
rect 11019 25846 12019 27661
rect 11019 25396 11079 25846
rect 11960 25396 12019 25846
rect 11019 -7940 12019 25396
rect 17475 27468 18475 27663
rect 17475 27018 17534 27468
rect 18415 27018 18475 27468
rect 17475 -7940 18475 27018
rect 22275 26744 23275 31996
rect 22275 26294 22335 26744
rect 23215 26294 23275 26744
rect 22275 23752 23275 26294
rect 22275 23302 22335 23752
rect 23215 23302 23275 23752
rect 22275 23242 23275 23302
use pa_nfet_w15_nf4  pa_nfet_w15_nf4_0
timestamp 1696585768
transform -1 0 26988 0 -1 26020
box -134 -318 1160 1588
use pa_nfet_w15_nf4  pa_nfet_w15_nf4_1
timestamp 1696585768
transform 1 0 2507 0 -1 26020
box -134 -318 1160 1588
use pa_nfet_w30_nf4  pa_nfet_w30_nf4_0
timestamp 1696592631
transform 1 0 4227 0 -1 26253
box -54 -85 2428 1821
use pa_nfet_w30_nf4  pa_nfet_w30_nf4_1
timestamp 1696592631
transform -1 0 25268 0 -1 26253
box -54 -85 2428 1821
use pa_nfet_w60_nf4  pa_nfet_w60_nf4_0
timestamp 1696592631
transform -1 0 22334 0 -1 26245
box 0 -93 4858 1813
use pa_nfet_w60_nf4  pa_nfet_w60_nf4_2
timestamp 1696592631
transform 1 0 7161 0 -1 26245
box 0 -93 4858 1813
use pa_nfet_w120_nf4  pa_nfet_w120_nf4_0
timestamp 1696592631
transform 1 0 17512 0 -1 23253
box 0 -93 9610 1813
use pa_nfet_w120_nf4  pa_nfet_w120_nf4_1
timestamp 1696592631
transform 1 0 2373 0 -1 23253
box 0 -93 9610 1813
use sky130_fd_pr__cap_mim_m3_1_H9ZJA7  sky130_fd_pr__cap_mim_m3_1_H9ZJA7_64
timestamp 1696250317
transform 0 1 18000 1 0 26432
box -686 -590 686 590
use sky130_fd_pr__cap_mim_m3_1_H9ZJA7  sky130_fd_pr__cap_mim_m3_1_H9ZJA7_65
timestamp 1696250317
transform 0 1 16570 -1 0 26432
box -686 -590 686 590
use sky130_fd_pr__cap_mim_m3_1_H9ZJA7  sky130_fd_pr__cap_mim_m3_1_H9ZJA7_70
timestamp 1696250317
transform 0 -1 11494 -1 0 26432
box -686 -590 686 590
use sky130_fd_pr__cap_mim_m3_1_H9ZJA7  sky130_fd_pr__cap_mim_m3_1_H9ZJA7_71
timestamp 1696250317
transform 0 1 12924 1 0 26432
box -686 -590 686 590
use sky130_fd_pr__nfet_01v8_SGMZ76  sky130_fd_pr__nfet_01v8_SGMZ76_0
timestamp 1696579262
transform 1 0 3920 0 -1 25457
box -359 -585 359 585
use sky130_fd_pr__nfet_01v8_SGMZ76  sky130_fd_pr__nfet_01v8_SGMZ76_1
timestamp 1696579262
transform 1 0 6908 0 -1 25457
box -359 -585 359 585
use sky130_fd_pr__nfet_01v8_SGMZ76  sky130_fd_pr__nfet_01v8_SGMZ76_2
timestamp 1696579262
transform -1 0 22587 0 -1 25457
box -359 -585 359 585
use sky130_fd_pr__nfet_01v8_SGMZ76  sky130_fd_pr__nfet_01v8_SGMZ76_3
timestamp 1696579262
transform -1 0 25575 0 -1 25457
box -359 -585 359 585
<< labels >>
flabel metal5 17475 32446 18475 35036 0 FreeSans 1600 0 0 0 inp_pa
port 1 nsew
flabel metal5 11019 31748 12019 35036 0 FreeSans 1600 0 0 0 inn_pa
port 2 nsew
flabel locali 14559 21329 14763 22090 0 FreeSans 1600 0 0 0 vss_pa
port 0 nsew
flabel metal2 27122 23098 27198 23194 0 FreeSans 320 0 0 0 en_pa[3]
port 3 nsew
flabel metal2 22334 26090 22412 26186 0 FreeSans 320 0 0 0 en_pa[2]
port 4 nsew
flabel metal2 25322 26090 25407 26186 0 FreeSans 320 0 0 0 en_pa[1]
port 5 nsew
flabel metal2 27122 26090 27207 26186 0 FreeSans 320 0 0 0 en_pa[0]
port 6 nsew
flabel metal5 17475 -7940 18475 -7176 0 FreeSans 1600 0 0 0 tunep_pa
port 7 nsew
flabel metal5 11019 -7940 12019 -7176 0 FreeSans 1600 0 0 0 tunen_pa
port 8 nsew
<< end >>
