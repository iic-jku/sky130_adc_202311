magic
tech sky130A
magscale 1 2
timestamp 1698999411
<< nwell >>
rect -38 261 682 582
<< pwell >>
rect 1 21 585 203
rect 30 -17 64 21
<< scnmos >>
rect 80 47 110 177
rect 179 47 209 177
rect 273 47 303 177
rect 369 47 399 177
rect 465 47 495 177
<< scpmoshvt >>
rect 80 297 110 497
rect 179 297 209 497
rect 273 297 303 497
rect 369 297 399 497
rect 465 297 495 497
<< ndiff >>
rect 27 162 80 177
rect 27 128 35 162
rect 69 128 80 162
rect 27 94 80 128
rect 27 60 35 94
rect 69 60 80 94
rect 27 47 80 60
rect 110 97 179 177
rect 110 63 135 97
rect 169 63 179 97
rect 110 47 179 63
rect 209 47 273 177
rect 303 47 369 177
rect 399 165 465 177
rect 399 131 411 165
rect 445 131 465 165
rect 399 97 465 131
rect 399 63 411 97
rect 445 63 465 97
rect 399 47 465 63
rect 495 97 559 177
rect 495 63 511 97
rect 545 63 559 97
rect 495 47 559 63
<< pdiff >>
rect 27 485 80 497
rect 27 451 35 485
rect 69 451 80 485
rect 27 417 80 451
rect 27 383 35 417
rect 69 383 80 417
rect 27 349 80 383
rect 27 315 35 349
rect 69 315 80 349
rect 27 297 80 315
rect 110 485 179 497
rect 110 451 127 485
rect 161 451 179 485
rect 110 417 179 451
rect 110 383 127 417
rect 161 383 179 417
rect 110 349 179 383
rect 110 315 127 349
rect 161 315 179 349
rect 110 297 179 315
rect 209 467 273 497
rect 209 433 223 467
rect 257 433 273 467
rect 209 399 273 433
rect 209 365 223 399
rect 257 365 273 399
rect 209 297 273 365
rect 303 467 369 497
rect 303 433 319 467
rect 353 433 369 467
rect 303 297 369 433
rect 399 467 465 497
rect 399 433 415 467
rect 449 433 465 467
rect 399 399 465 433
rect 399 365 415 399
rect 449 365 465 399
rect 399 297 465 365
rect 495 485 559 497
rect 495 451 517 485
rect 551 451 559 485
rect 495 399 559 451
rect 495 365 517 399
rect 551 365 559 399
rect 495 297 559 365
<< ndiffc >>
rect 35 128 69 162
rect 35 60 69 94
rect 135 63 169 97
rect 411 131 445 165
rect 411 63 445 97
rect 511 63 545 97
<< pdiffc >>
rect 35 451 69 485
rect 35 383 69 417
rect 35 315 69 349
rect 127 451 161 485
rect 127 383 161 417
rect 127 315 161 349
rect 223 433 257 467
rect 223 365 257 399
rect 319 433 353 467
rect 415 433 449 467
rect 415 365 449 399
rect 517 451 551 485
rect 517 365 551 399
<< poly >>
rect 80 497 110 523
rect 179 497 209 523
rect 273 497 303 523
rect 369 497 399 523
rect 465 497 495 523
rect 80 265 110 297
rect 179 265 209 297
rect 273 265 303 297
rect 369 265 399 297
rect 465 265 495 297
rect 80 249 135 265
rect 80 215 91 249
rect 125 215 135 249
rect 80 199 135 215
rect 177 249 231 265
rect 177 215 187 249
rect 221 215 231 249
rect 177 199 231 215
rect 273 249 327 265
rect 273 215 283 249
rect 317 215 327 249
rect 273 199 327 215
rect 369 249 423 265
rect 369 215 379 249
rect 413 215 423 249
rect 369 199 423 215
rect 465 249 519 265
rect 465 215 475 249
rect 509 215 519 249
rect 465 199 519 215
rect 80 177 110 199
rect 179 177 209 199
rect 273 177 303 199
rect 369 177 399 199
rect 465 177 495 199
rect 80 21 110 47
rect 179 21 209 47
rect 273 21 303 47
rect 369 21 399 47
rect 465 21 495 47
<< polycont >>
rect 91 215 125 249
rect 187 215 221 249
rect 283 215 317 249
rect 379 215 413 249
rect 475 215 509 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 644 561
rect 119 485 169 527
rect 19 451 35 485
rect 69 451 85 485
rect 19 417 85 451
rect 19 383 35 417
rect 69 383 85 417
rect 19 349 85 383
rect 19 315 35 349
rect 69 315 85 349
rect 119 451 127 485
rect 161 451 169 485
rect 119 417 169 451
rect 119 383 127 417
rect 161 383 169 417
rect 119 349 169 383
rect 207 467 257 483
rect 207 433 223 467
rect 303 467 369 527
rect 303 433 319 467
rect 353 433 369 467
rect 415 467 465 483
rect 449 433 465 467
rect 207 399 257 433
rect 415 399 465 433
rect 207 365 223 399
rect 257 365 415 399
rect 449 365 465 399
rect 501 451 517 485
rect 551 451 567 485
rect 501 399 567 451
rect 501 365 517 399
rect 551 365 592 399
rect 119 315 127 349
rect 161 315 169 349
rect 19 162 57 315
rect 119 299 169 315
rect 205 265 248 331
rect 91 249 153 265
rect 125 215 153 249
rect 91 199 153 215
rect 187 249 248 265
rect 221 215 248 249
rect 187 199 248 215
rect 283 249 340 331
rect 317 215 340 249
rect 283 199 340 215
rect 379 249 432 331
rect 413 215 432 249
rect 379 199 432 215
rect 475 249 524 331
rect 509 215 524 249
rect 475 199 524 215
rect 119 165 153 199
rect 558 165 592 365
rect 19 128 35 162
rect 69 128 85 162
rect 119 131 411 165
rect 445 131 592 165
rect 19 94 85 128
rect 395 97 461 131
rect 19 60 35 94
rect 69 60 85 94
rect 119 63 135 97
rect 169 63 185 97
rect 395 63 411 97
rect 445 63 461 97
rect 495 63 511 97
rect 545 63 561 97
rect 119 17 185 63
rect 495 17 561 63
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 644 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
<< metal1 >>
rect 0 561 644 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 644 561
rect 0 496 644 527
rect 0 17 644 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 644 17
rect 0 -48 644 -17
<< labels >>
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 1 nsew
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 2 nsew
flabel locali s 306 289 340 323 0 FreeSans 200 0 0 0 A2
port 5 nsew
flabel locali s 490 289 524 323 0 FreeSans 200 0 0 0 B1
port 7 nsew
flabel locali s 398 221 432 255 0 FreeSans 200 0 0 0 A1
port 6 nsew
flabel locali s 214 289 248 323 0 FreeSans 200 0 0 0 A3
port 4 nsew
flabel locali s 306 221 340 255 0 FreeSans 200 0 0 0 A2
port 5 nsew
flabel locali s 214 221 248 255 0 FreeSans 200 0 0 0 A3
port 4 nsew
flabel locali s 30 425 64 459 0 FreeSans 200 0 0 0 X
port 3 nsew
flabel locali s 398 289 432 323 0 FreeSans 200 0 0 0 A1
port 6 nsew
flabel locali s 30 357 64 391 0 FreeSans 200 0 0 0 X
port 3 nsew
flabel locali s 30 85 64 119 0 FreeSans 200 0 0 0 X
port 3 nsew
flabel locali s 490 221 524 255 0 FreeSans 200 0 0 0 B1
port 7 nsew
rlabel comment s 0 0 0 0 4 a31o_1
flabel nwell s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 9 nsew
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 10 nsew
<< properties >>
string FIXED_BBOX 0 0 644 544
string path 0.000 0.000 16.100 0.000 
<< end >>
