* Netlist for adc_top.mag
* Patrick Fath, IIC, JKU, 2023
* Netlist adapted for simulation, changes:
* -) Diodes removed
* -) Capmatrix replaced with PEX netlist of ADC capmatrix

.subckt sky130_fd_sc_hd__dfrtp_1 VGND VPWR CLK D RESET_B Q VPB VNB
X0 a_1217_47# a_27_47# a_1108_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X1 a_805_47# a_761_289# a_639_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.14 ps=1.1 w=0.42 l=0.15
X2 a_1108_47# a_193_47# a_761_289# VNB sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X3 a_1283_21# a_1108_47# a_1462_47# VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.064 ps=0.725 w=0.42 l=0.15
X4 a_651_413# a_27_47# a_543_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.116 pd=0.97 as=0.0724 ps=0.765 w=0.42 l=0.15
X5 VGND RESET_B a_805_47# VNB sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X6 Q a_1283_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.301 ps=2.66 w=1 l=0.15
X7 VPWR CLK a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X8 a_448_47# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.109 ps=1.36 w=0.42 l=0.15
X9 a_761_289# a_543_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.135 ps=1.15 w=0.64 l=0.15
X10 a_193_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X11 a_1108_47# a_27_47# a_761_289# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.129 ps=1.18 w=0.42 l=0.15
X12 a_543_47# a_27_47# a_448_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X13 a_1462_47# RESET_B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.064 pd=0.725 as=0.125 ps=1.01 w=0.42 l=0.15
X14 a_543_47# a_193_47# a_448_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0724 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X15 a_448_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.221 ps=1.89 w=0.42 l=0.15
X16 VPWR a_1283_21# a_1270_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X17 VPWR a_1108_47# a_1283_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X18 a_1270_413# a_193_47# a_1108_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X19 a_193_47# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X20 a_1283_21# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X21 VPWR a_761_289# a_651_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0703 pd=0.755 as=0.116 ps=0.97 w=0.42 l=0.15
X22 Q a_1283_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.209 ps=2.02 w=0.65 l=0.15
X23 a_639_47# a_193_47# a_543_47# VNB sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X24 VGND a_1283_21# a_1217_47# VNB sky130_fd_pr__nfet_01v8 ad=0.125 pd=1.01 as=0.0669 ps=0.75 w=0.42 l=0.15
X25 a_651_413# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0703 ps=0.755 w=0.42 l=0.15
X26 VGND CLK a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X27 a_761_289# a_543_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.129 pd=1.18 as=0.218 ps=2.2 w=0.84 l=0.15
.ends

.subckt sky130_fd_sc_hd__xor2_1 VPWR VGND A X B VPB VNB
X0 X a_35_297# a_285_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.26 ps=2.52 w=1 l=0.15
X1 X B a_285_47# VNB sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.42 as=0.0878 ps=0.92 w=0.65 l=0.15
X2 a_35_297# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3 a_117_297# B a_35_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4 VPWR B a_285_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5 VGND A a_35_297# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6 VGND a_35_297# X VNB sky130_fd_pr__nfet_01v8 ad=0.208 pd=1.94 as=0.25 ps=1.42 w=0.65 l=0.15
X7 a_285_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8 VPWR A a_117_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9 a_285_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__a221o_1 VPWR VGND A1 A2 X B1 B2 C1 VPB VNB
X0 a_465_47# A1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X1 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.157 ps=1.32 w=1 l=0.15
X2 a_109_297# B1 a_193_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3 a_193_297# B2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.102 ps=0.965 w=0.65 l=0.15
X5 a_205_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.86 as=0.107 ps=0.98 w=0.65 l=0.15
X6 VPWR A2 a_193_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.157 pd=1.32 as=0.165 ps=1.33 w=1 l=0.15
X7 a_193_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X8 a_27_47# B1 a_205_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0683 ps=0.86 w=0.65 l=0.15
X9 a_109_297# C1 a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X10 VGND C1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X11 VGND A2 a_465_47# VNB sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.965 as=0.107 ps=0.98 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__inv_2 VPWR VGND Y A VPB VNB
X0 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__clkbuf_2 VGND VPWR A X VPB VNB
X0 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.162 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X1 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.745 as=0.111 ps=1.37 w=0.42 l=0.15
X3 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.162 ps=1.33 w=1 l=0.15
X4 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0683 ps=0.745 w=0.42 l=0.15
X5 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__diode_2 VGND VPWR DIODE VPB VNB
C0 VNB DIODE 1f
.ends

.subckt sky130_fd_sc_hd__decap_6 VPWR VGND VPB VNB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=1.97
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.97
.ends

.subckt sky130_fd_sc_hd__decap_3 VPWR VGND VPB VNB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
.ends

.subckt sky130_fd_sc_hd__decap_8 VPWR VGND VPB VNB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
.ends

.subckt sky130_fd_sc_hd__decap_4 VGND VPWR VPB VNB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
.ends

.subckt sky130_fd_sc_hd__nand2_1 VGND VPWR A Y B VPB VNB
X0 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1 Y A a_113_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2 a_113_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__nor2_1 VGND VPWR A B Y VPB VNB
X0 VPWR A a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X1 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2 a_109_297# B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X3 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__o221a_2 VGND VPWR B1 B2 A2 A1 X C1 VPB VNB
X0 VPWR a_38_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1 VPWR A1 a_497_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.105 ps=1.21 w=1 l=0.15
X2 X a_38_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.165 ps=1.33 w=1 l=0.15
X3 a_141_47# B2 a_225_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4 a_497_297# A2 a_38_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.387 ps=1.77 w=1 l=0.15
X5 VGND A1 a_225_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6 VPWR C1 a_38_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.325 ps=2.65 w=1 l=0.15
X7 a_237_297# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.112 pd=1.23 as=0.165 ps=1.33 w=1 l=0.15
X8 a_38_47# B2 a_237_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.387 pd=1.77 as=0.112 ps=1.23 w=1 l=0.15
X9 a_225_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X10 X a_38_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X11 a_141_47# C1 a_38_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.237 ps=2.03 w=0.65 l=0.15
X12 VGND a_38_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X13 a_225_47# B1 a_141_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__clkbuf_1 VGND VPWR X A VPB VNB
X0 VPWR a_75_212# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X1 a_75_212# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X2 a_75_212# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X3 VGND a_75_212# X VNB sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
.ends

.subckt sky130_fd_sc_hd__nor2_2 VGND VPWR B Y A VPB VNB
X0 Y B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X5 VGND B Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X7 a_27_297# B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__nand2b_1 VGND VPWR A_N B Y VPB VNB
X0 VGND A_N a_27_93# VNB sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.985 as=0.109 ps=1.36 w=0.42 l=0.15
X1 Y a_27_93# a_206_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2 a_206_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.1 ps=0.985 w=0.65 l=0.15
X3 VPWR a_27_93# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X4 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.146 ps=1.34 w=1 l=0.15
X5 VPWR A_N a_27_93# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.146 pd=1.34 as=0.109 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_ef_sc_hd__decap_12 VGND VPWR VPB VNB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
.ends

.subckt sky130_fd_sc_hd__o21ai_1 VGND VPWR A2 B1 Y A1 VPB VNB
X0 Y A2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.39 as=0.105 ps=1.21 w=1 l=0.15
X1 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.182 pd=1.92 as=0.174 ps=1.39 w=0.7 l=0.15
X2 a_27_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.107 ps=0.98 w=0.65 l=0.15
X3 Y B1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4 a_109_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X5 VGND A1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__a211o_2 VGND VPWR X A2 A1 B1 C1 VPB VNB
X0 a_79_21# A1 a_348_47# VNB sky130_fd_pr__nfet_01v8 ad=0.115 pd=1 as=0.133 ps=1.06 w=0.65 l=0.15
X1 a_79_21# C1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.107 ps=0.98 w=0.65 l=0.15
X2 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.26 as=0.091 ps=0.93 w=0.65 l=0.15
X3 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4 a_79_21# C1 a_585_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X5 VPWR A2 a_299_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.26 ps=2.52 w=1 l=0.15
X6 a_299_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.195 ps=1.39 w=1 l=0.15
X7 a_585_297# B1 a_299_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.165 ps=1.33 w=1 l=0.15
X8 a_348_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.133 pd=1.06 as=0.2 ps=1.26 w=0.65 l=0.15
X9 X a_79_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X10 X a_79_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.169 ps=1.82 w=0.65 l=0.15
X11 VGND B1 a_79_21# VNB sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.115 ps=1 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__clkinv_2 VPWR VGND A Y VPB VNB
X0 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.111 ps=1.37 w=0.42 l=0.15
X1 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X3 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0588 ps=0.7 w=0.42 l=0.15
X4 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__a32o_1 VGND VPWR X A3 A2 A1 B1 B2 VPB VNB
X0 a_93_21# A1 a_346_47# VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.09 as=0.146 ps=1.1 w=0.65 l=0.15
X1 a_93_21# B1 a_250_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.185 ps=1.37 w=1 l=0.15
X2 a_584_47# B1 a_93_21# VNB sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.86 as=0.143 ps=1.09 w=0.65 l=0.15
X3 VPWR a_93_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.243 pd=1.49 as=0.33 ps=2.66 w=1 l=0.15
X4 VGND B2 a_584_47# VNB sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.0683 ps=0.86 w=0.65 l=0.15
X5 a_256_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0975 pd=0.95 as=0.167 ps=1.16 w=0.65 l=0.15
X6 a_250_297# B2 a_93_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X7 VGND a_93_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.167 pd=1.16 as=0.214 ps=1.96 w=0.65 l=0.15
X8 a_250_297# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.243 ps=1.49 w=1 l=0.15
X9 VPWR A2 a_250_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.45 as=0.165 ps=1.33 w=1 l=0.15
X10 a_250_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.185 pd=1.37 as=0.225 ps=1.45 w=1 l=0.15
X11 a_346_47# A2 a_256_47# VNB sky130_fd_pr__nfet_01v8 ad=0.146 pd=1.1 as=0.0975 ps=0.95 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__or3_1 VPWR VGND B C A X VPB VNB
X0 X a_29_53# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.148 ps=1.34 w=1 l=0.15
X1 a_111_297# C a_29_53# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X2 X a_29_53# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.102 ps=0.99 w=0.65 l=0.15
X3 a_183_297# B a_111_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X4 VPWR A a_183_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.148 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X5 a_29_53# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X6 VGND C a_29_53# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X7 VGND A a_29_53# VNB sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__a31o_1 VGND VPWR X A3 A2 A1 B1 VPB VNB
X0 VPWR a_80_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.172 pd=1.35 as=0.265 ps=2.53 w=1 l=0.15
X1 a_209_297# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.172 ps=1.35 w=1 l=0.15
X2 a_303_47# A2 a_209_47# VNB sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.104 ps=0.97 w=0.65 l=0.15
X3 a_209_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.104 pd=0.97 as=0.112 ps=0.995 w=0.65 l=0.15
X4 VGND a_80_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.112 pd=0.995 as=0.172 ps=1.83 w=0.65 l=0.15
X5 VGND B1 a_80_21# VNB sky130_fd_pr__nfet_01v8 ad=0.208 pd=1.94 as=0.107 ps=0.98 w=0.65 l=0.15
X6 a_80_21# A1 a_303_47# VNB sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.107 ps=0.98 w=0.65 l=0.15
X7 VPWR A2 a_209_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.16 ps=1.32 w=1 l=0.15
X8 a_80_21# B1 a_209_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.32 pd=2.64 as=0.165 ps=1.33 w=1 l=0.15
X9 a_209_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__or2_1 VPWR VGND X A B VPB VNB
X0 VGND A a_68_297# VNB sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X1 a_68_297# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X2 X a_68_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1 ps=0.985 w=0.65 l=0.15
X3 VPWR A a_150_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.146 pd=1.34 as=0.0441 ps=0.63 w=0.42 l=0.15
X4 X a_68_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.146 ps=1.34 w=1 l=0.15
X5 a_150_297# B a_68_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__buf_2 VPWR VGND X A VPB VNB
X0 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X1 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.33 w=1 l=0.15
X2 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.166 ps=1.8 w=0.64 l=0.15
X3 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X4 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.0878 ps=0.92 w=0.65 l=0.15
X5 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__nand3_1 VGND VPWR A B Y C VPB VNB
X0 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X1 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.165 ps=1.33 w=1 l=0.15
X2 a_193_47# B a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.0878 ps=0.92 w=0.65 l=0.15
X3 Y A a_193_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.107 ps=0.98 w=0.65 l=0.15
X4 Y C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5 a_109_47# C VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__and2_1 VPWR VGND X A B VPB VNB
X0 VPWR B a_59_75# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.167 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X1 X a_59_75# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.167 ps=1.39 w=1 l=0.15
X2 VGND B a_145_75# VNB sky130_fd_pr__nfet_01v8 ad=0.112 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X3 a_59_75# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
X4 X a_59_75# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.112 ps=1.04 w=0.65 l=0.15
X5 a_145_75# A a_59_75# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__a21oi_1 VPWR VGND A2 A1 B1 Y VPB VNB
X0 a_199_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.0959 pd=0.945 as=0.091 ps=0.93 w=0.65 l=0.15
X1 a_113_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.147 ps=1.29 w=1 l=0.15
X2 Y B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.172 ps=1.83 w=0.65 l=0.15
X3 VPWR A1 a_113_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.29 as=0.14 ps=1.28 w=1 l=0.15
X4 a_113_297# B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X5 VGND A2 a_199_47# VNB sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.0959 ps=0.945 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__a21oi_2 VGND VPWR A2 A1 Y B1 VPB VNB
X0 VGND A2 a_285_47# VNB sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.0683 ps=0.86 w=0.65 l=0.15
X1 VGND B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.26 pd=2.1 as=0.0878 ps=0.92 w=0.65 l=0.15
X2 Y A1 a_114_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.0894 ps=0.925 w=0.65 l=0.15
X3 a_114_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0894 pd=0.925 as=0.185 ps=1.87 w=0.65 l=0.15
X4 a_27_297# B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.36 pd=2.72 as=0.135 ps=1.27 w=1 l=0.15
X5 a_27_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6 Y B1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7 VPWR A2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.28 ps=2.56 w=1 l=0.15
X8 a_27_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9 VPWR A1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.14 ps=1.28 w=1 l=0.15
X10 a_285_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.86 as=0.091 ps=0.93 w=0.65 l=0.15
X11 Y B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.107 ps=0.98 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__dfrtp_2 VGND VPWR CLK D RESET_B Q VPB VNB
X0 a_1217_47# a_27_47# a_1108_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X1 a_805_47# a_761_289# a_639_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.14 ps=1.1 w=0.42 l=0.15
X2 VGND a_1283_21# Q VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3 a_1108_47# a_193_47# a_761_289# VNB sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X4 a_1283_21# a_1108_47# a_1462_47# VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.064 ps=0.725 w=0.42 l=0.15
X5 a_651_413# a_27_47# a_543_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.116 pd=0.97 as=0.0724 ps=0.765 w=0.42 l=0.15
X6 VPWR a_1283_21# Q VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7 VGND RESET_B a_805_47# VNB sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X8 Q a_1283_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.301 ps=2.66 w=1 l=0.15
X9 VPWR CLK a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X10 a_448_47# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.109 ps=1.36 w=0.42 l=0.15
X11 a_761_289# a_543_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.135 ps=1.15 w=0.64 l=0.15
X12 a_193_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X13 a_1108_47# a_27_47# a_761_289# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.129 ps=1.18 w=0.42 l=0.15
X14 a_543_47# a_27_47# a_448_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X15 a_1462_47# RESET_B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.064 pd=0.725 as=0.125 ps=1.01 w=0.42 l=0.15
X16 a_543_47# a_193_47# a_448_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0724 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X17 a_448_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.221 ps=1.89 w=0.42 l=0.15
X18 VPWR a_1283_21# a_1270_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X19 VPWR a_1108_47# a_1283_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X20 a_1270_413# a_193_47# a_1108_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X21 a_193_47# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X22 a_1283_21# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X23 VPWR a_761_289# a_651_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0703 pd=0.755 as=0.116 ps=0.97 w=0.42 l=0.15
X24 Q a_1283_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.209 ps=2.02 w=0.65 l=0.15
X25 a_639_47# a_193_47# a_543_47# VNB sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X26 VGND a_1283_21# a_1217_47# VNB sky130_fd_pr__nfet_01v8 ad=0.125 pd=1.01 as=0.0669 ps=0.75 w=0.42 l=0.15
X27 a_651_413# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0703 ps=0.755 w=0.42 l=0.15
X28 VGND CLK a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X29 a_761_289# a_543_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.129 pd=1.18 as=0.218 ps=2.2 w=0.84 l=0.15
.ends

.subckt sky130_fd_sc_hd__buf_6 VPWR VGND A X VPB VNB
X0 VPWR a_161_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1 a_161_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2 X a_161_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 VPWR a_161_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4 VGND A a_161_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5 X a_161_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6 VGND a_161_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X7 VGND a_161_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X8 VPWR a_161_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9 X a_161_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X10 X a_161_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X11 X a_161_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X12 X a_161_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X13 VPWR A a_161_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X14 VGND a_161_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X15 a_161_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__dlymetal6s2s_1 VPWR VGND X A VPB VNB
X0 a_558_47# a_381_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.141 ps=1.33 w=1 l=0.15
X1 VGND X a_381_47# VNB sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X2 a_841_47# a_664_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.141 ps=1.33 w=1 l=0.15
X3 VPWR A a_62_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.141 pd=1.33 as=0.109 ps=1.36 w=0.42 l=0.15
X4 VGND A a_62_47# VNB sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X5 a_558_47# a_381_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X6 X a_62_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.141 ps=1.33 w=1 l=0.15
X7 VPWR X a_381_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.141 pd=1.33 as=0.109 ps=1.36 w=0.42 l=0.15
X8 a_841_47# a_664_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X9 X a_62_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X10 VPWR a_558_47# a_664_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.141 pd=1.33 as=0.109 ps=1.36 w=0.42 l=0.15
X11 VGND a_558_47# a_664_47# VNB sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__or2b_1 VGND VPWR A X B_N VPB VNB
X0 a_219_297# a_27_53# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.157 ps=1.17 w=0.42 l=0.15
X1 VGND B_N a_27_53# VNB sky130_fd_pr__nfet_01v8 ad=0.157 pd=1.17 as=0.109 ps=1.36 w=0.42 l=0.15
X2 VPWR A a_301_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.148 pd=1.34 as=0.0441 ps=0.63 w=0.42 l=0.15
X3 X a_219_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.176 pd=1.84 as=0.102 ps=0.99 w=0.65 l=0.15
X4 a_301_297# a_27_53# a_219_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X5 X a_219_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.148 ps=1.34 w=1 l=0.15
X6 a_27_53# B_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.118 pd=1.4 as=0.109 ps=1.36 w=0.42 l=0.15
X7 VGND A a_219_297# VNB sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__o221a_1 VGND VPWR B1 B2 A2 A1 X C1 VPB VNB
X0 a_240_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1 X a_51_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.0878 ps=0.92 w=0.65 l=0.15
X2 VGND A1 a_240_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3 a_51_297# B2 a_245_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.412 pd=1.83 as=0.105 ps=1.21 w=1 l=0.15
X4 a_149_47# C1 a_51_297# VNB sky130_fd_pr__nfet_01v8 ad=0.0991 pd=0.955 as=0.201 ps=1.92 w=0.65 l=0.15
X5 a_240_47# B1 a_149_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0991 ps=0.955 w=0.65 l=0.15
X6 VPWR A1 a_512_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.105 ps=1.21 w=1 l=0.15
X7 X a_51_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.165 ps=1.33 w=1 l=0.15
X8 a_149_47# B2 a_240_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X9 a_245_297# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.165 ps=1.33 w=1 l=0.15
X10 VPWR C1 a_51_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.34 ps=2.68 w=1 l=0.15
X11 a_512_297# A2 a_51_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.412 ps=1.83 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__a21o_2 VGND VPWR A2 A1 B1 X VPB VNB
X0 VPWR a_80_199# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X1 X a_80_199# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X2 VGND a_80_199# X VNB sky130_fd_pr__nfet_01v8 ad=0.111 pd=0.99 as=0.091 ps=0.93 w=0.65 l=0.15
X3 a_386_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.157 ps=1.32 w=1 l=0.15
X4 X a_80_199# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.172 ps=1.83 w=0.65 l=0.15
X5 a_80_199# B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.162 pd=1.15 as=0.111 ps=0.99 w=0.65 l=0.15
X6 a_386_297# B1 a_80_199# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X7 a_458_47# A1 a_80_199# VNB sky130_fd_pr__nfet_01v8 ad=0.123 pd=1.03 as=0.162 ps=1.15 w=0.65 l=0.15
X8 VPWR A1 a_386_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.157 pd=1.32 as=0.14 ps=1.28 w=1 l=0.15
X9 VGND A2 a_458_47# VNB sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.123 ps=1.03 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__nand2_2 VGND VPWR Y A B VPB VNB
X0 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 a_27_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4 a_27_47# A Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5 Y A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7 VGND B a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__and3_1 VGND VPWR X C B A VPB VNB
X0 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1 VPWR C a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.0662 ps=0.735 w=0.42 l=0.15
X2 a_181_47# B a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X3 VGND C a_181_47# VNB sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X4 a_27_47# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X5 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142 ps=1.34 w=1 l=0.15
X6 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.132 ps=1.14 w=0.65 l=0.15
X7 a_109_47# A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__a221o_4 VPWR VGND A2 X A1 C1 B1 B2 VPB VNB
X0 VGND A2 a_445_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1 VGND B2 a_1053_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2 a_804_297# B1 a_445_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.345 pd=1.69 as=0.135 ps=1.27 w=1 l=0.15
X3 a_79_21# A1 a_445_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4 a_445_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5 a_804_297# C1 a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6 a_445_297# B1 a_804_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8 a_1053_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X9 a_79_21# C1 a_804_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X10 a_1053_47# B1 a_79_21# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X11 X a_79_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X12 a_445_47# A1 a_79_21# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X13 VGND C1 a_79_21# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X14 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X15 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X16 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X17 a_804_297# B2 a_445_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X18 a_79_21# B1 a_1053_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X19 a_79_21# C1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X20 a_445_297# B2 a_804_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.345 ps=1.69 w=1 l=0.15
X21 X a_79_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X22 a_445_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X23 a_445_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.138 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X24 VPWR A2 a_445_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X25 VPWR A1 a_445_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.138 ps=1.27 w=1 l=0.15
X26 X a_79_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X27 X a_79_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__nor3_1 VGND VPWR C B A Y VPB VNB
X0 VPWR A a_193_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1 a_193_297# B a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4 a_109_297# C Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5 VGND C Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__o21a_1 VGND VPWR A1 A2 B1 X VPB VNB
X0 VPWR A1 a_382_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.153 ps=1.3 w=1 l=0.15
X1 a_297_47# B1 a_79_21# VNB sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.169 ps=1.82 w=0.65 l=0.15
X2 a_297_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3 VGND A2 a_297_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.101 ps=0.96 w=0.65 l=0.15
X4 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.327 pd=1.65 as=0.28 ps=2.56 w=1 l=0.15
X5 a_79_21# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.327 ps=1.65 w=1 l=0.15
X6 a_382_297# A2 a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.153 pd=1.3 as=0.195 ps=1.39 w=1 l=0.15
X7 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__mux2_1 VGND VPWR X A1 S A0 VPB VNB
X0 VPWR a_505_21# a_535_374# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X1 a_505_21# S VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.118 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X2 a_218_374# S VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.158 ps=1.39 w=0.42 l=0.15
X3 VGND a_505_21# a_439_47# VNB sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X4 a_76_199# A0 a_218_374# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.193 pd=1.34 as=0.0767 ps=0.785 w=0.42 l=0.15
X5 a_505_21# S VGND VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.145 ps=1.11 w=0.42 l=0.15
X6 a_439_47# A0 a_76_199# VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0997 ps=0.895 w=0.42 l=0.15
X7 a_535_374# A1 a_76_199# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.193 ps=1.34 w=0.42 l=0.15
X8 a_76_199# A1 a_218_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0997 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X9 a_218_47# S VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.113 ps=1.04 w=0.42 l=0.15
X10 VPWR a_76_199# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.158 pd=1.39 as=0.26 ps=2.52 w=1 l=0.15
X11 VGND a_76_199# X VNB sky130_fd_pr__nfet_01v8 ad=0.113 pd=1.04 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__inv_1 VGND VPWR A Y VPB VNB
X0 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X1 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
.ends

.subckt pfet_01v8_w500_l500_nf2 a_n29_0# a_129_0# a_n129_n26# w_n224_n36# a_n187_0#
+ a_29_n26#
X0 a_129_0# a_29_n26# a_n29_0# w_n224_n36# sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.58 as=0.0725 ps=0.79 w=0.5 l=0.5
X1 a_n29_0# a_n129_n26# a_n187_0# w_n224_n36# sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.145 ps=1.58 w=0.5 l=0.5
.ends

.subckt sky130_fd_sc_hd__buf_4 VPWR VGND A X VPB VNB
X0 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X7 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X8 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X9 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__dlymetal6s6s_1 VPWR VGND X A VPB VNB
X0 X a_629_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X1 a_523_47# a_346_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X2 VGND a_240_47# a_346_47# VNB sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X3 a_240_47# a_63_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X4 VPWR a_240_47# a_346_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.141 pd=1.33 as=0.109 ps=1.36 w=0.42 l=0.15
X5 VGND A a_63_47# VNB sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X6 VPWR A a_63_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.141 pd=1.33 as=0.109 ps=1.36 w=0.42 l=0.15
X7 VPWR a_523_47# a_629_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.141 pd=1.33 as=0.109 ps=1.36 w=0.42 l=0.15
X8 VGND a_523_47# a_629_47# VNB sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X9 a_523_47# a_346_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.141 ps=1.33 w=1 l=0.15
X10 a_240_47# a_63_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.141 ps=1.33 w=1 l=0.15
X11 X a_629_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.141 ps=1.33 w=1 l=0.15
.ends

.subckt adc_noise_decoup_cell1 nmoscap_top nmoscap_bot pwell mimcap_top mimcap_bot
X0 nmoscap_top nmoscap_bot pwell sky130_fd_pr__cap_var_lvt w=16.4 l=16
X1 mimcap_top mimcap_bot sky130_fd_pr__cap_mim_m3_1 l=17.2 w=17.2
.ends

.subckt nfet_01v8_w500_l500_nf2 a_n129_n76# a_n29_n50# a_n187_n50# a_29_n76# a_129_n50#
+ VSUBS
X0 a_129_n50# a_29_n76# a_n29_n50# VSUBS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.0725 ps=0.79 w=0.5 l=0.5
X1 a_n29_n50# a_n129_n76# a_n187_n50# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.145 ps=1.58 w=0.5 l=0.5
.ends

.subckt adc_vcm_generator clk phi2 phi1_n phi1 phi2_n vcm VDD mimtop1 mimtop2 mimbot1
+ VSS
Xsky130_fd_sc_hd__inv_1_4 VSS VDD clk sky130_fd_sc_hd__inv_1_4/Y VDD VSS sky130_fd_sc_hd__inv_1
Xpfet_01v8_w500_l500_nf2_0 mimtop2 vcm phi1_n VDD vcm phi1_n pfet_01v8_w500_l500_nf2
Xpfet_01v8_w500_l500_nf2_1 mimtop1 vcm phi1_n VDD vcm phi1_n pfet_01v8_w500_l500_nf2
Xpfet_01v8_w500_l500_nf2_2 mimtop2 mimbot1 phi2_n VDD mimbot1 phi2_n pfet_01v8_w500_l500_nf2
Xsky130_fd_sc_hd__buf_4_0 VDD VSS sky130_fd_sc_hd__inv_1_2/A phi1 VDD VSS sky130_fd_sc_hd__buf_4
Xpfet_01v8_w500_l500_nf2_3 VDD mimtop1 phi2_n VDD mimtop1 phi2_n pfet_01v8_w500_l500_nf2
Xsky130_fd_sc_hd__buf_4_1 VDD VSS sky130_fd_sc_hd__inv_1_2/Y phi1_n VDD VSS sky130_fd_sc_hd__buf_4
Xsky130_fd_sc_hd__buf_4_2 VDD VSS sky130_fd_sc_hd__inv_1_3/A phi2 VDD VSS sky130_fd_sc_hd__buf_4
Xpfet_01v8_w500_l500_nf2_4 mimbot1 VSS phi1_n VDD VSS phi1_n pfet_01v8_w500_l500_nf2
Xsky130_fd_sc_hd__buf_4_3 VDD VSS sky130_fd_sc_hd__inv_1_3/Y phi2_n VDD VSS sky130_fd_sc_hd__buf_4
Xsky130_fd_sc_hd__dlymetal6s6s_1_0 VDD VSS sky130_fd_sc_hd__dlymetal6s6s_1_2/A sky130_fd_sc_hd__nand2_1_0/Y
+ VDD VSS sky130_fd_sc_hd__dlymetal6s6s_1
Xsky130_fd_sc_hd__dlymetal6s6s_1_1 VDD VSS sky130_fd_sc_hd__dlymetal6s6s_1_4/A sky130_fd_sc_hd__nand2_1_1/Y
+ VDD VSS sky130_fd_sc_hd__dlymetal6s6s_1
Xsky130_fd_sc_hd__dlymetal6s6s_1_2 VDD VSS sky130_fd_sc_hd__dlymetal6s6s_1_3/A sky130_fd_sc_hd__dlymetal6s6s_1_2/A
+ VDD VSS sky130_fd_sc_hd__dlymetal6s6s_1
Xsky130_fd_sc_hd__dlymetal6s6s_1_3 VDD VSS sky130_fd_sc_hd__inv_1_0/A sky130_fd_sc_hd__dlymetal6s6s_1_3/A
+ VDD VSS sky130_fd_sc_hd__dlymetal6s6s_1
Xsky130_fd_sc_hd__dlymetal6s6s_1_4 VDD VSS sky130_fd_sc_hd__dlymetal6s6s_1_5/A sky130_fd_sc_hd__dlymetal6s6s_1_4/A
+ VDD VSS sky130_fd_sc_hd__dlymetal6s6s_1
Xsky130_fd_sc_hd__dlymetal6s6s_1_5 VDD VSS sky130_fd_sc_hd__inv_1_1/A sky130_fd_sc_hd__dlymetal6s6s_1_5/A
+ VDD VSS sky130_fd_sc_hd__dlymetal6s6s_1
Xadc_noise_decoup_cell1_0[0] VDD VSS VSS VDD VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_0[1] VDD VSS VSS VDD VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_0[2] VDD VSS VSS VDD VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[0|0] vcm VSS VSS adc_noise_decoup_cell1_1[0|4]/mimcap_top
+ VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[1|0] vcm VSS VSS adc_noise_decoup_cell1_1[1|4]/mimcap_top
+ VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[2|0] vcm VSS VSS adc_noise_decoup_cell1_1[2|4]/mimcap_top
+ VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[3|0] vcm VSS VSS adc_noise_decoup_cell1_1[3|4]/mimcap_top
+ VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[4|0] vcm VSS VSS adc_noise_decoup_cell1_1[4|4]/mimcap_top
+ VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[5|0] vcm VSS VSS adc_noise_decoup_cell1_1[5|4]/mimcap_top
+ VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[6|0] vcm VSS VSS adc_noise_decoup_cell1_1[6|4]/mimcap_top
+ VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[7|0] vcm VSS VSS mimtop2 VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[0|1] vcm VSS VSS adc_noise_decoup_cell1_1[0|4]/mimcap_top
+ VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[1|1] vcm VSS VSS adc_noise_decoup_cell1_1[1|4]/mimcap_top
+ VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[2|1] vcm VSS VSS adc_noise_decoup_cell1_1[2|4]/mimcap_top
+ VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[3|1] vcm VSS VSS adc_noise_decoup_cell1_1[3|4]/mimcap_top
+ VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[4|1] vcm VSS VSS adc_noise_decoup_cell1_1[4|4]/mimcap_top
+ VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[5|1] vcm VSS VSS adc_noise_decoup_cell1_1[5|4]/mimcap_top
+ VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[6|1] vcm VSS VSS adc_noise_decoup_cell1_1[6|4]/mimcap_top
+ VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[7|1] vcm VSS VSS mimtop2 VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[0|2] vcm VSS VSS adc_noise_decoup_cell1_1[0|4]/mimcap_top
+ VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[1|2] vcm VSS VSS adc_noise_decoup_cell1_1[1|4]/mimcap_top
+ VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[2|2] vcm VSS VSS adc_noise_decoup_cell1_1[2|4]/mimcap_top
+ VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[3|2] vcm VSS VSS adc_noise_decoup_cell1_1[3|4]/mimcap_top
+ VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[4|2] vcm VSS VSS adc_noise_decoup_cell1_1[4|4]/mimcap_top
+ VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[5|2] vcm VSS VSS adc_noise_decoup_cell1_1[5|4]/mimcap_top
+ VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[6|2] vcm VSS VSS adc_noise_decoup_cell1_1[6|4]/mimcap_top
+ VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[7|2] vcm VSS VSS mimtop2 VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[0|3] vcm VSS VSS adc_noise_decoup_cell1_1[0|4]/mimcap_top
+ VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[1|3] vcm VSS VSS adc_noise_decoup_cell1_1[1|4]/mimcap_top
+ VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[2|3] vcm VSS VSS adc_noise_decoup_cell1_1[2|4]/mimcap_top
+ VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[3|3] vcm VSS VSS adc_noise_decoup_cell1_1[3|4]/mimcap_top
+ VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[4|3] vcm VSS VSS adc_noise_decoup_cell1_1[4|4]/mimcap_top
+ VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[5|3] vcm VSS VSS adc_noise_decoup_cell1_1[5|4]/mimcap_top
+ VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[6|3] vcm VSS VSS adc_noise_decoup_cell1_1[6|4]/mimcap_top
+ VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[7|3] vcm VSS VSS mimtop2 VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[0|4] vcm VSS VSS adc_noise_decoup_cell1_1[0|4]/mimcap_top
+ VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[1|4] vcm VSS VSS adc_noise_decoup_cell1_1[1|4]/mimcap_top
+ VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[2|4] vcm VSS VSS adc_noise_decoup_cell1_1[2|4]/mimcap_top
+ VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[3|4] vcm VSS VSS adc_noise_decoup_cell1_1[3|4]/mimcap_top
+ VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[4|4] vcm VSS VSS adc_noise_decoup_cell1_1[4|4]/mimcap_top
+ VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[5|4] vcm VSS VSS adc_noise_decoup_cell1_1[5|4]/mimcap_top
+ VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[6|4] vcm VSS VSS adc_noise_decoup_cell1_1[6|4]/mimcap_top
+ VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[7|4] vcm VSS VSS mimtop2 VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_3[0|0] vcm VSS VSS mimtop1 mimbot1 adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_3[1|0] vcm VSS VSS mimtop1 mimbot1 adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_3[2|0] vcm VSS VSS mimtop1 mimbot1 adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_3[3|0] vcm VSS VSS mimtop1 mimbot1 adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_3[4|0] vcm VSS VSS mimtop1 mimbot1 adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_3[5|0] vcm VSS VSS mimtop1 mimbot1 adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_3[6|0] vcm VSS VSS mimtop1 mimbot1 adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_3[7|0] vcm VSS VSS mimtop1 mimbot1 adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_3[0|1] vcm VSS VSS mimtop1 mimbot1 adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_3[1|1] vcm VSS VSS mimtop1 mimbot1 adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_3[2|1] vcm VSS VSS mimtop1 mimbot1 adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_3[3|1] vcm VSS VSS mimtop1 mimbot1 adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_3[4|1] vcm VSS VSS mimtop1 mimbot1 adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_3[5|1] vcm VSS VSS mimtop1 mimbot1 adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_3[6|1] vcm VSS VSS mimtop1 mimbot1 adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_3[7|1] vcm VSS VSS mimtop1 mimbot1 adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_3[0|2] vcm VSS VSS mimtop1 mimbot1 adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_3[1|2] vcm VSS VSS mimtop1 mimbot1 adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_3[2|2] vcm VSS VSS mimtop1 mimbot1 adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_3[3|2] vcm VSS VSS mimtop1 mimbot1 adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_3[4|2] vcm VSS VSS mimtop1 mimbot1 adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_3[5|2] vcm VSS VSS mimtop1 mimbot1 adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_3[6|2] vcm VSS VSS mimtop1 mimbot1 adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_3[7|2] vcm VSS VSS mimtop1 mimbot1 adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_3[0|3] vcm VSS VSS mimtop1 mimbot1 adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_3[1|3] vcm VSS VSS mimtop1 mimbot1 adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_3[2|3] vcm VSS VSS mimtop1 mimbot1 adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_3[3|3] vcm VSS VSS mimtop1 mimbot1 adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_3[4|3] vcm VSS VSS mimtop1 mimbot1 adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_3[5|3] vcm VSS VSS mimtop1 mimbot1 adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_3[6|3] vcm VSS VSS mimtop1 mimbot1 adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_3[7|3] vcm VSS VSS mimtop1 mimbot1 adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_3[0|4] vcm VSS VSS mimtop1 mimbot1 adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_3[1|4] vcm VSS VSS mimtop1 mimbot1 adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_3[2|4] vcm VSS VSS mimtop1 mimbot1 adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_3[3|4] vcm VSS VSS mimtop1 mimbot1 adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_3[4|4] vcm VSS VSS mimtop1 mimbot1 adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_3[5|4] vcm VSS VSS mimtop1 mimbot1 adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_3[6|4] vcm VSS VSS mimtop1 mimbot1 adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_3[7|4] vcm VSS VSS mimtop1 mimbot1 adc_noise_decoup_cell1
Xnfet_01v8_w500_l500_nf2_0 phi1 mimtop2 vcm phi1 vcm VSS nfet_01v8_w500_l500_nf2
Xsky130_fd_sc_hd__nand2_1_0 VSS VDD clk sky130_fd_sc_hd__nand2_1_0/Y sky130_fd_sc_hd__inv_1_3/Y
+ VDD VSS sky130_fd_sc_hd__nand2_1
Xnfet_01v8_w500_l500_nf2_1 phi1 mimtop1 vcm phi1 vcm VSS nfet_01v8_w500_l500_nf2
Xsky130_fd_sc_hd__nand2_1_1 VSS VDD sky130_fd_sc_hd__inv_1_2/Y sky130_fd_sc_hd__nand2_1_1/Y
+ sky130_fd_sc_hd__inv_1_4/Y VDD VSS sky130_fd_sc_hd__nand2_1
Xnfet_01v8_w500_l500_nf2_3 phi2 VDD mimtop1 phi2 mimtop1 VSS nfet_01v8_w500_l500_nf2
Xnfet_01v8_w500_l500_nf2_2 phi2 mimtop2 mimbot1 phi2 mimbot1 VSS nfet_01v8_w500_l500_nf2
Xnfet_01v8_w500_l500_nf2_4 phi1 mimbot1 VSS phi1 VSS VSS nfet_01v8_w500_l500_nf2
Xsky130_fd_sc_hd__inv_1_1 VSS VDD sky130_fd_sc_hd__inv_1_1/A sky130_fd_sc_hd__inv_1_3/A
+ VDD VSS sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_1_0 VSS VDD sky130_fd_sc_hd__inv_1_0/A sky130_fd_sc_hd__inv_1_2/A
+ VDD VSS sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_1_2 VSS VDD sky130_fd_sc_hd__inv_1_2/A sky130_fd_sc_hd__inv_1_2/Y
+ VDD VSS sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_1_3 VSS VDD sky130_fd_sc_hd__inv_1_3/A sky130_fd_sc_hd__inv_1_3/Y
+ VDD VSS sky130_fd_sc_hd__inv_1
.ends

.subckt sky130_fd_sc_hd__dfrtp_4 VGND VPWR CLK D RESET_B Q VPB VNB
X0 a_1217_47# a_27_47# a_1108_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X1 a_805_47# a_761_289# a_639_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.14 ps=1.1 w=0.42 l=0.15
X2 a_1108_47# a_193_47# a_761_289# VNB sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X3 a_1283_21# a_1108_47# a_1462_47# VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.064 ps=0.725 w=0.42 l=0.15
X4 a_651_413# a_27_47# a_543_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.116 pd=0.97 as=0.0724 ps=0.765 w=0.42 l=0.15
X5 VGND RESET_B a_805_47# VNB sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X6 VPWR a_1283_21# Q VPB sky130_fd_pr__pfet_01v8_hvt ad=0.305 pd=2.61 as=0.135 ps=1.27 w=1 l=0.15
X7 VPWR CLK a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X8 a_448_47# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.109 ps=1.36 w=0.42 l=0.15
X9 Q a_1283_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X10 VPWR a_1283_21# Q VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X11 a_761_289# a_543_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.135 ps=1.15 w=0.64 l=0.15
X12 Q a_1283_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X13 a_193_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X14 a_1108_47# a_27_47# a_761_289# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.129 ps=1.18 w=0.42 l=0.15
X15 a_543_47# a_27_47# a_448_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X16 a_1462_47# RESET_B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.064 pd=0.725 as=0.125 ps=1.01 w=0.42 l=0.15
X17 a_543_47# a_193_47# a_448_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0724 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X18 a_448_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.221 ps=1.89 w=0.42 l=0.15
X19 VPWR a_1283_21# a_1270_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X20 VPWR a_1108_47# a_1283_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X21 Q a_1283_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X22 a_1270_413# a_193_47# a_1108_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X23 a_193_47# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X24 a_1283_21# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X25 VGND a_1283_21# Q VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X26 VGND a_1283_21# Q VNB sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.0878 ps=0.92 w=0.65 l=0.15
X27 VPWR a_761_289# a_651_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0703 pd=0.755 as=0.116 ps=0.97 w=0.42 l=0.15
X28 a_639_47# a_193_47# a_543_47# VNB sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X29 VGND a_1283_21# a_1217_47# VNB sky130_fd_pr__nfet_01v8 ad=0.125 pd=1.01 as=0.0669 ps=0.75 w=0.42 l=0.15
X30 a_651_413# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0703 ps=0.755 w=0.42 l=0.15
X31 VGND CLK a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X32 a_761_289# a_543_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.129 pd=1.18 as=0.218 ps=2.2 w=0.84 l=0.15
X33 Q a_1283_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__o21ai_2 VGND VPWR B1 A1 Y A2 VPB VNB
X0 VGND A2 a_29_47# VNB sky130_fd_pr__nfet_01v8 ad=0.127 pd=1.04 as=0.091 ps=0.93 w=0.65 l=0.15
X1 Y B1 a_29_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X2 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X3 VPWR A1 a_112_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.175 ps=1.35 w=1 l=0.15
X4 a_29_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X5 Y A2 a_112_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6 VGND A1 a_29_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.172 ps=1.83 w=0.65 l=0.15
X7 a_112_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X8 a_112_297# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.175 pd=1.35 as=0.14 ps=1.28 w=1 l=0.15
X9 a_29_47# B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X10 Y B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.16 ps=1.32 w=1 l=0.15
X11 a_29_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.127 ps=1.04 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__a22o_1 VPWR VGND B1 A1 A2 X B2 VPB VNB
X0 VPWR A2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X1 a_27_297# B1 a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0747 ps=0.88 w=0.65 l=0.15
X2 VGND A2 a_373_47# VNB sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.114 ps=1 w=0.65 l=0.15
X3 X a_27_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X4 a_27_297# B1 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.253 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5 a_109_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.253 ps=2.52 w=1 l=0.15
X6 a_373_47# A1 a_27_297# VNB sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X7 X a_27_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.101 ps=0.96 w=0.65 l=0.15
X8 a_109_297# B2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X9 a_109_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0747 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__or4_1 VPWR VGND B D C A X VPB VNB
X0 a_27_297# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X1 a_27_297# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.109 ps=1.36 w=0.42 l=0.15
X2 a_277_297# B a_205_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X3 VPWR A a_277_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.148 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X4 X a_27_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.176 pd=1.84 as=0.102 ps=0.99 w=0.65 l=0.15
X5 a_205_297# C a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X6 X a_27_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.148 ps=1.34 w=1 l=0.15
X7 VGND C a_27_297# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0693 ps=0.75 w=0.42 l=0.15
X8 a_109_297# D a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.109 ps=1.36 w=0.42 l=0.15
X9 VGND A a_27_297# VNB sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__o221ai_1 VGND VPWR A1 A2 Y B2 C1 B1 VPB VNB
X0 a_109_47# B1 a_213_123# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.165 ps=1.82 w=0.65 l=0.15
X1 Y B2 a_295_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.45 as=0.12 ps=1.24 w=1 l=0.15
X2 VPWR A1 a_493_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X3 a_213_123# B2 a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0.117 pd=1.01 as=0.0878 ps=0.92 w=0.65 l=0.15
X4 a_295_297# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.12 pd=1.24 as=0.38 ps=1.76 w=1 l=0.15
X5 a_493_297# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.225 ps=1.45 w=1 l=0.15
X6 VPWR C1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.38 pd=1.76 as=0.28 ps=2.56 w=1 l=0.15
X7 VGND A2 a_213_123# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.117 ps=1.01 w=0.65 l=0.15
X8 a_213_123# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X9 a_109_47# C1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__nand3_2 VGND VPWR C A Y B VPB VNB
X0 VGND C a_277_47# VNB sky130_fd_pr__nfet_01v8 ad=0.201 pd=1.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2 a_277_47# C VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5 a_27_47# A Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6 a_27_47# B a_277_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7 VPWR C Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.31 pd=2.62 as=0.135 ps=1.27 w=1 l=0.15
X8 Y C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X9 a_277_47# B a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X10 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X11 Y A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__a21o_1 VPWR VGND A2 A1 B1 X VPB VNB
X0 a_81_21# B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0894 pd=0.925 as=0.257 ps=1.44 w=0.65 l=0.15
X1 a_299_297# B1 a_81_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.138 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2 VPWR a_81_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X3 VPWR A1 a_299_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.138 ps=1.27 w=1 l=0.15
X4 VGND a_81_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.257 pd=1.44 as=0.169 ps=1.82 w=0.65 l=0.15
X5 VGND A2 a_384_47# VNB sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X6 a_299_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X7 a_384_47# A1 a_81_21# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.0894 ps=0.925 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__mux2_2 VGND VPWR S A1 A0 X VPB VNB
X0 VPWR S a_591_369# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.0672 ps=0.85 w=0.64 l=0.15
X1 a_591_369# A0 a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0672 pd=0.85 as=0.131 ps=1.05 w=0.64 l=0.15
X2 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.178 pd=1.41 as=0.135 ps=1.27 w=1 l=0.15
X3 a_79_21# A1 a_306_369# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.131 pd=1.05 as=0.229 ps=1.36 w=0.64 l=0.15
X4 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.0878 ps=0.92 w=0.65 l=0.15
X5 VGND S a_578_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0578 ps=0.695 w=0.42 l=0.15
X6 a_306_369# a_257_199# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.229 pd=1.36 as=0.178 ps=1.41 w=0.64 l=0.15
X7 a_79_21# A0 a_288_47# VNB sky130_fd_pr__nfet_01v8 ad=0.173 pd=1.25 as=0.0683 ps=0.745 w=0.42 l=0.15
X8 a_288_47# a_257_199# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.745 as=0.097 ps=0.975 w=0.42 l=0.15
X9 a_257_199# S VGND VNB sky130_fd_pr__nfet_01v8 ad=0.113 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X10 a_578_47# A1 a_79_21# VNB sky130_fd_pr__nfet_01v8 ad=0.0578 pd=0.695 as=0.173 ps=1.25 w=0.42 l=0.15
X11 X a_79_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X12 a_257_199# S VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.173 pd=1.82 as=0.0864 ps=0.91 w=0.64 l=0.15
X13 X a_79_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__and4_1 VGND VPWR X D C B A VPB VNB
X0 a_27_47# C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0777 ps=0.79 w=0.42 l=0.15
X1 a_197_47# B a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0798 pd=0.8 as=0.0609 ps=0.71 w=0.42 l=0.15
X2 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.312 ps=1.68 w=1 l=0.15
X3 a_303_47# C a_197_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0798 ps=0.8 w=0.42 l=0.15
X4 a_27_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0735 pd=0.77 as=0.109 ps=1.36 w=0.42 l=0.15
X5 VPWR D a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.312 pd=1.68 as=0.0588 ps=0.7 w=0.42 l=0.15
X6 VGND D a_303_47# VNB sky130_fd_pr__nfet_01v8 ad=0.196 pd=1.33 as=0.0693 ps=0.75 w=0.42 l=0.15
X7 VPWR B a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0777 pd=0.79 as=0.0735 ps=0.77 w=0.42 l=0.15
X8 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.196 ps=1.33 w=0.65 l=0.15
X9 a_109_47# A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.109 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__and2b_1 VGND VPWR A_N X B VPB VNB
X0 VPWR B a_207_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.228 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X1 X a_207_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.228 ps=1.74 w=1 l=0.15
X2 a_297_47# a_27_413# a_207_413# VNB sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.109 ps=1.36 w=0.42 l=0.15
X3 X a_207_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.101 ps=0.99 w=0.65 l=0.15
X4 a_207_413# a_27_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X5 VPWR A_N a_27_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.109 ps=1.36 w=0.42 l=0.15
X6 VGND B a_297_47# VNB sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X7 a_27_413# A_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__clkinvlp_2 VGND VPWR A Y VPB VNB
X0 Y A a_150_67# VNB sky130_fd_pr__nfet_01v8 ad=0.157 pd=1.67 as=0.066 ps=0.79 w=0.55 l=0.15
X1 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.39 pd=2.78 as=0.14 ps=1.28 w=1 l=0.25
X2 a_150_67# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.79 as=0.157 ps=1.67 w=0.55 l=0.15
X3 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.25
.ends

.subckt sky130_fd_sc_hd__or3b_1 VGND VPWR B C_N A X VPB VNB
X0 a_109_93# C_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X1 a_215_53# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X2 VGND a_109_93# a_215_53# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X3 VGND A a_215_53# VNB sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X4 VPWR A a_369_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.148 pd=1.34 as=0.0683 ps=0.745 w=0.42 l=0.15
X5 a_369_297# B a_297_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0441 ps=0.63 w=0.42 l=0.15
X6 X a_215_53# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.275 pd=2.55 as=0.148 ps=1.34 w=1 l=0.15
X7 a_297_297# a_109_93# a_215_53# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X8 a_109_93# C_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X9 X a_215_53# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.179 pd=1.85 as=0.1 ps=0.985 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__clkbuf_16 VGND VPWR A X VPB VNB
X0 VPWR A a_110_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X6 a_110_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X7 a_110_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X8 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X9 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X10 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X11 a_110_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X12 VGND A a_110_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X13 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0578 pd=0.695 as=0.0588 ps=0.7 w=0.42 l=0.15
X14 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X15 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X16 VGND A a_110_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X17 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X18 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.138 pd=1.27 as=0.14 ps=1.28 w=1 l=0.15
X19 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X20 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.138 ps=1.27 w=1 l=0.15
X21 a_110_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.111 ps=1.37 w=0.42 l=0.15
X22 VPWR A a_110_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X23 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X24 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X25 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X26 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X27 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X28 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X29 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X30 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X31 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X32 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X33 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X34 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X35 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X36 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X37 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X38 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X39 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0578 ps=0.695 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__nand3b_1 VGND VPWR Y B C A_N VPB VNB
X0 Y a_53_93# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.192 ps=1.38 w=1 l=0.15
X1 a_232_47# C VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.1 ps=0.985 w=0.65 l=0.15
X2 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.192 pd=1.38 as=0.135 ps=1.27 w=1 l=0.15
X3 VPWR A_N a_53_93# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.146 pd=1.34 as=0.109 ps=1.36 w=0.42 l=0.15
X4 VGND A_N a_53_93# VNB sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.985 as=0.109 ps=1.36 w=0.42 l=0.15
X5 a_316_47# B a_232_47# VNB sky130_fd_pr__nfet_01v8 ad=0.125 pd=1.03 as=0.0878 ps=0.92 w=0.65 l=0.15
X6 Y a_53_93# a_316_47# VNB sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.125 ps=1.03 w=0.65 l=0.15
X7 Y C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.146 ps=1.34 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__a21boi_2 VPWR VGND B1_N A2 Y A1 VPB VNB
X0 Y a_61_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.183 ps=1.24 w=0.65 l=0.15
X1 VPWR A2 a_217_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2 a_217_297# a_61_47# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 a_479_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.86 as=0.107 ps=0.98 w=0.65 l=0.15
X4 a_217_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.285 pd=2.57 as=0.14 ps=1.28 w=1 l=0.15
X5 Y a_61_47# a_217_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6 VPWR A1 a_217_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X7 a_61_47# B1_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.111 ps=1.37 w=0.42 l=0.15
X8 VGND A2 a_637_47# VNB sky130_fd_pr__nfet_01v8 ad=0.185 pd=1.87 as=0.091 ps=0.93 w=0.65 l=0.15
X9 VGND a_61_47# Y VNB sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.0878 ps=0.92 w=0.65 l=0.15
X10 Y A1 a_479_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.0683 ps=0.86 w=0.65 l=0.15
X11 VGND B1_N a_61_47# VNB sky130_fd_pr__nfet_01v8 ad=0.183 pd=1.24 as=0.126 ps=1.44 w=0.42 l=0.15
X12 a_217_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.135 ps=1.27 w=1 l=0.15
X13 a_637_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__a21bo_1 VGND VPWR X A2 A1 B1_N VPB VNB
X0 a_298_297# a_27_413# a_215_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X1 a_215_297# a_27_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.136 ps=1.1 w=0.65 l=0.15
X2 a_298_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X3 X a_215_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.258 ps=1.45 w=0.65 l=0.15
X4 VPWR B1_N a_27_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X5 X a_215_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X6 a_382_47# A1 a_215_297# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.0878 ps=0.92 w=0.65 l=0.15
X7 VGND B1_N a_27_413# VNB sky130_fd_pr__nfet_01v8 ad=0.136 pd=1.1 as=0.111 ps=1.37 w=0.42 l=0.15
X8 VPWR A1 a_298_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.135 ps=1.27 w=1 l=0.15
X9 VGND A2 a_382_47# VNB sky130_fd_pr__nfet_01v8 ad=0.258 pd=1.45 as=0.091 ps=0.93 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__o22a_1 VGND VPWR B2 A2 A1 B1 X VPB VNB
X0 a_78_199# B1 a_215_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1 VPWR A1 a_493_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X2 a_493_297# A2 a_78_199# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.235 ps=1.47 w=1 l=0.15
X3 VPWR a_78_199# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.373 pd=1.75 as=0.28 ps=2.56 w=1 l=0.15
X4 VGND A2 a_215_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.114 ps=1 w=0.65 l=0.15
X5 a_78_199# B2 a_292_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.235 pd=1.47 as=0.117 ps=1.24 w=1 l=0.15
X6 a_215_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7 a_215_47# B2 a_78_199# VNB sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.0878 ps=0.92 w=0.65 l=0.15
X8 a_292_297# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.117 pd=1.24 as=0.373 ps=1.75 w=1 l=0.15
X9 VGND a_78_199# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__conb_1 VGND VPWR LO HI VPB VNB
R0 VPWR HI sky130_fd_pr__res_generic_po w=0.48 l=0.045
R1 LO VGND sky130_fd_pr__res_generic_po w=0.48 l=0.045
.ends

.subckt sky130_fd_sc_hd__nor2_4 VGND VPWR Y B A VPB VNB
X0 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4 a_27_297# B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X5 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X6 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X7 VGND B Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X8 VGND B Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X9 Y B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X10 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X11 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X12 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X13 a_27_297# B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X14 Y B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X15 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__a221oi_1 VGND VPWR Y B1 C1 A1 A2 B2 VPB VNB
X0 a_465_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.0991 pd=0.955 as=0.169 ps=1.82 w=0.65 l=0.15
X1 a_109_297# B1 a_193_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2 a_193_297# B2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 a_204_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0699 pd=0.865 as=0.106 ps=0.975 w=0.65 l=0.15
X4 VGND A2 a_465_47# VNB sky130_fd_pr__nfet_01v8 ad=0.198 pd=1.91 as=0.0991 ps=0.955 w=0.65 l=0.15
X5 a_193_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.153 pd=1.3 as=0.26 ps=2.52 w=1 l=0.15
X6 Y B1 a_204_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0699 ps=0.865 w=0.65 l=0.15
X7 VPWR A2 a_193_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.305 pd=2.61 as=0.153 ps=1.3 w=1 l=0.15
X8 a_109_297# C1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X9 VGND C1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.106 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__clkinv_4 VPWR VGND A Y VPB VNB
X0 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.63 as=0.0588 ps=0.7 w=0.42 l=0.15
X2 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.345 pd=2.69 as=0.14 ps=1.28 w=1 l=0.15
X5 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X6 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.305 ps=2.61 w=1 l=0.15
X7 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.139 ps=1.5 w=0.42 l=0.15
X8 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X9 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__buf_1 VGND VPWR X A VPB VNB
X0 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X1 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X2 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X3 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
.ends

.subckt adc_array_matrix_12bit row_n[0] row_n[1] row_n[2] row_n[3] row_n[4] row_n[5]
+ row_n[6] row_n[7] row_n[8] row_n[9] row_n[10] row_n[11] row_n[12] row_n[13] row_n[14]
+ row_n[15] rowon_n[0] rowon_n[1] rowon_n[2] rowon_n[3] rowon_n[4] rowon_n[5] rowon_n[6]
+ rowon_n[7] rowon_n[8] rowon_n[9] rowon_n[10] rowon_n[11] rowon_n[12] rowon_n[13]
+ rowon_n[14] rowon_n[15] rowoff_n[0] rowoff_n[1] rowoff_n[2] rowoff_n[3] rowoff_n[4]
+ rowoff_n[5] rowoff_n[6] rowoff_n[7] rowoff_n[8] rowoff_n[9] rowoff_n[10] rowoff_n[11]
+ rowoff_n[12] rowoff_n[13] rowoff_n[14] rowoff_n[15] vcm sample sample_n col_n[31]
+ col_n[30] col_n[29] col_n[28] col_n[27] col_n[26] col_n[25] col_n[24] col_n[23]
+ col_n[22] col_n[21] col_n[20] col_n[19] col_n[18] col_n[17] col_n[16] col_n[15]
+ col_n[14] col_n[13] col_n[12] col_n[11] col_n[10] col_n[9] col_n[8] col_n[7] col_n[6]
+ col_n[5] col_n[4] col_n[3] col_n[2] col_n[1] col_n[0] en_bit_n[2] en_bit_n[1] en_bit_n[0]
+ en_C0_n sw sw_n analog_in col[0] col[1] col[2] col[3] col[4] col[5] col[6] col[7]
+ col[8] col[9] col[10] col[11] col[12] col[13] col[14] col[15] col[16] col[17] col[18]
+ col[19] col[20] col[21] col[22] col[23] col[24] col[25] col[26] col[27] col[28]
+ col[29] col[30] col[31] VDD VSS ctop
X0 a_3970_15182# a_2475_15206# a_3878_15182# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X1 a_3878_9158# a_2275_9182# a_3970_9158# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2 VDD rowon_n[5] a_18938_7150# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3 a_30986_7150# row_n[5] a_31478_7512# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4 vcm a_2275_18218# a_32082_18194# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5 a_12002_2130# a_2475_2154# a_11910_2130# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X6 a_5374_4500# col_n[2] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X7 a_14410_15544# col_n[11] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X8 a_10906_12170# row_n[10] a_11398_12532# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X9 a_35398_9198# VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X10 a_17422_7512# col_n[14] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X11 a_18026_7150# a_2475_7174# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X12 VSS row_n[4] a_9294_6186# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X13 a_4370_15544# col_n[1] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X14 a_23046_11166# a_2475_11190# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X15 a_22346_10202# rowon_n[8] a_21950_10162# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X16 a_14922_11166# row_n[9] a_15414_11528# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X17 a_15414_2492# col_n[12] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X18 a_4882_11166# row_n[9] a_5374_11528# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X19 a_34394_2170# col_n[31] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X20 a_27062_12170# a_2475_12194# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X21 VSS row_n[6] a_26362_8194# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X22 a_1957_14202# VSS sample VDD sky130_fd_pr__pfet_01v8 ad=0.342 pd=2.97 as=0.342 ps=2.97 w=1.2 l=0.15
X23 a_34090_3134# a_2475_3158# a_33998_3134# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X24 a_1957_4162# VDD sample VSS sky130_fd_pr__nfet_01v8 ad=0.171 pd=1.77 as=0.171 ps=1.77 w=0.6 l=0.15
X25 a_26058_18194# a_2475_18218# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X26 a_21342_2170# rowon_n[0] a_20946_2130# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X27 a_35002_9158# row_n[7] a_35494_9520# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X28 a_23350_18234# VDD a_22954_18194# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X29 VSS row_n[13] a_20338_15222# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X30 a_26970_14178# a_2275_14202# a_27062_14178# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X31 a_11302_8194# rowon_n[6] a_10906_8154# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X32 a_29982_4138# a_2275_4162# a_30074_4138# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X33 a_12306_4178# rowon_n[2] a_11910_4138# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X34 vcm a_2275_2154# a_13006_2130# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X35 VDD rowon_n[3] a_22954_5142# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X36 VSS row_n[12] a_24354_14218# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X37 a_21342_11206# col_n[18] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X38 a_34394_10202# col_n[31] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X39 a_24962_17190# a_2275_17214# a_25054_17190# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X40 a_18938_7150# a_2275_7174# a_19030_7150# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X41 a_4274_13214# rowon_n[11] a_3878_13174# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X42 a_14314_13214# rowon_n[11] a_13918_13174# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X43 VSS row_n[8] a_11302_10202# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X44 a_20034_7150# a_2475_7174# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X45 a_21038_3134# a_2475_3158# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X46 a_19430_18556# col_n[16] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X47 a_19030_14178# a_2475_14202# a_18938_14178# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X48 a_11910_11166# a_2275_11190# a_12002_11166# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X49 VDD VSS VSS sky130_fd_pr__cap_var_lvt w=16.4 l=16
X50 VDD rowon_n[14] a_22954_16186# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X51 a_28978_14178# row_n[12] a_29470_14540# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X52 a_20434_13536# col_n[17] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X53 a_33486_12532# col_n[30] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X54 vcm a_2275_10186# a_29070_10162# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X55 a_20338_6186# col_n[17] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X56 a_15926_12170# a_2275_12194# a_16018_12170# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X57 a_3270_7190# rowon_n[5] a_2874_7150# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X58 VSS row_n[4] a_30378_6186# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X59 a_4274_3174# rowon_n[1] a_3878_3134# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X60 VDD rowon_n[2] a_11910_4138# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X61 a_5886_12170# a_2275_12194# a_5978_12170# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X62 VDD rowon_n[10] a_9902_12170# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X63 a_16322_6186# rowon_n[4] a_15926_6146# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X64 vcm a_2275_6170# a_24050_6146# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X65 a_35398_18234# VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X66 VDD rowon_n[9] a_3878_11166# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X67 VDD rowon_n[9] a_13918_11166# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X68 VDD rowon_n[4] a_5886_6146# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X69 VSS VDD a_12306_18234# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X70 a_30074_17190# a_2475_17214# a_29982_17190# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X71 a_16018_7150# a_2475_7174# a_15926_7150# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X72 a_26058_1126# a_2475_1150# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X73 a_25054_5142# a_2475_5166# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X74 a_13310_14218# col_n[10] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X75 VDD en_C0_n a_3878_1126# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X76 a_30986_17190# row_n[15] a_31478_17552# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X77 a_12002_16186# a_2475_16210# a_11910_16186# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X78 a_34090_16186# a_2475_16210# a_33998_16186# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X79 a_3270_14218# col_n[0] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X80 vcm a_2275_13198# a_31078_13174# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X81 a_25358_4178# col_n[22] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X82 a_35002_16186# row_n[14] a_35494_16548# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X83 a_10906_8154# row_n[6] a_11398_8516# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X84 VSS row_n[6] a_34394_8194# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X85 a_8290_5182# rowon_n[3] a_7894_5142# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X86 a_9294_1166# VSS a_8898_1126# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X87 VSS row_n[2] a_35398_4178# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X88 a_9994_9158# a_2475_9182# a_9902_9158# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X89 a_12402_16548# col_n[9] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X90 a_19334_16226# rowon_n[14] a_18938_16186# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X91 a_20338_11206# rowon_n[9] a_19942_11166# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X92 vcm a_2275_8178# a_28066_8154# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X93 vcm a_2275_4162# a_29070_4138# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X94 VSS a_2161_13198# a_2275_13198# VSS sky130_fd_pr__nfet_01v8 ad=0.124 pd=1.01 as=0.171 ps=1.77 w=0.6 l=0.15
X95 a_25358_7190# rowon_n[5] a_24962_7150# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X96 a_25054_13174# a_2475_13198# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X97 a_13310_7190# col_n[10] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X98 a_29070_7150# a_2475_7174# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X99 a_14314_3174# col_n[11] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X100 a_16018_12170# a_2475_12194# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X101 a_33998_9158# a_2275_9182# a_34090_9158# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X102 VDD rowon_n[1] a_7894_3134# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X103 a_24962_4138# row_n[2] a_25454_4500# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X104 a_5978_12170# a_2475_12194# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X105 a_2874_7150# row_n[5] a_3366_7512# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X106 vcm a_2275_7174# a_17022_7150# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X107 a_35494_4500# VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X108 a_19942_11166# a_2275_11190# a_20034_11166# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X109 a_32994_10162# a_2275_10186# a_33086_10162# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X110 a_15926_6146# row_n[4] a_16418_6508# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X111 a_34394_18234# VDD a_33998_18194# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X112 a_27366_17230# col_n[24] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X113 VSS row_n[13] a_31382_15222# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X114 a_13918_1126# VDD a_14410_1488# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X115 VSS row_n[12] a_35398_14218# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X116 a_32386_11206# col_n[29] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X117 a_6282_2170# col_n[3] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X118 a_22954_18194# a_2275_18218# a_23046_18194# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X119 a_12306_14218# rowon_n[12] a_11910_14178# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X120 a_18330_5182# col_n[15] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X121 a_19334_1166# en_bit_n[2] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X122 VDD VSS sky130_fd_pr__cap_mim_m3_1 l=17.2 w=17.2
X123 VDD rowon_n[15] a_29982_17190# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X124 a_26058_15182# a_2475_15206# a_25966_15182# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X125 VSS en_bit_n[0] a_20338_1166# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X126 vcm a_2275_11190# a_27062_11166# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X127 a_7894_5142# row_n[3] a_8386_5504# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X128 a_30378_1166# VSS a_29982_1126# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X129 VDD rowon_n[14] a_33998_16186# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X130 a_26970_15182# row_n[13] a_27462_15544# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X131 a_31478_13536# col_n[28] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X132 a_3878_13174# a_2275_13198# a_3970_13174# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X133 a_13918_13174# a_2275_13198# a_14010_13174# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X134 a_23046_5142# a_2475_5166# a_22954_5142# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X135 VDD rowon_n[6] a_30986_8154# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X136 a_17934_3134# row_n[1] a_18426_3496# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X137 a_29374_9198# col_n[26] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X138 a_29982_12170# row_n[10] a_30474_12532# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X139 VSS row_n[1] a_24354_3174# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X140 a_10394_7512# col_n[7] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X141 a_33390_7190# rowon_n[5] a_32994_7150# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X142 a_34394_3174# rowon_n[1] a_33998_3134# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X143 a_18330_11206# rowon_n[9] a_17934_11166# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X144 a_10998_7150# a_2475_7174# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X145 VSS row_n[7] a_14314_9198# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X146 a_27062_7150# a_2475_7174# a_26970_7150# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X147 a_28066_3134# a_2475_3158# a_27974_3134# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X148 vcm a_2275_9182# a_32082_9158# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X149 a_18938_18194# VDD a_19430_18556# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X150 vcm a_2275_14202# a_8990_14178# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X151 vcm a_2275_14202# a_19030_14178# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X152 a_4974_9158# a_2475_9182# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X153 a_28978_9158# row_n[7] a_29470_9520# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X154 a_8898_18194# VDD a_9390_18556# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X155 a_22954_8154# a_2275_8178# a_23046_8154# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X156 a_24450_1488# col_n[21] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X157 a_19030_2130# a_2475_2154# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X158 VSS row_n[0] a_13310_2170# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X159 a_23958_4138# a_2275_4162# a_24050_4138# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X160 a_33086_8154# a_2475_8178# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X161 a_23046_14178# a_2475_14202# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X162 VSS VDD a_29374_1166# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X163 a_14410_9520# col_n[11] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X164 a_15414_5504# col_n[12] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X165 VSS row_n[13] a_29374_15222# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X166 a_33390_13214# rowon_n[11] a_32994_13174# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X167 a_26362_12210# col_n[23] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X168 VSS row_n[8] a_30378_10202# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X169 a_16018_5142# a_2475_5166# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X170 VSS row_n[2] a_7286_4178# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X171 a_30986_11166# a_2275_11190# a_31078_11166# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X172 a_11910_7150# a_2275_7174# a_12002_7150# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X173 VDD rowon_n[15] a_27974_17190# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X174 a_25454_14540# col_n[22] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X175 a_35002_12170# a_2275_12194# a_35094_12170# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X176 a_25054_10162# a_2475_10186# a_24962_10162# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X177 a_27974_6146# a_2275_6170# a_28066_6146# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X178 a_32082_1126# a_2475_1150# a_31990_1126# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X179 a_5886_9158# a_2275_9182# a_5978_9158# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X180 a_33998_18194# a_2275_18218# a_34090_18194# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X181 a_29470_13536# col_n[26] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X182 VDD rowon_n[9] a_32994_11166# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X183 a_25966_10162# row_n[8] a_26458_10524# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X184 a_32994_7150# row_n[5] a_33486_7512# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X185 a_7382_4500# col_n[4] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X186 a_14010_2130# a_2475_2154# a_13918_2130# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X187 a_30986_2130# row_n[0] a_31478_2492# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X188 VDD rowon_n[0] a_18938_2130# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X189 a_11910_14178# a_2275_14202# a_12002_14178# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X190 VDD rowon_n[10] a_8898_12170# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X191 a_16930_5142# a_2275_5166# a_17022_5142# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X192 a_17422_2492# col_n[14] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X193 vcm a_2275_15206# a_23046_15182# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X194 VSS row_n[6] a_28370_8194# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X195 a_17022_17190# a_2475_17214# a_16930_17190# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X196 a_8290_15222# col_n[5] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X197 a_18330_15222# col_n[15] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X198 a_6982_17190# a_2475_17214# a_6890_17190# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X199 a_9902_17190# a_2275_17214# a_9994_17190# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X200 a_1957_8178# VSS sample VDD sky130_fd_pr__pfet_01v8 ad=0.342 pd=2.97 as=0.342 ps=2.97 w=1.2 l=0.15
X201 a_23350_2170# rowon_n[0] a_22954_2130# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X202 vcm a_2275_10186# a_14010_10162# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X203 a_2966_9158# a_2475_9182# a_2874_9158# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X204 a_2161_6170# sample VSS VSS sky130_fd_pr__nfet_01v8 ad=0.171 pd=1.77 as=0.171 ps=1.77 w=0.6 l=0.15
X205 a_7382_17552# col_n[4] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X206 a_17422_17552# col_n[14] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X207 a_3878_14178# row_n[12] a_4370_14540# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X208 a_13918_14178# row_n[12] a_14410_14540# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X209 a_25358_12210# rowon_n[10] a_24962_12170# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X210 vcm a_2275_10186# a_3970_10162# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X211 a_13310_8194# rowon_n[6] a_12914_8154# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X212 vcm a_2275_8178# a_21038_8154# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X213 vcm a_2275_4162# a_22042_4138# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X214 a_14314_4178# rowon_n[2] a_13918_4138# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X215 a_17934_13174# row_n[11] a_18426_13536# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X216 a_29374_11206# rowon_n[9] a_28978_11166# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X217 a_31078_8154# a_2475_8178# a_30986_8154# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X218 vcm a_2275_2154# a_15014_2130# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X219 a_7894_13174# row_n[11] a_8386_13536# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X220 VDD rowon_n[6] a_2874_8154# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X221 a_23046_3134# a_2475_3158# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X222 a_22042_7150# a_2475_7174# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X223 VDD rowon_n[8] a_24962_10162# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X224 VDD rowon_n[2] a_13918_4138# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X225 vcm a_2275_18218# a_4974_18194# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X226 vcm a_2275_18218# a_15014_18194# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X227 VSS row_n[15] a_23350_17230# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X228 VSS row_n[4] a_32386_6186# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X229 a_6282_3174# rowon_n[1] a_5886_3134# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X230 vcm a_2275_6170# a_26058_6146# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X231 VSS row_n[14] a_27366_16226# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X232 a_31382_14218# rowon_n[12] a_30986_14178# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X233 a_24354_13214# col_n[21] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X234 vcm a_2275_9182# a_3970_9158# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X235 VDD rowon_n[4] a_7894_6146# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X236 a_2475_4162# a_1957_4162# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.171 pd=1.77 as=0.124 ps=1.01 w=0.6 l=0.15
X237 a_32082_17190# a_2475_17214# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X238 a_17326_15222# rowon_n[13] a_16930_15182# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X239 a_11302_5182# col_n[8] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X240 a_12306_1166# col_n[9] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X241 a_28066_1126# a_2475_1150# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X242 a_7286_15222# rowon_n[13] a_6890_15182# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X243 a_19942_14178# a_2275_14202# a_20034_14178# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X244 a_32994_13174# a_2275_13198# a_33086_13174# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X245 a_18026_7150# a_2475_7174# a_17934_7150# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X246 a_27062_5142# a_2475_5166# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X247 VDD VDD a_25966_18194# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X248 a_3970_16186# a_2475_16210# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X249 a_14010_16186# a_2475_16210# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X250 a_23446_15544# col_n[20] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X251 VSS row_n[9] a_8290_11206# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X252 VSS row_n[9] a_18330_11206# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X253 a_23046_11166# a_2475_11190# a_22954_11166# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X254 VDD VSS a_5886_1126# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X255 a_23958_11166# row_n[9] a_24450_11528# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X256 a_12914_8154# row_n[6] a_13406_8516# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X257 VDD rowon_n[6] a_24962_8154# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X258 VDD rowon_n[11] a_6890_13174# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X259 VDD rowon_n[11] a_16930_13174# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X260 a_10906_3134# row_n[1] a_11398_3496# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X261 a_12306_17230# col_n[9] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X262 a_22346_9198# col_n[19] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X263 a_27366_7190# rowon_n[5] a_26970_7150# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X264 a_16322_3174# col_n[13] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X265 vcm a_2275_4162# a_30074_4138# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X266 a_16322_16226# col_n[13] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X267 vcm a_2275_16210# a_21038_16186# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X268 a_15318_7190# col_n[12] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X269 a_15014_18194# a_2475_18218# a_14922_18194# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X270 a_6282_16226# col_n[3] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X271 vcm a_2275_15206# a_34090_15182# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X272 a_4882_7150# row_n[5] a_5374_7512# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X273 a_4974_18194# a_2475_18218# a_4882_18194# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X274 vcm a_2275_7174# a_19030_7150# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X275 a_17934_6146# row_n[4] a_18426_6508# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X276 a_21038_3134# a_2475_3158# a_20946_3134# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X277 a_15414_18556# col_n[12] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X278 a_11910_15182# row_n[13] a_12402_15544# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X279 vcm a_2275_11190# a_12002_11166# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X280 a_20034_7150# a_2475_7174# a_19942_7150# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X281 a_2874_2130# row_n[0] a_3366_2492# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X282 a_5374_18556# col_n[2] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X283 a_21950_9158# row_n[7] a_22442_9520# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X284 a_15926_1126# VDD a_16418_1488# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X285 a_8290_2170# col_n[5] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X286 a_28066_15182# a_2475_15206# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X287 a_9902_2130# a_2275_2154# a_9994_2130# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X288 VSS row_n[10] a_22346_12210# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X289 VSS VDD a_22346_1166# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X290 a_32386_1166# VSS a_31990_1126# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X291 a_31382_5182# rowon_n[3] a_30986_5142# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X292 a_26058_1126# a_2475_1150# a_25966_1126# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X293 VSS VDD a_21342_18234# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X294 a_25054_5142# a_2475_5166# a_24962_5142# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X295 VDD rowon_n[12] a_20946_14178# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X296 a_22346_14218# col_n[19] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X297 a_16322_10202# rowon_n[8] a_15926_10162# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X298 VDD rowon_n[6] a_32994_8154# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X299 a_26970_7150# row_n[5] a_27462_7512# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X300 a_6282_10202# rowon_n[8] a_5886_10162# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X301 a_30074_18194# a_2475_18218# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X302 a_22442_10524# col_n[19] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X303 a_20946_6146# a_2275_6170# a_21038_6146# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X304 a_5278_16226# rowon_n[14] a_4882_16186# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X305 a_15318_16226# rowon_n[14] a_14922_16186# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X306 a_31078_6146# a_2475_6170# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X307 VDD rowon_n[1] a_30986_3134# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X308 a_20338_17230# col_n[17] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X309 a_21438_16548# col_n[18] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X310 a_30986_14178# a_2275_14202# a_31078_14178# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X311 a_18330_9198# rowon_n[7] a_17934_9158# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X312 a_30378_9198# col_n[27] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X313 a_12402_7512# col_n[9] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X314 a_13006_7150# a_2475_7174# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X315 VSS row_n[4] a_4274_6186# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X316 a_6890_15182# a_2275_15206# a_6982_15182# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X317 a_16930_15182# a_2275_15206# a_17022_15182# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X318 vcm a_2275_9182# a_34090_9158# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X319 a_29070_7150# a_2475_7174# a_28978_7150# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X320 a_10394_2492# col_n[7] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X321 VSS row_n[13] a_4274_15222# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X322 VSS row_n[13] a_14314_15222# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X323 a_11302_12210# col_n[8] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X324 a_19942_15182# row_n[13] a_20434_15544# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X325 a_15318_11206# col_n[12] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X326 vcm a_2275_11190# a_20034_11166# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X327 a_6982_9158# a_2475_9182# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X328 VSS row_n[6] a_21342_8194# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X329 VDD VSS sky130_fd_pr__cap_mim_m3_1 l=17.2 w=17.2
X330 a_32994_14178# row_n[12] a_33486_14540# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X331 a_14010_13174# a_2475_13198# a_13918_13174# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X332 a_5278_11206# col_n[2] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X333 vcm a_2275_10186# a_33086_10162# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X334 a_24962_8154# a_2275_8178# a_25054_8154# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X335 VSS row_n[0] a_15318_2170# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X336 a_25966_4138# a_2275_4162# a_26058_4138# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X337 a_3970_13174# a_2475_13198# a_3878_13174# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X338 VDD rowon_n[7] a_17934_9158# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X339 a_29982_9158# row_n[7] a_30474_9520# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X340 a_35094_8154# a_2475_8178# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X341 VDD rowon_n[3] a_18938_5142# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X342 a_30986_5142# row_n[3] a_31478_5504# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X343 VDD rowon_n[15] a_2874_17190# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X344 VDD rowon_n[15] a_12914_17190# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X345 vcm a_2275_16210# a_32082_16186# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X346 a_10394_14540# col_n[7] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X347 a_5978_2130# a_2475_2154# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X348 a_14410_13536# col_n[11] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X349 a_10906_10162# row_n[8] a_11398_10524# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X350 a_17422_5504# col_n[14] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X351 a_18026_5142# a_2475_5166# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X352 VSS row_n[2] a_9294_4178# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X353 a_4370_13536# col_n[1] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X354 VDD a_2161_7174# a_2275_7174# VDD sky130_fd_pr__pfet_01v8 ad=0.249 pd=1.62 as=0.342 ps=2.97 w=1.2 l=0.15
X355 a_13918_7150# a_2275_7174# a_14010_7150# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X356 VSS row_n[4] a_26362_6186# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X357 a_1957_2154# VDD sample VSS sky130_fd_pr__nfet_01v8 ad=0.171 pd=1.77 as=0.171 ps=1.77 w=0.6 l=0.15
X358 a_26058_16186# a_2475_16210# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X359 a_7894_9158# a_2275_9182# a_7986_9158# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X360 a_35002_7150# row_n[5] a_35494_7512# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X361 a_9390_4500# col_n[6] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X362 VSS VDD a_19334_18234# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X363 a_23350_16226# rowon_n[14] a_22954_16186# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X364 VSS row_n[11] a_20338_13214# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X365 a_11302_6186# rowon_n[4] a_10906_6146# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X366 VSS row_n[10] a_33390_12210# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X367 a_32994_2130# row_n[0] a_33486_2492# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X368 a_6890_2130# a_2275_2154# a_6982_2130# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X369 a_10298_12210# rowon_n[10] a_9902_12170# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X370 a_24962_15182# a_2275_15206# a_25054_15182# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X371 a_18938_5142# a_2275_5166# a_19030_5142# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X372 a_28066_12170# a_2475_12194# a_27974_12170# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X373 a_4274_11206# rowon_n[9] a_3878_11166# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X374 a_14314_11206# rowon_n[9] a_13918_11166# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X375 a_10998_7150# a_2475_7174# a_10906_7150# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X376 a_21038_1126# a_2475_1150# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X377 a_20034_5142# a_2475_5166# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X378 a_8990_17190# a_2475_17214# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X379 a_19430_16548# col_n[16] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X380 VDD rowon_n[12] a_31990_14178# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X381 a_28978_12170# row_n[10] a_29470_12532# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X382 a_20434_11528# col_n[17] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X383 a_33486_10524# col_n[30] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X384 a_20338_4178# col_n[17] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X385 a_3270_5182# rowon_n[3] a_2874_5142# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X386 a_4274_1166# en_C0_n a_3878_1126# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X387 VSS row_n[2] a_30378_4178# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X388 a_31382_17230# col_n[28] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X389 VDD rowon_n[8] a_9902_10162# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X390 a_4974_9158# a_2475_9182# a_4882_9158# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X391 a_19030_2130# a_2475_2154# a_18938_2130# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X392 a_16322_4178# rowon_n[2] a_15926_4138# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X393 vcm a_2275_8178# a_23046_8154# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X394 vcm a_2275_4162# a_24050_4138# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X395 a_35398_16226# VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X396 a_33086_8154# a_2475_8178# a_32994_8154# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X397 VSS row_n[14] a_12306_16226# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X398 a_20338_7190# rowon_n[5] a_19942_7150# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X399 vcm a_2275_17214# a_26058_17190# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X400 a_30074_15182# a_2475_15206# a_29982_15182# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X401 a_24050_7150# a_2475_7174# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X402 a_16018_5142# a_2475_5166# a_15926_5142# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X403 a_25054_3134# a_2475_3158# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X404 a_34090_14178# a_2475_14202# a_33998_14178# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X405 VDD rowon_n[1] a_2874_3134# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X406 a_19942_4138# row_n[2] a_20434_4500# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X407 a_34490_18556# col_n[31] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X408 a_30986_15182# row_n[13] a_31478_15544# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X409 a_12002_14178# a_2475_14202# a_11910_14178# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X410 vcm a_2275_11190# a_31078_11166# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X411 vcm a_2275_7174# a_12002_7150# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X412 a_30474_4500# col_n[27] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X413 VDD VDD a_10906_18194# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X414 vcm a_2275_12194# a_17022_12170# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X415 a_10906_6146# row_n[4] a_11398_6508# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X416 VSS row_n[4] a_34394_6186# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X417 a_8290_3174# rowon_n[1] a_7894_3134# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X418 VDD rowon_n[2] a_15926_4138# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X419 vcm a_2275_12194# a_6982_12170# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X420 a_19334_14218# rowon_n[12] a_18938_14178# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X421 vcm a_2275_6170# a_28066_6146# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X422 vcm a_2275_9182# a_5978_9158# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X423 a_21038_12170# a_2475_12194# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X424 a_2475_8178# a_1957_8178# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.342 pd=2.97 as=0.249 ps=1.62 w=1.2 l=0.15
X425 a_25358_5182# rowon_n[3] a_24962_5142# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X426 a_13310_5182# col_n[10] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X427 a_14314_1166# col_n[11] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X428 a_29070_5142# a_2475_5166# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X429 VDD VSS a_7894_1126# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X430 VDD rowon_n[6] a_26970_8154# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X431 a_2874_5142# row_n[3] a_3366_5504# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X432 vcm a_2275_5166# a_17022_5142# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X433 a_30378_17230# rowon_n[15] a_29982_17190# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X434 a_14922_8154# row_n[6] a_15414_8516# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X435 a_3970_11166# a_2475_11190# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X436 a_14010_11166# a_2475_11190# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X437 a_34394_16226# rowon_n[14] a_33998_16186# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X438 a_27366_15222# col_n[24] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X439 VSS row_n[11] a_31382_13214# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X440 VDD rowon_n[1] a_24962_3134# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X441 a_12914_3134# row_n[1] a_13406_3496# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X442 a_24354_9198# col_n[21] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X443 VSS row_n[5] a_19334_7190# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X444 a_29374_7190# rowon_n[5] a_28978_7150# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X445 a_22954_16186# a_2275_16210# a_23046_16186# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X446 a_18330_3174# col_n[15] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X447 a_6982_18194# a_2475_18218# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X448 a_17022_18194# a_2475_18218# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X449 a_26458_17552# col_n[23] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X450 VDD rowon_n[13] a_29982_15182# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X451 a_26058_13174# a_2475_13198# a_25966_13174# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X452 VDD VSS VSS sky130_fd_pr__cap_var_lvt w=16.4 l=16
X453 a_30378_12210# col_n[27] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X454 a_26970_13174# row_n[11] a_27462_13536# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X455 a_31478_11528# col_n[28] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X456 a_22042_7150# a_2475_7174# a_21950_7150# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X457 a_23046_3134# a_2475_3158# a_22954_3134# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X458 VDD rowon_n[4] a_30986_6146# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X459 a_4882_2130# row_n[0] a_5374_2492# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X460 vcm a_2275_12194# a_25054_12170# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X461 a_23958_9158# row_n[7] a_24450_9520# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X462 a_17934_1126# en_bit_n[1] a_18426_1488# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X463 a_19334_18234# col_n[16] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X464 vcm a_2275_18218# a_24050_18194# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X465 a_29982_10162# row_n[8] a_30474_10524# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X466 a_9294_18234# col_n[6] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X467 VSS VDD a_24354_1166# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X468 a_9390_14540# col_n[6] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X469 a_10394_5504# col_n[7] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X470 a_33390_5182# rowon_n[3] a_32994_5142# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X471 a_28066_10162# a_2475_10186# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X472 a_10998_5142# a_2475_5166# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X473 a_28066_1126# a_2475_1150# a_27974_1126# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X474 a_27062_5142# a_2475_5166# a_26970_5142# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X475 a_19030_12170# a_2475_12194# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X476 a_18938_16186# row_n[14] a_19430_16548# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X477 a_28978_7150# row_n[5] a_29470_7512# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X478 a_8898_16186# row_n[14] a_9390_16548# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X479 a_22954_6146# a_2275_6170# a_23046_6146# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X480 a_33086_6146# a_2475_6170# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X481 a_26970_2130# row_n[0] a_27462_2492# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X482 VDD rowon_n[1] a_32994_3134# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X483 a_28370_17230# rowon_n[15] a_27974_17190# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X484 a_14410_7512# col_n[11] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X485 VSS row_n[11] a_29374_13214# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X486 a_33390_11206# rowon_n[9] a_32994_11166# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X487 a_26362_10202# col_n[23] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X488 a_15014_7150# a_2475_7174# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X489 VSS a_2161_1150# a_2275_1150# VSS sky130_fd_pr__nfet_01v8 ad=0.124 pd=1.01 as=0.171 ps=1.77 w=0.6 l=0.15
X490 a_16018_3134# a_2475_3158# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X491 a_11910_5142# a_2275_5166# a_12002_5142# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X492 a_12402_2492# col_n[9] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X493 a_9294_12210# rowon_n[10] a_8898_12170# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X494 a_16930_10162# a_2275_10186# a_17022_10162# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X495 a_8990_9158# a_2475_9182# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X496 VSS row_n[6] a_23350_8194# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X497 a_31382_2170# col_n[28] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X498 a_19334_2170# rowon_n[0] a_18938_2130# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X499 VDD rowon_n[13] a_27974_15182# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X500 a_25454_12532# col_n[22] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X501 a_6890_10162# a_2275_10186# a_6982_10162# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X502 VSS row_n[0] a_17326_2170# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X503 a_27974_4138# a_2275_4162# a_28066_4138# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X504 a_33998_16186# a_2275_16210# a_34090_16186# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X505 a_29470_11528# col_n[26] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X506 a_32994_5142# row_n[3] a_33486_5504# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X507 a_7986_2130# a_2475_2154# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X508 VDD rowon_n[8] a_8898_10162# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X509 vcm a_2275_2154# a_9994_2130# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X510 VSS row_n[15] a_7286_17230# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X511 VSS row_n[15] a_17326_17230# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X512 a_22042_17190# a_2475_17214# a_21950_17190# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X513 a_15926_7150# a_2275_7174# a_16018_7150# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X514 a_16930_3134# a_2275_3158# a_17022_3134# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X515 a_18330_13214# col_n[15] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X516 vcm a_2275_13198# a_23046_13174# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X517 VSS row_n[4] a_28370_6186# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X518 a_22954_17190# row_n[15] a_23446_17552# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X519 a_17022_15182# a_2475_15206# a_16930_15182# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X520 a_8290_13214# col_n[5] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X521 VSS row_n[7] a_6282_9198# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X522 a_6982_15182# a_2475_15206# a_6890_15182# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X523 a_9902_15182# a_2275_15206# a_9994_15182# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X524 a_1957_6170# VSS sample VDD sky130_fd_pr__pfet_01v8 ad=0.342 pd=2.97 as=0.342 ps=2.97 w=1.2 l=0.15
X525 a_17422_15544# col_n[14] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X526 a_2161_4162# sample VSS VSS sky130_fd_pr__nfet_01v8 ad=0.171 pd=1.77 as=0.171 ps=1.77 w=0.6 l=0.15
X527 a_7382_15544# col_n[4] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X528 a_3878_12170# row_n[10] a_4370_12532# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X529 a_13918_12170# row_n[10] a_14410_12532# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X530 a_26058_11166# a_2475_11190# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X531 a_25358_10202# rowon_n[8] a_24962_10162# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X532 a_13310_6186# rowon_n[4] a_12914_6146# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X533 vcm a_2275_6170# a_21038_6146# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X534 a_17934_11166# row_n[9] a_18426_11528# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X535 a_31078_6146# a_2475_6170# a_30986_6146# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X536 a_35002_2130# row_n[0] a_35494_2492# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X537 a_8898_2130# a_2275_2154# a_8990_2130# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X538 a_7894_11166# row_n[9] a_8386_11528# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X539 VDD rowon_n[4] a_2874_6146# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X540 a_6378_9520# col_n[3] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X541 a_23046_1126# a_2475_1150# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X542 a_13006_7150# a_2475_7174# a_12914_7150# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X543 a_22042_5142# a_2475_5166# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X544 vcm a_2275_17214# a_10998_17190# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X545 a_24962_10162# a_2275_10186# a_25054_10162# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X546 VDD rowon_n[6] a_19942_8154# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X547 a_26362_18234# VDD a_25966_18194# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X548 vcm a_2275_16210# a_4974_16186# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X549 vcm a_2275_16210# a_15014_16186# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X550 VSS row_n[13] a_23350_15222# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X551 a_6982_9158# a_2475_9182# a_6890_9158# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X552 a_6282_1166# VSS a_5886_1126# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X553 VSS row_n[2] a_32386_4178# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X554 vcm a_2275_8178# a_25054_8154# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X555 vcm a_2275_4162# a_26058_4138# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X556 VSS row_n[12] a_27366_14218# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X557 a_24354_11206# col_n[21] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X558 a_35094_8154# a_2475_8178# a_35002_8154# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X559 a_27974_17190# a_2275_17214# a_28066_17190# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X560 a_5978_2130# a_2475_2154# a_5886_2130# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X561 a_2475_2154# a_1957_2154# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.171 pd=1.77 as=0.124 ps=1.01 w=0.6 l=0.15
X562 VDD rowon_n[15] a_21950_17190# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X563 a_32082_15182# a_2475_15206# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X564 a_17326_13214# rowon_n[11] a_16930_13174# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X565 a_22346_7190# rowon_n[5] a_21950_7150# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X566 a_11302_3174# col_n[8] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X567 a_7286_13214# rowon_n[11] a_6890_13174# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X568 a_30986_9158# a_2275_9182# a_31078_9158# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X569 a_10298_7190# col_n[7] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X570 a_18026_5142# a_2475_5166# a_17934_5142# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X571 a_27062_3134# a_2475_3158# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X572 VDD rowon_n[14] a_25966_16186# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X573 a_3970_14178# a_2475_14202# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X574 a_14010_14178# a_2475_14202# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X575 a_23446_13536# col_n[20] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X576 a_32482_4500# col_n[29] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X577 a_18938_12170# a_2275_12194# a_19030_12170# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X578 vcm a_2275_7174# a_14010_7150# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X579 a_12914_6146# row_n[4] a_13406_6508# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X580 VDD rowon_n[4] a_24962_6146# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X581 a_8898_12170# a_2275_12194# a_8990_12170# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X582 VDD rowon_n[9] a_6890_11166# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X583 VDD rowon_n[9] a_16930_11166# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X584 a_10906_1126# VDD a_11398_1488# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X585 VSS VDD a_15318_18234# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X586 a_20034_18194# a_2475_18218# a_19942_18194# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X587 a_12306_15222# col_n[9] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X588 vcm a_2275_9182# a_7986_9158# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X589 a_3270_2170# col_n[0] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X590 VSS VDD a_5278_18234# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X591 a_10998_17190# a_2475_17214# a_10906_17190# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X592 a_33086_17190# a_2475_17214# a_32994_17190# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X593 a_16322_1166# col_n[13] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X594 a_27366_5182# rowon_n[3] a_26970_5142# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X595 a_20946_18194# VDD a_21438_18556# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X596 a_16322_14218# col_n[13] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X597 vcm a_2275_14202# a_21038_14178# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X598 a_5278_8194# rowon_n[6] a_4882_8154# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X599 a_15318_5182# col_n[12] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X600 a_33998_17190# row_n[15] a_34490_17552# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X601 a_15014_16186# a_2475_16210# a_14922_16186# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X602 a_6282_14218# col_n[3] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X603 vcm a_2275_13198# a_34090_13174# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X604 a_19430_8516# col_n[16] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X605 a_4882_5142# row_n[3] a_5374_5504# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X606 vcm a_2275_2154# a_6982_2130# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X607 a_11398_17552# col_n[8] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X608 a_4974_16186# a_2475_16210# a_4882_16186# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X609 VDD rowon_n[6] a_28978_8154# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X610 vcm a_2275_5166# a_19030_5142# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X611 a_21038_1126# a_2475_1150# a_20946_1126# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X612 a_20034_5142# a_2475_5166# a_19942_5142# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X613 a_15414_16548# col_n[12] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X614 a_11910_13174# row_n[11] a_12402_13536# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X615 VDD rowon_n[1] a_26970_3134# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X616 a_5374_16548# col_n[2] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X617 a_21950_7150# row_n[5] a_22442_7512# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X618 a_14922_3134# row_n[1] a_15414_3496# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X619 a_2475_16210# a_1957_16210# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.171 pd=1.77 as=0.124 ps=1.01 w=0.6 l=0.15
X620 a_28066_13174# a_2475_13198# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X621 vcm a_2275_12194# a_9994_12170# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X622 a_26362_9198# col_n[23] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X623 VSS row_n[8] a_22346_10202# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X624 a_22954_11166# a_2275_11190# a_23046_11166# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X625 a_31382_3174# rowon_n[1] a_30986_3134# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X626 a_25054_3134# a_2475_3158# a_24962_3134# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X627 VSS row_n[14] a_21342_16226# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X628 a_24050_7150# a_2475_7174# a_23958_7150# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X629 VDD rowon_n[10] a_20946_12170# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X630 a_25966_9158# row_n[7] a_26458_9520# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X631 VDD rowon_n[4] a_32994_6146# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X632 a_26970_5142# row_n[3] a_27462_5504# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X633 a_25966_18194# a_2275_18218# a_26058_18194# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X634 a_30074_16186# a_2475_16210# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X635 a_19942_8154# a_2275_8178# a_20034_8154# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X636 VDD VSS a_30986_1126# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X637 VSS row_n[0] a_10298_2170# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X638 a_31078_4138# a_2475_4162# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X639 a_20946_4138# a_2275_4162# a_21038_4138# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X640 VDD VDD a_19942_18194# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X641 a_5278_14218# rowon_n[12] a_4882_14178# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X642 a_15318_14218# rowon_n[12] a_14922_14178# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X643 a_30074_8154# a_2475_8178# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X644 a_20338_15222# col_n[17] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X645 a_2475_17214# a_1957_17214# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.342 pd=2.97 as=0.249 ps=1.62 w=1.2 l=0.15
X646 a_12402_5504# col_n[9] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X647 a_13006_5142# a_2475_5166# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X648 VSS row_n[2] a_4274_4178# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X649 a_13310_17230# rowon_n[15] a_12914_17190# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X650 a_6890_13174# a_2275_13198# a_6982_13174# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X651 a_16930_13174# a_2275_13198# a_17022_13174# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X652 a_7286_7190# col_n[4] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X653 a_3270_17230# rowon_n[15] a_2874_17190# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X654 a_29070_5142# a_2475_5166# a_28978_5142# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X655 VSS row_n[11] a_4274_13214# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X656 VSS row_n[11] a_14314_13214# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X657 a_32082_12170# a_2475_12194# a_31990_12170# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X658 a_11302_10202# col_n[8] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X659 a_19942_13174# row_n[11] a_20434_13536# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X660 VSS row_n[4] a_21342_6186# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X661 a_32994_12170# row_n[10] a_33486_12532# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X662 a_14010_11166# a_2475_11190# a_13918_11166# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X663 a_24962_6146# a_2275_6170# a_25054_6146# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X664 a_31078_18194# a_2475_18218# a_30986_18194# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X665 a_3970_11166# a_2475_11190# a_3878_11166# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X666 a_2874_9158# a_2275_9182# a_2966_9158# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X667 VDD rowon_n[5] a_17934_7150# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X668 a_29982_7150# row_n[5] a_30474_7512# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X669 a_35094_6146# a_2475_6170# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X670 a_28978_2130# row_n[0] a_29470_2492# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X671 a_31990_18194# VDD a_32482_18556# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X672 VDD rowon_n[13] a_2874_15182# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X673 VDD rowon_n[13] a_12914_15182# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X674 vcm a_2275_14202# a_32082_14178# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X675 a_10394_12532# col_n[7] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X676 a_4370_4500# col_n[1] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X677 a_14410_11528# col_n[11] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X678 a_18026_3134# a_2475_3158# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X679 a_4370_11528# col_n[1] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X680 a_17022_7150# a_2475_7174# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X681 VDD a_2161_5166# a_2275_5166# VDD sky130_fd_pr__pfet_01v8 ad=0.249 pd=1.62 as=0.342 ps=2.97 w=1.2 l=0.15
X682 vcm a_2275_17214# a_30074_17190# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X683 a_13918_5142# a_2275_5166# a_14010_5142# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X684 a_33390_2170# col_n[30] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X685 a_14410_2492# col_n[11] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X686 VSS row_n[6] a_25358_8194# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X687 VSS row_n[2] a_26362_4178# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X688 a_35398_8194# rowon_n[6] a_35002_8154# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X689 a_26058_14178# a_2475_14202# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X690 a_35002_5142# row_n[3] a_35494_5504# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X691 a_9994_2130# a_2475_2154# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X692 VSS row_n[14] a_19334_16226# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X693 a_23350_14218# rowon_n[12] a_22954_14178# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X694 a_29374_12210# col_n[26] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X695 VSS row_n[9] a_20338_11206# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X696 VSS row_n[8] a_33390_10202# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X697 a_11302_4178# rowon_n[2] a_10906_4138# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X698 a_24050_17190# a_2475_17214# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X699 a_33998_11166# a_2275_11190# a_34090_11166# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X700 a_10298_10202# rowon_n[8] a_9902_10162# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X701 a_26458_4500# col_n[23] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X702 a_24962_13174# a_2275_13198# a_25054_13174# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X703 a_17934_7150# a_2275_7174# a_18026_7150# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X704 a_18938_3134# a_2275_3158# a_19030_3134# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X705 VDD VDD a_17934_18194# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X706 a_28466_14540# col_n[25] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X707 VDD rowon_n[10] a_31990_12170# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X708 a_28066_10162# a_2475_10186# a_27974_10162# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X709 a_10998_5142# a_2475_5166# a_10906_5142# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X710 a_20034_3134# a_2475_3158# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X711 a_8990_15182# a_2475_15206# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X712 VSS row_n[7] a_8290_9198# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X713 a_28978_10162# row_n[8] a_29470_10524# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X714 VDD VSS sky130_fd_pr__cap_mim_m3_1 l=17.2 w=17.2
X715 a_3270_3174# rowon_n[1] a_2874_3134# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X716 VDD rowon_n[2] a_10906_4138# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X717 VSS VDD a_34394_18234# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X718 a_31382_15222# col_n[28] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X719 a_9902_10162# a_2275_10186# a_9994_10162# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X720 a_2161_8178# sample VDD VDD sky130_fd_pr__pfet_01v8 ad=0.342 pd=2.97 as=0.342 ps=2.97 w=1.2 l=0.15
X721 vcm a_2275_6170# a_23046_6146# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X722 a_11302_18234# VDD a_10906_18194# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X723 a_35398_14218# VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X724 a_33086_6146# a_2475_6170# a_32994_6146# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X725 a_29070_18194# a_2475_18218# a_28978_18194# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X726 VSS row_n[12] a_12306_14218# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X727 a_20338_5182# rowon_n[3] a_19942_5142# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X728 a_30474_17552# col_n[27] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X729 vcm a_2275_15206# a_26058_15182# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X730 a_30074_13174# a_2475_13198# a_29982_13174# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X731 a_8386_9520# col_n[5] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X732 a_15014_7150# a_2475_7174# a_14922_7150# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X733 a_25054_1126# a_2475_1150# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X734 a_16018_3134# a_2475_3158# a_15926_3134# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X735 a_24050_5142# a_2475_5166# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X736 a_2874_17190# a_2275_17214# a_2966_17190# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X737 a_9994_17190# a_2475_17214# a_9902_17190# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X738 a_12914_17190# a_2275_17214# a_13006_17190# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X739 VDD VSS a_2874_1126# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X740 a_34490_16548# col_n[31] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X741 a_30986_13174# row_n[11] a_31478_13536# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X742 VDD rowon_n[6] a_21950_8154# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X743 vcm a_2275_5166# a_12002_5142# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X744 VDD rowon_n[14] a_10906_16186# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X745 vcm a_2275_10186# a_17022_10162# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X746 a_9902_8154# row_n[6] a_10394_8516# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X747 a_8290_1166# VSS a_7894_1126# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X748 VSS row_n[2] a_34394_4178# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X749 a_6890_14178# row_n[12] a_7382_14540# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X750 a_16930_14178# row_n[12] a_17422_14540# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X751 vcm a_2275_10186# a_6982_10162# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X752 a_8990_9158# a_2475_9182# a_8898_9158# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X753 VDD rowon_n[1] a_19942_3134# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X754 vcm a_2275_4162# a_28066_4138# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X755 a_24354_7190# rowon_n[5] a_23958_7150# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X756 a_2475_6170# a_1957_6170# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.342 pd=2.97 as=0.249 ps=1.62 w=1.2 l=0.15
X757 a_7986_2130# a_2475_2154# a_7894_2130# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X758 a_25358_3174# rowon_n[1] a_24962_3134# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X759 a_29070_3134# a_2475_3158# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X760 a_13310_3174# col_n[10] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X761 a_15318_9198# rowon_n[7] a_14922_9158# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X762 a_32994_9158# a_2275_9182# a_33086_9158# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X763 a_32082_10162# a_2475_10186# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X764 VDD rowon_n[4] a_26970_6146# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X765 vcm a_2275_3158# a_17022_3134# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X766 a_34490_4500# col_n[31] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X767 vcm a_2275_18218# a_7986_18194# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X768 vcm a_2275_18218# a_18026_18194# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X769 VSS row_n[15] a_26362_17230# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X770 a_30378_15222# rowon_n[13] a_29982_15182# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X771 vcm a_2275_7174# a_16018_7150# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X772 a_14922_6146# row_n[4] a_15414_6508# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X773 a_31990_2130# a_2275_2154# a_32082_2130# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X774 a_34394_14218# rowon_n[12] a_33998_14178# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X775 a_27366_13214# col_n[24] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X776 VSS row_n[9] a_31382_11206# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X777 VDD VSS a_24962_1126# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X778 a_22042_18194# a_2475_18218# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X779 a_12914_1126# VDD a_13406_1488# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X780 VSS row_n[3] a_19334_5182# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X781 a_13006_17190# a_2475_17214# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X782 a_35094_17190# a_2475_17214# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X783 a_5278_2170# col_n[2] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X784 a_29374_5182# rowon_n[3] a_28978_5142# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X785 a_2966_17190# a_2475_17214# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X786 a_22954_14178# a_2275_14202# a_23046_14178# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X787 VDD rowon_n[7] a_14922_9158# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X788 a_7286_8194# rowon_n[6] a_6890_8154# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X789 a_18330_1166# en_bit_n[1] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X790 VDD VDD a_28978_18194# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X791 a_6982_16186# a_2475_16210# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X792 a_17022_16186# a_2475_16210# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X793 a_26458_15544# col_n[23] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X794 VDD rowon_n[11] a_29982_13174# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X795 a_26058_11166# a_2475_11190# a_25966_11166# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X796 vcm a_2275_2154# a_8990_2130# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X797 a_30378_10202# col_n[27] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X798 VDD a_2161_12194# a_2275_12194# VDD sky130_fd_pr__pfet_01v8 ad=0.249 pd=1.62 as=0.342 ps=2.97 w=1.2 l=0.15
X799 a_26970_11166# row_n[9] a_27462_11528# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X800 a_23046_1126# a_2475_1150# a_22954_1126# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X801 a_19430_3496# col_n[16] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X802 a_22042_5142# a_2475_5166# a_21950_5142# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X803 VDD rowon_n[1] a_28978_3134# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X804 a_24962_14178# row_n[12] a_25454_14540# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X805 vcm a_2275_10186# a_25054_10162# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X806 a_23958_7150# row_n[5] a_24450_7512# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X807 a_8990_12170# a_2475_12194# a_8898_12170# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X808 a_28370_9198# col_n[25] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X809 a_19334_16226# col_n[16] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X810 vcm a_2275_16210# a_24050_16186# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X811 a_21950_2130# row_n[0] a_22442_2492# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X812 a_10906_18194# a_2275_18218# a_10998_18194# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X813 a_18026_18194# a_2475_18218# a_17934_18194# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X814 a_9294_16226# col_n[6] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X815 a_7986_18194# a_2475_18218# a_7894_18194# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X816 a_9390_12532# col_n[6] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X817 a_2475_11190# a_1957_11190# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.171 pd=1.77 as=0.124 ps=1.01 w=0.6 l=0.15
X818 a_27366_2170# col_n[24] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X819 a_33390_3174# rowon_n[1] a_32994_3134# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X820 a_10998_3134# a_2475_3158# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X821 a_18426_18556# col_n[15] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X822 a_27062_3134# a_2475_3158# a_26970_3134# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X823 a_8386_18556# col_n[5] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X824 vcm a_2275_9182# a_31078_9158# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X825 a_17326_8194# col_n[14] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X826 a_3970_9158# a_2475_9182# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X827 a_27974_9158# row_n[7] a_28466_9520# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X828 a_28978_5142# row_n[3] a_29470_5504# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X829 a_6890_8154# row_n[6] a_7382_8516# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X830 VSS row_n[0] a_12306_2170# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X831 a_22954_4138# a_2275_4162# a_23046_4138# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X832 a_32082_8154# a_2475_8178# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X833 VDD VSS a_32994_1126# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X834 a_33086_4138# a_2475_4162# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X835 a_2161_17214# sample VSS VSS sky130_fd_pr__nfet_01v8 ad=0.171 pd=1.77 as=0.171 ps=1.77 w=0.6 l=0.15
X836 a_28370_15222# rowon_n[13] a_27974_15182# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X837 VSS row_n[10] a_25358_12210# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X838 a_30074_11166# a_2475_11190# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X839 a_14410_5504# col_n[11] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X840 a_2966_2130# a_2475_2154# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X841 VSS row_n[9] a_29374_11206# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X842 a_15014_5142# a_2475_5166# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X843 a_16018_1126# a_2475_1150# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X844 a_9294_7190# col_n[6] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X845 VDD rowon_n[12] a_23958_14178# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X846 a_12002_12170# a_2475_12194# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X847 a_34090_12170# a_2475_12194# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X848 a_10906_7150# a_2275_7174# a_10998_7150# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X849 a_11910_3134# a_2275_3158# a_12002_3134# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X850 a_9294_10202# rowon_n[8] a_8898_10162# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X851 VSS row_n[4] a_23350_6186# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X852 a_33086_18194# a_2475_18218# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X853 VDD rowon_n[11] a_27974_13174# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X854 a_25454_10524# col_n[22] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X855 a_10998_18194# a_2475_18218# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X856 a_23350_17230# col_n[20] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X857 a_33998_14178# a_2275_14202# a_34090_14178# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X858 a_4882_9158# a_2275_9182# a_4974_9158# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X859 VDD rowon_n[0] a_17934_2130# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X860 a_2161_18218# sample VDD VDD sky130_fd_pr__pfet_01v8 ad=0.342 pd=2.97 as=0.342 ps=2.97 w=1.2 l=0.15
X861 a_29982_2130# row_n[0] a_30474_2492# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X862 a_3878_2130# a_2275_2154# a_3970_2130# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X863 VSS row_n[13] a_7286_15222# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X864 VSS row_n[13] a_17326_15222# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X865 a_22042_15182# a_2475_15206# a_21950_15182# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X866 a_4274_12210# col_n[1] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X867 a_14314_12210# col_n[11] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X868 a_15926_5142# a_2275_5166# a_16018_5142# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X869 a_16930_1126# a_2275_1150# a_17022_1126# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X870 a_18330_11206# col_n[15] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X871 vcm a_2275_11190# a_23046_11166# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X872 a_35398_2170# VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X873 VSS row_n[2] a_28370_4178# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X874 a_22954_15182# row_n[13] a_23446_15544# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X875 a_17022_13174# a_2475_13198# a_16930_13174# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X876 a_8290_11206# col_n[5] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X877 VSS row_n[6] a_27366_8194# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X878 a_6982_13174# a_2475_13198# a_6890_13174# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X879 a_9902_13174# a_2275_13198# a_9994_13174# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X880 a_1957_4162# VSS sample VDD sky130_fd_pr__pfet_01v8 ad=0.342 pd=2.97 as=0.342 ps=2.97 w=1.2 l=0.15
X881 VDD rowon_n[15] a_5886_17190# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X882 VDD rowon_n[15] a_15926_17190# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X883 a_3366_14540# col_n[0] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X884 a_13406_14540# col_n[10] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X885 a_17422_13536# col_n[14] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X886 a_13918_10162# row_n[8] a_14410_10524# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X887 a_2161_2154# sample VSS VSS sky130_fd_pr__nfet_01v8 ad=0.171 pd=1.77 as=0.171 ps=1.77 w=0.6 l=0.15
X888 a_7382_13536# col_n[4] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X889 a_3878_10162# row_n[8] a_4370_10524# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X890 vcm a_2275_8178# a_20034_8154# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X891 vcm a_2275_4162# a_21038_4138# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X892 a_13310_4178# rowon_n[2] a_12914_4138# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X893 a_26970_9158# a_2275_9182# a_27062_9158# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X894 a_30074_8154# a_2475_8178# a_29982_8154# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X895 VSS row_n[5] a_16322_7190# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X896 a_31078_4138# a_2475_4162# a_30986_4138# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X897 a_28466_4500# col_n[25] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X898 a_6378_7512# col_n[3] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X899 a_13006_5142# a_2475_5166# a_12914_5142# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X900 a_22042_3134# a_2475_3158# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X901 a_22346_17230# rowon_n[15] a_21950_17190# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X902 vcm a_2275_15206# a_10998_15182# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X903 VDD rowon_n[4] a_19942_6146# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X904 a_4882_18194# VDD a_5374_18556# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X905 a_14922_18194# VDD a_15414_18556# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X906 a_26362_16226# rowon_n[14] a_25966_16186# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X907 vcm a_2275_14202# a_4974_14178# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X908 vcm a_2275_14202# a_15014_14178# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X909 VSS row_n[11] a_23350_13214# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X910 a_8990_10162# a_2475_10186# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X911 VDD rowon_n[2] a_12914_4138# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X912 vcm a_2275_6170# a_25054_6146# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X913 a_35094_6146# a_2475_6170# a_35002_6146# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X914 a_27974_15182# a_2275_15206# a_28066_15182# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X915 a_32082_13174# a_2475_13198# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X916 vcm a_2275_9182# a_2966_9158# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X917 VDD rowon_n[13] a_21950_15182# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X918 a_17326_11206# rowon_n[9] a_16930_11166# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X919 a_11302_1166# col_n[8] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X920 a_22346_5182# rowon_n[3] a_21950_5142# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X921 VDD rowon_n[12] a_35002_14178# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X922 a_7286_11206# rowon_n[9] a_6890_11166# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X923 a_17022_7150# a_2475_7174# a_16930_7150# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X924 a_10298_5182# col_n[7] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X925 a_27062_1126# a_2475_1150# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X926 a_18026_3134# a_2475_3158# a_17934_3134# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X927 a_23446_11528# col_n[20] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X928 VDD VSS VSS sky130_fd_pr__cap_var_lvt w=16.4 l=16
X929 a_21342_18234# col_n[18] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X930 VDD rowon_n[6] a_23958_8154# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X931 vcm a_2275_5166# a_14010_5142# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X932 a_34394_17230# col_n[31] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X933 VDD rowon_n[1] a_21950_3134# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X934 VSS row_n[15] a_11302_17230# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X935 a_9902_3134# row_n[1] a_10394_3496# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X936 a_29982_18194# a_2275_18218# a_30074_18194# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X937 VSS row_n[14] a_15318_16226# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X938 a_20034_16186# a_2475_16210# a_19942_16186# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X939 a_12306_13214# col_n[9] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X940 vcm a_2275_17214# a_29070_17190# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X941 VSS row_n[14] a_5278_16226# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X942 a_10998_15182# a_2475_15206# a_10906_15182# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X943 a_33086_15182# a_2475_15206# a_32994_15182# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X944 a_21342_9198# col_n[18] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X945 VSS row_n[7] a_31382_9198# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X946 a_26362_7190# rowon_n[5] a_25966_7150# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X947 a_9994_2130# a_2475_2154# a_9902_2130# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X948 a_27366_3174# rowon_n[1] a_26970_3134# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X949 a_15318_3174# col_n[12] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X950 a_20946_16186# row_n[14] a_21438_16548# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X951 a_5278_6186# rowon_n[4] a_4882_6146# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X952 a_33998_15182# row_n[13] a_34490_15544# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X953 a_15014_14178# a_2475_14202# a_14922_14178# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X954 vcm a_2275_11190# a_34090_11166# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X955 a_17326_9198# rowon_n[7] a_16930_9158# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X956 a_35002_9158# a_2275_9182# a_35094_9158# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X957 a_19430_6508# col_n[16] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X958 VDD VDD a_13918_18194# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X959 a_11398_15544# col_n[8] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X960 a_4974_14178# a_2475_14202# a_4882_14178# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X961 vcm a_2275_7174# a_18026_7150# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X962 VDD rowon_n[4] a_28978_6146# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X963 vcm a_2275_3158# a_19030_3134# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X964 VDD VDD a_3878_18194# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X965 a_20034_3134# a_2475_3158# a_19942_3134# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X966 a_11910_11166# row_n[9] a_12402_11528# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X967 a_33998_2130# a_2275_2154# a_34090_2130# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X968 VDD VSS a_26970_1126# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X969 a_20946_9158# row_n[7] a_21438_9520# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X970 a_26058_8154# a_2475_8178# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X971 a_14922_1126# VDD a_15414_1488# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X972 a_21950_5142# row_n[3] a_22442_5504# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X973 a_31478_9520# col_n[28] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X974 a_2475_14202# a_1957_14202# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.171 pd=1.77 as=0.124 ps=1.01 w=0.6 l=0.15
X975 a_9902_14178# row_n[12] a_10394_14540# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X976 vcm a_2275_10186# a_9994_10162# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X977 a_21342_12210# rowon_n[10] a_20946_12170# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X978 VDD rowon_n[7] a_16930_9158# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X979 a_9294_8194# rowon_n[6] a_8898_8154# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X980 a_20338_18234# VDD a_19942_18194# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X981 a_31382_1166# VSS a_30986_1126# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X982 a_17022_11166# a_2475_11190# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X983 a_25054_1126# a_2475_1150# a_24962_1126# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X984 VSS row_n[12] a_21342_14218# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X985 a_6982_11166# a_2475_11190# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X986 a_24050_5142# a_2475_5166# a_23958_5142# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X987 a_21950_17190# a_2275_17214# a_22042_17190# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X988 VDD rowon_n[8] a_20946_10162# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X989 a_25966_7150# row_n[5] a_26458_7512# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X990 VDD VSS VSS sky130_fd_pr__cap_var_lvt w=16.4 l=16
X991 a_25966_16186# a_2275_16210# a_26058_16186# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X992 a_30074_14178# a_2475_14202# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X993 a_19942_6146# a_2275_6170# a_20034_6146# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X994 a_9994_18194# a_2475_18218# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X995 VDD rowon_n[14] a_19942_16186# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X996 a_30074_6146# a_2475_6170# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X997 a_23958_2130# row_n[0] a_24450_2492# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X998 a_20338_13214# col_n[17] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X999 a_33390_12210# col_n[30] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1000 a_2475_15206# a_1957_15206# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.342 pd=2.97 as=0.249 ps=1.62 w=1.2 l=0.15
X1001 a_12002_7150# a_2475_7174# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1002 a_29374_2170# col_n[26] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1003 a_13006_3134# a_2475_3158# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1004 a_3270_15222# rowon_n[13] a_2874_15182# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X1005 a_13310_15222# rowon_n[13] a_12914_15182# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X1006 VSS row_n[10] a_10298_12210# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1007 a_7286_5182# col_n[4] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1008 a_32386_18234# col_n[29] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1009 a_19334_8194# col_n[16] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1010 a_29070_3134# a_2475_3158# a_28978_3134# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X1011 a_32482_14540# col_n[29] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X1012 vcm a_2275_12194# a_28066_12170# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1013 VSS row_n[9] a_4274_11206# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1014 VSS row_n[9] a_14314_11206# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1015 a_32082_10162# a_2475_10186# a_31990_10162# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X1016 vcm a_2275_9182# a_33086_9158# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1017 a_19942_11166# row_n[9] a_20434_11528# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1018 a_8898_8154# row_n[6] a_9390_8516# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1019 VSS row_n[6] a_20338_8194# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1020 VSS row_n[2] a_21342_4178# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1021 vcm a_2275_18218# a_27062_18194# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1022 a_31078_16186# a_2475_16210# a_30986_16186# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X1023 a_32994_10162# row_n[8] a_33486_10524# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1024 a_30378_8194# rowon_n[6] a_29982_8154# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X1025 VSS row_n[0] a_14314_2170# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1026 a_24962_4138# a_2275_4162# a_25054_4138# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1027 a_34090_8154# a_2475_8178# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1028 VDD rowon_n[3] a_17934_5142# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1029 vcm a_2275_2154# a_32082_2130# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1030 a_35094_4138# a_2475_4162# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1031 a_29982_5142# row_n[3] a_30474_5504# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1032 a_31990_16186# row_n[14] a_32482_16548# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1033 VDD rowon_n[11] a_2874_13174# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1034 VDD rowon_n[11] a_12914_13174# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1035 a_10394_10524# col_n[7] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X1036 a_4974_2130# a_2475_2154# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1037 a_6890_3134# row_n[1] a_7382_3496# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1038 a_17022_5142# a_2475_5166# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1039 a_18026_1126# a_2475_1150# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1040 a_2161_12194# sample VSS VSS sky130_fd_pr__nfet_01v8 ad=0.171 pd=1.77 as=0.171 ps=1.77 w=0.6 l=0.15
X1041 VDD a_2161_3158# a_2275_3158# VDD sky130_fd_pr__pfet_01v8 ad=0.249 pd=1.62 as=0.342 ps=2.97 w=1.2 l=0.15
X1042 a_13918_3134# a_2275_3158# a_14010_3134# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1043 a_21438_4500# col_n[18] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X1044 vcm a_2275_15206# a_30074_15182# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1045 a_12914_7150# a_2275_7174# a_13006_7150# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1046 VSS row_n[4] a_25358_6186# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1047 VSS row_n[7] a_3270_9198# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1048 a_35398_6186# rowon_n[4] a_35002_6146# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X1049 a_18330_18234# VDD a_17934_18194# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X1050 a_32386_12210# rowon_n[10] a_31990_12170# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X1051 VSS row_n[12] a_19334_14218# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1052 a_29374_10202# col_n[26] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1053 ctop sw ctop VDD sky130_fd_pr__pfet_01v8 ad=0.275 pd=2.19 as=2.71 ps=21.9 w=1.9 l=0.22
X1054 a_24050_15182# a_2475_15206# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1055 a_20946_12170# a_2275_12194# a_21038_12170# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1056 a_5886_2130# a_2275_2154# a_5978_2130# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1057 a_18938_1126# a_2275_1150# a_19030_1126# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1058 a_17934_5142# a_2275_5166# a_18026_5142# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1059 VDD rowon_n[14] a_17934_16186# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1060 a_28466_12532# col_n[25] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X1061 VDD rowon_n[8] a_31990_10162# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1062 a_3366_9520# col_n[0] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X1063 VSS row_n[6] a_29374_8194# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1064 a_20034_1126# a_2475_1150# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1065 a_10998_3134# a_2475_3158# a_10906_3134# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X1066 a_8990_13174# a_2475_13198# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1067 a_16418_8516# col_n[13] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X1068 VSS row_n[15] a_30378_17230# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1069 a_3270_1166# VSS a_2874_1126# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X1070 VSS row_n[14] a_34394_16226# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1071 a_31382_13214# col_n[28] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1072 a_3970_9158# a_2475_9182# a_3878_9158# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X1073 a_32386_7190# col_n[29] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1074 a_2161_6170# sample VDD VDD sky130_fd_pr__pfet_01v8 ad=0.342 pd=2.97 as=0.342 ps=2.97 w=1.2 l=0.15
X1075 a_11302_16226# rowon_n[14] a_10906_16186# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X1076 vcm a_2275_4162# a_23046_4138# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1077 a_25054_17190# a_2475_17214# a_24962_17190# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X1078 a_28978_9158# a_2275_9182# a_29070_9158# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1079 a_32082_8154# a_2475_8178# a_31990_8154# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X1080 VSS row_n[5] a_18330_7190# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1081 a_33086_4138# a_2475_4162# a_32994_4138# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X1082 a_29070_16186# a_2475_16210# a_28978_16186# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X1083 vcm a_2275_13198# a_26058_13174# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1084 a_2966_2130# a_2475_2154# a_2874_2130# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X1085 a_20338_3174# rowon_n[1] a_19942_3134# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X1086 VDD VDD a_32994_18194# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1087 a_25966_17190# row_n[15] a_26458_17552# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1088 a_30474_15544# col_n[27] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X1089 a_30074_11166# a_2475_11190# a_29982_11166# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X1090 a_8386_7512# col_n[5] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X1091 a_15014_5142# a_2475_5166# a_14922_5142# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X1092 a_16018_1126# a_2475_1150# a_15926_1126# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X1093 a_24050_3134# a_2475_3158# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1094 a_2874_15182# a_2275_15206# a_2966_15182# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1095 a_9994_15182# a_2475_15206# a_9902_15182# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X1096 a_12914_15182# a_2275_15206# a_13006_15182# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1097 a_10298_9198# rowon_n[7] a_9902_9158# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X1098 a_30986_11166# row_n[9] a_31478_11528# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1099 VDD rowon_n[4] a_21950_6146# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1100 a_6378_2492# col_n[3] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X1101 vcm a_2275_3158# a_12002_3134# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1102 vcm a_2275_7174# a_10998_7150# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1103 a_9902_6146# row_n[4] a_10394_6508# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1104 a_6890_12170# row_n[10] a_7382_12532# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1105 a_16930_12170# row_n[10] a_17422_12532# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1106 VDD en_bit_n[0] a_19942_1126# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1107 vcm a_2275_9182# a_4974_9158# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1108 a_25358_1166# VSS a_24962_1126# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X1109 a_2475_4162# a_1957_4162# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.342 pd=2.97 as=0.249 ps=1.62 w=1.2 l=0.15
X1110 a_24354_5182# rowon_n[3] a_23958_5142# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X1111 VDD rowon_n[7] a_9902_9158# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1112 a_13310_1166# col_n[10] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1113 a_29070_1126# a_2475_1150# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1114 vcm a_2275_17214# a_14010_17190# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1115 a_27974_10162# a_2275_10186# a_28066_10162# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1116 vcm a_2275_2154# a_3970_2130# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1117 vcm a_2275_17214# a_3970_17190# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1118 VDD rowon_n[6] a_25966_8154# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1119 vcm a_2275_1150# a_17022_1126# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1120 a_29374_18234# VDD a_28978_18194# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X1121 vcm a_2275_16210# a_7986_16186# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1122 vcm a_2275_16210# a_18026_16186# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1123 VSS row_n[13] a_26362_15222# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1124 a_30378_13214# rowon_n[11] a_29982_13174# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X1125 vcm a_2275_5166# a_16018_5142# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1126 a_27366_11206# col_n[24] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1127 VDD rowon_n[1] a_23958_3134# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1128 a_22042_16186# a_2475_16210# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1129 VSS row_n[1] a_19334_3174# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1130 VDD rowon_n[15] a_24962_17190# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1131 a_13006_15182# a_2475_15206# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1132 a_35094_15182# a_2475_15206# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1133 a_31990_12170# a_2275_12194# a_32082_12170# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1134 a_23350_9198# col_n[20] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1135 a_28370_7190# rowon_n[5] a_27974_7150# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X1136 a_29374_3174# rowon_n[1] a_28978_3134# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X1137 a_2966_15182# a_2475_15206# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1138 VSS row_n[7] a_33390_9198# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1139 VDD rowon_n[5] a_14922_7150# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1140 a_7286_6186# rowon_n[4] a_6890_6146# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X1141 VDD rowon_n[14] a_28978_16186# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1142 a_6982_14178# a_2475_14202# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1143 a_17022_14178# a_2475_14202# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1144 a_26458_13536# col_n[23] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X1145 VDD rowon_n[9] a_29982_11166# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1146 vcm a_2275_9182# a_27062_9158# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1147 a_22346_2170# col_n[19] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1148 VDD a_2161_10186# a_2275_10186# VDD sky130_fd_pr__pfet_01v8 ad=0.249 pd=1.62 as=0.342 ps=2.97 w=1.2 l=0.15
X1149 a_24050_12170# a_2475_12194# a_23958_12170# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X1150 a_19430_1488# en_bit_n[2] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X1151 a_22042_3134# a_2475_3158# a_21950_3134# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X1152 VSS row_n[10] a_9294_12210# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1153 a_12306_8194# col_n[9] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1154 a_28066_8154# a_2475_8178# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1155 VDD VSS a_28978_1126# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1156 VSS VDD a_18330_18234# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1157 a_23046_18194# a_2475_18218# a_22954_18194# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X1158 a_24962_12170# row_n[10] a_25454_12532# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1159 a_22954_9158# row_n[7] a_23446_9520# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1160 a_23958_5142# row_n[3] a_24450_5504# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1161 VSS VDD a_8290_18234# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1162 a_8990_10162# a_2475_10186# a_8898_10162# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X1163 a_33486_9520# col_n[30] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X1164 a_23958_18194# VDD a_24450_18556# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1165 a_19334_14218# col_n[16] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1166 vcm a_2275_14202# a_24050_14178# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1167 a_10906_16186# a_2275_16210# a_10998_16186# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1168 a_18026_16186# a_2475_16210# a_17934_16186# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X1169 VDD rowon_n[12] a_7894_14178# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1170 a_9294_14218# col_n[6] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1171 a_7986_16186# a_2475_16210# a_7894_16186# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X1172 a_9390_10524# col_n[6] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X1173 a_33390_1166# VSS a_32994_1126# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X1174 a_10998_1126# a_2475_1150# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1175 a_18426_16548# col_n[15] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X1176 a_4274_7190# col_n[1] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1177 a_27062_1126# a_2475_1150# a_26970_1126# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X1178 a_8386_16548# col_n[5] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X1179 a_17326_6186# col_n[14] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1180 VDD VSS sky130_fd_pr__cap_mim_m3_1 l=17.2 w=17.2
X1181 a_27974_7150# row_n[5] a_28466_7512# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1182 vcm a_2275_12194# a_13006_12170# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1183 a_6890_6146# row_n[4] a_7382_6508# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1184 vcm a_2275_12194# a_2966_12170# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1185 a_32082_6146# a_2475_6170# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1186 a_25966_2130# row_n[0] a_26458_2492# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1187 a_2161_15206# sample VSS VSS sky130_fd_pr__nfet_01v8 ad=0.171 pd=1.77 as=0.171 ps=1.77 w=0.6 l=0.15
X1188 a_28370_13214# rowon_n[11] a_27974_13174# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X1189 VSS row_n[8] a_25358_10202# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1190 vcm a_2275_18218# a_12002_18194# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1191 a_25966_11166# a_2275_11190# a_26058_11166# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1192 a_14010_7150# a_2475_7174# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1193 a_15014_3134# a_2475_3158# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1194 a_9294_5182# col_n[6] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1195 VDD rowon_n[10] a_23958_12170# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1196 vcm a_2275_9182# a_35094_9158# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1197 a_10906_5142# a_2275_5166# a_10998_5142# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1198 a_11910_1126# a_2275_1150# a_12002_1126# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1199 a_30378_2170# col_n[27] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1200 a_18330_2170# rowon_n[0] a_17934_2130# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X1201 VSS row_n[2] a_23350_4178# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1202 a_28978_18194# a_2275_18218# a_29070_18194# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1203 a_33086_16186# a_2475_16210# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1204 VDD rowon_n[9] a_27974_11166# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1205 VSS row_n[6] a_22346_8194# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1206 a_32386_8194# rowon_n[6] a_31990_8154# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X1207 a_10998_16186# a_2475_16210# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1208 vcm a_2275_2154# a_34090_2130# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1209 a_23350_15222# col_n[20] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1210 a_26058_8154# a_2475_8178# a_25966_8154# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X1211 a_8898_3134# row_n[1] a_9390_3496# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1212 a_6982_2130# a_2475_2154# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1213 a_16322_17230# rowon_n[15] a_15926_17190# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X1214 a_6282_17230# rowon_n[15] a_5886_17190# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X1215 a_2161_16210# sample VDD VDD sky130_fd_pr__pfet_01v8 ad=0.342 pd=2.97 as=0.342 ps=2.97 w=1.2 l=0.15
X1216 a_21950_9158# a_2275_9182# a_22042_9158# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1217 VSS row_n[5] a_11302_7190# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1218 a_22442_17552# col_n[19] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X1219 VSS row_n[11] a_7286_13214# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1220 VSS row_n[11] a_17326_13214# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1221 a_22042_13174# a_2475_13198# a_21950_13174# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X1222 a_35094_12170# a_2475_12194# a_35002_12170# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X1223 a_4274_10202# col_n[1] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1224 a_14314_10202# col_n[11] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1225 a_14922_7150# a_2275_7174# a_15014_7150# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1226 a_15926_3134# a_2275_3158# a_16018_3134# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1227 a_23446_4500# col_n[20] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X1228 a_2966_12170# a_2475_12194# a_2874_12170# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X1229 a_13006_12170# a_2475_12194# a_12914_12170# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X1230 a_22954_13174# row_n[11] a_23446_13536# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1231 a_17022_11166# a_2475_11190# a_16930_11166# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X1232 VSS row_n[4] a_27366_6186# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1233 a_6982_11166# a_2475_11190# a_6890_11166# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X1234 VSS row_n[7] a_5278_9198# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1235 a_1957_18218# VDD sample VSS sky130_fd_pr__nfet_01v8 ad=0.171 pd=1.77 as=0.171 ps=1.77 w=0.6 l=0.15
X1236 VDD rowon_n[13] a_5886_15182# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1237 VDD rowon_n[13] a_15926_15182# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1238 a_3366_12532# col_n[0] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X1239 a_13406_12532# col_n[10] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X1240 a_17422_11528# col_n[14] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X1241 a_7382_11528# col_n[4] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X1242 vcm a_2275_6170# a_20034_6146# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1243 a_15318_18234# col_n[12] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1244 vcm a_2275_18218# a_20034_18194# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1245 a_30074_6146# a_2475_6170# a_29982_6146# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X1246 VSS row_n[3] a_16322_5182# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1247 a_7894_2130# a_2275_2154# a_7986_2130# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1248 a_5278_18234# col_n[2] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1249 vcm a_2275_17214# a_33086_17190# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1250 a_5374_9520# col_n[2] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X1251 a_31990_8154# row_n[6] a_32482_8516# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1252 a_6378_5504# col_n[3] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X1253 a_24050_10162# a_2475_10186# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1254 a_18426_8516# col_n[15] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X1255 a_12002_7150# a_2475_7174# a_11910_7150# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X1256 a_22042_1126# a_2475_1150# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1257 a_13006_3134# a_2475_3158# a_12914_3134# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X1258 a_10906_17190# row_n[15] a_11398_17552# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1259 a_22346_15222# rowon_n[13] a_21950_15182# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X1260 vcm a_2275_13198# a_10998_13174# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1261 a_4882_16186# row_n[14] a_5374_16548# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1262 a_14922_16186# row_n[14] a_15414_16548# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1263 a_26362_14218# rowon_n[12] a_25966_14178# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X1264 VSS row_n[9] a_23350_11206# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1265 a_16418_3496# col_n[13] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X1266 a_34394_7190# col_n[31] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1267 vcm a_2275_4162# a_25054_4138# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1268 a_27062_17190# a_2475_17214# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1269 a_34090_8154# a_2475_8178# a_33998_8154# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X1270 a_35094_4138# a_2475_4162# a_35002_4138# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X1271 a_27974_13174# a_2275_13198# a_28066_13174# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1272 a_1957_9182# VDD sample VSS sky130_fd_pr__nfet_01v8 ad=0.171 pd=1.77 as=0.171 ps=1.77 w=0.6 l=0.15
X1273 VDD rowon_n[11] a_21950_13174# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1274 a_21342_7190# rowon_n[5] a_20946_7150# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X1275 a_4974_2130# a_2475_2154# a_4882_2130# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X1276 a_22346_3174# rowon_n[1] a_21950_3134# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X1277 a_10298_3174# col_n[7] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1278 VDD rowon_n[10] a_35002_12170# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1279 a_17022_5142# a_2475_5166# a_16930_5142# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X1280 a_18026_1126# a_2475_1150# a_17934_1126# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X1281 a_12306_9198# rowon_n[7] a_11910_9158# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X1282 a_29982_9158# a_2275_9182# a_30074_9158# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1283 a_21342_16226# col_n[18] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1284 vcm a_2275_7174# a_13006_7150# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1285 VDD rowon_n[4] a_23958_6146# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1286 a_8386_2492# col_n[5] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X1287 vcm a_2275_3158# a_14010_3134# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1288 a_34394_15222# col_n[31] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1289 a_12914_10162# a_2275_10186# a_13006_10162# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1290 VDD VSS sky130_fd_pr__cap_mim_m3_1 l=17.2 w=17.2
X1291 a_2874_10162# a_2275_10186# a_2966_10162# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1292 VDD VSS a_21950_1126# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1293 a_4274_18234# VDD a_3878_18194# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X1294 a_14314_18234# VDD a_13918_18194# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X1295 VSS row_n[13] a_11302_15222# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1296 a_21038_8154# a_2475_8178# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1297 a_9902_1126# VDD a_10394_1488# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1298 a_20434_18556# col_n[17] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X1299 a_29982_16186# a_2275_16210# a_30074_16186# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1300 VSS row_n[12] a_15318_14218# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1301 a_20034_14178# a_2475_14202# a_19942_14178# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X1302 a_12306_11206# col_n[9] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1303 a_33486_17552# col_n[30] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X1304 vcm a_2275_15206# a_29070_15182# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1305 VSS row_n[12] a_5278_14218# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1306 a_10998_13174# a_2475_13198# a_10906_13174# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X1307 a_33086_13174# a_2475_13198# a_32994_13174# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X1308 a_15318_1166# col_n[12] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1309 a_27366_1166# VSS a_26970_1126# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X1310 a_26362_5182# rowon_n[3] a_25966_5142# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X1311 a_5886_17190# a_2275_17214# a_5978_17190# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1312 a_15926_17190# a_2275_17214# a_16018_17190# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1313 VDD rowon_n[7] a_11910_9158# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1314 a_4274_8194# rowon_n[6] a_3878_8154# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X1315 a_5278_4178# rowon_n[2] a_4882_4138# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X1316 VDD rowon_n[15] a_9902_17190# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1317 a_33998_13174# row_n[11] a_34490_13536# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1318 vcm a_2275_2154# a_5978_2130# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1319 VDD rowon_n[14] a_13918_16186# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1320 a_11398_13536# col_n[8] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X1321 VDD rowon_n[6] a_27974_8154# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1322 vcm a_2275_5166# a_18026_5142# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1323 vcm a_2275_1150# a_19030_1126# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1324 VDD rowon_n[14] a_3878_16186# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1325 a_20034_1126# a_2475_1150# a_19942_1126# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X1326 a_20946_7150# row_n[5] a_21438_7512# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1327 a_26058_6146# a_2475_6170# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1328 VDD rowon_n[1] a_25966_3134# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1329 vcm a_2275_18218# a_31078_18194# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1330 a_31478_7512# col_n[28] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X1331 VDD rowon_n[2] a_4882_4138# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1332 a_9902_12170# row_n[10] a_10394_12532# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1333 a_21342_10202# rowon_n[8] a_20946_10162# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X1334 a_25358_9198# col_n[22] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1335 a_22042_11166# a_2475_11190# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1336 VSS row_n[7] a_35398_9198# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1337 VDD rowon_n[5] a_16930_7150# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1338 a_9294_6186# rowon_n[4] a_8898_6146# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X1339 a_13006_10162# a_2475_10186# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1340 a_35094_10162# a_2475_10186# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1341 vcm a_2275_9182# a_29070_9158# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1342 a_20338_16226# rowon_n[14] a_19942_16186# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X1343 a_2966_10162# a_2475_10186# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1344 a_24354_2170# col_n[21] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1345 VDD rowon_n[0] a_14922_2130# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1346 a_14314_8194# col_n[11] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1347 a_24050_3134# a_2475_3158# a_23958_3134# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X1348 a_25054_18194# a_2475_18218# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1349 a_21950_15182# a_2275_15206# a_22042_15182# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1350 a_24962_9158# row_n[7] a_25454_9520# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1351 a_25966_5142# row_n[3] a_26458_5504# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1352 a_16018_17190# a_2475_17214# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1353 a_35494_9520# VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X1354 a_3878_8154# row_n[6] a_4370_8516# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1355 a_5978_17190# a_2475_17214# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1356 a_25966_14178# a_2275_14202# a_26058_14178# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1357 a_19942_4138# a_2275_4162# a_20034_4138# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1358 a_9994_16186# a_2475_16210# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1359 a_30074_4138# a_2475_4162# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1360 a_20338_11206# col_n[17] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1361 a_33390_10202# col_n[30] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1362 a_2475_13198# a_1957_13198# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.342 pd=2.97 as=0.249 ps=1.62 w=1.2 l=0.15
X1363 a_12002_5142# a_2475_5166# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1364 a_13006_1126# a_2475_1150# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1365 a_3270_13214# rowon_n[11] a_2874_13174# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X1366 a_13310_13214# rowon_n[11] a_12914_13174# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X1367 VSS row_n[8] a_10298_10202# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1368 a_6282_7190# col_n[3] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1369 a_7286_3174# col_n[4] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1370 a_32386_16226# col_n[29] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1371 a_10906_11166# a_2275_11190# a_10998_11166# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1372 a_19334_6186# col_n[16] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1373 a_29070_1126# a_2475_1150# a_28978_1126# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X1374 a_27974_14178# row_n[12] a_28466_14540# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1375 a_32482_12532# col_n[29] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X1376 vcm a_2275_10186# a_28066_10162# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1377 a_14922_12170# a_2275_12194# a_15014_12170# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1378 a_8898_6146# row_n[4] a_9390_6508# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1379 VSS row_n[4] a_20338_6186# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1380 vcm a_2275_16210# a_27062_16186# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1381 a_31078_14178# a_2475_14202# a_30986_14178# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X1382 a_4882_12170# a_2275_12194# a_4974_12170# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1383 a_30378_6186# rowon_n[4] a_29982_6146# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X1384 a_13918_18194# a_2275_18218# a_14010_18194# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1385 a_31478_18556# col_n[28] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X1386 a_34090_6146# a_2475_6170# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1387 a_27974_2130# row_n[0] a_28466_2492# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1388 a_3878_18194# a_2275_18218# a_3970_18194# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1389 VDD rowon_n[9] a_2874_11166# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1390 VDD rowon_n[9] a_12914_11166# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1391 a_6890_1126# VDD a_7382_1488# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1392 a_17022_3134# a_2475_3158# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1393 a_2161_10186# sample VSS VSS sky130_fd_pr__nfet_01v8 ad=0.171 pd=1.77 as=0.171 ps=1.77 w=0.6 l=0.15
X1394 VDD a_2161_1150# a_2275_1150# VDD sky130_fd_pr__pfet_01v8 ad=0.249 pd=1.62 as=0.342 ps=2.97 w=1.2 l=0.15
X1395 a_13918_1126# a_2275_1150# a_14010_1126# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1396 a_29982_17190# row_n[15] a_30474_17552# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1397 vcm a_2275_13198# a_30074_13174# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1398 a_12914_5142# a_2275_5166# a_13006_5142# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1399 VSS row_n[6] a_24354_8194# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1400 VSS row_n[2] a_25358_4178# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1401 a_11398_8516# col_n[8] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X1402 a_34394_8194# rowon_n[6] a_33998_8154# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X1403 a_35398_4178# rowon_n[2] a_35002_4138# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X1404 a_18330_16226# rowon_n[14] a_17934_16186# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X1405 VSS row_n[10] a_28370_12210# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1406 a_33086_11166# a_2475_11190# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1407 a_32386_10202# rowon_n[8] a_31990_10162# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X1408 a_28066_8154# a_2475_8178# a_27974_8154# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X1409 a_8990_2130# a_2475_2154# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1410 a_10998_11166# a_2475_11190# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1411 a_24050_13174# a_2475_13198# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1412 a_19030_7150# a_2475_7174# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1413 VDD rowon_n[12] a_26970_14178# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1414 a_15014_12170# a_2475_12194# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1415 a_23958_9158# a_2275_9182# a_24050_9158# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1416 VSS row_n[5] a_13310_7190# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1417 a_4974_12170# a_2475_12194# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1418 a_17934_3134# a_2275_3158# a_18026_3134# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1419 VDD rowon_n[2] a_35002_4138# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1420 a_25454_4500# col_n[22] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X1421 a_28466_10524# col_n[25] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X1422 a_3366_7512# col_n[0] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X1423 VSS row_n[4] a_29374_6186# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1424 a_10998_1126# a_2475_1150# a_10906_1126# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X1425 VSS row_n[7] a_7286_9198# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1426 a_16418_6508# col_n[13] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X1427 a_33390_18234# VDD a_32994_18194# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X1428 a_26362_17230# col_n[23] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1429 VSS row_n[13] a_30378_15222# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1430 VSS row_n[12] a_34394_14218# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1431 a_31382_11206# col_n[28] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1432 VSS row_n[0] a_6282_2170# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1433 a_2161_4162# sample VDD VDD sky130_fd_pr__pfet_01v8 ad=0.342 pd=2.97 as=0.342 ps=2.97 w=1.2 l=0.15
X1434 a_32386_5182# col_n[29] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1435 a_35002_17190# a_2275_17214# a_35094_17190# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1436 a_11302_14218# rowon_n[12] a_10906_14178# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X1437 a_1957_13198# VDD sample VSS sky130_fd_pr__nfet_01v8 ad=0.171 pd=1.77 as=0.171 ps=1.77 w=0.6 l=0.15
X1438 a_25054_15182# a_2475_15206# a_24962_15182# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X1439 a_7286_12210# col_n[4] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1440 a_17326_12210# col_n[14] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1441 vcm a_2275_12194# a_22042_12170# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1442 a_32082_6146# a_2475_6170# a_31990_6146# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X1443 VSS row_n[3] a_18330_5182# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1444 a_29070_14178# a_2475_14202# a_28978_14178# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X1445 vcm a_2275_11190# a_26058_11166# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1446 a_33998_8154# row_n[6] a_34490_8516# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1447 a_20338_1166# en_bit_n[0] a_19942_1126# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X1448 a_29470_18556# col_n[26] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X1449 VDD rowon_n[14] a_32994_16186# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1450 a_25966_15182# row_n[13] a_26458_15544# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1451 a_30474_13536# col_n[27] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X1452 a_7382_9520# col_n[4] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X1453 a_8386_5504# col_n[5] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X1454 a_24050_1126# a_2475_1150# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1455 a_15014_3134# a_2475_3158# a_14922_3134# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X1456 a_2874_13174# a_2275_13198# a_2966_13174# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1457 a_9994_13174# a_2475_13198# a_9902_13174# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X1458 a_12914_13174# a_2275_13198# a_13006_13174# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1459 a_14010_7150# a_2475_7174# a_13918_7150# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X1460 VDD rowon_n[15] a_8898_17190# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1461 a_6378_14540# col_n[3] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X1462 a_16418_14540# col_n[13] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X1463 VDD rowon_n[6] a_20946_8154# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1464 vcm a_2275_1150# a_12002_1126# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1465 a_31990_3134# row_n[1] a_32482_3496# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1466 vcm a_2275_5166# a_10998_5142# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1467 a_18426_3496# col_n[15] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X1468 a_6890_10162# row_n[8] a_7382_10524# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1469 a_16930_10162# row_n[8] a_17422_10524# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1470 a_23350_7190# rowon_n[5] a_22954_7150# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X1471 a_6982_2130# a_2475_2154# a_6890_2130# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X1472 a_24354_3174# rowon_n[1] a_23958_3134# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X1473 VDD rowon_n[5] a_9902_7150# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1474 a_25358_17230# rowon_n[15] a_24962_17190# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X1475 vcm a_2275_15206# a_14010_15182# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1476 vcm a_2275_15206# a_3970_15182# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1477 a_14314_9198# rowon_n[7] a_13918_9158# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X1478 vcm a_2275_9182# a_22042_9158# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1479 VDD rowon_n[4] a_25966_6146# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1480 a_17934_18194# VDD a_18426_18556# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1481 a_29374_16226# rowon_n[14] a_28978_16186# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X1482 vcm a_2275_14202# a_7986_14178# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1483 vcm a_2275_14202# a_18026_14178# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1484 VSS row_n[11] a_26362_13214# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1485 a_30378_11206# rowon_n[9] a_29982_11166# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X1486 vcm a_2275_7174# a_15014_7150# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1487 vcm a_2275_3158# a_16018_3134# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1488 a_7894_18194# VDD a_8386_18556# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1489 a_30986_2130# a_2275_2154# a_31078_2130# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1490 a_23046_8154# a_2475_8178# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1491 VDD VSS a_23958_1126# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1492 a_22042_14178# a_2475_14202# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1493 VSS en_bit_n[2] a_19334_1166# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1494 VDD rowon_n[13] a_24962_15182# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1495 a_13006_13174# a_2475_13198# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1496 a_35094_13174# a_2475_13198# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1497 a_29374_1166# VSS a_28978_1126# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X1498 a_28370_5182# rowon_n[3] a_27974_5142# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X1499 a_2966_13174# a_2475_13198# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1500 a_25358_12210# col_n[22] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1501 VDD rowon_n[7] a_13918_9158# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1502 VDD rowon_n[3] a_14922_5142# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1503 a_7286_4178# rowon_n[2] a_6890_4138# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X1504 a_26458_11528# col_n[23] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X1505 a_29982_11166# a_2275_11190# a_30074_11166# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1506 a_6282_8194# rowon_n[6] a_5886_8154# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X1507 vcm a_2275_2154# a_7986_2130# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1508 a_24354_18234# col_n[21] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1509 a_24450_14540# col_n[21] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X1510 a_24050_10162# a_2475_10186# a_23958_10162# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X1511 a_2475_9182# a_1957_9182# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.171 pd=1.77 as=0.124 ps=1.01 w=0.6 l=0.15
X1512 a_22042_1126# a_2475_1150# a_21950_1126# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X1513 VSS row_n[8] a_9294_10202# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1514 a_12306_6186# col_n[9] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1515 a_28066_6146# a_2475_6170# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1516 VDD rowon_n[1] a_27974_3134# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1517 a_32994_18194# a_2275_18218# a_33086_18194# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1518 VSS row_n[14] a_18330_16226# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1519 a_23046_16186# a_2475_16210# a_22954_16186# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X1520 a_24962_10162# row_n[8] a_25454_10524# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1521 a_22954_7150# row_n[5] a_23446_7512# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1522 VSS row_n[14] a_8290_16226# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1523 a_33486_7512# col_n[30] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X1524 VDD rowon_n[2] a_6890_4138# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1525 a_23958_16186# row_n[14] a_24450_16548# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1526 a_20946_2130# row_n[0] a_21438_2492# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1527 a_10906_14178# a_2275_14202# a_10998_14178# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1528 a_18026_14178# a_2475_14202# a_17934_14178# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X1529 VDD rowon_n[10] a_7894_12170# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1530 a_31478_2492# col_n[28] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X1531 VDD VDD a_16930_18194# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1532 a_7986_14178# a_2475_14202# a_7894_14178# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X1533 VDD VDD a_6890_18194# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1534 a_26362_2170# col_n[23] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1535 VDD rowon_n[0] a_16930_2130# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1536 a_4274_5182# col_n[1] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1537 vcm a_2275_9182# a_30074_9158# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1538 a_16322_8194# col_n[13] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1539 a_17326_4178# col_n[14] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1540 a_27974_5142# row_n[3] a_28466_5504# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1541 vcm a_2275_10186# a_13006_10162# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1542 a_5886_8154# row_n[6] a_6378_8516# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1543 a_2874_14178# row_n[12] a_3366_14540# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1544 a_12914_14178# row_n[12] a_13406_14540# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1545 a_24354_12210# rowon_n[10] a_23958_12170# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X1546 vcm a_2275_10186# a_2966_10162# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1547 a_21950_10162# a_2275_10186# a_22042_10162# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1548 a_32082_4138# a_2475_4162# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1549 a_28370_11206# rowon_n[9] a_27974_11166# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X1550 a_21038_8154# a_2475_8178# a_20946_8154# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X1551 a_3878_3134# row_n[1] a_4370_3496# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1552 vcm a_2275_16210# a_12002_16186# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1553 a_14010_5142# a_2475_5166# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1554 a_15014_1126# a_2475_1150# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1555 a_16930_4138# row_n[2] a_17422_4500# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1556 a_9994_11166# a_2475_11190# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1557 a_8290_7190# col_n[5] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1558 a_9294_3174# col_n[6] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1559 VDD rowon_n[8] a_23958_10162# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1560 a_9902_7150# a_2275_7174# a_9994_7150# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1561 a_10906_3134# a_2275_3158# a_10998_3134# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1562 VSS row_n[15] a_22346_17230# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1563 a_28978_16186# a_2275_16210# a_29070_16186# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1564 a_33086_14178# a_2475_14202# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1565 VSS row_n[4] a_22346_6186# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1566 a_32386_6186# rowon_n[4] a_31990_6146# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X1567 a_10998_14178# a_2475_14202# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1568 a_23350_13214# col_n[20] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1569 a_26058_6146# a_2475_6170# a_25966_6146# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X1570 a_8898_1126# VDD a_9390_1488# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1571 a_16322_15222# rowon_n[13] a_15926_15182# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X1572 VSS row_n[10] a_13310_12210# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1573 a_6282_15222# rowon_n[13] a_5886_15182# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X1574 a_2161_14202# sample VDD VDD sky130_fd_pr__pfet_01v8 ad=0.342 pd=2.97 as=0.342 ps=2.97 w=1.2 l=0.15
X1575 VSS row_n[10] a_3270_12210# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1576 VSS row_n[3] a_11302_5182# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1577 a_2874_2130# a_2275_2154# a_2966_2130# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1578 a_22442_15544# col_n[19] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X1579 a_35494_14540# VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X1580 VSS row_n[9] a_7286_11206# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1581 VSS row_n[9] a_17326_11206# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1582 a_22042_11166# a_2475_11190# a_21950_11166# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X1583 a_35094_10162# a_2475_10186# a_35002_10162# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X1584 a_14922_5142# a_2275_5166# a_15014_5142# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1585 a_15926_1126# a_2275_1150# a_16018_1126# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1586 a_22954_11166# row_n[9] a_23446_11528# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1587 a_2966_10162# a_2475_10186# a_2874_10162# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X1588 a_13006_10162# a_2475_10186# a_12914_10162# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X1589 VDD VSS sky130_fd_pr__cap_mim_m3_1 l=17.2 w=17.2
X1590 VSS row_n[2] a_27366_4178# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1591 VDD rowon_n[12] a_11910_14178# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1592 a_13406_8516# col_n[10] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X1593 VDD rowon_n[11] a_5886_13174# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1594 VDD rowon_n[11] a_15926_13174# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1595 a_3366_10524# col_n[0] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X1596 a_13406_10524# col_n[10] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X1597 a_11302_17230# col_n[8] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1598 a_11398_3496# col_n[8] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X1599 vcm a_2275_4162# a_20034_4138# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1600 a_15318_16226# col_n[12] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1601 vcm a_2275_16210# a_20034_16186# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1602 a_25966_9158# a_2275_9182# a_26058_9158# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1603 VSS row_n[5] a_15318_7190# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1604 VSS row_n[1] a_16322_3174# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1605 a_30074_4138# a_2475_4162# a_29982_4138# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X1606 a_14010_18194# a_2475_18218# a_13918_18194# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X1607 a_5278_16226# col_n[2] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1608 vcm a_2275_15206# a_33086_15182# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1609 a_27462_4500# col_n[24] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X1610 a_3970_18194# a_2475_18218# a_3878_18194# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X1611 a_5374_7512# col_n[2] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X1612 a_31990_6146# row_n[4] a_32482_6508# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1613 a_5978_7150# a_2475_7174# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1614 a_18426_6508# col_n[15] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X1615 a_12002_5142# a_2475_5166# a_11910_5142# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X1616 a_13006_1126# a_2475_1150# a_12914_1126# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X1617 a_14410_18556# col_n[11] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X1618 a_10906_15182# row_n[13] a_11398_15544# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1619 a_22346_13214# rowon_n[11] a_21950_13174# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X1620 vcm a_2275_11190# a_10998_11166# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1621 VSS row_n[7] a_9294_9198# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1622 a_4370_18556# col_n[1] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X1623 a_35398_12210# rowon_n[10] a_35002_12170# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X1624 a_3366_2492# col_n[0] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X1625 a_16418_1488# col_n[13] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X1626 a_27062_15182# a_2475_15206# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1627 a_23958_12170# a_2275_12194# a_24050_12170# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1628 VSS row_n[0] a_8290_2170# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1629 a_34394_5182# col_n[31] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1630 a_34090_6146# a_2475_6170# a_33998_6146# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X1631 a_1957_7174# VDD sample VSS sky130_fd_pr__nfet_01v8 ad=0.171 pd=1.77 as=0.171 ps=1.77 w=0.6 l=0.15
X1632 VDD rowon_n[9] a_21950_11166# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1633 a_9390_9520# col_n[6] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X1634 a_10298_1166# col_n[7] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1635 a_22346_1166# VSS a_21950_1126# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X1636 a_21342_5182# rowon_n[3] a_20946_5142# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X1637 VDD rowon_n[8] a_35002_10162# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1638 a_17022_3134# a_2475_3158# a_16930_3134# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X1639 VSS VDD a_20338_18234# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1640 VSS row_n[15] a_33390_17230# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1641 a_33998_3134# row_n[1] a_34490_3496# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1642 a_21342_14218# col_n[18] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1643 VDD rowon_n[6] a_22954_8154# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1644 a_6890_7150# a_2275_7174# a_6982_7150# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1645 vcm a_2275_5166# a_13006_5142# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1646 vcm a_2275_1150# a_14010_1126# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1647 a_10298_17230# rowon_n[15] a_9902_17190# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X1648 a_34394_13214# col_n[31] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1649 a_28066_17190# a_2475_17214# a_27974_17190# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X1650 a_4274_16226# rowon_n[14] a_3878_16186# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X1651 a_14314_16226# rowon_n[14] a_13918_16186# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X1652 VSS row_n[11] a_11302_13214# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1653 a_21038_6146# a_2475_6170# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1654 VDD rowon_n[1] a_20946_3134# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1655 a_20434_16548# col_n[17] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X1656 a_29982_14178# a_2275_14202# a_30074_14178# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1657 a_28978_17190# row_n[15] a_29470_17552# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1658 a_33486_15544# col_n[30] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X1659 vcm a_2275_13198# a_29070_13174# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1660 a_10998_11166# a_2475_11190# a_10906_11166# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X1661 a_33086_11166# a_2475_11190# a_32994_11166# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X1662 a_20338_9198# col_n[17] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1663 a_8990_2130# a_2475_2154# a_8898_2130# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X1664 a_26362_3174# rowon_n[1] a_25966_3134# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X1665 a_5886_15182# a_2275_15206# a_5978_15182# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1666 a_15926_15182# a_2275_15206# a_16018_15182# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1667 VSS row_n[7] a_30378_9198# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1668 VDD rowon_n[5] a_11910_7150# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1669 a_4274_6186# rowon_n[4] a_3878_6146# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X1670 VDD rowon_n[13] a_9902_15182# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1671 a_33998_11166# row_n[9] a_34490_11528# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1672 a_16322_9198# rowon_n[7] a_15926_9158# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X1673 vcm a_2275_9182# a_24050_9158# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1674 a_19030_7150# a_2475_7174# a_18938_7150# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X1675 a_10298_12210# col_n[7] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1676 a_11398_11528# col_n[8] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X1677 VDD rowon_n[4] a_27974_6146# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1678 VDD rowon_n[0] a_9902_2130# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1679 vcm a_2275_3158# a_18026_3134# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1680 VDD VSS a_25966_1126# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1681 a_32994_2130# a_2275_2154# a_33086_2130# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1682 a_15318_2170# rowon_n[0] a_14922_2130# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X1683 a_26058_4138# a_2475_4162# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1684 a_19942_9158# row_n[7] a_20434_9520# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1685 a_25054_8154# a_2475_8178# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1686 a_20946_5142# row_n[3] a_21438_5504# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1687 vcm a_2275_16210# a_31078_16186# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1688 a_30474_9520# col_n[27] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X1689 a_31478_5504# col_n[28] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X1690 a_9902_10162# row_n[8] a_10394_10524# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1691 vcm a_2275_17214# a_17022_17190# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1692 VDD rowon_n[7] a_15926_9158# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1693 a_8290_8194# rowon_n[6] a_7894_8154# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X1694 VDD rowon_n[3] a_16930_5142# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1695 a_9294_4178# rowon_n[2] a_8898_4138# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X1696 vcm a_2275_17214# a_6982_17190# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1697 a_20338_14218# rowon_n[12] a_19942_14178# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X1698 a_21038_17190# a_2475_17214# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1699 a_14314_6186# col_n[11] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1700 a_24050_1126# a_2475_1150# a_23958_1126# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X1701 a_25054_16186# a_2475_16210# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1702 a_21950_13174# a_2275_13198# a_22042_13174# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1703 a_24962_7150# row_n[5] a_25454_7512# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1704 a_16018_15182# a_2475_15206# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1705 a_35494_7512# VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X1706 a_3878_6146# row_n[4] a_4370_6508# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1707 a_5978_15182# a_2475_15206# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1708 VDD rowon_n[2] a_8898_4138# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1709 a_9994_14178# a_2475_14202# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1710 VSS row_n[10] a_32386_12210# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1711 a_22954_2130# row_n[0] a_23446_2492# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1712 a_33486_2492# col_n[30] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X1713 VSS VDD a_31382_18234# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1714 a_2475_11190# a_1957_11190# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.342 pd=2.97 as=0.249 ps=1.62 w=1.2 l=0.15
X1715 a_28370_2170# col_n[25] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1716 a_12002_3134# a_2475_3158# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1717 VDD rowon_n[12] a_30986_14178# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1718 a_27062_12170# a_2475_12194# a_26970_12170# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X1719 a_3270_11206# rowon_n[9] a_2874_11166# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X1720 a_13310_11206# rowon_n[9] a_12914_11166# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X1721 a_6282_5182# col_n[3] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1722 a_7286_1166# col_n[4] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1723 a_32386_14218# col_n[29] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1724 a_19334_4178# col_n[16] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1725 a_26058_18194# a_2475_18218# a_25966_18194# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X1726 a_27974_12170# row_n[10] a_28466_12532# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1727 a_32482_10524# col_n[29] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X1728 a_18330_8194# col_n[15] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1729 VSS row_n[2] a_20338_4178# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1730 a_26970_18194# VDD a_27462_18556# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1731 a_30378_17230# col_n[27] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1732 vcm a_2275_14202# a_27062_14178# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1733 a_7894_8154# row_n[6] a_8386_8516# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1734 a_30378_4178# rowon_n[2] a_29982_4138# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X1735 a_13918_16186# a_2275_16210# a_14010_16186# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1736 a_31478_16548# col_n[28] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X1737 vcm a_2275_2154# a_31078_2130# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1738 a_34090_4138# a_2475_4162# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1739 a_3878_16186# a_2275_16210# a_3970_16186# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1740 a_23046_8154# a_2475_8178# a_22954_8154# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X1741 a_3970_2130# a_2475_2154# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1742 a_5886_3134# row_n[1] a_6378_3496# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1743 a_17022_1126# a_2475_1150# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1744 vcm a_2275_17214# a_25054_17190# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1745 a_18938_4138# row_n[2] a_19430_4500# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1746 vcm a_2275_11190# a_30074_11166# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1747 a_20434_4500# col_n[17] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X1748 a_29982_15182# row_n[13] a_30474_15544# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1749 a_12914_3134# a_2275_3158# a_13006_3134# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1750 VDD rowon_n[2] a_29982_4138# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1751 vcm a_2275_12194# a_16018_12170# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1752 VSS row_n[4] a_24354_6186# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1753 vcm a_2275_12194# a_5978_12170# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1754 a_11398_6508# col_n[8] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X1755 a_34394_6186# rowon_n[4] a_33998_6146# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X1756 a_18330_14218# rowon_n[12] a_17934_14178# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X1757 VSS row_n[8] a_28370_10202# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1758 a_19030_17190# a_2475_17214# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1759 a_28978_11166# a_2275_11190# a_29070_11166# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1760 a_28066_6146# a_2475_6170# a_27974_6146# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X1761 a_20034_12170# a_2475_12194# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1762 a_19030_5142# a_2475_5166# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1763 VDD rowon_n[10] a_26970_12170# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1764 VSS row_n[3] a_13310_5182# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1765 a_4882_2130# a_2275_2154# a_4974_2130# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1766 a_17934_1126# a_2275_1150# a_18026_1126# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1767 a_3366_5504# col_n[0] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X1768 VSS row_n[2] a_29374_4178# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1769 a_15414_8516# col_n[12] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X1770 a_16018_8154# a_2475_8178# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1771 VSS VDD a_29374_18234# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1772 a_33390_16226# rowon_n[14] a_32994_16186# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X1773 a_26362_15222# col_n[23] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1774 VSS row_n[11] a_30378_13214# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1775 VSS a_2161_6170# a_2275_6170# VSS sky130_fd_pr__nfet_01v8 ad=0.124 pd=1.01 as=0.171 ps=1.77 w=0.6 l=0.15
X1776 a_13406_3496# col_n[10] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X1777 a_19334_7190# rowon_n[5] a_18938_7150# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X1778 a_31382_7190# col_n[28] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1779 a_32386_3174# col_n[29] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1780 a_9294_17230# rowon_n[15] a_8898_17190# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X1781 a_35002_15182# a_2275_15206# a_35094_15182# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1782 a_25454_17552# col_n[22] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X1783 a_21950_14178# row_n[12] a_22442_14540# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1784 a_25054_13174# a_2475_13198# a_24962_13174# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X1785 a_7286_10202# col_n[4] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1786 a_17326_10202# col_n[14] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1787 vcm a_2275_10186# a_22042_10162# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1788 a_27974_9158# a_2275_9182# a_28066_9158# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1789 VSS row_n[5] a_17326_7190# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1790 VSS row_n[1] a_18330_3174# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1791 a_32082_4138# a_2475_4162# a_31990_4138# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X1792 a_5978_12170# a_2475_12194# a_5886_12170# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X1793 a_16018_12170# a_2475_12194# a_15926_12170# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X1794 a_33998_6146# row_n[4] a_34490_6508# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1795 a_29470_4500# col_n[26] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X1796 a_29470_16548# col_n[26] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X1797 a_25966_13174# row_n[11] a_26458_13536# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1798 a_30474_11528# col_n[27] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X1799 a_7382_7512# col_n[4] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X1800 a_7986_7150# a_2475_7174# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1801 a_14010_5142# a_2475_5166# a_13918_5142# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X1802 a_15014_1126# a_2475_1150# a_14922_1126# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X1803 a_9994_11166# a_2475_11190# a_9902_11166# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X1804 a_26970_2130# a_2275_2154# a_27062_2130# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1805 VDD rowon_n[13] a_8898_15182# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1806 a_6378_12532# col_n[3] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X1807 a_16418_12532# col_n[13] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X1808 VDD rowon_n[4] a_20946_6146# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1809 a_31990_1126# VDD a_32482_1488# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1810 a_5374_2492# col_n[2] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X1811 vcm a_2275_3158# a_10998_3134# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1812 vcm a_2275_7174# a_9994_7150# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1813 a_18426_1488# en_bit_n[1] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X1814 a_16930_8154# a_2275_8178# a_17022_8154# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1815 a_18330_18234# col_n[15] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1816 vcm a_2275_18218# a_23046_18194# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1817 VDD VSS VSS sky130_fd_pr__cap_var_lvt w=16.4 l=16
X1818 a_8290_18234# col_n[5] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1819 a_24354_1166# VSS a_23958_1126# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X1820 a_23350_5182# rowon_n[3] a_22954_5142# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X1821 a_27062_10162# a_2475_10186# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1822 VDD rowon_n[3] a_9902_5142# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1823 a_13918_17190# row_n[15] a_14410_17552# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1824 a_25358_15222# rowon_n[13] a_24962_15182# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X1825 vcm a_2275_13198# a_14010_13174# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1826 a_2161_9182# sample VSS VSS sky130_fd_pr__nfet_01v8 ad=0.171 pd=1.77 as=0.171 ps=1.77 w=0.6 l=0.15
X1827 vcm a_2275_2154# a_2966_2130# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1828 a_3878_17190# row_n[15] a_4370_17552# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1829 vcm a_2275_13198# a_3970_13174# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1830 vcm a_2275_1150# a_16018_1126# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1831 a_17934_16186# row_n[14] a_18426_16548# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1832 a_29374_14218# rowon_n[12] a_28978_14178# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X1833 VSS row_n[9] a_26362_11206# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1834 a_8898_7150# a_2275_7174# a_8990_7150# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1835 vcm a_2275_5166# a_15014_5142# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1836 a_7894_16186# row_n[14] a_8386_16548# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1837 a_31078_12170# a_2475_12194# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1838 a_23046_6146# a_2475_6170# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1839 VDD rowon_n[1] a_22954_3134# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1840 VDD rowon_n[11] a_24962_13174# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1841 a_28370_3174# rowon_n[1] a_27974_3134# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X1842 a_25358_10202# col_n[22] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1843 VSS row_n[7] a_32386_9198# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1844 VDD rowon_n[5] a_13918_7150# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1845 a_6282_6186# rowon_n[4] a_5886_6146# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X1846 a_24354_16226# col_n[21] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1847 vcm a_2275_9182# a_26058_9158# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1848 a_8290_12210# rowon_n[10] a_7894_12170# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X1849 a_15926_10162# a_2275_10186# a_16018_10162# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1850 VSS row_n[0] a_31382_2170# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1851 a_21342_2170# col_n[18] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1852 VDD rowon_n[0] a_11910_2130# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1853 a_24450_12532# col_n[21] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X1854 a_5886_10162# a_2275_10186# a_5978_10162# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1855 a_2475_7174# a_1957_7174# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.171 pd=1.77 as=0.124 ps=1.01 w=0.6 l=0.15
X1856 a_5978_7150# a_2475_7174# a_5886_7150# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X1857 a_7286_18234# VDD a_6890_18194# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X1858 a_17326_18234# VDD a_16930_18194# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X1859 a_11302_8194# col_n[8] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1860 a_27062_8154# a_2475_8178# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1861 a_35002_2130# a_2275_2154# a_35094_2130# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1862 VDD VSS a_27974_1126# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1863 a_17326_2170# rowon_n[0] a_16930_2130# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X1864 a_28066_4138# a_2475_4162# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1865 a_12306_4178# col_n[9] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1866 a_23446_18556# col_n[20] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X1867 a_32994_16186# a_2275_16210# a_33086_16186# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1868 VSS row_n[12] a_18330_14218# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1869 a_23046_14178# a_2475_14202# a_22954_14178# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X1870 a_22954_5142# row_n[3] a_23446_5504# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1871 VSS row_n[12] a_8290_14218# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1872 a_32482_9520# col_n[29] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X1873 a_33486_5504# col_n[30] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X1874 a_18938_17190# a_2275_17214# a_19030_17190# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1875 a_8898_17190# a_2275_17214# a_8990_17190# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1876 VDD rowon_n[8] a_7894_10162# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1877 VDD VSS sky130_fd_pr__cap_mim_m3_1 l=17.2 w=17.2
X1878 VDD rowon_n[14] a_16930_16186# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1879 VDD rowon_n[14] a_6890_16186# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1880 a_11910_4138# row_n[2] a_12402_4500# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1881 vcm a_2275_12194# a_35094_12170# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1882 a_3270_7190# col_n[0] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1883 a_4274_3174# col_n[1] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1884 a_16322_6186# col_n[13] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1885 vcm a_2275_18218# a_34090_18194# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1886 vcm a_2275_7174# a_6982_7150# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1887 a_12914_12170# row_n[10] a_13406_12532# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1888 a_5886_6146# row_n[4] a_6378_6508# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1889 a_2874_12170# row_n[10] a_3366_12532# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1890 a_25054_11166# a_2475_11190# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1891 a_24354_10202# rowon_n[8] a_23958_10162# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X1892 a_16018_10162# a_2475_10186# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1893 a_21038_6146# a_2475_6170# a_20946_6146# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X1894 a_35494_2492# VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X1895 a_3878_1126# en_C0_n a_4370_1488# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1896 a_24962_2130# row_n[0] a_25454_2492# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1897 a_11910_18194# VDD a_12402_18556# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1898 vcm a_2275_14202# a_12002_14178# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1899 a_5978_10162# a_2475_10186# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1900 VDD rowon_n[12] a_18938_14178# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1901 a_29070_12170# a_2475_12194# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1902 a_14010_3134# a_2475_3158# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1903 a_8290_5182# col_n[5] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1904 a_9294_1166# col_n[6] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1905 a_28066_18194# a_2475_18218# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1906 vcm a_2275_17214# a_9994_17190# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1907 a_9902_5142# a_2275_5166# a_9994_5142# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1908 a_10906_1126# a_2275_1150# a_10998_1126# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1909 VSS row_n[2] a_22346_4178# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1910 VSS row_n[13] a_22346_15222# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1911 a_28978_14178# a_2275_14202# a_29070_14178# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1912 a_32386_4178# rowon_n[2] a_31990_4138# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X1913 a_31382_8194# rowon_n[6] a_30986_8154# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X1914 vcm a_2275_2154# a_33086_2130# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1915 a_23350_11206# col_n[20] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1916 a_25054_8154# a_2475_8178# a_24962_8154# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X1917 a_26058_4138# a_2475_4162# a_25966_4138# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X1918 a_7894_3134# row_n[1] a_8386_3496# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1919 VDD rowon_n[15] a_20946_17190# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1920 a_16322_13214# rowon_n[11] a_15926_13174# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X1921 VSS row_n[8] a_13310_10202# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1922 a_6282_13214# rowon_n[11] a_5886_13174# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X1923 a_3878_11166# a_2275_11190# a_3970_11166# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1924 a_13918_11166# a_2275_11190# a_14010_11166# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1925 VSS row_n[8] a_3270_10202# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1926 a_20946_9158# a_2275_9182# a_21038_9158# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1927 VSS row_n[5] a_10298_7190# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1928 VSS row_n[1] a_11302_3174# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1929 a_22442_13536# col_n[19] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X1930 a_35494_12532# VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X1931 a_31078_9158# a_2475_9182# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1932 a_14922_3134# a_2275_3158# a_15014_3134# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1933 a_22442_4500# col_n[19] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X1934 a_17934_12170# a_2275_12194# a_18026_12170# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1935 VDD rowon_n[2] a_31990_4138# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1936 a_7894_12170# a_2275_12194# a_7986_12170# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1937 VDD rowon_n[10] a_11910_12170# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1938 a_13406_6508# col_n[10] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X1939 VSS row_n[7] a_4274_9198# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1940 a_6890_18194# a_2275_18218# a_6982_18194# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1941 a_16930_18194# a_2275_18218# a_17022_18194# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1942 VDD rowon_n[9] a_5886_11166# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1943 VDD rowon_n[9] a_15926_11166# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1944 VSS VDD a_14314_18234# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1945 a_11302_15222# col_n[8] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1946 a_11398_1488# col_n[8] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X1947 VSS VDD a_4274_18234# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1948 a_32082_17190# a_2475_17214# a_31990_17190# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X1949 VSS row_n[0] a_3270_2170# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1950 a_19942_18194# VDD a_20434_18556# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1951 a_15318_14218# col_n[12] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1952 vcm a_2275_14202# a_20034_14178# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1953 VSS row_n[3] a_15318_5182# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1954 VSS VDD a_16322_1166# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1955 a_32994_17190# row_n[15] a_33486_17552# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1956 a_14010_16186# a_2475_16210# a_13918_16186# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X1957 a_5278_14218# col_n[2] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1958 vcm a_2275_13198# a_33086_13174# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1959 a_10394_17552# col_n[7] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X1960 a_3970_16186# a_2475_16210# a_3878_16186# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X1961 a_4370_9520# col_n[1] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X1962 VDD rowon_n[6] a_18938_8154# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1963 a_30986_8154# row_n[6] a_31478_8516# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1964 a_5374_5504# col_n[2] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X1965 a_17422_8516# col_n[14] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X1966 a_5978_5142# a_2475_5166# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1967 a_12002_3134# a_2475_3158# a_11910_3134# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X1968 a_14410_16548# col_n[11] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X1969 a_10906_13174# row_n[11] a_11398_13536# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1970 a_22346_11206# rowon_n[9] a_21950_11166# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X1971 a_18026_8154# a_2475_8178# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1972 analog_in sw ctop VSS sky130_fd_pr__nfet_01v8 ad=0.275 pd=2.19 as=0.551 ps=4.38 w=1.9 l=0.22
X1973 a_4370_16548# col_n[1] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X1974 a_35398_10202# rowon_n[8] a_35002_10162# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X1975 a_15414_3496# col_n[12] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X1976 a_27062_13174# a_2475_13198# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1977 VSS row_n[7] a_26362_9198# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1978 a_33390_7190# col_n[30] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1979 a_34394_3174# col_n[31] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1980 a_18026_12170# a_2475_12194# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1981 a_34090_4138# a_2475_4162# a_33998_4138# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X1982 a_7986_12170# a_2475_12194# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1983 a_1957_5166# VDD sample VSS sky130_fd_pr__nfet_01v8 ad=0.171 pd=1.77 as=0.171 ps=1.77 w=0.6 l=0.15
X1984 a_9390_7512# col_n[6] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X1985 a_3970_2130# a_2475_2154# a_3878_2130# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X1986 a_21342_3174# rowon_n[1] a_20946_3134# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X1987 a_35002_10162# a_2275_10186# a_35094_10162# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1988 a_9994_7150# a_2475_7174# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1989 a_17022_1126# a_2475_1150# a_16930_1126# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X1990 a_29374_17230# col_n[26] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1991 VSS row_n[14] a_20338_16226# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1992 VSS row_n[13] a_33390_15222# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1993 a_11302_9198# rowon_n[7] a_10906_9158# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X1994 a_28978_2130# a_2275_2154# a_29070_2130# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1995 VDD rowon_n[4] a_22954_6146# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1996 a_6890_5142# a_2275_5166# a_6982_5142# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X1997 a_7382_2492# col_n[4] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X1998 vcm a_2275_3158# a_13006_3134# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1999 a_10298_15222# rowon_n[13] a_9902_15182# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X2000 a_34394_11206# col_n[31] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2001 a_26458_9520# col_n[23] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X2002 a_18938_8154# a_2275_8178# a_19030_8154# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2003 a_24962_18194# a_2275_18218# a_25054_18194# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2004 VDD VSS a_20946_1126# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2005 a_10298_2170# rowon_n[0] a_9902_2130# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X2006 a_21038_4138# a_2475_4162# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2007 VDD rowon_n[15] a_31990_17190# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2008 a_28066_15182# a_2475_15206# a_27974_15182# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X2009 a_4274_14218# rowon_n[12] a_3878_14178# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X2010 a_14314_14218# rowon_n[12] a_13918_14178# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X2011 VSS row_n[9] a_11302_11206# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X2012 a_20034_8154# a_2475_8178# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2013 a_28978_15182# row_n[13] a_29470_15544# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2014 a_33486_13536# col_n[30] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X2015 vcm a_2275_11190# a_29070_11166# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2016 VDD rowon_n[3] a_11910_5142# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2017 a_26362_1166# VSS a_25966_1126# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X2018 a_5886_13174# a_2275_13198# a_5978_13174# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2019 a_15926_13174# a_2275_13198# a_16018_13174# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2020 VDD rowon_n[7] a_10906_9158# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2021 a_3270_8194# rowon_n[6] a_2874_8154# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X2022 a_4274_4178# rowon_n[2] a_3878_4138# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X2023 VDD rowon_n[11] a_9902_13174# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2024 vcm a_2275_2154# a_4974_2130# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2025 a_19030_5142# a_2475_5166# a_18938_5142# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X2026 a_10298_10202# col_n[7] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2027 vcm a_2275_1150# a_18026_1126# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2028 a_30074_18194# a_2475_18218# a_29982_18194# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X2029 a_16018_8154# a_2475_8178# a_15926_8154# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X2030 a_19942_7150# row_n[5] a_20434_7512# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2031 a_25054_6146# a_2475_6170# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2032 a_30986_18194# VDD a_31478_18556# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2033 vcm a_2275_14202# a_31078_14178# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2034 a_30474_7512# col_n[27] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X2035 VDD rowon_n[2] a_3878_4138# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2036 vcm a_2275_15206# a_17022_15182# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2037 VSS row_n[7] a_34394_9198# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X2038 VDD rowon_n[5] a_15926_7150# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2039 a_8290_6186# rowon_n[4] a_7894_6146# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X2040 vcm a_2275_15206# a_6982_15182# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2041 vcm a_2275_9182# a_28066_9158# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2042 a_23350_2170# col_n[20] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2043 VDD rowon_n[0] a_13918_2130# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2044 a_21038_15182# a_2475_15206# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2045 VSS row_n[0] a_33390_2170# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X2046 a_25358_8194# rowon_n[6] a_24962_8154# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X2047 a_7986_7150# a_2475_7174# a_7894_7150# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X2048 a_14314_4178# col_n[11] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2049 VSS a_2161_16210# a_2275_16210# VSS sky130_fd_pr__nfet_01v8 ad=0.124 pd=1.01 as=0.171 ps=1.77 w=0.6 l=0.15
X2050 a_25054_14178# a_2475_14202# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2051 a_13310_8194# col_n[10] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2052 a_29070_8154# a_2475_8178# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2053 vcm a_2275_2154# a_27062_2130# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2054 a_24962_5142# row_n[3] a_25454_5504# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2055 a_16018_13174# a_2475_13198# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2056 a_34490_9520# col_n[31] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X2057 a_35494_5504# VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X2058 a_5978_13174# a_2475_13198# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2059 a_28370_12210# col_n[25] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2060 VSS row_n[8] a_32386_10202# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X2061 a_2874_8154# row_n[6] a_3366_8516# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2062 vcm a_2275_8178# a_17022_8154# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2063 a_32994_11166# a_2275_11190# a_33086_11166# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2064 a_31990_7150# a_2275_7174# a_32082_7150# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2065 a_27366_18234# col_n[24] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2066 VSS row_n[14] a_31382_16226# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X2067 a_12002_1126# a_2475_1150# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2068 a_27462_14540# col_n[24] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X2069 VDD rowon_n[10] a_30986_12170# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2070 a_27062_10162# a_2475_10186# a_26970_10162# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X2071 a_6282_3174# col_n[3] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2072 a_13918_4138# row_n[2] a_14410_4500# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2073 a_5278_7190# col_n[2] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2074 a_26058_16186# a_2475_16210# a_25966_16186# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X2075 a_27974_10162# row_n[8] a_28466_10524# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2076 a_18330_6186# col_n[15] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2077 VDD VDD a_29982_18194# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2078 vcm a_2275_7174# a_8990_7150# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2079 a_26970_16186# row_n[14] a_27462_16548# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2080 a_30378_15222# col_n[27] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2081 a_7894_6146# row_n[4] a_8386_6508# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2082 VDD a_2161_17214# a_2275_17214# VDD sky130_fd_pr__pfet_01v8 ad=0.249 pd=1.62 as=0.342 ps=2.97 w=1.2 l=0.15
X2083 a_13918_14178# a_2275_14202# a_14010_14178# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2084 a_3878_14178# a_2275_14202# a_3970_14178# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2085 a_23046_6146# a_2475_6170# a_22954_6146# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X2086 a_5886_1126# VDD a_6378_1488# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2087 vcm a_2275_15206# a_25054_15182# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2088 a_8990_17190# a_2475_17214# a_8898_17190# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X2089 a_29982_13174# row_n[11] a_30474_13536# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2090 a_12914_1126# a_2275_1150# a_13006_1126# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2091 vcm a_2275_10186# a_16018_10162# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2092 VSS row_n[2] a_24354_4178# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X2093 a_9390_17552# col_n[6] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X2094 a_5886_14178# row_n[12] a_6378_14540# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2095 a_15926_14178# row_n[12] a_16418_14540# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2096 a_27366_12210# rowon_n[10] a_26970_12170# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X2097 vcm a_2275_10186# a_5978_10162# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2098 a_10394_8516# col_n[7] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X2099 a_10998_8154# a_2475_8178# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2100 a_33390_8194# rowon_n[6] a_32994_8154# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X2101 a_27366_7190# col_n[24] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2102 a_34394_4178# rowon_n[2] a_33998_4138# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X2103 vcm a_2275_2154# a_35094_2130# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2104 a_19030_15182# a_2475_15206# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2105 a_27062_8154# a_2475_8178# a_26970_8154# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X2106 a_28066_4138# a_2475_4162# a_27974_4138# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X2107 a_19030_3134# a_2475_3158# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2108 VDD rowon_n[8] a_26970_10162# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2109 a_22954_9158# a_2275_9182# a_23046_9158# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2110 VSS row_n[5] a_12306_7190# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X2111 VSS row_n[1] a_13310_3174# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X2112 a_33086_9158# a_2475_9182# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2113 VDD rowon_n[2] a_33998_4138# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2114 a_24450_4500# col_n[21] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X2115 VSS row_n[15] a_25358_17230# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X2116 a_2966_7150# a_2475_7174# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2117 a_15414_6508# col_n[12] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X2118 a_16018_6146# a_2475_6170# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2119 a_21950_2130# a_2275_2154# a_22042_2130# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2120 VSS row_n[14] a_29374_16226# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X2121 a_33390_14218# rowon_n[12] a_32994_14178# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X2122 a_26362_13214# col_n[23] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2123 VSS row_n[9] a_30378_11206# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X2124 VSS a_2161_4162# a_2275_4162# VSS sky130_fd_pr__nfet_01v8 ad=0.124 pd=1.01 as=0.171 ps=1.77 w=0.6 l=0.15
X2125 a_13406_1488# col_n[10] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X2126 a_12002_17190# a_2475_17214# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2127 a_34090_17190# a_2475_17214# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2128 VSS row_n[10] a_16322_12210# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X2129 a_21038_12170# a_2475_12194# a_20946_12170# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X2130 a_11910_8154# a_2275_8178# a_12002_8154# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2131 a_32386_1166# col_n[29] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2132 a_31382_5182# col_n[28] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2133 a_19334_5182# rowon_n[3] a_18938_5142# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X2134 a_9294_15222# rowon_n[13] a_8898_15182# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X2135 a_35002_13174# a_2275_13198# a_35094_13174# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2136 VSS row_n[10] a_6282_12210# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X2137 VSS row_n[0] a_5278_2170# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X2138 VDD VDD a_27974_18194# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2139 a_25454_15544# col_n[22] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X2140 a_21950_12170# row_n[10] a_22442_12532# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2141 a_25054_11166# a_2475_11190# a_24962_11166# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X2142 VSS row_n[3] a_17326_5182# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X2143 VSS en_bit_n[1] a_18330_1166# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X2144 a_5978_10162# a_2475_10186# a_5886_10162# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X2145 a_16018_10162# a_2475_10186# a_15926_10162# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X2146 VDD rowon_n[12] a_14922_14178# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2147 a_25966_11166# row_n[9] a_26458_11528# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2148 a_32994_8154# row_n[6] a_33486_8516# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2149 a_7382_5504# col_n[4] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X2150 a_7986_5142# a_2475_5166# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2151 a_14010_3134# a_2475_3158# a_13918_3134# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X2152 VDD rowon_n[12] a_4882_14178# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2153 VDD rowon_n[11] a_8898_13174# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2154 a_6378_10524# col_n[3] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X2155 a_16418_10524# col_n[13] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X2156 vcm a_2275_1150# a_10998_1126# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2157 a_30986_3134# row_n[1] a_31478_3496# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2158 VDD rowon_n[1] a_18938_3134# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2159 a_14314_17230# col_n[11] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2160 a_3878_7150# a_2275_7174# a_3970_7150# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2161 vcm a_2275_5166# a_9994_5142# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2162 a_4274_17230# col_n[1] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2163 a_16930_6146# a_2275_6170# a_17022_6146# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2164 a_17422_3496# col_n[14] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X2165 a_18330_16226# col_n[15] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2166 vcm a_2275_16210# a_23046_16186# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2167 VSS row_n[7] a_28370_9198# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X2168 a_35398_7190# VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2169 a_9902_18194# a_2275_18218# a_9994_18194# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2170 a_17022_18194# a_2475_18218# a_16930_18194# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X2171 a_8290_16226# col_n[5] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2172 a_1957_9182# VSS sample VDD sky130_fd_pr__pfet_01v8 ad=0.342 pd=2.97 as=0.342 ps=2.97 w=1.2 l=0.15
X2173 a_6982_18194# a_2475_18218# a_6890_18194# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X2174 a_23350_3174# rowon_n[1] a_22954_3134# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X2175 a_17422_18556# col_n[14] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X2176 a_13918_15182# row_n[13] a_14410_15544# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2177 a_25358_13214# rowon_n[11] a_24962_13174# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X2178 a_1957_12194# VSS sample VDD sky130_fd_pr__pfet_01v8 ad=0.342 pd=2.97 as=0.342 ps=2.97 w=1.2 l=0.15
X2179 vcm a_2275_11190# a_14010_11166# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2180 a_2161_7174# sample VSS VSS sky130_fd_pr__nfet_01v8 ad=0.171 pd=1.77 as=0.171 ps=1.77 w=0.6 l=0.15
X2181 a_7382_18556# col_n[4] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X2182 a_3878_15182# row_n[13] a_4370_15544# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2183 vcm a_2275_11190# a_3970_11166# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2184 a_13310_9198# rowon_n[7] a_12914_9158# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X2185 vcm a_2275_9182# a_21038_9158# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2186 a_31078_9158# a_2475_9182# a_30986_9158# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X2187 a_8898_5142# a_2275_5166# a_8990_5142# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2188 a_9390_2492# col_n[6] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X2189 vcm a_2275_3158# a_15014_3134# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2190 a_28466_9520# col_n[25] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X2191 a_26970_12170# a_2275_12194# a_27062_12170# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2192 a_22042_8154# a_2475_8178# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2193 VDD VSS a_22954_1126# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2194 a_29982_2130# a_2275_2154# a_30074_2130# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2195 a_12306_2170# rowon_n[0] a_11910_2130# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X2196 a_23046_4138# a_2475_4162# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2197 VSS row_n[10] a_24354_12210# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X2198 VDD rowon_n[9] a_24962_11166# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2199 a_28370_1166# VSS a_27974_1126# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X2200 VDD rowon_n[7] a_12914_9158# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2201 VDD rowon_n[3] a_13918_5142# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2202 a_6282_4178# rowon_n[2] a_5886_4138# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X2203 VSS VDD a_23350_18234# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X2204 VDD rowon_n[12] a_22954_14178# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2205 a_24354_14218# col_n[21] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2206 a_19030_12170# a_2475_12194# a_18938_12170# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X2207 a_8290_10202# rowon_n[8] a_7894_10162# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X2208 a_32082_18194# a_2475_18218# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2209 a_24450_10524# col_n[21] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X2210 a_2475_5166# a_1957_5166# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.171 pd=1.77 as=0.124 ps=1.01 w=0.6 l=0.15
X2211 a_5978_5142# a_2475_5166# a_5886_5142# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X2212 a_7286_16226# rowon_n[14] a_6890_16186# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X2213 a_17326_16226# rowon_n[14] a_16930_16186# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X2214 a_18026_8154# a_2475_8178# a_17934_8154# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X2215 a_11302_6186# col_n[8] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2216 a_27062_6146# a_2475_6170# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2217 a_23446_16548# col_n[20] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X2218 a_32994_14178# a_2275_14202# a_33086_14178# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2219 a_32482_7512# col_n[29] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X2220 VDD rowon_n[2] a_5886_4138# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2221 a_18938_15182# a_2275_15206# a_19030_15182# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2222 a_8898_15182# a_2275_15206# a_8990_15182# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2223 a_30474_2492# col_n[27] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X2224 a_19942_2130# row_n[0] a_20434_2492# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2225 a_3270_12210# col_n[0] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2226 a_13310_12210# col_n[10] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2227 a_25358_2170# col_n[22] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2228 VDD rowon_n[0] a_15926_2130# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2229 a_12306_18234# col_n[9] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2230 a_35002_14178# row_n[12] a_35494_14540# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2231 vcm a_2275_10186# a_35094_10162# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2232 a_27366_8194# rowon_n[6] a_26970_8154# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X2233 a_9994_7150# a_2475_7174# a_9902_7150# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X2234 a_3270_5182# col_n[0] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2235 VSS row_n[0] a_35398_2170# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X2236 a_4274_1166# en_C0_n VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2237 a_15318_8194# col_n[12] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2238 vcm a_2275_2154# a_29070_2130# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2239 a_16322_4178# col_n[13] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2240 vcm a_2275_16210# a_34090_16186# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2241 a_12402_14540# col_n[9] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X2242 a_21038_10162# a_2475_10186# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2243 vcm a_2275_5166# a_6982_5142# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2244 a_12914_10162# row_n[8] a_13406_10524# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2245 a_4882_8154# row_n[6] a_5374_8516# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2246 VSS a_2161_11190# a_2275_11190# VSS sky130_fd_pr__nfet_01v8 ad=0.124 pd=1.01 as=0.171 ps=1.77 w=0.6 l=0.15
X2247 a_2874_10162# row_n[8] a_3366_10524# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2248 vcm a_2275_8178# a_19030_8154# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2249 a_20034_8154# a_2475_8178# a_19942_8154# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X2250 a_21038_4138# a_2475_4162# a_20946_4138# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X2251 a_11910_16186# row_n[14] a_12402_16548# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2252 a_33998_7150# a_2275_7174# a_34090_7150# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2253 a_2874_3134# row_n[1] a_3366_3496# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2254 VDD rowon_n[10] a_18938_12170# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2255 a_14010_1126# a_2475_1150# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2256 a_8290_3174# col_n[5] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2257 a_15926_4138# row_n[2] a_16418_4500# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2258 a_21342_17230# rowon_n[15] a_20946_17190# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X2259 a_28066_16186# a_2475_16210# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2260 vcm a_2275_15206# a_9994_15182# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2261 a_9902_3134# a_2275_3158# a_9994_3134# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2262 VSS row_n[11] a_22346_13214# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X2263 a_31382_6186# rowon_n[4] a_30986_6146# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X2264 VSS row_n[10] a_35398_12210# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X2265 a_12306_12210# rowon_n[10] a_11910_12170# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X2266 a_25054_6146# a_2475_6170# a_24962_6146# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X2267 a_7894_1126# VDD a_8386_1488# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2268 VDD rowon_n[13] a_20946_15182# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2269 a_6282_11206# rowon_n[9] a_5886_11166# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X2270 a_16322_11206# rowon_n[9] a_15926_11166# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X2271 a_26970_8154# row_n[6] a_27462_8516# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2272 VDD rowon_n[12] a_33998_14178# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2273 VSS row_n[3] a_10298_5182# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X2274 VSS VDD a_11302_1166# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X2275 a_22442_11528# col_n[19] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X2276 a_35494_10524# VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X2277 a_14922_1126# a_2275_1150# a_15014_1126# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2278 a_20338_18234# col_n[17] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2279 a_33390_17230# col_n[30] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2280 VDD rowon_n[8] a_11910_10162# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2281 a_12402_8516# col_n[9] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X2282 a_13006_8154# a_2475_8178# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2283 a_29374_7190# col_n[26] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2284 VSS row_n[15] a_10298_17230# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X2285 a_6890_16186# a_2275_16210# a_6982_16186# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2286 a_16930_16186# a_2275_16210# a_17022_16186# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2287 a_29070_8154# a_2475_8178# a_28978_8154# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X2288 VSS row_n[14] a_14314_16226# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X2289 a_11302_13214# col_n[8] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2290 a_10394_3496# col_n[7] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X2291 vcm a_2275_17214# a_28066_17190# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2292 VSS row_n[14] a_4274_16226# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X2293 a_32082_15182# a_2475_15206# a_31990_15182# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X2294 VSS row_n[7] a_21342_9198# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X2295 a_19942_16186# row_n[14] a_20434_16548# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2296 a_19030_10162# a_2475_10186# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2297 VSS row_n[1] a_15318_3174# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X2298 a_32994_15182# row_n[13] a_33486_15544# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2299 a_14010_14178# a_2475_14202# a_13918_14178# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X2300 vcm a_2275_11190# a_33086_11166# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2301 a_24962_9158# a_2275_9182# a_25054_9158# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2302 a_35094_9158# a_2475_9182# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2303 VSS row_n[5] a_14314_7190# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X2304 vcm a_2275_7174# a_32082_7150# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2305 VDD VDD a_12914_18194# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2306 a_10394_15544# col_n[7] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X2307 a_3970_14178# a_2475_14202# a_3878_14178# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X2308 a_4370_7512# col_n[1] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X2309 VDD rowon_n[4] a_18938_6146# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2310 a_30986_6146# row_n[4] a_31478_6508# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2311 VDD VDD a_2874_18194# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2312 vcm a_2275_12194# a_8990_12170# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2313 vcm a_2275_12194# a_19030_12170# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2314 a_4974_7150# a_2475_7174# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2315 a_17422_6508# col_n[14] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X2316 a_12002_1126# a_2475_1150# a_11910_1126# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X2317 a_5978_3134# a_2475_3158# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2318 a_10906_11166# row_n[9] a_11398_11528# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2319 VDD a_2161_8178# a_2275_8178# VDD sky130_fd_pr__pfet_01v8 ad=0.249 pd=1.62 as=0.342 ps=2.97 w=1.2 l=0.15
X2320 a_18026_6146# a_2475_6170# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2321 a_23958_2130# a_2275_2154# a_24050_2130# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2322 ctop sw analog_in VSS sky130_fd_pr__nfet_01v8 ad=0.275 pd=2.19 as=0.275 ps=2.19 w=1.9 l=0.22
X2323 a_23046_12170# a_2475_12194# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2324 a_21438_9520# col_n[18] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X2325 a_13918_8154# a_2275_8178# a_14010_8154# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2326 a_15414_1488# col_n[12] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X2327 VSS row_n[0] a_7286_2170# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X2328 a_33390_5182# col_n[30] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2329 a_1957_3158# VDD sample VSS sky130_fd_pr__nfet_01v8 ad=0.171 pd=1.77 as=0.171 ps=1.77 w=0.6 l=0.15
X2330 a_32386_17230# rowon_n[15] a_31990_17190# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X2331 a_35002_8154# row_n[6] a_35494_8516# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2332 a_9390_5504# col_n[6] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X2333 a_21342_1166# VSS a_20946_1126# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X2334 a_9994_5142# a_2475_5166# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2335 a_29374_15222# col_n[26] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2336 VSS row_n[12] a_20338_14218# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X2337 VSS row_n[11] a_33390_13214# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X2338 a_20946_17190# a_2275_17214# a_21038_17190# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2339 a_5886_7150# a_2275_7174# a_5978_7150# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2340 vcm a_2275_1150# a_13006_1126# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2341 a_32994_3134# row_n[1] a_33486_3496# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2342 a_6890_3134# a_2275_3158# a_6982_3134# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2343 a_10298_13214# rowon_n[11] a_9902_13174# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X2344 a_26458_7512# col_n[23] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X2345 a_18938_6146# a_2275_6170# a_19030_6146# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2346 a_24962_16186# a_2275_16210# a_25054_16186# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2347 a_8990_18194# a_2475_18218# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2348 a_28466_17552# col_n[25] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X2349 VDD rowon_n[13] a_31990_15182# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2350 a_28066_13174# a_2475_13198# a_27974_13174# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X2351 a_10998_8154# a_2475_8178# a_10906_8154# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X2352 a_20034_6146# a_2475_6170# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2353 a_11910_12170# a_2275_12194# a_12002_12170# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2354 a_28978_13174# row_n[11] a_29470_13536# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2355 a_33486_11528# col_n[30] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X2356 VDD rowon_n[9] a_9902_11166# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2357 VDD rowon_n[5] a_10906_7150# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2358 a_3270_6186# rowon_n[4] a_2874_6146# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X2359 a_31382_18234# col_n[28] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2360 vcm a_2275_9182# a_23046_9158# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2361 a_19030_3134# a_2475_3158# a_18938_3134# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X2362 a_33086_9158# a_2475_9182# a_32994_9158# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X2363 vcm a_2275_18218# a_26058_18194# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2364 a_30074_16186# a_2475_16210# a_29982_16186# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X2365 a_20338_8194# rowon_n[6] a_19942_8154# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X2366 a_2966_7150# a_2475_7174# a_2874_7150# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X2367 a_24050_8154# a_2475_8178# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2368 a_16018_6146# a_2475_6170# a_15926_6146# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X2369 vcm a_2275_2154# a_22042_2130# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2370 a_14314_2170# rowon_n[0] a_13918_2130# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X2371 a_25054_4138# a_2475_4162# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2372 a_19942_5142# row_n[3] a_20434_5504# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2373 a_30986_16186# row_n[14] a_31478_16548# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2374 a_30474_5504# col_n[27] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X2375 vcm a_2275_8178# a_12002_8154# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2376 a_16930_17190# row_n[15] a_17422_17552# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2377 vcm a_2275_13198# a_17022_13174# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2378 VDD rowon_n[3] a_15926_5142# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2379 a_8290_4178# rowon_n[2] a_7894_4138# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X2380 a_6890_17190# row_n[15] a_7382_17552# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2381 vcm a_2275_13198# a_6982_13174# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2382 a_21038_13174# a_2475_13198# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2383 a_2475_9182# a_1957_9182# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.342 pd=2.97 as=0.249 ps=1.62 w=1.2 l=0.15
X2384 a_25358_6186# rowon_n[4] a_24962_6146# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X2385 a_7986_5142# a_2475_5166# a_7894_5142# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X2386 VSS a_2161_14202# a_2275_14202# VSS sky130_fd_pr__nfet_01v8 ad=0.124 pd=1.01 as=0.171 ps=1.77 w=0.6 l=0.15
X2387 a_13310_6186# col_n[10] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2388 a_29070_6146# a_2475_6170# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2389 a_31382_12210# rowon_n[10] a_30986_12170# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X2390 vcm a_2275_7174# a_3970_7150# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2391 a_34490_7512# col_n[31] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X2392 a_2874_6146# row_n[4] a_3366_6508# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2393 a_28370_10202# col_n[25] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2394 vcm a_2275_6170# a_17022_6146# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2395 VDD rowon_n[2] a_7894_4138# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2396 a_30378_18234# VDD a_29982_18194# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X2397 a_19942_12170# a_2275_12194# a_20034_12170# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2398 a_32482_2492# col_n[29] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X2399 a_31990_5142# a_2275_5166# a_32082_5142# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2400 a_27366_16226# col_n[24] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2401 VSS row_n[12] a_31382_14218# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X2402 a_18938_10162# a_2275_10186# a_19030_10162# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2403 a_31990_17190# a_2275_17214# a_32082_17190# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2404 a_27462_12532# col_n[24] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X2405 a_8898_10162# a_2275_10186# a_8990_10162# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2406 VDD rowon_n[8] a_30986_10162# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2407 VSS row_n[6] a_19334_8194# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X2408 a_6282_1166# col_n[3] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2409 a_29374_8194# rowon_n[6] a_28978_8154# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X2410 a_5278_5182# col_n[2] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2411 a_26058_14178# a_2475_14202# a_25966_14178# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X2412 a_18330_4178# col_n[15] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2413 a_26458_18556# col_n[23] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X2414 VDD rowon_n[14] a_29982_16186# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2415 vcm a_2275_5166# a_8990_5142# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2416 a_30378_13214# col_n[27] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2417 a_22346_7190# col_n[19] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2418 VDD a_2161_15206# a_2275_15206# VDD sky130_fd_pr__pfet_01v8 ad=0.249 pd=1.62 as=0.342 ps=2.97 w=1.2 l=0.15
X2419 vcm a_2275_2154# a_30074_2130# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2420 VSS row_n[15] a_9294_17230# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X2421 a_24050_17190# a_2475_17214# a_23958_17190# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X2422 a_22042_8154# a_2475_8178# a_21950_8154# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X2423 a_4882_3134# row_n[1] a_5374_3496# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2424 a_23046_4138# a_2475_4162# a_22954_4138# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X2425 vcm a_2275_13198# a_25054_13174# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2426 a_24962_17190# row_n[15] a_25454_17552# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2427 a_17934_4138# row_n[2] a_18426_4500# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2428 a_8990_15182# a_2475_15206# a_8898_15182# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X2429 a_29982_11166# row_n[9] a_30474_11528# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2430 a_9390_15544# col_n[6] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X2431 a_5886_12170# row_n[10] a_6378_12532# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2432 a_15926_12170# row_n[10] a_16418_12532# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2433 a_28066_11166# a_2475_11190# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2434 a_27366_10202# rowon_n[8] a_26970_10162# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X2435 a_10394_6508# col_n[7] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X2436 a_10998_6146# a_2475_6170# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2437 a_33390_6186# rowon_n[4] a_32994_6146# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X2438 a_27366_5182# col_n[24] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2439 a_19030_13174# a_2475_13198# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2440 a_27062_6146# a_2475_6170# a_26970_6146# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X2441 a_28978_8154# row_n[6] a_29470_8516# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2442 a_19030_1126# a_2475_1150# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2443 vcm a_2275_17214# a_13006_17190# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2444 VSS row_n[3] a_12306_5182# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X2445 VSS VDD a_13310_1166# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X2446 vcm a_2275_17214# a_2966_17190# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2447 a_26970_3134# row_n[1] a_27462_3496# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2448 a_28370_18234# VDD a_27974_18194# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X2449 VSS row_n[13] a_25358_15222# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X2450 a_22346_12210# col_n[19] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2451 a_2966_5142# a_2475_5166# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2452 a_14410_8516# col_n[11] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X2453 a_16018_4138# a_2475_4162# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2454 VSS row_n[12] a_29374_14218# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X2455 a_26362_11206# col_n[23] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2456 a_15014_8154# a_2475_8178# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2457 VSS a_2161_2154# a_2275_2154# VSS sky130_fd_pr__nfet_01v8 ad=0.124 pd=1.01 as=0.171 ps=1.77 w=0.6 l=0.15
X2458 VDD rowon_n[15] a_23958_17190# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2459 a_12002_15182# a_2475_15206# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2460 a_34090_15182# a_2475_15206# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2461 a_21438_14540# col_n[18] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X2462 a_30986_12170# a_2275_12194# a_31078_12170# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2463 VSS row_n[8] a_16322_10202# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X2464 a_21038_10162# a_2475_10186# a_20946_10162# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X2465 a_18330_7190# rowon_n[5] a_17934_7150# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X2466 a_11910_6146# a_2275_6170# a_12002_6146# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2467 a_31382_3174# col_n[28] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2468 a_19334_3174# rowon_n[1] a_18938_3134# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X2469 a_12402_3496# col_n[9] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X2470 a_9294_13214# rowon_n[11] a_8898_13174# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X2471 a_6890_11166# a_2275_11190# a_6982_11166# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2472 a_16930_11166# a_2275_11190# a_17022_11166# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2473 VSS row_n[8] a_6282_10202# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X2474 VSS row_n[7] a_23350_9198# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X2475 a_30378_7190# col_n[27] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2476 VDD rowon_n[14] a_27974_16186# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2477 a_25454_13536# col_n[22] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X2478 a_21950_10162# row_n[8] a_22442_10524# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2479 VSS row_n[1] a_17326_3174# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X2480 vcm a_2275_7174# a_34090_7150# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2481 a_32994_6146# row_n[4] a_33486_6508# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2482 VDD rowon_n[10] a_14922_12170# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2483 a_14010_1126# a_2475_1150# a_13918_1126# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X2484 a_7986_3134# a_2475_3158# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2485 VDD rowon_n[10] a_4882_12170# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2486 a_6982_7150# a_2475_7174# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2487 a_25966_2130# a_2275_2154# a_26058_2130# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2488 VDD rowon_n[9] a_8898_11166# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2489 VDD en_bit_n[2] a_18938_1126# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2490 a_30986_1126# VDD a_31478_1488# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2491 VSS VDD a_17326_18234# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X2492 a_22042_18194# a_2475_18218# a_21950_18194# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X2493 a_14314_15222# col_n[11] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2494 a_3878_5142# a_2275_5166# a_3970_5142# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2495 a_4370_2492# col_n[1] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X2496 vcm a_2275_3158# a_9994_3134# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2497 VSS VDD a_7286_18234# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X2498 a_13006_17190# a_2475_17214# a_12914_17190# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X2499 a_35094_17190# a_2475_17214# a_35002_17190# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X2500 a_4274_15222# col_n[1] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2501 a_23446_9520# col_n[20] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X2502 a_15926_8154# a_2275_8178# a_16018_8154# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2503 a_17422_1488# col_n[14] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X2504 a_16930_4138# a_2275_4162# a_17022_4138# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2505 a_22954_18194# VDD a_23446_18556# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2506 a_2966_17190# a_2475_17214# a_2874_17190# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X2507 a_18330_14218# col_n[15] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2508 vcm a_2275_14202# a_23046_14178# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2509 VSS row_n[0] a_9294_2170# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X2510 a_35398_5182# VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2511 a_9902_16186# a_2275_16210# a_9994_16186# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2512 a_17022_16186# a_2475_16210# a_16930_16186# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X2513 a_8290_14218# col_n[5] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2514 a_13406_17552# col_n[10] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X2515 a_6982_16186# a_2475_16210# a_6890_16186# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X2516 a_23350_1166# VSS a_22954_1126# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X2517 a_3366_17552# col_n[0] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X2518 a_17422_16548# col_n[14] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X2519 a_13918_13174# row_n[11] a_14410_13536# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2520 a_25358_11206# rowon_n[9] a_24962_11166# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X2521 a_1957_10186# VSS sample VDD sky130_fd_pr__pfet_01v8 ad=0.342 pd=2.97 as=0.342 ps=2.97 w=1.2 l=0.15
X2522 a_2161_5166# sample VSS VSS sky130_fd_pr__nfet_01v8 ad=0.171 pd=1.77 as=0.171 ps=1.77 w=0.6 l=0.15
X2523 a_7382_16548# col_n[4] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X2524 a_3878_13174# row_n[11] a_4370_13536# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2525 a_35002_3134# row_n[1] a_35494_3496# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2526 a_7894_7150# a_2275_7174# a_7986_7150# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2527 vcm a_2275_1150# a_15014_1126# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2528 a_8898_3134# a_2275_3158# a_8990_3134# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2529 a_28466_7512# col_n[25] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X2530 a_13006_8154# a_2475_8178# a_12914_8154# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X2531 a_22042_6146# a_2475_6170# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2532 ctop sw_n analog_in VDD sky130_fd_pr__pfet_01v8 ad=0.551 pd=4.38 as=0.275 ps=2.19 w=1.9 l=0.22
X2533 VSS row_n[8] a_24354_10202# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X2534 a_26458_2492# col_n[23] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X2535 vcm a_2275_18218# a_10998_18194# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2536 a_24962_11166# a_2275_11190# a_25054_11166# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2537 VDD rowon_n[5] a_12914_7150# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2538 VSS row_n[14] a_23350_16226# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X2539 a_19430_14540# col_n[16] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X2540 VDD rowon_n[10] a_22954_12170# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2541 a_19030_10162# a_2475_10186# a_18938_10162# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X2542 vcm a_2275_9182# a_25054_9158# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2543 a_35094_9158# a_2475_9182# a_35002_9158# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X2544 a_20338_2170# col_n[17] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2545 VDD rowon_n[0] a_10906_2130# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2546 a_27974_18194# a_2275_18218# a_28066_18194# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2547 a_32082_16186# a_2475_16210# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2548 a_22346_8194# rowon_n[6] a_21950_8154# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X2549 a_4974_7150# a_2475_7174# a_4882_7150# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X2550 VSS row_n[0] a_30378_2170# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X2551 a_5978_3134# a_2475_3158# a_5886_3134# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X2552 a_2475_3158# a_1957_3158# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.171 pd=1.77 as=0.124 ps=1.01 w=0.6 l=0.15
X2553 VDD VDD a_21950_18194# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2554 VDD rowon_n[15] a_35002_17190# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2555 a_7286_14218# rowon_n[12] a_6890_14178# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X2556 a_17326_14218# rowon_n[12] a_16930_14178# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X2557 a_10298_8194# col_n[7] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2558 a_18026_6146# a_2475_6170# a_17934_6146# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X2559 vcm a_2275_2154# a_24050_2130# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2560 a_16322_2170# rowon_n[0] a_15926_2130# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X2561 a_27062_4138# a_2475_4162# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2562 a_11302_4178# col_n[8] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2563 analog_in sw_n ctop VDD sky130_fd_pr__pfet_01v8 ad=0.275 pd=2.19 as=0.275 ps=2.19 w=1.9 l=0.22
X2564 a_32482_5504# col_n[29] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X2565 a_8898_13174# a_2275_13198# a_8990_13174# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2566 a_18938_13174# a_2275_13198# a_19030_13174# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2567 vcm a_2275_8178# a_14010_8154# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2568 a_34090_12170# a_2475_12194# a_33998_12170# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X2569 a_3270_10202# col_n[0] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2570 a_13310_10202# col_n[10] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2571 a_12002_12170# a_2475_12194# a_11910_12170# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X2572 a_12306_16226# col_n[9] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2573 a_35002_12170# row_n[10] a_35494_12532# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2574 a_27366_6186# rowon_n[4] a_26970_6146# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X2575 a_9994_5142# a_2475_5166# a_9902_5142# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X2576 a_3270_3174# col_n[0] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2577 a_10906_4138# row_n[2] a_11398_4500# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2578 a_10998_18194# a_2475_18218# a_10906_18194# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X2579 a_33086_18194# a_2475_18218# a_32994_18194# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X2580 a_5278_9198# rowon_n[7] a_4882_9158# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X2581 a_15318_6186# col_n[12] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2582 a_33998_18194# VDD a_34490_18556# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2583 vcm a_2275_14202# a_34090_14178# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2584 a_12402_12532# col_n[9] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X2585 a_19334_12210# rowon_n[10] a_18938_12170# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X2586 vcm a_2275_3158# a_6982_3134# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2587 vcm a_2275_7174# a_5978_7150# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2588 a_4882_6146# row_n[4] a_5374_6508# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2589 a_11398_18556# col_n[8] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X2590 vcm a_2275_6170# a_19030_6146# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2591 a_20034_6146# a_2475_6170# a_19942_6146# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X2592 a_34490_2492# col_n[31] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X2593 a_2874_1126# VDD a_3366_1488# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2594 a_33998_5142# a_2275_5166# a_34090_5142# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2595 VDD rowon_n[8] a_18938_10162# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2596 a_21950_8154# row_n[6] a_22442_8516# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2597 a_2475_17214# a_1957_17214# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.171 pd=1.77 as=0.124 ps=1.01 w=0.6 l=0.15
X2598 VDD rowon_n[7] a_4882_9158# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2599 a_8290_1166# col_n[5] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2600 a_9902_17190# row_n[15] a_10394_17552# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2601 a_21342_15222# rowon_n[13] a_20946_15182# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X2602 a_28066_14178# a_2475_14202# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2603 vcm a_2275_13198# a_9994_13174# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2604 a_9902_1126# a_2275_1150# a_9994_1126# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2605 VSS row_n[9] a_22346_11206# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X2606 a_31382_4178# rowon_n[2] a_30986_4138# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X2607 VSS row_n[8] a_35398_10202# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X2608 a_24354_7190# col_n[21] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2609 a_12306_10202# rowon_n[8] a_11910_10162# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X2610 a_24050_8154# a_2475_8178# a_23958_8154# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X2611 a_25054_4138# a_2475_4162# a_24962_4138# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X2612 VDD rowon_n[11] a_20946_13174# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2613 a_26970_6146# row_n[4] a_27462_6508# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2614 VDD rowon_n[10] a_33998_12170# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2615 VSS row_n[1] a_10298_3174# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X2616 a_19942_9158# a_2275_9182# a_20034_9158# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2617 a_30074_9158# a_2475_9182# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2618 a_20338_16226# col_n[17] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2619 VDD rowon_n[2] a_30986_4138# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2620 a_2475_18218# a_1957_18218# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.342 pd=2.97 as=0.249 ps=1.62 w=1.2 l=0.15
X2621 a_33390_15222# col_n[30] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2622 a_12402_6508# col_n[9] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X2623 a_16930_14178# a_2275_14202# a_17022_14178# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2624 a_13006_6146# a_2475_6170# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2625 a_29374_5182# col_n[26] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2626 a_3270_18234# VDD a_2874_18194# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X2627 a_13310_18234# VDD a_12914_18194# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X2628 VSS row_n[13] a_10298_15222# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X2629 a_6890_14178# a_2275_14202# a_6982_14178# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2630 a_7286_8194# col_n[4] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2631 a_29070_6146# a_2475_6170# a_28978_6146# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X2632 VSS row_n[12] a_14314_14218# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X2633 a_11302_11206# col_n[8] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2634 a_10394_1488# col_n[7] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X2635 a_32482_17552# col_n[29] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X2636 vcm a_2275_15206# a_28066_15182# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2637 VSS row_n[12] a_4274_14218# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X2638 a_32082_13174# a_2475_13198# a_31990_13174# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X2639 a_4882_17190# a_2275_17214# a_4974_17190# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2640 a_14922_17190# a_2275_17214# a_15014_17190# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2641 VSS row_n[3] a_14314_5182# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X2642 VSS VDD a_15318_1166# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X2643 a_32994_13174# row_n[11] a_33486_13536# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2644 a_28978_3134# row_n[1] a_29470_3496# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2645 vcm a_2275_5166# a_32082_5142# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2646 VDD rowon_n[14] a_12914_16186# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2647 a_10394_13536# col_n[7] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X2648 vcm a_2275_10186# a_19030_10162# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2649 VDD rowon_n[6] a_17934_8154# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2650 a_29982_8154# row_n[6] a_30474_8516# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2651 a_4370_5504# col_n[1] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X2652 VDD rowon_n[14] a_2874_16186# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2653 a_8898_14178# row_n[12] a_9390_14540# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2654 a_18938_14178# row_n[12] a_19430_14540# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2655 vcm a_2275_10186# a_8990_10162# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2656 a_4974_5142# a_2475_5166# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2657 a_5978_1126# a_2475_1150# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2658 a_17022_8154# a_2475_8178# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2659 VDD a_2161_6170# a_2275_6170# VDD sky130_fd_pr__pfet_01v8 ad=0.249 pd=1.62 as=0.342 ps=2.97 w=1.2 l=0.15
X2660 a_18026_4138# a_2475_4162# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2661 vcm a_2275_18218# a_30074_18194# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2662 a_21438_7512# col_n[18] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X2663 a_13918_6146# a_2275_6170# a_14010_6146# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2664 analog_in sw ctop VSS sky130_fd_pr__nfet_01v8 ad=0.275 pd=2.19 as=0.275 ps=2.19 w=1.9 l=0.22
X2665 a_14410_3496# col_n[11] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X2666 a_33390_3174# col_n[30] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2667 VSS row_n[7] a_25358_9198# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X2668 a_35398_9198# rowon_n[7] a_35002_9158# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X2669 a_12002_10162# a_2475_10186# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2670 a_34090_10162# a_2475_10186# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2671 VSS row_n[15] a_28370_17230# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X2672 a_32386_15222# rowon_n[13] a_31990_15182# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X2673 a_35002_6146# row_n[4] a_35494_6508# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2674 a_8990_7150# a_2475_7174# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2675 a_9994_3134# a_2475_3158# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2676 a_29374_13214# col_n[26] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2677 VSS row_n[9] a_33390_11206# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X2678 a_27974_2130# a_2275_2154# a_28066_2130# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2679 a_24050_18194# a_2475_18218# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2680 a_20946_15182# a_2275_15206# a_21038_15182# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2681 a_5886_5142# a_2275_5166# a_5978_5142# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2682 a_6890_1126# a_2275_1150# a_6982_1126# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2683 a_32994_1126# VDD a_33486_1488# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2684 a_15014_17190# a_2475_17214# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2685 a_10298_11206# rowon_n[9] a_9902_11166# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X2686 a_25454_9520# col_n[22] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X2687 a_17934_8154# a_2275_8178# a_18026_8154# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2688 a_18938_4138# a_2275_4162# a_19030_4138# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2689 a_26458_5504# col_n[23] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X2690 a_4974_17190# a_2475_17214# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2691 a_24962_14178# a_2275_14202# a_25054_14178# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2692 VDD rowon_n[7] a_35002_9158# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2693 a_8990_16186# a_2475_16210# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2694 a_28466_15544# col_n[25] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X2695 VDD rowon_n[11] a_31990_13174# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2696 a_28066_11166# a_2475_11190# a_27974_11166# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X2697 a_10998_6146# a_2475_6170# a_10906_6146# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X2698 a_20034_4138# a_2475_4162# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2699 a_28978_11166# row_n[9] a_29470_11528# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2700 a_9902_11166# a_2275_11190# a_9994_11166# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2701 a_2161_9182# sample VDD VDD sky130_fd_pr__pfet_01v8 ad=0.342 pd=2.97 as=0.342 ps=2.97 w=1.2 l=0.15
X2702 VDD rowon_n[3] a_10906_5142# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2703 a_3270_4178# rowon_n[2] a_2874_4138# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X2704 a_31382_16226# col_n[28] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2705 VSS row_n[5] a_6282_7190# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X2706 a_19030_1126# a_2475_1150# a_18938_1126# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X2707 vcm a_2275_17214# a_22042_17190# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2708 a_7286_17230# col_n[4] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2709 a_17326_17230# col_n[14] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2710 vcm a_2275_16210# a_26058_16186# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2711 a_30074_14178# a_2475_14202# a_29982_14178# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X2712 a_20338_6186# rowon_n[4] a_19942_6146# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X2713 a_2966_5142# a_2475_5166# a_2874_5142# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X2714 a_12914_18194# a_2275_18218# a_13006_18194# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2715 a_30474_18556# col_n[27] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X2716 a_15014_8154# a_2475_8178# a_14922_8154# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X2717 a_24050_6146# a_2475_6170# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2718 a_16018_4138# a_2475_4162# a_15926_4138# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X2719 a_2874_18194# a_2275_18218# a_2966_18194# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2720 a_9994_18194# a_2475_18218# a_9902_18194# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X2721 a_28466_2492# col_n[25] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X2722 vcm a_2275_6170# a_12002_6146# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2723 VDD rowon_n[2] a_2874_4138# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2724 a_16930_15182# row_n[13] a_17422_15544# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2725 vcm a_2275_11190# a_17022_11166# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2726 a_6890_15182# row_n[13] a_7382_15544# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2727 vcm a_2275_11190# a_6982_11166# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2728 VDD rowon_n[0] a_12914_2130# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2729 VSS row_n[0] a_32386_2170# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X2730 a_24354_8194# rowon_n[6] a_23958_8154# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X2731 a_6982_7150# a_2475_7174# a_6890_7150# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X2732 a_7986_3134# a_2475_3158# a_7894_3134# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X2733 a_25358_4178# rowon_n[2] a_24962_4138# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X2734 VSS row_n[10] a_27366_12210# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X2735 vcm a_2275_2154# a_26058_2130# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2736 a_29070_4138# a_2475_4162# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2737 a_13310_4178# col_n[10] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2738 a_32082_11166# a_2475_11190# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2739 a_31382_10202# rowon_n[8] a_30986_10162# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X2740 vcm a_2275_5166# a_3970_5142# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2741 a_34490_5504# col_n[31] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X2742 vcm a_2275_8178# a_16018_8154# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2743 vcm a_2275_4162# a_17022_4138# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2744 VSS VDD a_26362_18234# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X2745 a_30378_16226# rowon_n[14] a_29982_16186# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X2746 VDD rowon_n[12] a_25966_14178# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2747 a_14010_12170# a_2475_12194# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2748 a_30986_7150# a_2275_7174# a_31078_7150# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2749 a_31990_3134# a_2275_3158# a_32082_3134# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2750 a_27366_14218# col_n[24] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2751 a_3970_12170# a_2475_12194# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2752 VDD rowon_n[2] a_24962_4138# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2753 a_35094_18194# a_2475_18218# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2754 a_31990_15182# a_2275_15206# a_32082_15182# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2755 a_27462_10524# col_n[24] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X2756 VSS row_n[4] a_19334_6186# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X2757 a_12914_4138# row_n[2] a_13406_4500# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2758 a_2966_18194# a_2475_18218# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2759 a_13006_18194# a_2475_18218# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2760 a_29374_6186# rowon_n[4] a_28978_6146# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X2761 a_5278_3174# col_n[2] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2762 a_25358_17230# col_n[22] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2763 a_26458_16548# col_n[23] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X2764 a_7286_9198# rowon_n[7] a_6890_9158# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X2765 vcm a_2275_7174# a_7986_7150# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2766 vcm a_2275_3158# a_8990_3134# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2767 a_30378_11206# col_n[27] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2768 ctop sw analog_in VSS sky130_fd_pr__nfet_01v8 ad=0.275 pd=2.19 as=0.275 ps=2.19 w=1.9 l=0.22
X2769 a_22346_5182# col_n[19] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2770 VDD a_2161_13198# a_2275_13198# VDD sky130_fd_pr__pfet_01v8 ad=0.249 pd=1.62 as=0.342 ps=2.97 w=1.2 l=0.15
X2771 VSS row_n[13] a_9294_15222# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X2772 a_24050_15182# a_2475_15206# a_23958_15182# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X2773 a_6282_12210# col_n[3] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2774 a_16322_12210# col_n[13] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2775 vcm a_2275_12194# a_21038_12170# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2776 a_22042_6146# a_2475_6170# a_21950_6146# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X2777 a_4882_1126# VDD a_5374_1488# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2778 vcm a_2275_11190# a_25054_11166# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2779 a_23958_8154# row_n[6] a_24450_8516# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2780 a_24962_15182# row_n[13] a_25454_15544# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2781 a_8990_13174# a_2475_13198# a_8898_13174# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X2782 VDD rowon_n[7] a_6890_9158# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2783 VDD rowon_n[15] a_7894_17190# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2784 a_5374_14540# col_n[2] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X2785 a_15414_14540# col_n[12] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X2786 a_21950_3134# row_n[1] a_22442_3496# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2787 a_9390_13536# col_n[6] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X2788 a_2475_12194# a_1957_12194# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.171 pd=1.77 as=0.124 ps=1.01 w=0.6 l=0.15
X2789 a_5886_10162# row_n[8] a_6378_10524# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2790 a_15926_10162# row_n[8] a_16418_10524# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2791 a_26362_7190# col_n[23] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2792 a_27366_3174# col_n[24] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2793 a_33390_4178# rowon_n[2] a_32994_4138# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X2794 a_10998_4138# a_2475_4162# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2795 a_17326_9198# col_n[14] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2796 a_27062_4138# a_2475_4162# a_26970_4138# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X2797 a_28978_6146# row_n[4] a_29470_6508# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2798 a_24354_17230# rowon_n[15] a_23958_17190# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X2799 vcm a_2275_15206# a_13006_15182# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2800 VDD VSS VSS sky130_fd_pr__cap_var_lvt w=16.4 l=16
X2801 VSS row_n[1] a_12306_3174# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X2802 vcm a_2275_15206# a_2966_15182# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2803 a_32082_9158# a_2475_9182# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2804 a_26970_1126# VDD a_27462_1488# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2805 a_2161_18218# sample VSS VSS sky130_fd_pr__nfet_01v8 ad=0.171 pd=1.77 as=0.171 ps=1.77 w=0.6 l=0.15
X2806 a_28370_16226# rowon_n[14] a_27974_16186# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X2807 VSS row_n[11] a_25358_13214# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X2808 a_22346_10202# col_n[19] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2809 a_2966_3134# a_2475_3158# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2810 VDD rowon_n[2] a_32994_4138# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2811 a_14410_6508# col_n[11] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X2812 a_20946_2130# a_2275_2154# a_21038_2130# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2813 a_15318_12210# rowon_n[10] a_14922_12170# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X2814 a_16930_9158# row_n[7] a_17422_9520# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2815 a_9294_8194# col_n[6] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2816 a_15014_6146# a_2475_6170# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2817 a_31078_2130# a_2475_2154# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2818 a_5278_12210# rowon_n[10] a_4882_12170# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X2819 VDD rowon_n[13] a_23958_15182# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2820 a_12002_13174# a_2475_13198# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2821 a_34090_13174# a_2475_13198# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2822 a_21438_12532# col_n[18] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X2823 a_10906_8154# a_2275_8178# a_10998_8154# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2824 a_18330_5182# rowon_n[3] a_17934_5142# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X2825 a_12402_1488# col_n[9] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X2826 a_19334_1166# en_bit_n[2] a_18938_1126# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X2827 a_31382_1166# col_n[28] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2828 a_11910_4138# a_2275_4162# a_12002_4138# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2829 a_9294_11206# rowon_n[9] a_8898_11166# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X2830 VSS row_n[0] a_4274_2170# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X2831 a_30378_5182# col_n[27] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2832 a_25454_11528# col_n[22] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X2833 VSS VDD a_17326_1166# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X2834 a_23350_18234# col_n[20] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2835 vcm a_2275_5166# a_34090_5142# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2836 VDD rowon_n[8] a_14922_10162# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2837 a_7986_1126# a_2475_1150# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2838 VDD rowon_n[8] a_4882_10162# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2839 a_6982_5142# a_2475_5166# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2840 VSS row_n[15] a_3270_17230# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X2841 VSS row_n[15] a_13310_17230# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X2842 a_29982_3134# row_n[1] a_30474_3496# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2843 VDD rowon_n[1] a_17934_3134# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2844 VSS row_n[14] a_17326_16226# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X2845 a_22042_16186# a_2475_16210# a_21950_16186# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X2846 a_14314_13214# col_n[11] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2847 a_2874_7150# a_2275_7174# a_2966_7150# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2848 vcm a_2275_1150# a_9994_1126# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2849 a_3878_3134# a_2275_3158# a_3970_3134# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2850 VSS row_n[14] a_7286_16226# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X2851 a_13006_15182# a_2475_15206# a_12914_15182# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X2852 a_35094_15182# a_2475_15206# a_35002_15182# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X2853 a_4274_13214# col_n[1] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2854 vcm a_2275_12194# a_32082_12170# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2855 a_23446_7512# col_n[20] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X2856 a_15926_6146# a_2275_6170# a_16018_6146# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2857 a_22954_16186# row_n[14] a_23446_16548# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2858 a_2966_15182# a_2475_15206# a_2874_15182# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X2859 VSS row_n[7] a_27366_9198# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X2860 a_35398_3174# VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2861 a_9902_14178# a_2275_14202# a_9994_14178# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2862 a_17022_14178# a_2475_14202# a_16930_14178# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X2863 a_21438_2492# col_n[18] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X2864 VDD VDD a_15926_18194# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2865 a_13406_15544# col_n[10] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X2866 a_6982_14178# a_2475_14202# a_6890_14178# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X2867 VDD VDD a_5886_18194# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2868 a_3366_15544# col_n[0] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X2869 VSS row_n[0] a_26362_2170# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X2870 a_2161_3158# sample VSS VSS sky130_fd_pr__nfet_01v8 ad=0.171 pd=1.77 as=0.171 ps=1.77 w=0.6 l=0.15
X2871 a_13918_11166# row_n[9] a_14410_11528# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2872 a_3878_11166# row_n[9] a_4370_11528# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2873 vcm a_2275_9182# a_20034_9158# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2874 a_35002_1126# VDD a_35494_1488# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2875 a_26058_12170# a_2475_12194# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2876 a_30074_9158# a_2475_9182# a_29982_9158# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X2877 VSS row_n[6] a_16322_8194# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X2878 a_7894_5142# a_2275_5166# a_7986_5142# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2879 a_8898_1126# a_2275_1150# a_8990_1126# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2880 a_27462_9520# col_n[24] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X2881 a_28466_5504# col_n[25] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X2882 a_23350_12210# rowon_n[10] a_22954_12170# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X2883 a_20946_10162# a_2275_10186# a_21038_10162# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2884 a_6378_8516# col_n[3] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X2885 a_13006_6146# a_2475_6170# a_12914_6146# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X2886 a_11302_2170# rowon_n[0] a_10906_2130# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X2887 a_22042_4138# a_2475_4162# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2888 a_22346_18234# VDD a_21950_18194# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X2889 vcm a_2275_16210# a_10998_16186# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2890 a_35398_17230# rowon_n[15] a_35002_17190# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X2891 VDD rowon_n[3] a_12914_5142# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2892 VSS row_n[12] a_23350_14218# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X2893 a_8990_11166# a_2475_11190# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2894 a_23958_17190# a_2275_17214# a_24050_17190# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2895 a_19430_12532# col_n[16] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X2896 VDD rowon_n[8] a_22954_10162# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2897 VSS row_n[5] a_8290_7190# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X2898 a_27974_16186# a_2275_16210# a_28066_16186# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2899 a_32082_14178# a_2475_14202# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2900 a_22346_6186# rowon_n[4] a_21950_6146# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X2901 a_4974_5142# a_2475_5166# a_4882_5142# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X2902 a_5978_1126# a_2475_1150# a_5886_1126# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X2903 VDD rowon_n[14] a_21950_16186# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2904 VDD rowon_n[13] a_35002_15182# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2905 a_10298_6186# col_n[7] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2906 a_18026_4138# a_2475_4162# a_17934_4138# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X2907 a_35398_12210# VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2908 a_17022_8154# a_2475_8178# a_16930_8154# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X2909 VSS row_n[10] a_12306_12210# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X2910 vcm a_2275_6170# a_14010_6146# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2911 a_34394_18234# col_n[31] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2912 VSS VDD a_11302_18234# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X2913 a_34490_14540# col_n[31] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X2914 a_34090_10162# a_2475_10186# a_33998_10162# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X2915 a_12002_10162# a_2475_10186# a_11910_10162# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X2916 vcm a_2275_18218# a_29070_18194# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2917 VDD rowon_n[12] a_10906_14178# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2918 a_12306_14218# col_n[9] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2919 a_35002_10162# row_n[8] a_35494_10524# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2920 VSS row_n[0] a_34394_2170# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X2921 a_3270_1166# col_n[0] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2922 a_9994_3134# a_2475_3158# a_9902_3134# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X2923 a_27366_4178# rowon_n[2] a_26970_4138# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X2924 a_10998_16186# a_2475_16210# a_10906_16186# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X2925 a_33086_16186# a_2475_16210# a_32994_16186# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X2926 a_19334_10202# rowon_n[8] a_18938_10162# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X2927 a_26362_8194# rowon_n[6] a_25966_8154# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X2928 a_8990_7150# a_2475_7174# a_8898_7150# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X2929 vcm a_2275_2154# a_28066_2130# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2930 a_15318_4178# col_n[12] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2931 a_33998_16186# row_n[14] a_34490_16548# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2932 a_12402_10524# col_n[9] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X2933 vcm a_2275_1150# a_6982_1126# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2934 VDD VSS sky130_fd_pr__cap_mim_m3_1 l=17.2 w=17.2
X2935 a_10298_17230# col_n[7] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2936 vcm a_2275_5166# a_5978_5142# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2937 a_11398_16548# col_n[8] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X2938 vcm a_2275_8178# a_18026_8154# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2939 vcm a_2275_4162# a_19030_4138# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2940 a_20034_4138# a_2475_4162# a_19942_4138# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X2941 a_26058_9158# a_2475_9182# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2942 a_15318_7190# rowon_n[5] a_14922_7150# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X2943 a_32994_7150# a_2275_7174# a_33086_7150# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2944 a_33998_3134# a_2275_3158# a_34090_3134# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2945 a_21950_6146# row_n[4] a_22442_6508# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2946 VDD rowon_n[2] a_26970_4138# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2947 a_2475_15206# a_1957_15206# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.171 pd=1.77 as=0.124 ps=1.01 w=0.6 l=0.15
X2948 VDD rowon_n[5] a_4882_7150# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2949 a_14922_4138# row_n[2] a_15414_4500# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2950 a_9902_15182# row_n[13] a_10394_15544# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2951 a_21342_13214# rowon_n[11] a_20946_13174# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X2952 vcm a_2275_11190# a_9994_11166# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2953 a_34394_12210# rowon_n[10] a_33998_12170# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X2954 a_31990_10162# a_2275_10186# a_32082_10162# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2955 a_9294_9198# rowon_n[7] a_8898_9158# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X2956 a_22954_12170# a_2275_12194# a_23046_12170# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2957 a_24354_5182# col_n[21] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2958 a_24050_6146# a_2475_6170# a_23958_6146# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X2959 a_21950_18194# a_2275_18218# a_22042_18194# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2960 VDD rowon_n[9] a_20946_11166# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2961 VDD rowon_n[8] a_33998_10162# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2962 a_25966_8154# row_n[6] a_26458_8516# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2963 VDD rowon_n[7] a_8898_9158# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2964 VSS VDD a_10298_1166# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X2965 VSS row_n[15] a_32386_17230# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X2966 a_23958_3134# row_n[1] a_24450_3496# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2967 a_20338_14218# col_n[17] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2968 a_2475_16210# a_1957_16210# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.342 pd=2.97 as=0.249 ps=1.62 w=1.2 l=0.15
X2969 a_33390_13214# col_n[30] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2970 a_12002_8154# a_2475_8178# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2971 a_28370_7190# col_n[25] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2972 a_29374_3174# col_n[26] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2973 a_13006_4138# a_2475_4162# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2974 a_27062_17190# a_2475_17214# a_26970_17190# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X2975 a_3270_16226# rowon_n[14] a_2874_16186# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X2976 a_13310_16226# rowon_n[14] a_12914_16186# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X2977 VSS row_n[11] a_10298_13214# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X2978 a_7286_6186# col_n[4] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2979 a_29070_4138# a_2475_4162# a_28978_4138# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X2980 a_19334_9198# col_n[16] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2981 a_27974_17190# row_n[15] a_28466_17552# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2982 a_32482_15544# col_n[29] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X2983 vcm a_2275_13198# a_28066_13174# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2984 a_32082_11166# a_2475_11190# a_31990_11166# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X2985 a_4882_15182# a_2275_15206# a_4974_15182# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2986 a_14922_15182# a_2275_15206# a_15014_15182# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2987 VSS row_n[7] a_20338_9198# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X2988 a_30378_9198# rowon_n[7] a_29982_9158# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X2989 VSS row_n[1] a_14314_3174# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X2990 a_32994_11166# row_n[9] a_33486_11528# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2991 a_28978_1126# VDD a_29470_1488# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2992 vcm a_2275_3158# a_32082_3134# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2993 a_10394_11528# col_n[7] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X2994 a_34090_9158# a_2475_9182# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2995 vcm a_2275_7174# a_31078_7150# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2996 VDD rowon_n[4] a_17934_6146# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X2997 a_29982_6146# row_n[4] a_30474_6508# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2998 a_8898_12170# row_n[10] a_9390_12532# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X2999 a_18938_12170# row_n[10] a_19430_12532# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3000 a_3970_7150# a_2475_7174# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3001 VDD VSS sky130_fd_pr__cap_mim_m3_1 l=17.2 w=17.2
X3002 a_4974_3134# a_2475_3158# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3003 a_17022_6146# a_2475_6170# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3004 a_22954_2130# a_2275_2154# a_23046_2130# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3005 VDD a_2161_4162# a_2275_4162# VDD sky130_fd_pr__pfet_01v8 ad=0.249 pd=1.62 as=0.342 ps=2.97 w=1.2 l=0.15
X3006 a_2161_13198# sample VSS VSS sky130_fd_pr__nfet_01v8 ad=0.171 pd=1.77 as=0.171 ps=1.77 w=0.6 l=0.15
X3007 a_18938_9158# row_n[7] a_19430_9520# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3008 a_33086_2130# a_2475_2154# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3009 vcm a_2275_16210# a_30074_16186# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3010 a_20434_9520# col_n[17] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X3011 a_12914_8154# a_2275_8178# a_13006_8154# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3012 a_14410_1488# col_n[11] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X3013 a_13918_4138# a_2275_4162# a_14010_4138# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3014 a_21438_5504# col_n[18] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X3015 VDD rowon_n[7] a_29982_9158# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3016 a_33390_1166# col_n[30] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3017 vcm a_2275_17214# a_16018_17190# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3018 vcm a_2275_17214# a_5978_17190# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3019 VSS row_n[13] a_28370_15222# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3020 a_32386_13214# rowon_n[11] a_31990_13174# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X3021 a_20034_17190# a_2475_17214# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3022 a_8990_5142# a_2475_5166# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3023 a_9994_1126# a_2475_1150# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3024 a_29374_11206# col_n[26] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3025 a_24050_16186# a_2475_16210# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3026 a_20946_13174# a_2275_13198# a_21038_13174# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3027 a_4882_7150# a_2275_7174# a_4974_7150# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3028 a_5886_3134# a_2275_3158# a_5978_3134# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3029 VDD rowon_n[15] a_26970_17190# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3030 a_15014_15182# a_2475_15206# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3031 a_33998_12170# a_2275_12194# a_34090_12170# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3032 a_25454_7512# col_n[22] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X3033 a_17934_6146# a_2275_6170# a_18026_6146# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3034 a_4974_15182# a_2475_15206# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3035 VDD rowon_n[5] a_35002_7150# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3036 a_8990_14178# a_2475_14202# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3037 a_28466_13536# col_n[25] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X3038 VDD rowon_n[9] a_31990_11166# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3039 VSS row_n[7] a_29374_9198# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3040 a_10998_4138# a_2475_4162# a_10906_4138# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X3041 a_23446_2492# col_n[20] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X3042 VSS VDD a_30378_18234# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3043 VSS row_n[0] a_28370_2170# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3044 a_31382_14218# col_n[28] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3045 a_32386_8194# col_n[29] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3046 VSS row_n[3] a_6282_5182# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3047 a_1957_2154# VSS sample VDD sky130_fd_pr__pfet_01v8 ad=0.342 pd=2.97 as=0.342 ps=2.97 w=1.2 l=0.15
X3048 a_25054_18194# a_2475_18218# a_24962_18194# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X3049 vcm a_2275_15206# a_22042_15182# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3050 a_32082_9158# a_2475_9182# a_31990_9158# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X3051 VSS row_n[6] a_18330_8194# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3052 a_16018_17190# a_2475_17214# a_15926_17190# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X3053 a_7286_15222# col_n[4] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3054 a_17326_15222# col_n[14] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3055 a_29470_9520# col_n[26] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X3056 a_25966_18194# VDD a_26458_18556# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3057 a_5978_17190# a_2475_17214# a_5886_17190# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X3058 vcm a_2275_14202# a_26058_14178# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3059 a_8386_8516# col_n[5] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X3060 a_2966_3134# a_2475_3158# a_2874_3134# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X3061 a_20338_4178# rowon_n[2] a_19942_4138# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X3062 a_12914_16186# a_2275_16210# a_13006_16186# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3063 a_30474_16548# col_n[27] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X3064 a_15014_6146# a_2475_6170# a_14922_6146# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X3065 vcm a_2275_2154# a_21038_2130# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3066 a_13310_2170# rowon_n[0] a_12914_2130# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X3067 a_24050_4138# a_2475_4162# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3068 a_2874_16186# a_2275_16210# a_2966_16186# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3069 a_9994_16186# a_2475_16210# a_9902_16186# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X3070 a_26970_7150# a_2275_7174# a_27062_7150# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3071 a_31078_2130# a_2475_2154# a_30986_2130# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X3072 a_6378_17552# col_n[3] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X3073 a_16418_17552# col_n[13] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X3074 vcm a_2275_8178# a_10998_8154# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3075 a_6378_3496# col_n[3] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X3076 vcm a_2275_4162# a_12002_4138# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3077 a_16930_13174# row_n[11] a_17422_13536# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3078 a_6890_13174# row_n[11] a_7382_13536# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3079 VDD rowon_n[2] a_19942_4138# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3080 vcm a_2275_12194# a_15014_12170# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3081 vcm a_2275_12194# a_4974_12170# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3082 a_24354_6186# rowon_n[4] a_23958_6146# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X3083 a_6982_5142# a_2475_5166# a_6890_5142# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X3084 a_7986_1126# a_2475_1150# a_7894_1126# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X3085 VSS row_n[8] a_27366_10202# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3086 vcm a_2275_18218# a_3970_18194# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3087 vcm a_2275_18218# a_14010_18194# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3088 a_27974_11166# a_2275_11190# a_28066_11166# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3089 vcm a_2275_7174# a_2966_7150# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3090 vcm a_2275_3158# a_3970_3134# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3091 vcm a_2275_6170# a_16018_6146# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3092 VSS row_n[14] a_26362_16226# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3093 a_30378_14218# rowon_n[12] a_29982_14178# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X3094 VDD rowon_n[10] a_25966_12170# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3095 a_31990_1126# a_2275_1150# a_32082_1126# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3096 a_30986_5142# a_2275_5166# a_31078_5142# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3097 a_31078_17190# a_2475_17214# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3098 a_35094_16186# a_2475_16210# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3099 a_31990_13174# a_2275_13198# a_32082_13174# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3100 a_5278_1166# col_n[2] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3101 VSS row_n[2] a_19334_4178# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3102 VDD VDD a_24962_18194# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3103 a_2966_16186# a_2475_16210# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3104 a_13006_16186# a_2475_16210# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3105 a_28370_8194# rowon_n[6] a_27974_8154# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X3106 a_29374_4178# rowon_n[2] a_28978_4138# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X3107 a_25358_15222# col_n[22] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3108 VDD rowon_n[6] a_14922_8154# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3109 vcm a_2275_5166# a_7986_5142# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3110 vcm a_2275_1150# a_8990_1126# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3111 a_21342_7190# col_n[18] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3112 a_22346_3174# col_n[19] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3113 a_8290_17230# rowon_n[15] a_7894_17190# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X3114 VDD a_2161_11190# a_2275_11190# VDD sky130_fd_pr__pfet_01v8 ad=0.249 pd=1.62 as=0.342 ps=2.97 w=1.2 l=0.15
X3115 VSS row_n[5] a_31382_7190# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3116 ctop sw_n ctop VSS sky130_fd_pr__nfet_01v8 ad=0.275 pd=2.19 as=2.76 ps=21.9 w=1.9 l=0.22
X3117 a_24450_17552# col_n[21] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X3118 a_20946_14178# row_n[12] a_21438_14540# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3119 VSS row_n[11] a_9294_13214# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3120 a_24050_13174# a_2475_13198# a_23958_13174# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X3121 a_6282_10202# col_n[3] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3122 a_16322_10202# col_n[13] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3123 vcm a_2275_10186# a_21038_10162# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3124 a_12306_9198# col_n[9] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3125 a_35002_7150# a_2275_7174# a_35094_7150# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3126 a_22042_4138# a_2475_4162# a_21950_4138# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X3127 a_4974_12170# a_2475_12194# a_4882_12170# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X3128 a_15014_12170# a_2475_12194# a_14922_12170# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X3129 a_28066_9158# a_2475_9182# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3130 a_17326_7190# rowon_n[5] a_16930_7150# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X3131 a_23958_6146# row_n[4] a_24450_6508# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3132 VDD rowon_n[2] a_28978_4138# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3133 a_19430_4500# col_n[16] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X3134 a_24962_13174# row_n[11] a_25454_13536# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3135 a_8990_11166# a_2475_11190# a_8898_11166# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X3136 VDD rowon_n[5] a_6890_7150# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3137 VDD rowon_n[13] a_7894_15182# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3138 a_5374_12532# col_n[2] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X3139 a_15414_12532# col_n[12] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X3140 a_21950_1126# VDD a_22442_1488# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3141 VDD rowon_n[0] a_4882_2130# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3142 a_9390_11528# col_n[6] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X3143 a_2475_10186# a_1957_10186# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.171 pd=1.77 as=0.124 ps=1.01 w=0.6 l=0.15
X3144 a_27366_1166# col_n[24] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3145 a_26362_5182# col_n[23] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3146 a_11910_9158# row_n[7] a_12402_9520# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3147 a_4274_8194# col_n[1] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3148 vcm a_2275_17214# a_35094_17190# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3149 a_27974_8154# row_n[6] a_28466_8516# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3150 a_12914_17190# row_n[15] a_13406_17552# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3151 a_24354_15222# rowon_n[13] a_23958_15182# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X3152 vcm a_2275_13198# a_13006_13174# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3153 VSS row_n[10] a_21342_12210# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3154 VSS VDD a_12306_1166# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3155 a_2874_17190# row_n[15] a_3366_17552# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3156 vcm a_2275_13198# a_2966_13174# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3157 a_25966_3134# row_n[1] a_26458_3496# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3158 a_28370_14218# rowon_n[12] a_27974_14178# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X3159 VSS row_n[9] a_25358_11206# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3160 a_2966_1126# a_2475_1150# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3161 a_15014_4138# a_2475_4162# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3162 a_29070_17190# a_2475_17214# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3163 VDD rowon_n[12] a_19942_14178# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3164 a_30074_12170# a_2475_12194# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3165 a_15318_10202# rowon_n[8] a_14922_10162# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X3166 a_14010_8154# a_2475_8178# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3167 a_16930_7150# row_n[5] a_17422_7512# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3168 a_9294_6186# col_n[6] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3169 a_5278_10202# rowon_n[8] a_4882_10162# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X3170 VDD rowon_n[11] a_23958_13174# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3171 a_21438_10524# col_n[18] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X3172 a_10906_6146# a_2275_6170# a_10998_6146# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3173 a_18330_3174# rowon_n[1] a_17934_3134# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X3174 VSS row_n[7] a_22346_9198# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3175 a_30378_3174# col_n[27] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3176 a_32386_9198# rowon_n[7] a_31990_9158# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X3177 a_23350_16226# col_n[20] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3178 vcm a_2275_7174# a_33086_7150# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3179 vcm a_2275_3158# a_34090_3134# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3180 a_14922_10162# a_2275_10186# a_15014_10162# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3181 a_26058_9158# a_2475_9182# a_25966_9158# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X3182 VSS row_n[0] a_21342_2170# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3183 a_6982_3134# a_2475_3158# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3184 a_4882_10162# a_2275_10186# a_4974_10162# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3185 a_6282_18234# VDD a_5886_18194# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X3186 a_16322_18234# VDD a_15926_18194# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X3187 VSS row_n[13] a_3270_15222# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3188 VSS row_n[13] a_13310_15222# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3189 a_35094_2130# a_2475_2154# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3190 a_3878_1126# a_2275_1150# a_3970_1126# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3191 VDD en_bit_n[1] a_17934_1126# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3192 a_29982_1126# VDD a_30474_1488# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3193 a_24962_2130# a_2275_2154# a_25054_2130# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3194 a_22442_18556# col_n[19] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X3195 VSS row_n[12] a_17326_14218# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3196 a_22042_14178# a_2475_14202# a_21950_14178# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X3197 a_14314_11206# col_n[11] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3198 VSS row_n[6] a_11302_8194# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3199 a_2874_5142# a_2275_5166# a_2966_5142# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3200 a_35494_17552# VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X3201 VSS row_n[12] a_7286_14218# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3202 a_31990_14178# row_n[12] a_32482_14540# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3203 a_13006_13174# a_2475_13198# a_12914_13174# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X3204 a_35094_13174# a_2475_13198# a_35002_13174# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X3205 a_4274_11206# col_n[1] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3206 vcm a_2275_10186# a_32082_10162# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3207 a_22442_9520# col_n[19] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X3208 a_14922_8154# a_2275_8178# a_15014_8154# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3209 a_35398_1166# VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3210 a_15926_4138# a_2275_4162# a_16018_4138# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3211 a_23446_5504# col_n[20] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X3212 a_17934_17190# a_2275_17214# a_18026_17190# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3213 a_2966_13174# a_2475_13198# a_2874_13174# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X3214 VDD rowon_n[7] a_31990_9158# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3215 a_7894_17190# a_2275_17214# a_7986_17190# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3216 VDD rowon_n[15] a_11910_17190# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3217 VDD rowon_n[14] a_15926_16186# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3218 a_13406_13536# col_n[10] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X3219 VDD rowon_n[14] a_5886_16186# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3220 a_3366_13536# col_n[0] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X3221 VSS row_n[5] a_3270_7190# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3222 vcm a_2275_18218# a_33086_18194# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3223 VSS row_n[4] a_16322_6186# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3224 a_7894_3134# a_2275_3158# a_7986_3134# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3225 VSS row_n[10] a_19334_12210# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3226 a_27462_7512# col_n[24] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X3227 a_24050_11166# a_2475_11190# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3228 a_23350_10202# rowon_n[8] a_22954_10162# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X3229 a_6378_6508# col_n[3] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X3230 a_13006_4138# a_2475_4162# a_12914_4138# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X3231 a_15014_10162# a_2475_10186# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3232 a_12002_8154# a_2475_8178# a_11910_8154# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X3233 a_25454_2492# col_n[22] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X3234 a_10906_18194# VDD a_11398_18556# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3235 a_22346_16226# rowon_n[14] a_21950_16186# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X3236 a_35398_15222# rowon_n[13] a_35002_15182# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X3237 vcm a_2275_14202# a_10998_14178# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3238 a_4974_10162# a_2475_10186# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3239 VDD rowon_n[0] a_35002_2130# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3240 VDD rowon_n[12] a_17934_14178# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3241 a_34394_8194# col_n[31] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3242 a_27062_18194# a_2475_18218# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3243 a_23958_15182# a_2275_15206# a_24050_15182# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3244 a_19430_10524# col_n[16] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X3245 VSS row_n[3] a_8290_5182# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3246 a_18026_17190# a_2475_17214# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3247 a_34090_9158# a_2475_9182# a_33998_9158# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X3248 a_7986_17190# a_2475_17214# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3249 a_27974_14178# a_2275_14202# a_28066_14178# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3250 a_21342_8194# rowon_n[6] a_20946_8154# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X3251 a_4974_3134# a_2475_3158# a_4882_3134# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X3252 a_22346_4178# rowon_n[2] a_21950_4138# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X3253 VDD rowon_n[11] a_35002_13174# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3254 a_3970_7150# a_2475_7174# a_3878_7150# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X3255 vcm a_2275_2154# a_23046_2130# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3256 a_10298_4178# col_n[7] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3257 a_35398_10202# VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3258 a_17022_6146# a_2475_6170# a_16930_6146# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X3259 a_33086_2130# a_2475_2154# a_32994_2130# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X3260 a_28978_7150# a_2275_7174# a_29070_7150# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3261 a_8386_3496# col_n[5] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X3262 VSS row_n[8] a_12306_10202# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3263 vcm a_2275_8178# a_13006_8154# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3264 vcm a_2275_4162# a_14010_4138# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3265 a_34394_16226# col_n[31] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3266 a_2874_11166# a_2275_11190# a_2966_11166# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3267 a_12914_11166# a_2275_11190# a_13006_11166# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3268 VSS row_n[14] a_11302_16226# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3269 a_34490_12532# col_n[31] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X3270 a_21038_9158# a_2475_9182# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3271 a_10298_7190# rowon_n[5] a_9902_7150# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X3272 VDD rowon_n[2] a_21950_4138# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3273 vcm a_2275_16210# a_29070_16186# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3274 a_33086_14178# a_2475_14202# a_32994_14178# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X3275 VDD rowon_n[10] a_10906_12170# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3276 a_26362_6186# rowon_n[4] a_25966_6146# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X3277 a_9994_1126# a_2475_1150# a_9902_1126# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X3278 a_9902_4138# row_n[2] a_10394_4500# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3279 a_33486_18556# col_n[30] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X3280 a_10998_14178# a_2475_14202# a_10906_14178# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X3281 a_8990_5142# a_2475_5166# a_8898_5142# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X3282 a_5886_18194# a_2275_18218# a_5978_18194# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3283 VDD VDD a_9902_18194# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3284 a_15926_18194# a_2275_18218# a_16018_18194# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3285 a_4274_9198# rowon_n[7] a_3878_9158# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X3286 a_10298_15222# col_n[7] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3287 vcm a_2275_7174# a_4974_7150# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3288 vcm a_2275_3158# a_5978_3134# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3289 vcm a_2275_6170# a_18026_6146# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3290 a_2475_2154# a_1957_2154# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.342 pd=2.97 as=0.249 ps=1.62 w=1.2 l=0.15
X3291 a_15318_5182# rowon_n[3] a_14922_5142# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X3292 a_32994_5142# a_2275_5166# a_33086_5142# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3293 a_20946_8154# row_n[6] a_21438_8516# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3294 VDD rowon_n[7] a_3878_9158# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3295 a_31478_8516# col_n[28] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X3296 VDD rowon_n[3] a_4882_5142# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3297 a_9902_13174# row_n[11] a_10394_13536# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3298 a_21342_11206# rowon_n[9] a_20946_11166# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X3299 VDD rowon_n[6] a_16930_8154# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3300 a_35094_11166# a_2475_11190# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3301 a_34394_10202# rowon_n[8] a_33998_10162# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X3302 a_2966_11166# a_2475_11190# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3303 a_13006_11166# a_2475_11190# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3304 a_23350_7190# col_n[20] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3305 a_24354_3174# col_n[21] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3306 VDD rowon_n[1] a_14922_3134# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3307 VDD rowon_n[12] a_28978_14178# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3308 a_17022_12170# a_2475_12194# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3309 VSS row_n[5] a_33390_7190# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3310 a_24050_4138# a_2475_4162# a_23958_4138# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X3311 a_6982_12170# a_2475_12194# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3312 a_14314_9198# col_n[11] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3313 vcm a_2275_7174# a_27062_7150# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3314 a_21950_16186# a_2275_16210# a_22042_16186# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3315 a_25966_6146# row_n[4] a_26458_6508# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3316 a_5978_18194# a_2475_18218# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3317 a_16018_18194# a_2475_18218# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3318 VDD rowon_n[5] a_8898_7150# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3319 a_28370_17230# col_n[25] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3320 VSS row_n[13] a_32386_15222# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3321 a_23958_1126# VDD a_24450_1488# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3322 a_2475_14202# a_1957_14202# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.342 pd=2.97 as=0.249 ps=1.62 w=1.2 l=0.15
X3323 a_33390_11206# col_n[30] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3324 VDD rowon_n[0] a_6890_2130# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3325 a_13310_14218# rowon_n[12] a_12914_14178# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X3326 a_12002_6146# a_2475_6170# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3327 a_29374_1166# col_n[26] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3328 a_28370_5182# col_n[25] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3329 VDD rowon_n[15] a_30986_17190# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3330 a_27062_15182# a_2475_15206# a_26970_15182# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X3331 a_3270_14218# rowon_n[12] a_2874_14178# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X3332 a_9294_12210# col_n[6] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3333 a_19334_12210# col_n[16] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3334 vcm a_2275_12194# a_24050_12170# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3335 VSS row_n[9] a_10298_11206# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3336 a_13918_9158# row_n[7] a_14410_9520# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3337 a_6282_8194# col_n[3] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3338 a_7286_4178# col_n[4] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3339 vcm a_2275_11190# a_28066_11166# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3340 a_27974_15182# row_n[13] a_28466_15544# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3341 a_32482_13536# col_n[29] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X3342 a_4882_13174# a_2275_13198# a_4974_13174# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3343 a_14922_13174# a_2275_13198# a_15014_13174# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3344 VSS VDD a_14314_1166# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3345 a_8386_14540# col_n[5] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X3346 a_18426_14540# col_n[15] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X3347 vcm a_2275_1150# a_32082_1126# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3348 a_27974_3134# row_n[1] a_28466_3496# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3349 vcm a_2275_5166# a_31078_5142# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3350 a_8898_10162# row_n[8] a_9390_10524# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3351 a_18938_10162# row_n[8] a_19430_10524# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3352 a_3970_5142# a_2475_5166# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3353 a_4974_1126# a_2475_1150# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3354 a_6890_4138# row_n[2] a_7382_4500# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3355 a_17022_4138# a_2475_4162# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3356 a_18938_7150# row_n[5] a_19430_7512# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3357 a_29982_18194# VDD a_30474_18556# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3358 vcm a_2275_14202# a_30074_14178# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3359 a_20434_7512# col_n[17] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X3360 a_12914_6146# a_2275_6170# a_13006_6146# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3361 VDD rowon_n[5] a_29982_7150# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3362 a_16930_2130# row_n[0] a_17422_2492# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3363 a_27366_17230# rowon_n[15] a_26970_17190# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X3364 vcm a_2275_15206# a_16018_15182# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3365 VSS row_n[7] a_24354_9198# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3366 vcm a_2275_15206# a_5978_15182# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3367 a_34394_9198# rowon_n[7] a_33998_9158# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X3368 VSS row_n[11] a_28370_13214# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3369 a_32386_11206# rowon_n[9] a_31990_11166# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X3370 a_28066_9158# a_2475_9182# a_27974_9158# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X3371 vcm a_2275_7174# a_35094_7150# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3372 a_20034_15182# a_2475_15206# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3373 VSS row_n[0] a_23350_2170# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3374 a_8990_3134# a_2475_3158# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3375 a_24050_14178# a_2475_14202# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3376 VSS row_n[6] a_13310_8194# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3377 a_19030_8154# a_2475_8178# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3378 a_4882_5142# a_2275_5166# a_4974_5142# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3379 a_5886_1126# a_2275_1150# a_5978_1126# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3380 VDD rowon_n[13] a_26970_15182# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3381 a_15014_13174# a_2475_13198# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3382 a_24450_9520# col_n[21] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X3383 a_17934_4138# a_2275_4162# a_18026_4138# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3384 a_25454_5504# col_n[22] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X3385 a_4974_13174# a_2475_13198# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3386 VDD rowon_n[7] a_33998_9158# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3387 a_3366_8516# col_n[0] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X3388 VDD rowon_n[3] a_35002_5142# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3389 a_28466_11528# col_n[25] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X3390 VSS a_2161_9182# a_2275_9182# VSS sky130_fd_pr__nfet_01v8 ad=0.124 pd=1.01 as=0.171 ps=1.77 w=0.6 l=0.15
X3391 a_21950_7150# a_2275_7174# a_22042_7150# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3392 a_26362_18234# col_n[23] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3393 VSS row_n[14] a_30378_16226# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3394 VSS row_n[15] a_6282_17230# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3395 VSS row_n[15] a_16322_17230# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3396 a_21038_17190# a_2475_17214# a_20946_17190# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X3397 VSS row_n[5] a_5278_7190# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3398 a_32386_6186# col_n[29] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3399 VSS row_n[1] a_6282_3174# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3400 a_35002_18194# a_2275_18218# a_35094_18194# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3401 a_25054_16186# a_2475_16210# a_24962_16186# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X3402 a_17326_13214# col_n[14] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3403 vcm a_2275_13198# a_22042_13174# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3404 VSS row_n[4] a_18330_6186# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3405 a_21950_17190# row_n[15] a_22442_17552# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3406 a_1957_16210# VDD sample VSS sky130_fd_pr__nfet_01v8 ad=0.171 pd=1.77 as=0.171 ps=1.77 w=0.6 l=0.15
X3407 a_16018_15182# a_2475_15206# a_15926_15182# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X3408 a_7286_13214# col_n[4] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3409 a_29470_7512# col_n[26] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X3410 a_25966_16186# row_n[14] a_26458_16548# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3411 a_5978_15182# a_2475_15206# a_5886_15182# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X3412 a_8386_6508# col_n[5] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X3413 a_2966_1126# a_2475_1150# a_2874_1126# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X3414 a_12914_14178# a_2275_14202# a_13006_14178# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3415 a_14010_8154# a_2475_8178# a_13918_8154# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X3416 a_15014_4138# a_2475_4162# a_14922_4138# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X3417 a_16418_15544# col_n[13] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X3418 a_2874_14178# a_2275_14202# a_2966_14178# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3419 a_9994_14178# a_2475_14202# a_9902_14178# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X3420 a_27462_2492# col_n[24] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X3421 a_26970_5142# a_2275_5166# a_27062_5142# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3422 VDD VDD a_8898_18194# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3423 a_6378_15544# col_n[3] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X3424 vcm a_2275_6170# a_10998_6146# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3425 a_6378_1488# col_n[3] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X3426 a_16930_11166# row_n[9] a_17422_11528# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3427 a_6890_11166# row_n[9] a_7382_11528# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3428 vcm a_2275_10186# a_15014_10162# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3429 a_4882_14178# row_n[12] a_5374_14540# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3430 a_14922_14178# row_n[12] a_15414_14540# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3431 a_26362_12210# rowon_n[10] a_25966_12170# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X3432 vcm a_2275_10186# a_4974_10162# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3433 a_23958_10162# a_2275_10186# a_24050_10162# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3434 a_23350_8194# rowon_n[6] a_22954_8154# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X3435 a_6982_3134# a_2475_3158# a_6890_3134# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X3436 a_24354_4178# rowon_n[2] a_23958_4138# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X3437 VDD rowon_n[6] a_9902_8154# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3438 vcm a_2275_2154# a_25054_2130# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3439 a_25358_18234# VDD a_24962_18194# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X3440 a_1957_17214# VSS sample VDD sky130_fd_pr__pfet_01v8 ad=0.342 pd=2.97 as=0.342 ps=2.97 w=1.2 l=0.15
X3441 vcm a_2275_16210# a_3970_16186# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3442 vcm a_2275_16210# a_14010_16186# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3443 vcm a_2275_5166# a_2966_5142# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3444 a_35094_2130# a_2475_2154# a_35002_2130# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X3445 vcm a_2275_1150# a_3970_1126# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3446 vcm a_2275_8178# a_15014_8154# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3447 vcm a_2275_4162# a_16018_4138# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3448 VSS row_n[12] a_26362_14218# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3449 a_26970_17190# a_2275_17214# a_27062_17190# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3450 VDD rowon_n[8] a_25966_10162# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3451 a_29982_7150# a_2275_7174# a_30074_7150# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3452 a_30986_3134# a_2275_3158# a_31078_3134# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3453 a_31078_15182# a_2475_15206# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3454 a_23046_9158# a_2475_9182# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3455 a_12306_7190# rowon_n[5] a_11910_7150# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X3456 VDD rowon_n[2] a_23958_4138# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3457 VSS row_n[15] a_24354_17230# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3458 a_35094_14178# a_2475_14202# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3459 VDD rowon_n[14] a_24962_16186# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3460 a_2966_14178# a_2475_14202# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3461 a_13006_14178# a_2475_14202# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3462 a_28370_6186# rowon_n[4] a_27974_6146# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X3463 a_25358_13214# col_n[22] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3464 a_6282_9198# rowon_n[7] a_5886_9158# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X3465 VDD rowon_n[4] a_14922_6146# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3466 vcm a_2275_3158# a_7986_3134# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3467 a_19030_17190# a_2475_17214# a_18938_17190# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X3468 VSS row_n[10] a_15318_12210# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3469 a_20034_12170# a_2475_12194# a_19942_12170# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X3470 a_22346_1166# col_n[19] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3471 a_21342_5182# col_n[18] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3472 a_8290_15222# rowon_n[13] a_7894_15182# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X3473 VSS row_n[10] a_5278_12210# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3474 a_5278_2170# rowon_n[0] a_4882_2130# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X3475 VSS row_n[3] a_31382_5182# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3476 a_24450_15544# col_n[21] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X3477 a_20946_12170# row_n[10] a_21438_12532# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3478 VSS row_n[9] a_9294_11206# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3479 a_24050_11166# a_2475_11190# a_23958_11166# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X3480 ctop sw_n ctop VSS sky130_fd_pr__nfet_01v8 ad=0.275 pd=2.19 as=0 ps=0 w=1.9 l=0.22
X3481 a_35002_5142# a_2275_5166# a_35094_5142# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3482 a_4974_10162# a_2475_10186# a_4882_10162# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X3483 a_15014_10162# a_2475_10186# a_14922_10162# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X3484 a_22954_8154# row_n[6] a_23446_8516# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3485 a_17326_5182# rowon_n[3] a_16930_5142# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X3486 VDD rowon_n[12] a_13918_14178# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3487 a_24962_11166# row_n[9] a_25454_11528# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3488 a_33486_8516# col_n[30] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X3489 VDD rowon_n[12] a_3878_14178# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3490 VDD rowon_n[7] a_5886_9158# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3491 VDD rowon_n[3] a_6890_5142# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3492 VDD rowon_n[11] a_7894_13174# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3493 a_5374_10524# col_n[2] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X3494 a_15414_10524# col_n[12] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X3495 a_20946_3134# row_n[1] a_21438_3496# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3496 a_13310_17230# col_n[10] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3497 a_31478_3496# col_n[28] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X3498 a_3270_17230# col_n[0] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3499 a_26362_3174# col_n[23] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3500 VDD rowon_n[1] a_16930_3134# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3501 a_11910_7150# row_n[5] a_12402_7512# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3502 a_25358_7190# col_n[22] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3503 VSS row_n[5] a_35398_7190# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3504 a_4274_6186# col_n[1] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3505 vcm a_2275_15206# a_35094_15182# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3506 a_16322_9198# col_n[13] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3507 vcm a_2275_7174# a_29070_7150# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3508 a_27974_6146# row_n[4] a_28466_6508# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3509 a_12914_15182# row_n[13] a_13406_15544# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3510 a_24354_13214# rowon_n[11] a_23958_13174# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X3511 vcm a_2275_11190# a_13006_11166# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3512 VSS row_n[8] a_21342_10202# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3513 a_2874_15182# row_n[13] a_3366_15544# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3514 vcm a_2275_11190# a_2966_11166# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3515 a_21950_11166# a_2275_11190# a_22042_11166# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3516 a_25966_1126# VDD a_26458_1488# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3517 a_21038_9158# a_2475_9182# a_20946_9158# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X3518 VDD rowon_n[0] a_8898_2130# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3519 VDD rowon_n[15] a_18938_17190# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3520 a_29070_15182# a_2475_15206# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3521 VDD rowon_n[10] a_19942_12170# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3522 a_25966_12170# a_2275_12194# a_26058_12170# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3523 a_15926_9158# row_n[7] a_16418_9520# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3524 a_14010_6146# a_2475_6170# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3525 a_16930_5142# row_n[3] a_17422_5504# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3526 a_30074_2130# a_2475_2154# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3527 a_19942_2130# a_2275_2154# a_20034_2130# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3528 a_9294_4178# col_n[6] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3529 a_8290_8194# col_n[5] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3530 VDD rowon_n[9] a_23958_11166# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3531 a_9902_8154# a_2275_8178# a_9994_8154# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3532 a_18330_1166# en_bit_n[1] a_17934_1126# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X3533 a_30378_1166# col_n[27] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3534 a_10906_4138# a_2275_4162# a_10998_4138# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3535 VSS VDD a_22346_18234# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3536 VSS row_n[15] a_35398_17230# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3537 a_23350_14218# col_n[20] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3538 vcm a_2275_5166# a_33086_5142# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3539 a_12306_17230# rowon_n[15] a_11910_17190# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X3540 a_6982_1126# a_2475_1150# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3541 a_8898_4138# row_n[2] a_9390_4500# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3542 a_6282_16226# rowon_n[14] a_5886_16186# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X3543 a_16322_16226# rowon_n[14] a_15926_16186# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X3544 VSS row_n[11] a_3270_13214# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3545 VSS row_n[11] a_13310_13214# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3546 a_31078_12170# a_2475_12194# a_30986_12170# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X3547 a_22442_16548# col_n[19] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X3548 VSS row_n[4] a_11302_6186# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3549 a_2874_3134# a_2275_3158# a_2966_3134# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3550 a_35494_15544# VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X3551 a_31990_12170# row_n[10] a_32482_12532# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3552 a_13006_11166# a_2475_11190# a_12914_11166# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X3553 a_35094_11166# a_2475_11190# a_35002_11166# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X3554 a_22442_7512# col_n[19] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X3555 a_14922_6146# a_2275_6170# a_15014_6146# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3556 a_7894_15182# a_2275_15206# a_7986_15182# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3557 a_17934_15182# a_2275_15206# a_18026_15182# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3558 a_2966_11166# a_2475_11190# a_2874_11166# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X3559 VDD rowon_n[5] a_31990_7150# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3560 a_18938_2130# row_n[0] a_19430_2492# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3561 VDD rowon_n[13] a_11910_15182# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3562 a_20434_2492# col_n[17] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X3563 a_13406_11528# col_n[10] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X3564 VDD rowon_n[0] a_29982_2130# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3565 a_3366_11528# col_n[0] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X3566 a_11302_18234# col_n[8] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3567 a_35398_2170# rowon_n[0] a_35002_2130# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X3568 VSS row_n[0] a_25358_2170# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3569 VSS row_n[3] a_3270_5182# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3570 vcm a_2275_16210# a_33086_16186# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3571 a_20034_10162# a_2475_10186# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3572 VSS row_n[6] a_15318_8194# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3573 a_7894_1126# a_2275_1150# a_7986_1126# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3574 VSS row_n[2] a_16322_4178# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3575 VSS row_n[8] a_19334_10202# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3576 a_27462_5504# col_n[24] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X3577 vcm a_2275_17214# a_19030_17190# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3578 a_5374_8516# col_n[2] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X3579 a_5978_8154# a_2475_8178# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3580 vcm a_2275_17214# a_8990_17190# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3581 a_12002_6146# a_2475_6170# a_11910_6146# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X3582 a_10906_16186# row_n[14] a_11398_16548# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3583 a_22346_14218# rowon_n[12] a_21950_14178# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X3584 a_35398_13214# rowon_n[11] a_35002_13174# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X3585 a_23958_7150# a_2275_7174# a_24050_7150# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3586 a_3366_3496# col_n[0] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X3587 a_23046_17190# a_2475_17214# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3588 VDD rowon_n[10] a_17934_12170# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3589 a_34394_6186# col_n[31] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3590 a_16418_4500# col_n[13] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X3591 a_27062_16186# a_2475_16210# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3592 a_23958_13174# a_2275_13198# a_24050_13174# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3593 VSS row_n[5] a_7286_7190# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3594 VSS row_n[1] a_8290_3174# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3595 a_18026_15182# a_2475_15206# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3596 a_1957_8178# VDD sample VSS sky130_fd_pr__nfet_01v8 ad=0.171 pd=1.77 as=0.171 ps=1.77 w=0.6 l=0.15
X3597 a_7986_15182# a_2475_15206# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3598 a_21342_6186# rowon_n[4] a_20946_6146# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X3599 a_4974_1126# a_2475_1150# a_4882_1126# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X3600 a_2161_2154# sample VDD VDD sky130_fd_pr__pfet_01v8 ad=0.342 pd=2.97 as=0.342 ps=2.97 w=1.2 l=0.15
X3601 VSS row_n[10] a_34394_12210# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3602 VDD rowon_n[9] a_35002_11166# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3603 a_3970_5142# a_2475_5166# a_3878_5142# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X3604 a_11302_12210# rowon_n[10] a_10906_12170# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X3605 a_1957_11190# VDD sample VSS sky130_fd_pr__nfet_01v8 ad=0.171 pd=1.77 as=0.171 ps=1.77 w=0.6 l=0.15
X3606 a_17022_4138# a_2475_4162# a_16930_4138# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X3607 VSS VDD a_33390_18234# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3608 a_8386_1488# col_n[5] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X3609 a_29470_2492# col_n[26] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X3610 a_28978_5142# a_2275_5166# a_29070_5142# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3611 a_29070_12170# a_2475_12194# a_28978_12170# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X3612 a_6890_8154# a_2275_8178# a_6982_8154# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3613 vcm a_2275_6170# a_13006_6146# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3614 a_10298_18234# VDD a_9902_18194# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X3615 VDD rowon_n[12] a_32994_14178# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3616 a_34394_14218# col_n[31] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3617 a_28066_18194# a_2475_18218# a_27974_18194# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X3618 VSS row_n[12] a_11302_14218# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3619 a_34490_10524# col_n[31] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X3620 a_10298_5182# rowon_n[3] a_9902_5142# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X3621 a_28978_18194# VDD a_29470_18556# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3622 a_11910_17190# a_2275_17214# a_12002_17190# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3623 vcm a_2275_14202# a_29070_14178# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3624 VDD rowon_n[8] a_10906_10162# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3625 a_26362_4178# rowon_n[2] a_25966_4138# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X3626 a_15926_16186# a_2275_16210# a_16018_16186# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3627 a_33486_16548# col_n[30] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X3628 VDD rowon_n[6] a_11910_8154# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3629 a_8990_3134# a_2475_3158# a_8898_3134# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X3630 a_5886_16186# a_2275_16210# a_5978_16186# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3631 VDD rowon_n[14] a_9902_16186# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3632 a_19030_8154# a_2475_8178# a_18938_8154# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X3633 a_10298_13214# col_n[7] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3634 vcm a_2275_5166# a_4974_5142# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3635 vcm a_2275_1150# a_5978_1126# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3636 VDD rowon_n[1] a_9902_3134# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3637 vcm a_2275_4162# a_18026_4138# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3638 a_25054_9158# a_2475_9182# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3639 a_14314_7190# rowon_n[5] a_13918_7150# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X3640 vcm a_2275_7174# a_22042_7150# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3641 a_32994_3134# a_2275_3158# a_33086_3134# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3642 a_15318_3174# rowon_n[1] a_14922_3134# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X3643 vcm a_2275_12194# a_18026_12170# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3644 a_20946_6146# row_n[4] a_21438_6508# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3645 VDD rowon_n[2] a_25966_4138# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3646 vcm a_2275_12194# a_7986_12170# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3647 VDD rowon_n[5] a_3878_7150# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3648 a_31478_6508# col_n[28] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X3649 a_9902_11166# row_n[9] a_10394_11528# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3650 a_31078_10162# a_2475_10186# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3651 VDD rowon_n[4] a_16930_6146# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3652 vcm a_2275_18218# a_6982_18194# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3653 vcm a_2275_18218# a_17022_18194# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3654 a_8290_9198# rowon_n[7] a_7894_9158# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X3655 a_22042_12170# a_2475_12194# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3656 VDD VSS a_14922_1126# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3657 a_24354_1166# col_n[21] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3658 a_23350_5182# col_n[20] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3659 a_21038_18194# a_2475_18218# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3660 VDD rowon_n[10] a_28978_12170# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3661 a_7286_2170# rowon_n[0] a_6890_2130# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X3662 VSS row_n[3] a_33390_5182# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3663 vcm a_2275_5166# a_27062_5142# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3664 a_31382_17230# rowon_n[15] a_30986_17190# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X3665 a_21950_14178# a_2275_14202# a_22042_14178# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3666 a_24962_8154# row_n[6] a_25454_8516# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3667 a_5978_16186# a_2475_16210# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3668 a_16018_16186# a_2475_16210# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3669 VDD rowon_n[7] a_7894_9158# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3670 a_35494_8516# VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X3671 VDD rowon_n[3] a_8898_5142# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3672 a_28370_15222# col_n[25] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3673 VSS row_n[11] a_32386_13214# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3674 a_19942_17190# a_2275_17214# a_20034_17190# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3675 a_33486_3496# col_n[30] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X3676 a_22954_3134# row_n[1] a_23446_3496# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3677 a_28370_3174# col_n[25] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3678 a_12002_4138# a_2475_4162# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3679 a_27462_17552# col_n[24] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X3680 VDD rowon_n[13] a_30986_15182# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3681 a_23958_14178# row_n[12] a_24450_14540# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3682 a_27062_13174# a_2475_13198# a_26970_13174# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X3683 a_9294_10202# col_n[6] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3684 a_19334_10202# col_n[16] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3685 vcm a_2275_10186# a_24050_10162# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3686 a_13918_7150# row_n[5] a_14410_7512# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3687 a_6282_6186# col_n[3] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3688 a_7986_12170# a_2475_12194# a_7894_12170# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X3689 a_10906_12170# a_2275_12194# a_10998_12170# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3690 a_18026_12170# a_2475_12194# a_17934_12170# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X3691 a_18330_9198# col_n[15] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3692 a_27974_13174# row_n[11] a_28466_13536# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3693 a_32482_11528# col_n[29] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X3694 a_11910_2130# row_n[0] a_12402_2492# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3695 a_30378_18234# col_n[27] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3696 a_8386_12532# col_n[5] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X3697 a_18426_12532# col_n[15] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X3698 a_17326_2170# col_n[14] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3699 a_23046_9158# a_2475_9182# a_22954_9158# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X3700 vcm a_2275_7174# a_30074_7150# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3701 a_27974_1126# VDD a_28466_1488# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3702 vcm a_2275_3158# a_31078_3134# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3703 VDD VSS sky130_fd_pr__cap_mim_m3_1 l=17.2 w=17.2
X3704 a_3970_3134# a_2475_3158# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3705 vcm a_2275_18218# a_25054_18194# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3706 a_17934_9158# row_n[7] a_18426_9520# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3707 a_18938_5142# row_n[3] a_19430_5504# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3708 a_32082_2130# a_2475_2154# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3709 a_29982_16186# row_n[14] a_30474_16548# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3710 a_12914_4138# a_2275_4162# a_13006_4138# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3711 a_20434_5504# col_n[17] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X3712 a_29070_10162# a_2475_10186# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3713 VDD rowon_n[3] a_29982_5142# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3714 a_15926_17190# row_n[15] a_16418_17552# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3715 a_27366_15222# rowon_n[13] a_26970_15182# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X3716 vcm a_2275_13198# a_16018_13174# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3717 a_5886_17190# row_n[15] a_6378_17552# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3718 vcm a_2275_13198# a_5978_13174# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3719 VSS row_n[9] a_28370_11206# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3720 vcm a_2275_5166# a_35094_5142# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3721 a_19030_18194# a_2475_18218# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3722 a_20034_13174# a_2475_13198# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3723 a_8990_1126# a_2475_1150# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3724 a_10998_12170# a_2475_12194# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3725 a_33086_12170# a_2475_12194# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3726 VSS row_n[4] a_13310_6186# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3727 a_19030_6146# a_2475_6170# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3728 a_4882_3134# a_2275_3158# a_4974_3134# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3729 VDD rowon_n[11] a_26970_13174# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3730 a_24450_7512# col_n[21] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X3731 VDD rowon_n[5] a_33998_7150# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3732 a_3366_6508# col_n[0] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X3733 a_22346_17230# col_n[19] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3734 a_2161_12194# sample VDD VDD sky130_fd_pr__pfet_01v8 ad=0.342 pd=2.97 as=0.342 ps=2.97 w=1.2 l=0.15
X3735 a_16018_9158# a_2475_9182# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3736 VSS a_2161_7174# a_2275_7174# VSS sky130_fd_pr__nfet_01v8 ad=0.124 pd=1.01 as=0.171 ps=1.77 w=0.6 l=0.15
X3737 a_22442_2492# col_n[19] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X3738 a_21950_5142# a_2275_5166# a_22042_5142# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3739 a_26362_16226# col_n[23] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3740 VSS row_n[12] a_30378_14218# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3741 a_17934_10162# a_2275_10186# a_18026_10162# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3742 VDD rowon_n[0] a_31990_2130# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3743 a_30986_17190# a_2275_17214# a_31078_17190# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3744 a_7894_10162# a_2275_10186# a_7986_10162# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3745 VSS row_n[0] a_27366_2170# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3746 a_9294_18234# VDD a_8898_18194# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X3747 VSS row_n[13] a_6282_15222# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3748 VSS row_n[13] a_16322_15222# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3749 a_21038_15182# a_2475_15206# a_20946_15182# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X3750 a_19334_8194# rowon_n[6] a_18938_8154# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X3751 a_31382_8194# col_n[28] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3752 VSS row_n[3] a_5278_5182# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3753 VSS VDD a_6282_1166# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3754 a_32386_4178# col_n[29] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3755 a_35002_16186# a_2275_16210# a_35094_16186# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3756 a_25054_14178# a_2475_14202# a_24962_14178# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X3757 a_17326_11206# col_n[14] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3758 vcm a_2275_11190# a_22042_11166# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3759 VSS row_n[2] a_18330_4178# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3760 a_25454_18556# col_n[22] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X3761 a_21950_15182# row_n[13] a_22442_15544# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3762 a_1957_14202# VDD sample VSS sky130_fd_pr__nfet_01v8 ad=0.171 pd=1.77 as=0.171 ps=1.77 w=0.6 l=0.15
X3763 a_16018_13174# a_2475_13198# a_15926_13174# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X3764 a_7286_11206# col_n[4] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3765 VSS row_n[6] a_17326_8194# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3766 a_29470_5504# col_n[26] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X3767 a_5978_13174# a_2475_13198# a_5886_13174# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X3768 a_7382_8516# col_n[4] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X3769 VDD rowon_n[15] a_4882_17190# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3770 VDD rowon_n[15] a_14922_17190# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3771 a_7986_8154# a_2475_8178# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3772 a_14010_6146# a_2475_6170# a_13918_6146# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X3773 vcm a_2275_2154# a_20034_2130# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3774 a_16418_13536# col_n[13] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X3775 a_25966_7150# a_2275_7174# a_26058_7150# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3776 a_30074_2130# a_2475_2154# a_29982_2130# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X3777 a_26970_3134# a_2275_3158# a_27062_3134# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3778 VDD rowon_n[14] a_8898_16186# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3779 a_6378_13536# col_n[3] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X3780 vcm a_2275_8178# a_9994_8154# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3781 a_5374_3496# col_n[2] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X3782 a_31990_4138# row_n[2] a_32482_4500# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3783 vcm a_2275_4162# a_10998_4138# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3784 a_16930_9158# a_2275_9182# a_17022_9158# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3785 a_18426_4500# col_n[15] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X3786 VSS row_n[5] a_9294_7190# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3787 a_4882_12170# row_n[10] a_5374_12532# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3788 a_14922_12170# row_n[10] a_15414_12532# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3789 a_27062_11166# a_2475_11190# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3790 a_26362_10202# rowon_n[8] a_25966_10162# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X3791 a_23350_6186# rowon_n[4] a_22954_6146# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X3792 a_6982_1126# a_2475_1150# a_6890_1126# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X3793 a_18026_10162# a_2475_10186# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3794 VDD rowon_n[4] a_9902_6146# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3795 a_3878_18194# VDD a_4370_18556# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3796 a_13918_18194# VDD a_14410_18556# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3797 a_25358_16226# rowon_n[14] a_24962_16186# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X3798 a_1957_15206# VSS sample VDD sky130_fd_pr__pfet_01v8 ad=0.342 pd=2.97 as=0.342 ps=2.97 w=1.2 l=0.15
X3799 vcm a_2275_14202# a_3970_14178# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3800 vcm a_2275_14202# a_14010_14178# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3801 a_7986_10162# a_2475_10186# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3802 vcm a_2275_3158# a_2966_3134# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3803 a_8898_8154# a_2275_8178# a_8990_8154# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3804 vcm a_2275_6170# a_15014_6146# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3805 a_26970_15182# a_2275_15206# a_27062_15182# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3806 a_31078_13174# a_2475_13198# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3807 a_30986_1126# a_2275_1150# a_31078_1126# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3808 a_29982_5142# a_2275_5166# a_30074_5142# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3809 a_12306_5182# rowon_n[3] a_11910_5142# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X3810 VSS row_n[13] a_24354_15222# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3811 a_21342_12210# col_n[18] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3812 a_28370_4178# rowon_n[2] a_27974_4138# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X3813 a_25358_11206# col_n[22] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3814 VDD rowon_n[6] a_13918_8154# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3815 vcm a_2275_1150# a_7986_1126# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3816 VDD rowon_n[15] a_22954_17190# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3817 a_19030_15182# a_2475_15206# a_18938_15182# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X3818 a_20434_14540# col_n[17] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X3819 a_29982_12170# a_2275_12194# a_30074_12170# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3820 VSS row_n[8] a_15318_10202# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3821 a_20034_10162# a_2475_10186# a_19942_10162# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X3822 a_21342_3174# col_n[18] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3823 VDD rowon_n[1] a_11910_3134# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3824 a_8290_13214# rowon_n[11] a_7894_13174# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X3825 a_5886_11166# a_2275_11190# a_5978_11166# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3826 a_15926_11166# a_2275_11190# a_16018_11166# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3827 VSS row_n[8] a_5278_10202# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3828 a_20338_7190# col_n[17] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3829 VSS row_n[5] a_30378_7190# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3830 VSS row_n[1] a_31382_3174# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3831 a_24450_13536# col_n[21] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X3832 a_20946_10162# row_n[8] a_21438_10524# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3833 a_2475_8178# a_1957_8178# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.171 pd=1.77 as=0.124 ps=1.01 w=0.6 l=0.15
X3834 a_5978_8154# a_2475_8178# a_5886_8154# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X3835 a_35002_3134# a_2275_3158# a_35094_3134# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3836 a_11302_9198# col_n[8] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3837 a_27062_9158# a_2475_9182# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3838 a_16322_7190# rowon_n[5] a_15926_7150# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X3839 vcm a_2275_7174# a_24050_7150# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3840 a_22954_6146# row_n[4] a_23446_6508# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3841 a_17326_3174# rowon_n[1] a_16930_3134# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X3842 VDD rowon_n[10] a_13918_12170# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3843 a_33486_6508# col_n[30] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X3844 VDD rowon_n[2] a_27974_4138# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3845 VDD rowon_n[10] a_3878_12170# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3846 VDD rowon_n[5] a_5886_7150# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3847 a_8898_18194# a_2275_18218# a_8990_18194# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3848 a_18938_18194# a_2275_18218# a_19030_18194# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3849 VDD rowon_n[9] a_7894_11166# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3850 a_20946_1126# VDD a_21438_1488# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3851 a_26058_2130# a_2475_2154# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3852 a_13310_15222# col_n[10] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3853 a_31478_1488# col_n[28] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X3854 VDD rowon_n[0] a_3878_2130# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3855 a_12002_17190# a_2475_17214# a_11910_17190# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X3856 a_34090_17190# a_2475_17214# a_33998_17190# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X3857 a_3270_15222# col_n[0] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3858 VDD VSS a_16930_1126# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3859 a_26362_1166# col_n[23] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3860 a_10906_9158# row_n[7] a_11398_9520# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3861 a_11910_5142# row_n[3] a_12402_5504# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3862 a_4274_4178# col_n[1] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3863 VSS row_n[3] a_35398_5182# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3864 a_25358_5182# col_n[22] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3865 a_35002_17190# row_n[15] a_35494_17552# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3866 vcm a_2275_13198# a_35094_13174# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3867 a_3270_8194# col_n[0] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3868 a_9294_2170# rowon_n[0] a_8898_2130# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X3869 a_12402_17552# col_n[9] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X3870 a_19334_17230# rowon_n[15] a_18938_17190# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X3871 vcm a_2275_5166# a_29070_5142# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3872 a_20338_12210# rowon_n[10] a_19942_12170# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X3873 vcm a_2275_8178# a_6982_8154# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3874 a_12914_13174# row_n[11] a_13406_13536# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3875 a_24354_11206# rowon_n[9] a_23958_11166# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X3876 a_2874_13174# row_n[11] a_3366_13536# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3877 a_24962_3134# row_n[1] a_25454_3496# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3878 a_5978_11166# a_2475_11190# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3879 a_16018_11166# a_2475_11190# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3880 a_35494_3496# VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X3881 a_29070_13174# a_2475_13198# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3882 a_3878_4138# row_n[2] a_4370_4500# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3883 VDD rowon_n[13] a_18938_15182# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3884 VDD rowon_n[8] a_19942_10162# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3885 a_15926_7150# row_n[5] a_16418_7512# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3886 a_14010_4138# a_2475_4162# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3887 a_9994_12170# a_2475_12194# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3888 a_8290_6186# col_n[5] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3889 vcm a_2275_18218# a_9994_18194# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3890 a_9902_6146# a_2275_6170# a_9994_6146# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3891 a_13918_2130# row_n[0] a_14410_2492# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3892 VSS row_n[14] a_22346_16226# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3893 VSS row_n[13] a_35398_15222# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3894 a_32386_12210# col_n[29] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3895 a_31382_9198# rowon_n[7] a_30986_9158# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X3896 a_19334_2170# col_n[16] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3897 vcm a_2275_3158# a_33086_3134# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3898 a_12306_15222# rowon_n[13] a_11910_15182# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X3899 a_25054_9158# a_2475_9182# a_24962_9158# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X3900 a_30378_2170# rowon_n[0] a_29982_2130# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X3901 VSS row_n[0] a_20338_2170# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3902 VDD VDD a_20946_18194# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3903 VDD rowon_n[15] a_33998_17190# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3904 a_6282_14218# rowon_n[12] a_5886_14178# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X3905 a_16322_14218# rowon_n[12] a_15926_14178# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X3906 a_31478_14540# col_n[28] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X3907 vcm a_2275_12194# a_27062_12170# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3908 VSS row_n[9] a_3270_11206# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3909 VSS row_n[9] a_13310_11206# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3910 a_31078_10162# a_2475_10186# a_30986_10162# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X3911 VSS row_n[6] a_10298_8194# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3912 a_34090_2130# a_2475_2154# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3913 a_2874_1126# a_2275_1150# a_2966_1126# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3914 VSS row_n[2] a_11302_4178# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3915 a_35494_13536# VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X3916 a_31990_10162# row_n[8] a_32482_10524# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3917 a_14922_4138# a_2275_4162# a_15014_4138# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3918 a_22442_5504# col_n[19] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X3919 a_7894_13174# a_2275_13198# a_7986_13174# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3920 a_17934_13174# a_2275_13198# a_18026_13174# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3921 VDD rowon_n[7] a_30986_9158# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3922 VDD rowon_n[3] a_31990_5142# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3923 VDD rowon_n[11] a_11910_13174# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3924 a_11302_16226# col_n[8] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3925 a_11398_4500# col_n[8] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X3926 a_32082_18194# a_2475_18218# a_31990_18194# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X3927 VSS row_n[1] a_3270_3174# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3928 a_32994_18194# VDD a_33486_18556# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3929 vcm a_2275_14202# a_33086_14178# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3930 a_18330_12210# rowon_n[10] a_17934_12170# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X3931 VSS row_n[4] a_15318_6186# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3932 a_10394_18556# col_n[7] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X3933 vcm a_2275_15206# a_19030_15182# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3934 a_5374_6508# col_n[2] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X3935 a_5978_6146# a_2475_6170# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3936 a_12002_4138# a_2475_4162# a_11910_4138# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X3937 vcm a_2275_15206# a_8990_15182# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3938 a_35398_11206# rowon_n[9] a_35002_11166# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X3939 a_18026_9158# a_2475_9182# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3940 VDD rowon_n[0] a_33998_2130# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3941 a_3366_1488# col_n[0] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X3942 VDD VSS sky130_fd_pr__cap_mim_m3_1 l=17.2 w=17.2
X3943 a_24450_2492# col_n[21] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X3944 a_23958_5142# a_2275_5166# a_24050_5142# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3945 a_23046_15182# a_2475_15206# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3946 VDD rowon_n[8] a_17934_10162# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3947 VSS row_n[0] a_29374_2170# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3948 a_34394_4178# col_n[31] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3949 a_27062_14178# a_2475_14202# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3950 a_33390_8194# col_n[30] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3951 VSS row_n[3] a_7286_5182# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3952 VSS VDD a_8290_1166# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3953 a_18026_13174# a_2475_13198# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3954 a_7986_13174# a_2475_13198# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3955 a_3970_3134# a_2475_3158# a_3878_3134# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X3956 a_21342_4178# rowon_n[2] a_20946_4138# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X3957 a_35002_11166# a_2275_11190# a_35094_11166# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3958 VSS row_n[8] a_34394_10202# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3959 a_9390_8516# col_n[6] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X3960 a_11302_10202# rowon_n[8] a_10906_10162# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X3961 a_9994_8154# a_2475_8178# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3962 a_32082_2130# a_2475_2154# a_31990_2130# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X3963 a_29374_18234# col_n[26] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3964 VSS row_n[14] a_33390_16226# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3965 a_27974_7150# a_2275_7174# a_28066_7150# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3966 a_28978_3134# a_2275_3158# a_29070_3134# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3967 a_10298_16226# rowon_n[14] a_9902_16186# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X3968 a_29470_14540# col_n[26] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X3969 VDD rowon_n[10] a_32994_12170# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3970 a_29070_10162# a_2475_10186# a_28978_10162# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X3971 a_6890_6146# a_2275_6170# a_6982_6146# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3972 a_7382_3496# col_n[4] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X3973 a_33998_4138# row_n[2] a_34490_4500# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3974 vcm a_2275_4162# a_13006_4138# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3975 a_18938_9158# a_2275_9182# a_19030_9158# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3976 a_28066_16186# a_2475_16210# a_27974_16186# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X3977 a_20034_9158# a_2475_9182# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3978 a_10298_3174# rowon_n[1] a_9902_3134# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X3979 VDD VDD a_31990_18194# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3980 VDD rowon_n[2] a_20946_4138# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3981 a_28978_16186# row_n[14] a_29470_16548# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3982 a_11910_15182# a_2275_15206# a_12002_15182# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3983 a_8990_1126# a_2475_1150# a_8898_1126# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X3984 VDD VSS VSS sky130_fd_pr__cap_var_lvt w=16.4 l=16
X3985 a_15926_14178# a_2275_14202# a_16018_14178# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3986 VDD rowon_n[4] a_11910_6146# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3987 a_5886_14178# a_2275_14202# a_5978_14178# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3988 a_3270_9198# rowon_n[7] a_2874_9158# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X3989 a_19030_6146# a_2475_6170# a_18938_6146# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X3990 a_10298_11206# col_n[7] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3991 vcm a_2275_3158# a_4974_3134# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3992 VDD VSS a_9902_1126# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X3993 a_16018_9158# a_2475_9182# a_15926_9158# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X3994 a_14314_5182# rowon_n[3] a_13918_5142# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X3995 a_15318_1166# VSS a_14922_1126# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X3996 a_32994_1126# a_2275_1150# a_33086_1126# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X3997 vcm a_2275_5166# a_22042_5142# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3998 vcm a_2275_10186# a_18026_10162# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3999 a_19942_8154# row_n[6] a_20434_8516# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4000 a_7894_14178# row_n[12] a_8386_14540# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4001 a_17934_14178# row_n[12] a_18426_14540# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4002 a_29374_12210# rowon_n[10] a_28978_12170# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X4003 vcm a_2275_10186# a_7986_10162# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4004 a_26970_10162# a_2275_10186# a_27062_10162# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4005 VDD rowon_n[7] a_2874_9158# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4006 a_30474_8516# col_n[27] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X4007 VDD rowon_n[3] a_3878_5142# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4008 VDD rowon_n[6] a_15926_8154# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4009 vcm a_2275_16210# a_6982_16186# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4010 vcm a_2275_16210# a_17022_16186# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4011 a_23350_3174# col_n[20] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4012 VDD rowon_n[1] a_13918_3134# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4013 a_21038_16186# a_2475_16210# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4014 VDD rowon_n[8] a_28978_10162# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4015 a_25358_9198# rowon_n[7] a_24962_9158# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X4016 a_7986_8154# a_2475_8178# a_7894_8154# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X4017 VSS row_n[5] a_32386_7190# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4018 VSS row_n[1] a_33390_3174# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4019 a_13310_9198# col_n[10] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4020 vcm a_2275_3158# a_27062_3134# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4021 VSS a_2161_17214# a_2275_17214# VSS sky130_fd_pr__nfet_01v8 ad=0.124 pd=1.01 as=0.171 ps=1.77 w=0.6 l=0.15
X4022 VSS row_n[15] a_27366_17230# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4023 a_31382_15222# rowon_n[13] a_30986_15182# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X4024 a_29070_9158# a_2475_9182# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4025 vcm a_2275_7174# a_26058_7150# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4026 a_24962_6146# row_n[4] a_25454_6508# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4027 a_5978_14178# a_2475_14202# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4028 a_16018_14178# a_2475_14202# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4029 VDD rowon_n[5] a_7894_7150# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4030 a_35494_6508# VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X4031 a_28370_13214# col_n[25] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4032 VSS row_n[9] a_32386_11206# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4033 vcm a_2275_9182# a_17022_9158# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4034 a_12306_2170# col_n[9] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4035 a_19942_15182# a_2275_15206# a_20034_15182# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4036 a_22954_1126# VDD a_23446_1488# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4037 a_33486_1488# col_n[30] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X4038 a_28066_2130# a_2475_2154# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4039 a_14010_17190# a_2475_17214# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4040 VSS row_n[10] a_18330_12210# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4041 a_23046_12170# a_2475_12194# a_22954_12170# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X4042 a_31990_8154# a_2275_8178# a_32082_8154# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4043 VDD rowon_n[0] a_5886_2130# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4044 a_3970_17190# a_2475_17214# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4045 VSS row_n[10] a_8290_12210# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4046 VDD rowon_n[7] a_24962_9158# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4047 a_28370_1166# col_n[25] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4048 a_27462_15544# col_n[24] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X4049 VDD rowon_n[11] a_30986_13174# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4050 a_23958_12170# row_n[10] a_24450_12532# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4051 a_27062_11166# a_2475_11190# a_26970_11166# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X4052 a_12914_9158# row_n[7] a_13406_9520# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4053 a_5278_8194# col_n[2] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4054 a_13918_5142# row_n[3] a_14410_5504# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4055 a_6282_4178# col_n[3] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4056 a_7986_10162# a_2475_10186# a_7894_10162# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X4057 a_18026_10162# a_2475_10186# a_17934_10162# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X4058 VDD rowon_n[12] a_16930_14178# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4059 a_27974_11166# row_n[9] a_28466_11528# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4060 VDD rowon_n[12] a_6890_14178# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4061 vcm a_2275_8178# a_8990_8154# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4062 a_30378_16226# col_n[27] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4063 a_8386_10524# col_n[5] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X4064 a_18426_10524# col_n[15] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X4065 vcm a_2275_1150# a_31078_1126# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4066 VDD a_2161_18218# a_2275_18218# VDD sky130_fd_pr__pfet_01v8 ad=0.249 pd=1.62 as=0.342 ps=2.97 w=1.2 l=0.15
X4067 vcm a_2275_17214# a_21038_17190# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4068 vcm a_2275_5166# a_30074_5142# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4069 a_6282_17230# col_n[3] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4070 a_16322_17230# col_n[13] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4071 a_3970_1126# a_2475_1150# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4072 vcm a_2275_16210# a_25054_16186# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4073 a_5886_4138# row_n[2] a_6378_4500# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4074 a_17934_7150# row_n[5] a_18426_7512# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4075 ctop sw_n analog_in VDD sky130_fd_pr__pfet_01v8 ad=0.275 pd=2.19 as=0.275 ps=2.19 w=1.9 l=0.22
X4076 a_8990_18194# a_2475_18218# a_8898_18194# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X4077 vcm a_2275_12194# a_12002_12170# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4078 a_15926_2130# row_n[0] a_16418_2492# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4079 a_15926_15182# row_n[13] a_16418_15544# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4080 a_27366_13214# rowon_n[11] a_26970_13174# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X4081 vcm a_2275_11190# a_16018_11166# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4082 a_9390_18556# col_n[6] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X4083 a_5886_15182# row_n[13] a_6378_15544# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4084 vcm a_2275_11190# a_5978_11166# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4085 a_10998_9158# a_2475_9182# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4086 a_33390_9198# rowon_n[7] a_32994_9158# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X4087 a_27366_8194# col_n[24] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4088 a_27062_9158# a_2475_9182# a_26970_9158# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X4089 vcm a_2275_3158# a_35094_3134# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4090 VDD VSS VSS sky130_fd_pr__cap_var_lvt w=16.4 l=16
X4091 a_19030_16186# a_2475_16210# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4092 VSS row_n[0] a_22346_2170# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4093 a_28978_12170# a_2275_12194# a_29070_12170# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4094 a_32386_2170# rowon_n[0] a_31990_2130# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X4095 a_4882_1126# a_2275_1150# a_4974_1126# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4096 a_19030_4138# a_2475_4162# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4097 VSS row_n[2] a_13310_4178# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4098 VDD rowon_n[9] a_26970_11166# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4099 VSS row_n[6] a_12306_8194# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4100 a_26058_2130# a_2475_2154# a_25966_2130# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X4101 a_24450_5504# col_n[21] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X4102 VDD rowon_n[7] a_32994_9158# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4103 VDD rowon_n[3] a_33998_5142# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4104 VSS VDD a_25358_18234# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4105 a_22346_15222# col_n[19] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4106 a_2966_8154# a_2475_8178# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4107 a_26362_14218# col_n[23] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4108 a_2161_10186# sample VDD VDD sky130_fd_pr__pfet_01v8 ad=0.342 pd=2.97 as=0.342 ps=2.97 w=1.2 l=0.15
X4109 a_20946_7150# a_2275_7174# a_21038_7150# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4110 VSS a_2161_5166# a_2275_5166# VSS sky130_fd_pr__nfet_01v8 ad=0.124 pd=1.01 as=0.171 ps=1.77 w=0.6 l=0.15
X4111 a_21950_3134# a_2275_3158# a_22042_3134# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4112 a_15318_17230# rowon_n[15] a_14922_17190# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X4113 a_31078_7150# a_2475_7174# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4114 a_34090_18194# a_2475_18218# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4115 a_5278_17230# rowon_n[15] a_4882_17190# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X4116 a_30986_15182# a_2275_15206# a_31078_15182# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4117 a_11910_9158# a_2275_9182# a_12002_9158# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4118 a_12002_18194# a_2475_18218# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4119 a_21438_17552# col_n[18] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X4120 a_9294_16226# rowon_n[14] a_8898_16186# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X4121 VSS row_n[11] a_6282_13214# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4122 VSS row_n[11] a_16322_13214# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4123 a_21038_13174# a_2475_13198# a_20946_13174# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X4124 a_19334_6186# rowon_n[4] a_18938_6146# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X4125 a_31382_6186# col_n[28] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4126 VSS row_n[1] a_5278_3174# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4127 a_13406_4500# col_n[10] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X4128 a_25454_16548# col_n[22] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X4129 a_35002_14178# a_2275_14202# a_35094_14178# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4130 a_21950_13174# row_n[11] a_22442_13536# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4131 VSS row_n[5] a_4274_7190# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4132 a_16018_11166# a_2475_11190# a_15926_11166# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X4133 VSS row_n[4] a_17326_6186# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4134 a_5978_11166# a_2475_11190# a_5886_11166# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X4135 a_7382_6508# col_n[4] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X4136 VDD rowon_n[13] a_4882_15182# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4137 VDD rowon_n[13] a_14922_15182# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4138 a_7986_6146# a_2475_6170# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4139 a_14010_4138# a_2475_4162# a_13918_4138# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X4140 a_5278_12210# col_n[2] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4141 a_15318_12210# col_n[12] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4142 vcm a_2275_12194# a_20034_12170# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4143 a_16418_11528# col_n[13] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X4144 a_26970_1126# a_2275_1150# a_27062_1126# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4145 a_25966_5142# a_2275_5166# a_26058_5142# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4146 a_6378_11528# col_n[3] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X4147 a_3878_8154# a_2275_8178# a_3970_8154# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4148 vcm a_2275_6170# a_9994_6146# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4149 a_5374_1488# col_n[2] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X4150 a_14314_18234# col_n[11] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4151 a_4274_18234# col_n[1] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4152 vcm a_2275_17214# a_32082_17190# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4153 a_35398_8194# VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4154 a_4370_14540# col_n[1] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X4155 a_14410_14540# col_n[11] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X4156 VSS row_n[3] a_9294_5182# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4157 a_14922_10162# row_n[8] a_15414_10524# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4158 a_23046_10162# a_2475_10186# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4159 a_4882_10162# row_n[8] a_5374_10524# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4160 a_23350_4178# rowon_n[2] a_22954_4138# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X4161 a_2161_8178# sample VSS VSS sky130_fd_pr__nfet_01v8 ad=0.171 pd=1.77 as=0.171 ps=1.77 w=0.6 l=0.15
X4162 VSS row_n[5] a_26362_7190# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4163 a_3878_16186# row_n[14] a_4370_16548# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4164 a_13918_16186# row_n[14] a_14410_16548# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4165 a_25358_14218# rowon_n[12] a_24962_14178# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X4166 a_1957_13198# VSS sample VDD sky130_fd_pr__pfet_01v8 ad=0.342 pd=2.97 as=0.342 ps=2.97 w=1.2 l=0.15
X4167 a_34090_2130# a_2475_2154# a_33998_2130# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X4168 vcm a_2275_1150# a_2966_1126# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4169 a_8898_6146# a_2275_6170# a_8990_6146# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4170 a_9390_3496# col_n[6] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X4171 vcm a_2275_4162# a_15014_4138# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4172 a_26058_17190# a_2475_17214# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4173 a_23350_17230# rowon_n[15] a_22954_17190# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X4174 a_26970_13174# a_2275_13198# a_27062_13174# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4175 a_29982_3134# a_2275_3158# a_30074_3134# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4176 a_22042_9158# a_2475_9182# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4177 a_11302_7190# rowon_n[5] a_10906_7150# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X4178 a_12306_3174# rowon_n[1] a_11910_3134# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X4179 VSS row_n[11] a_24354_13214# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4180 a_21342_10202# col_n[18] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4181 VDD rowon_n[2] a_22954_4138# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4182 a_14314_12210# rowon_n[10] a_13918_12170# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X4183 VDD rowon_n[4] a_13918_6146# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4184 a_21038_2130# a_2475_2154# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4185 a_4274_12210# rowon_n[10] a_3878_12170# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X4186 a_11910_10162# a_2275_10186# a_12002_10162# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4187 a_19430_17552# col_n[16] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X4188 VDD VSS VSS sky130_fd_pr__cap_var_lvt w=16.4 l=16
X4189 VDD rowon_n[13] a_22954_15182# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4190 a_19030_13174# a_2475_13198# a_18938_13174# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X4191 a_20434_12532# col_n[17] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X4192 VDD VSS a_11910_1126# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4193 a_21342_1166# col_n[18] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4194 a_8290_11206# rowon_n[9] a_7894_11166# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X4195 VSS VDD a_31382_1166# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4196 VSS row_n[3] a_30378_5182# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4197 a_20338_5182# col_n[17] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4198 a_24450_11528# col_n[21] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X4199 a_5978_6146# a_2475_6170# a_5886_6146# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X4200 a_35002_1126# a_2275_1150# a_35094_1126# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4201 a_4274_2170# rowon_n[0] a_3878_2130# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X4202 a_18026_9158# a_2475_9182# a_17934_9158# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X4203 a_16322_5182# rowon_n[3] a_15926_5142# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X4204 a_17326_1166# VSS a_16930_1126# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X4205 vcm a_2275_5166# a_24050_5142# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4206 a_35398_17230# VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4207 VDD rowon_n[8] a_13918_10162# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4208 a_32482_8516# col_n[29] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X4209 VDD rowon_n[8] a_3878_10162# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4210 VDD rowon_n[3] a_5886_5142# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4211 VSS row_n[15] a_12306_17230# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4212 a_8898_16186# a_2275_16210# a_8990_16186# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4213 a_18938_16186# a_2275_16210# a_19030_16186# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4214 a_19942_3134# row_n[1] a_20434_3496# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4215 a_13310_13214# col_n[10] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4216 a_30474_3496# col_n[27] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X4217 a_12002_15182# a_2475_15206# a_11910_15182# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X4218 a_34090_15182# a_2475_15206# a_33998_15182# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X4219 a_3270_13214# col_n[0] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4220 vcm a_2275_12194# a_31078_12170# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4221 a_25358_3174# col_n[22] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4222 a_10906_7150# row_n[5] a_11398_7512# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4223 VSS row_n[1] a_35398_3174# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4224 VDD rowon_n[1] a_15926_3134# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4225 a_35002_15182# row_n[13] a_35494_15544# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4226 vcm a_2275_11190# a_35094_11166# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4227 a_27366_9198# rowon_n[7] a_26970_9158# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X4228 a_9994_8154# a_2475_8178# a_9902_8154# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X4229 VSS row_n[5] a_34394_7190# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4230 a_3270_6186# col_n[0] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4231 a_12402_15544# col_n[9] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X4232 a_19334_15222# rowon_n[13] a_18938_15182# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X4233 a_20338_10202# rowon_n[8] a_19942_10162# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X4234 a_15318_9198# col_n[12] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4235 vcm a_2275_7174# a_28066_7150# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4236 vcm a_2275_3158# a_29070_3134# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4237 a_21038_11166# a_2475_11190# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4238 vcm a_2275_6170# a_6982_6146# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4239 a_12914_11166# row_n[9] a_13406_11528# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4240 vcm a_2275_9182# a_19030_9158# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4241 VSS a_2161_12194# a_2275_12194# VSS sky130_fd_pr__nfet_01v8 ad=0.124 pd=1.01 as=0.171 ps=1.77 w=0.6 l=0.15
X4242 a_2874_11166# row_n[9] a_3366_11528# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4243 a_24962_1126# VDD a_25454_1488# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4244 a_14314_2170# col_n[11] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4245 a_25054_12170# a_2475_12194# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4246 a_20034_9158# a_2475_9182# a_19942_9158# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X4247 a_33998_8154# a_2275_8178# a_34090_8154# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4248 a_35494_1488# VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X4249 VDD rowon_n[0] a_7894_2130# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4250 VDD rowon_n[11] a_18938_13174# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4251 a_19942_10162# a_2275_10186# a_20034_10162# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4252 a_14922_9158# row_n[7] a_15414_9520# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4253 VDD rowon_n[7] a_26970_9158# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4254 a_15926_5142# row_n[3] a_16418_5504# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4255 a_8290_4178# col_n[5] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4256 a_21342_18234# VDD a_20946_18194# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X4257 vcm a_2275_16210# a_9994_16186# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4258 a_9902_4138# a_2275_4162# a_9994_4138# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4259 a_34394_17230# rowon_n[15] a_33998_17190# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X4260 VSS row_n[12] a_22346_14218# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4261 VSS row_n[11] a_35398_13214# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4262 a_32386_10202# col_n[29] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4263 a_22954_17190# a_2275_17214# a_23046_17190# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4264 vcm a_2275_1150# a_33086_1126# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4265 a_12306_13214# rowon_n[11] a_11910_13174# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X4266 a_7894_4138# row_n[2] a_8386_4500# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4267 VDD rowon_n[14] a_20946_16186# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4268 VDD rowon_n[13] a_33998_15182# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4269 a_26970_14178# row_n[12] a_27462_14540# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4270 a_31478_12532# col_n[28] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X4271 vcm a_2275_10186# a_27062_10162# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4272 a_13918_12170# a_2275_12194# a_14010_12170# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4273 VSS row_n[4] a_10298_6186# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4274 a_3878_12170# a_2275_12194# a_3970_12170# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4275 a_35494_11528# VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X4276 VDD rowon_n[5] a_30986_7150# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4277 a_17934_2130# row_n[0] a_18426_2492# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4278 a_33390_18234# col_n[30] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4279 VDD rowon_n[9] a_11910_11166# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4280 a_29374_8194# col_n[26] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4281 VSS VDD a_10298_18234# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4282 a_13006_9158# a_2475_9182# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4283 a_29070_9158# a_2475_9182# a_28978_9158# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X4284 vcm a_2275_18218# a_28066_18194# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4285 a_32082_16186# a_2475_16210# a_31990_16186# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X4286 a_11302_14218# col_n[8] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4287 VSS row_n[0] a_24354_2170# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4288 a_18330_10202# rowon_n[8] a_17934_10162# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X4289 a_34394_2170# rowon_n[0] a_33998_2130# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X4290 VSS VDD a_3270_1166# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4291 a_32994_16186# row_n[14] a_33486_16548# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4292 a_19030_11166# a_2475_11190# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4293 VSS row_n[6] a_14314_8194# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4294 a_28066_2130# a_2475_2154# a_27974_2130# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X4295 VSS row_n[2] a_15318_4178# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4296 vcm a_2275_8178# a_32082_8154# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4297 a_18938_17190# row_n[15] a_19430_17552# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4298 a_10394_16548# col_n[7] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X4299 vcm a_2275_13198# a_19030_13174# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4300 a_4370_8516# col_n[1] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X4301 a_5978_4138# a_2475_4162# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4302 a_8898_17190# row_n[15] a_9390_17552# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4303 vcm a_2275_13198# a_8990_13174# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4304 a_4974_8154# a_2475_8178# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4305 a_23958_3134# a_2275_3158# a_24050_3134# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4306 VDD a_2161_9182# a_2275_9182# VDD sky130_fd_pr__pfet_01v8 ad=0.249 pd=1.62 as=0.342 ps=2.97 w=1.2 l=0.15
X4307 a_22954_7150# a_2275_7174# a_23046_7150# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4308 a_23046_13174# a_2475_13198# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4309 a_33086_7150# a_2475_7174# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4310 a_13918_9158# a_2275_9182# a_14010_9158# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4311 a_33390_6186# col_n[30] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4312 VSS row_n[1] a_7286_3174# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4313 a_15414_4500# col_n[12] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X4314 a_33390_12210# rowon_n[10] a_32994_12170# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X4315 a_30986_10162# a_2275_10186# a_31078_10162# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4316 a_3970_1126# a_2475_1150# a_3878_1126# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X4317 a_32386_18234# VDD a_31990_18194# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X4318 a_9390_6508# col_n[6] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X4319 a_9994_6146# a_2475_6170# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4320 a_28978_1126# a_2275_1150# a_29070_1126# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4321 a_29374_16226# col_n[26] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4322 VSS row_n[12] a_33390_14218# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4323 a_27974_5142# a_2275_5166# a_28066_5142# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4324 a_20946_18194# a_2275_18218# a_21038_18194# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4325 a_33998_17190# a_2275_17214# a_34090_17190# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4326 a_10298_14218# rowon_n[12] a_9902_14178# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X4327 a_29470_12532# col_n[26] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X4328 VDD rowon_n[8] a_32994_10162# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4329 a_5886_8154# a_2275_8178# a_5978_8154# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4330 a_7382_1488# col_n[4] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X4331 a_6890_4138# a_2275_4162# a_6982_4138# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4332 a_26458_8516# col_n[23] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X4333 a_28066_14178# a_2475_14202# a_27974_14178# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X4334 a_10998_9158# a_2475_9182# a_10906_9158# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X4335 a_10298_1166# VSS a_9902_1126# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X4336 a_28466_18556# col_n[25] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X4337 VDD rowon_n[14] a_31990_16186# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4338 a_11910_13174# a_2275_13198# a_12002_13174# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4339 VDD rowon_n[6] a_10906_8154# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4340 VSS row_n[5] a_28370_7190# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4341 a_19030_4138# a_2475_4162# a_18938_4138# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X4342 a_1957_7174# VSS sample VDD sky130_fd_pr__pfet_01v8 ad=0.342 pd=2.97 as=0.342 ps=2.97 w=1.2 l=0.15
X4343 vcm a_2275_1150# a_4974_1126# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4344 a_20338_9198# rowon_n[7] a_19942_9158# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X4345 a_2966_8154# a_2475_8178# a_2874_8154# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X4346 a_13310_7190# rowon_n[5] a_12914_7150# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X4347 vcm a_2275_3158# a_22042_3134# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4348 a_14314_3174# rowon_n[1] a_13918_3134# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X4349 a_24050_9158# a_2475_9182# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4350 vcm a_2275_7174# a_21038_7150# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4351 a_31078_7150# a_2475_7174# a_30986_7150# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X4352 a_19942_6146# row_n[4] a_20434_6508# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4353 a_7894_12170# row_n[10] a_8386_12532# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4354 a_17934_12170# row_n[10] a_18426_12532# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4355 a_29374_10202# rowon_n[8] a_28978_10162# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X4356 VDD rowon_n[5] a_2874_7150# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4357 a_30474_6508# col_n[27] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X4358 vcm a_2275_9182# a_12002_9158# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4359 VDD rowon_n[4] a_15926_6146# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4360 a_16930_18194# VDD a_17422_18556# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4361 vcm a_2275_14202# a_6982_14178# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4362 vcm a_2275_14202# a_17022_14178# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4363 a_23046_2130# a_2475_2154# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4364 a_6890_18194# VDD a_7382_18556# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4365 VDD rowon_n[7] a_19942_9158# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4366 VDD VSS a_13918_1126# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4367 a_23350_1166# col_n[20] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4368 vcm a_2275_17214# a_15014_17190# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4369 a_21038_14178# a_2475_14202# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4370 a_7986_6146# a_2475_6170# a_7894_6146# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X4371 VSS VDD a_33390_1166# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4372 a_6282_2170# rowon_n[0] a_5886_2130# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X4373 VSS row_n[3] a_32386_5182# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4374 vcm a_2275_17214# a_4974_17190# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4375 vcm a_2275_1150# a_27062_1126# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4376 VSS a_2161_15206# a_2275_15206# VSS sky130_fd_pr__nfet_01v8 ad=0.124 pd=1.01 as=0.171 ps=1.77 w=0.6 l=0.15
X4377 VSS row_n[13] a_27366_15222# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4378 a_31382_13214# rowon_n[11] a_30986_13174# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X4379 a_24354_12210# col_n[21] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4380 vcm a_2275_5166# a_26058_5142# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4381 vcm a_2275_8178# a_3970_8154# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4382 a_34490_8516# col_n[31] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X4383 VDD rowon_n[3] a_7894_5142# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4384 a_28370_11206# col_n[25] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4385 a_19942_13174# a_2275_13198# a_20034_13174# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4386 VDD rowon_n[15] a_25966_17190# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4387 a_14010_15182# a_2475_15206# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4388 a_23446_14540# col_n[20] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X4389 a_32994_12170# a_2275_12194# a_33086_12170# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4390 VSS row_n[8] a_18330_10202# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4391 a_23046_10162# a_2475_10186# a_22954_10162# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X4392 a_31990_6146# a_2275_6170# a_32082_6146# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4393 a_32482_3496# col_n[29] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X4394 a_3970_15182# a_2475_15206# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4395 a_8898_11166# a_2275_11190# a_8990_11166# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4396 a_18938_11166# a_2275_11190# a_19030_11166# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4397 VSS row_n[8] a_8290_10202# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4398 VDD rowon_n[5] a_24962_7150# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4399 a_31990_18194# a_2275_18218# a_32082_18194# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4400 a_27462_13536# col_n[24] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X4401 VDD rowon_n[9] a_30986_11166# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4402 a_23958_10162# row_n[8] a_24450_10524# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4403 VSS row_n[7] a_19334_9198# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4404 a_12914_7150# row_n[5] a_13406_7512# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4405 a_5278_6186# col_n[2] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4406 a_29374_9198# rowon_n[7] a_28978_9158# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X4407 VDD rowon_n[10] a_16930_12170# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4408 a_10906_2130# row_n[0] a_11398_2492# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4409 VDD rowon_n[10] a_6890_12170# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4410 vcm a_2275_6170# a_8990_6146# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4411 a_30378_14218# col_n[27] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4412 a_22346_8194# col_n[19] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4413 a_24050_18194# a_2475_18218# a_23958_18194# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X4414 VDD a_2161_16210# a_2275_16210# VDD sky130_fd_pr__pfet_01v8 ad=0.249 pd=1.62 as=0.342 ps=2.97 w=1.2 l=0.15
X4415 a_16322_15222# col_n[13] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4416 vcm a_2275_15206# a_21038_15182# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4417 a_22042_9158# a_2475_9182# a_21950_9158# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X4418 a_16322_2170# col_n[13] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4419 vcm a_2275_3158# a_30074_3134# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4420 VSS VDD a_9294_18234# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4421 a_15014_17190# a_2475_17214# a_14922_17190# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X4422 a_6282_15222# col_n[3] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4423 a_19430_9520# col_n[16] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X4424 a_24962_18194# VDD a_25454_18556# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4425 a_4974_17190# a_2475_17214# a_4882_17190# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X4426 vcm a_2275_14202# a_25054_14178# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4427 VDD rowon_n[7] a_28978_9158# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4428 a_17934_5142# row_n[3] a_18426_5504# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4429 a_15414_17552# col_n[12] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X4430 a_8990_16186# a_2475_16210# a_8898_16186# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X4431 vcm a_2275_10186# a_12002_10162# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4432 a_21038_2130# a_2475_2154# a_20946_2130# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X4433 a_5374_17552# col_n[2] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X4434 a_11910_14178# row_n[12] a_12402_14540# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4435 a_15926_13174# row_n[11] a_16418_13536# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4436 a_27366_11206# rowon_n[9] a_26970_11166# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X4437 a_9390_16548# col_n[6] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X4438 a_5886_13174# row_n[11] a_6378_13536# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4439 a_27366_6186# col_n[24] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4440 vcm a_2275_1150# a_35094_1126# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4441 a_19030_14178# a_2475_14202# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4442 vcm a_2275_18218# a_2966_18194# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4443 vcm a_2275_18218# a_13006_18194# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4444 VSS row_n[15] a_21342_17230# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4445 VSS row_n[4] a_12306_6186# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4446 VDD rowon_n[5] a_32994_7150# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4447 VSS row_n[14] a_25358_16226# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4448 a_22346_13214# col_n[19] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4449 a_2966_6146# a_2475_6170# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4450 a_15014_9158# a_2475_9182# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4451 a_21950_1126# a_2275_1150# a_22042_1126# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4452 VSS a_2161_3158# a_2275_3158# VSS sky130_fd_pr__nfet_01v8 ad=0.124 pd=1.01 as=0.171 ps=1.77 w=0.6 l=0.15
X4453 a_20946_5142# a_2275_5166# a_21038_5142# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4454 a_30074_17190# a_2475_17214# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4455 a_15318_15222# rowon_n[13] a_14922_15182# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X4456 VDD rowon_n[0] a_30986_2130# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4457 a_31078_5142# a_2475_5166# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4458 a_34090_16186# a_2475_16210# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4459 a_5278_15222# rowon_n[13] a_4882_15182# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X4460 a_30986_13174# a_2275_13198# a_31078_13174# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4461 VDD VDD a_23958_18194# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4462 a_12002_16186# a_2475_16210# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4463 a_21438_15544# col_n[18] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X4464 a_9294_14218# rowon_n[12] a_8898_14178# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X4465 VSS row_n[9] a_6282_11206# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4466 VSS row_n[9] a_16322_11206# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4467 a_21038_11166# a_2475_11190# a_20946_11166# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X4468 a_18330_8194# rowon_n[6] a_17934_8154# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X4469 a_30378_8194# col_n[27] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4470 VSS VDD a_5278_1166# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4471 a_31382_4178# col_n[28] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4472 a_19334_4178# rowon_n[2] a_18938_4138# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X4473 a_21950_11166# row_n[9] a_22442_11528# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4474 VSS row_n[3] a_4274_5182# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4475 VSS row_n[2] a_17326_4178# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4476 vcm a_2275_8178# a_34090_8154# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4477 VDD rowon_n[11] a_4882_13174# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4478 VDD rowon_n[11] a_14922_13174# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4479 a_6982_8154# a_2475_8178# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4480 VSS row_n[5] a_21342_7190# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4481 a_7986_4138# a_2475_4162# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4482 a_19942_14178# row_n[12] a_20434_14540# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4483 a_5278_10202# col_n[2] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4484 a_15318_10202# col_n[12] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4485 vcm a_2275_10186# a_20034_10162# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4486 a_24962_7150# a_2275_7174# a_25054_7150# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4487 a_25966_3134# a_2275_3158# a_26058_3134# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4488 a_3970_12170# a_2475_12194# a_3878_12170# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X4489 a_14010_12170# a_2475_12194# a_13918_12170# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X4490 a_35094_7150# a_2475_7174# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4491 a_3878_6146# a_2275_6170# a_3970_6146# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4492 a_4370_3496# col_n[1] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X4493 VDD rowon_n[2] a_18938_4138# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4494 vcm a_2275_4162# a_9994_4138# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4495 a_14314_16226# col_n[11] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4496 a_15926_9158# a_2275_9182# a_16018_9158# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4497 a_30986_4138# row_n[2] a_31478_4500# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4498 a_13006_18194# a_2475_18218# a_12914_18194# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X4499 a_35094_18194# a_2475_18218# a_35002_18194# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X4500 a_4274_16226# col_n[1] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4501 vcm a_2275_15206# a_32082_15182# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4502 a_35398_6186# VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4503 VSS row_n[1] a_9294_3174# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4504 a_17422_4500# col_n[14] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X4505 a_2966_18194# a_2475_18218# a_2874_18194# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X4506 a_4370_12532# col_n[1] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X4507 a_14410_12532# col_n[11] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X4508 a_13406_18556# col_n[10] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X4509 a_3366_18556# col_n[0] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X4510 VSS row_n[3] a_26362_5182# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4511 a_1957_11190# VSS sample VDD sky130_fd_pr__pfet_01v8 ad=0.342 pd=2.97 as=0.342 ps=2.97 w=1.2 l=0.15
X4512 a_1957_1150# VDD sample VSS sky130_fd_pr__nfet_01v8 ad=0.171 pd=1.77 as=0.171 ps=1.77 w=0.6 l=0.15
X4513 a_26058_15182# a_2475_15206# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4514 a_7894_8154# a_2275_8178# a_7986_8154# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4515 a_9390_1488# col_n[6] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X4516 a_8898_4138# a_2275_4162# a_8990_4138# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4517 a_28466_8516# col_n[25] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X4518 VSS row_n[15] a_19334_17230# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4519 a_23350_15222# rowon_n[13] a_22954_15182# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X4520 VSS row_n[10] a_20338_12210# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4521 a_29982_1126# a_2275_1150# a_30074_1126# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4522 a_13006_9158# a_2475_9182# a_12914_9158# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X4523 a_11302_5182# rowon_n[3] a_10906_5142# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X4524 a_12306_1166# VSS a_11910_1126# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X4525 VSS row_n[9] a_24354_11206# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4526 a_26458_3496# col_n[23] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X4527 a_14314_10202# rowon_n[8] a_13918_10162# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X4528 VDD rowon_n[6] a_12914_8154# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4529 a_4274_10202# rowon_n[8] a_3878_10162# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X4530 a_19430_15544# col_n[16] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X4531 VDD rowon_n[11] a_22954_13174# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4532 a_19030_11166# a_2475_11190# a_18938_11166# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X4533 a_20434_10524# col_n[17] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X4534 a_20338_3174# col_n[17] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4535 VSS row_n[1] a_30378_3174# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4536 VDD rowon_n[1] a_10906_3134# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4537 VDD VSS VSS sky130_fd_pr__cap_var_lvt w=16.4 l=16
X4538 a_22346_9198# rowon_n[7] a_21950_9158# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X4539 a_4974_8154# a_2475_8178# a_4882_8154# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X4540 a_5978_4138# a_2475_4162# a_5886_4138# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X4541 VDD VDD a_35002_18194# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4542 a_10298_9198# col_n[7] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4543 vcm a_2275_7174# a_23046_7150# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4544 vcm a_2275_3158# a_24050_3134# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4545 a_16322_3174# rowon_n[1] a_15926_3134# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X4546 a_35398_15222# VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4547 a_33086_7150# a_2475_7174# a_32994_7150# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X4548 a_32482_6508# col_n[29] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X4549 vcm a_2275_9182# a_14010_9158# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4550 VSS row_n[13] a_12306_15222# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4551 a_8898_14178# a_2275_14202# a_8990_14178# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4552 a_18938_14178# a_2275_14202# a_19030_14178# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4553 a_19942_1126# en_bit_n[0] a_20434_1488# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4554 a_25054_2130# a_2475_2154# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4555 a_13310_11206# col_n[10] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4556 a_30474_1488# col_n[27] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X4557 a_34490_17552# col_n[31] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X4558 a_30986_14178# row_n[12] a_31478_14540# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4559 a_12002_13174# a_2475_13198# a_11910_13174# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X4560 a_34090_13174# a_2475_13198# a_33998_13174# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X4561 a_3270_11206# col_n[0] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4562 vcm a_2275_10186# a_31078_10162# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4563 VDD VSS a_15926_1126# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4564 a_25358_1166# col_n[22] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4565 VDD rowon_n[0] a_2874_2130# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4566 a_9902_9158# row_n[7] a_10394_9520# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4567 VDD rowon_n[7] a_21950_9158# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4568 a_10906_5142# row_n[3] a_11398_5504# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4569 VSS VDD a_35398_1166# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4570 VDD rowon_n[15] a_10906_17190# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4571 a_35002_13174# row_n[11] a_35494_13536# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4572 a_9994_6146# a_2475_6170# a_9902_6146# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X4573 a_8290_2170# rowon_n[0] a_7894_2130# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X4574 a_3270_4178# col_n[0] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4575 VSS row_n[3] a_34394_5182# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4576 a_12402_13536# col_n[9] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X4577 a_19334_13214# rowon_n[11] a_18938_13174# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X4578 vcm a_2275_1150# a_29070_1126# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4579 vcm a_2275_5166# a_28066_5142# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4580 vcm a_2275_8178# a_5978_8154# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4581 vcm a_2275_4162# a_6982_4138# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4582 a_2475_7174# a_1957_7174# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.342 pd=2.97 as=0.249 ps=1.62 w=1.2 l=0.15
X4583 VSS a_2161_10186# a_2275_10186# VSS sky130_fd_pr__nfet_01v8 ad=0.124 pd=1.01 as=0.171 ps=1.77 w=0.6 l=0.15
X4584 a_33998_6146# a_2275_6170# a_34090_6146# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4585 a_34490_3496# col_n[31] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X4586 a_2874_4138# row_n[2] a_3366_4500# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4587 VDD rowon_n[9] a_18938_11166# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4588 a_14922_7150# row_n[5] a_15414_7512# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4589 VDD rowon_n[5] a_26970_7150# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4590 a_2475_18218# a_1957_18218# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.171 pd=1.77 as=0.124 ps=1.01 w=0.6 l=0.15
X4591 a_14010_10162# a_2475_10186# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4592 a_9902_18194# VDD a_10394_18556# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4593 a_21342_16226# rowon_n[14] a_20946_16186# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X4594 a_34394_15222# rowon_n[13] a_33998_15182# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X4595 vcm a_2275_14202# a_9994_14178# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4596 VSS row_n[10] a_31382_12210# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4597 a_3970_10162# a_2475_10186# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4598 VDD rowon_n[0] a_24962_2130# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4599 a_12914_2130# row_n[0] a_13406_2492# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4600 VSS row_n[9] a_35398_11206# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4601 a_24354_8194# col_n[21] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4602 a_22954_15182# a_2275_15206# a_23046_15182# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4603 a_18330_2170# col_n[15] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4604 a_17022_17190# a_2475_17214# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4605 VDD rowon_n[12] a_29982_14178# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4606 a_26058_12170# a_2475_12194# a_25966_12170# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X4607 a_12306_11206# rowon_n[9] a_11910_11166# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X4608 a_24050_9158# a_2475_9182# a_23958_9158# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X4609 a_6982_17190# a_2475_17214# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4610 VDD rowon_n[11] a_33998_13174# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4611 a_26970_12170# row_n[10] a_27462_12532# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4612 a_31478_10524# col_n[28] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X4613 a_23046_2130# a_2475_2154# a_22954_2130# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X4614 VSS row_n[2] a_10298_4178# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4615 VDD rowon_n[3] a_30986_5142# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4616 a_33390_16226# col_n[30] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4617 a_29374_6186# col_n[26] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4618 VSS row_n[14] a_10298_16226# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4619 a_9294_17230# col_n[6] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4620 a_19334_17230# col_n[16] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4621 vcm a_2275_17214# a_24050_17190# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4622 a_7286_9198# col_n[4] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4623 vcm a_2275_16210# a_28066_16186# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4624 a_32082_14178# a_2475_14202# a_31990_14178# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X4625 a_10394_4500# col_n[7] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X4626 a_14922_18194# a_2275_18218# a_15014_18194# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4627 a_32482_18556# col_n[29] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X4628 a_4882_18194# a_2275_18218# a_4974_18194# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4629 VSS row_n[4] a_14314_6186# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4630 VDD VSS VSS sky130_fd_pr__cap_var_lvt w=16.4 l=16
X4631 vcm a_2275_6170# a_32082_6146# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4632 a_18938_15182# row_n[13] a_19430_15544# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4633 vcm a_2275_11190# a_19030_11166# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4634 a_4370_6508# col_n[1] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X4635 a_8898_15182# row_n[13] a_9390_15544# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4636 vcm a_2275_11190# a_8990_11166# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4637 a_6890_9158# row_n[7] a_7382_9520# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4638 a_4974_6146# a_2475_6170# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4639 a_23958_1126# a_2275_1150# a_24050_1126# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4640 a_17022_9158# a_2475_9182# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4641 a_33086_5142# a_2475_5166# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4642 a_22954_5142# a_2275_5166# a_23046_5142# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4643 VDD rowon_n[0] a_32994_2130# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4644 a_21438_8516# col_n[18] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X4645 VSS row_n[10] a_29374_12210# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4646 VSS VDD a_7286_1166# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4647 a_16018_2130# a_2475_2154# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4648 a_33390_4178# col_n[30] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4649 a_34090_11166# a_2475_11190# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4650 a_33390_10202# rowon_n[8] a_32994_10162# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X4651 a_12002_11166# a_2475_11190# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4652 VSS VDD a_28370_18234# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4653 a_32386_16226# rowon_n[14] a_31990_16186# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X4654 VDD rowon_n[12] a_27974_14178# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4655 a_8990_8154# a_2475_8178# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4656 VSS row_n[5] a_23350_7190# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4657 a_9994_4138# a_2475_4162# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4658 a_29374_14218# col_n[26] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4659 a_27974_3134# a_2275_3158# a_28066_3134# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4660 a_20946_16186# a_2275_16210# a_21038_16186# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4661 a_33998_15182# a_2275_15206# a_34090_15182# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4662 a_29470_10524# col_n[26] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X4663 a_5886_6146# a_2275_6170# a_5978_6146# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4664 a_32994_4138# row_n[2] a_33486_4500# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4665 a_4974_18194# a_2475_18218# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4666 a_15014_18194# a_2475_18218# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4667 a_17934_9158# a_2275_9182# a_18026_9158# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4668 a_26458_6508# col_n[23] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X4669 a_28466_16548# col_n[25] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X4670 a_16930_2130# a_2275_2154# a_17022_2130# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4671 VDD rowon_n[4] a_10906_6146# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4672 a_8290_12210# col_n[5] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4673 a_18330_12210# col_n[15] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4674 vcm a_2275_12194# a_23046_12170# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4675 VSS row_n[3] a_28370_5182# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4676 VSS row_n[6] a_6282_8194# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4677 a_1957_5166# VSS sample VDD sky130_fd_pr__pfet_01v8 ad=0.342 pd=2.97 as=0.342 ps=2.97 w=1.2 l=0.15
X4678 a_17326_18234# col_n[14] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4679 vcm a_2275_18218# a_22042_18194# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4680 a_7286_18234# col_n[4] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4681 a_2966_6146# a_2475_6170# a_2874_6146# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X4682 a_7382_14540# col_n[4] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X4683 a_17422_14540# col_n[14] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X4684 a_13310_5182# rowon_n[3] a_12914_5142# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X4685 a_14314_1166# VSS a_13918_1126# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X4686 vcm a_2275_1150# a_22042_1126# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4687 a_26058_10162# a_2475_10186# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4688 a_15014_9158# a_2475_9182# a_14922_9158# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X4689 a_28466_3496# col_n[25] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X4690 a_31078_5142# a_2475_5166# a_30986_5142# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X4691 vcm a_2275_5166# a_21038_5142# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4692 a_7894_10162# row_n[8] a_8386_10524# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4693 a_17934_10162# row_n[8] a_18426_10524# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4694 VDD rowon_n[3] a_2874_5142# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4695 a_16930_16186# row_n[14] a_17422_16548# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4696 a_6890_16186# row_n[14] a_7382_16548# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4697 VDD rowon_n[5] a_19942_7150# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4698 VDD rowon_n[1] a_12914_3134# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4699 a_26362_17230# rowon_n[15] a_25966_17190# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X4700 vcm a_2275_15206# a_15014_15182# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4701 VSS row_n[1] a_32386_3174# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4702 a_7986_4138# a_2475_4162# a_7894_4138# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X4703 vcm a_2275_15206# a_4974_15182# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4704 a_24354_9198# rowon_n[7] a_23958_9158# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X4705 a_6982_8154# a_2475_8178# a_6890_8154# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X4706 VSS row_n[11] a_27366_13214# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4707 a_31382_11206# rowon_n[9] a_30986_11166# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X4708 a_24354_10202# col_n[21] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4709 vcm a_2275_7174# a_25054_7150# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4710 vcm a_2275_3158# a_26058_3134# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4711 a_35094_7150# a_2475_7174# a_35002_7150# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X4712 vcm a_2275_6170# a_3970_6146# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4713 a_34490_6508# col_n[31] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X4714 a_17326_12210# rowon_n[10] a_16930_12170# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X4715 vcm a_2275_9182# a_16018_9158# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4716 a_2475_1150# a_1957_1150# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.171 pd=1.77 as=0.124 ps=1.01 w=0.6 l=0.15
X4717 a_7286_12210# rowon_n[10] a_6890_12170# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X4718 a_27062_2130# a_2475_2154# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4719 a_11302_2170# col_n[8] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4720 VDD rowon_n[13] a_25966_15182# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4721 a_14010_13174# a_2475_13198# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4722 a_23446_12532# col_n[20] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X4723 a_30986_8154# a_2275_8178# a_31078_8154# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4724 a_32482_1488# col_n[29] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X4725 a_31990_4138# a_2275_4162# a_32082_4138# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4726 a_3970_13174# a_2475_13198# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4727 VDD rowon_n[7] a_23958_9158# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4728 VDD rowon_n[3] a_24962_5142# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4729 a_31990_16186# a_2275_16210# a_32082_16186# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4730 a_27462_11528# col_n[24] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X4731 a_12914_5142# row_n[3] a_13406_5504# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4732 a_5278_4178# col_n[2] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4733 a_25358_18234# col_n[22] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4734 VDD rowon_n[8] a_16930_10162# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4735 VDD rowon_n[8] a_6890_10162# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4736 vcm a_2275_8178# a_7986_8154# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4737 vcm a_2275_4162# a_8990_4138# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4738 VSS row_n[15] a_5278_17230# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4739 VSS row_n[15] a_15318_17230# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4740 a_20034_17190# a_2475_17214# a_19942_17190# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X4741 a_22346_6186# col_n[19] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4742 a_24050_16186# a_2475_16210# a_23958_16186# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X4743 VDD a_2161_14202# a_2275_14202# VDD sky130_fd_pr__pfet_01v8 ad=0.249 pd=1.62 as=0.342 ps=2.97 w=1.2 l=0.15
X4744 a_16322_13214# col_n[13] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4745 vcm a_2275_13198# a_21038_13174# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4746 a_5278_7190# rowon_n[5] a_4882_7150# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X4747 vcm a_2275_1150# a_30074_1126# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4748 a_20946_17190# row_n[15] a_21438_17552# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4749 VSS row_n[14] a_9294_16226# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4750 a_15014_15182# a_2475_15206# a_14922_15182# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X4751 a_6282_13214# col_n[3] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4752 vcm a_2275_12194# a_34090_12170# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4753 a_19430_7512# col_n[16] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X4754 a_24962_16186# row_n[14] a_25454_16548# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4755 a_4974_15182# a_2475_15206# a_4882_15182# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X4756 VDD rowon_n[5] a_28978_7150# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4757 a_4882_4138# row_n[2] a_5374_4500# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4758 a_15414_15544# col_n[12] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X4759 a_8990_14178# a_2475_14202# a_8898_14178# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X4760 a_11910_12170# row_n[10] a_12402_12532# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4761 VDD VDD a_7894_18194# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4762 a_5374_15544# col_n[2] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X4763 VDD rowon_n[0] a_26970_2130# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4764 a_2475_13198# a_1957_13198# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.171 pd=1.77 as=0.124 ps=1.01 w=0.6 l=0.15
X4765 a_15926_11166# row_n[9] a_16418_11528# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4766 a_14922_2130# row_n[0] a_15414_2492# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4767 a_5886_11166# row_n[9] a_6378_11528# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4768 a_26362_8194# col_n[23] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4769 a_27366_4178# col_n[24] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4770 a_28066_12170# a_2475_12194# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4771 a_22954_10162# a_2275_10186# a_23046_10162# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4772 a_31382_2170# rowon_n[0] a_30986_2130# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X4773 VSS row_n[2] a_12306_4178# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4774 a_24354_18234# VDD a_23958_18194# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X4775 vcm a_2275_16210# a_2966_16186# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4776 vcm a_2275_16210# a_13006_16186# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4777 VSS row_n[13] a_21342_15222# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4778 a_25054_2130# a_2475_2154# a_24962_2130# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X4779 a_26970_4138# row_n[2] a_27462_4500# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4780 VDD rowon_n[3] a_32994_5142# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4781 VSS row_n[12] a_25358_14218# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4782 a_22346_11206# col_n[19] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4783 a_2966_4138# a_2475_4162# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4784 a_25966_17190# a_2275_17214# a_26058_17190# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4785 a_30074_15182# a_2475_15206# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4786 a_19942_7150# a_2275_7174# a_20034_7150# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4787 a_20946_3134# a_2275_3158# a_21038_3134# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4788 VDD rowon_n[15] a_19942_17190# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4789 a_15318_13214# rowon_n[11] a_14922_13174# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X4790 a_9294_9198# col_n[6] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4791 a_30074_7150# a_2475_7174# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4792 a_31078_3134# a_2475_3158# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4793 a_34090_14178# a_2475_14202# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4794 a_5278_13214# rowon_n[11] a_4882_13174# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X4795 a_10906_9158# a_2275_9182# a_10998_9158# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4796 VDD rowon_n[14] a_23958_16186# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4797 a_12002_14178# a_2475_14202# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4798 a_21438_13536# col_n[18] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X4799 a_18330_6186# rowon_n[4] a_17934_6146# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X4800 a_30378_6186# col_n[27] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4801 VSS row_n[1] a_4274_3174# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4802 a_12402_4500# col_n[9] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X4803 a_16930_12170# a_2275_12194# a_17022_12170# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4804 a_6890_12170# a_2275_12194# a_6982_12170# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4805 VSS row_n[10] a_14314_12210# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4806 vcm a_2275_6170# a_34090_6146# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4807 VSS row_n[10] a_4274_12210# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4808 VDD rowon_n[9] a_4882_11166# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4809 VDD rowon_n[9] a_14922_11166# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4810 a_6982_6146# a_2475_6170# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4811 VSS row_n[3] a_21342_5182# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4812 VSS VDD a_13310_18234# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4813 a_19942_12170# row_n[10] a_20434_12532# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4814 a_8898_9158# row_n[7] a_9390_9520# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4815 a_25966_1126# a_2275_1150# a_26058_1126# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4816 a_24962_5142# a_2275_5166# a_25054_5142# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4817 VSS VDD a_3270_18234# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4818 a_31078_17190# a_2475_17214# a_30986_17190# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X4819 a_3970_10162# a_2475_10186# a_3878_10162# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X4820 a_14010_10162# a_2475_10186# a_13918_10162# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X4821 a_2874_8154# a_2275_8178# a_2966_8154# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4822 a_4370_1488# en_C0_n VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X4823 a_3878_4138# a_2275_4162# a_3970_4138# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4824 a_35094_5142# a_2475_5166# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4825 VDD rowon_n[12] a_12914_14178# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4826 a_14314_14218# col_n[11] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4827 a_23446_8516# col_n[20] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X4828 a_31990_17190# row_n[15] a_32482_17552# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4829 a_13006_16186# a_2475_16210# a_12914_16186# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X4830 a_35094_16186# a_2475_16210# a_35002_16186# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X4831 VDD rowon_n[12] a_2874_14178# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4832 a_4274_14218# col_n[1] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4833 vcm a_2275_13198# a_32082_13174# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4834 VSS VDD a_9294_1166# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4835 a_35398_4178# VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4836 a_2966_16186# a_2475_16210# a_2874_16186# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X4837 a_4370_10524# col_n[1] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X4838 a_14410_10524# col_n[11] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X4839 a_18026_2130# a_2475_2154# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4840 a_21438_3496# col_n[18] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X4841 a_13406_16548# col_n[10] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X4842 a_3366_16548# col_n[0] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X4843 VSS row_n[5] a_25358_7190# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4844 VSS row_n[1] a_26362_3174# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4845 a_35398_7190# rowon_n[5] a_35002_7150# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X4846 VDD VSS sky130_fd_pr__cap_mim_m3_1 l=17.2 w=17.2
X4847 a_26058_13174# a_2475_13198# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4848 VSS row_n[7] a_16322_9198# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4849 a_7894_6146# a_2275_6170# a_7986_6146# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4850 a_28466_6508# col_n[25] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X4851 a_35002_4138# row_n[2] a_35494_4500# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4852 VSS row_n[13] a_19334_15222# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4853 a_23350_13214# rowon_n[11] a_22954_13174# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X4854 VSS row_n[8] a_20338_10202# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4855 a_20946_11166# a_2275_11190# a_21038_11166# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4856 a_11302_3174# rowon_n[1] a_10906_3134# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X4857 a_33998_10162# a_2275_10186# a_34090_10162# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4858 a_26458_1488# col_n[23] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X4859 a_35398_18234# VDD a_35002_18194# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X4860 a_18938_2130# a_2275_2154# a_19030_2130# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4861 VDD rowon_n[15] a_17934_17190# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4862 a_24962_12170# a_2275_12194# a_25054_12170# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4863 VDD rowon_n[4] a_12914_6146# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4864 a_20034_2130# a_2475_2154# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4865 a_16418_9520# col_n[13] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X4866 VSS row_n[6] a_8290_8194# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4867 a_23958_18194# a_2275_18218# a_24050_18194# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4868 a_19430_13536# col_n[16] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X4869 VDD rowon_n[9] a_22954_11166# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4870 VDD VSS a_10906_1126# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4871 a_20338_1166# en_bit_n[0] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4872 VSS VDD a_30378_1166# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4873 VSS row_n[15] a_34394_17230# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4874 a_2161_7174# sample VDD VDD sky130_fd_pr__pfet_01v8 ad=0.342 pd=2.97 as=0.342 ps=2.97 w=1.2 l=0.15
X4875 a_4974_6146# a_2475_6170# a_4882_6146# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X4876 a_3270_2170# rowon_n[0] a_2874_2130# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X4877 VDD rowon_n[14] a_35002_16186# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4878 a_17022_9158# a_2475_9182# a_16930_9158# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X4879 a_16322_1166# VSS a_15926_1126# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X4880 vcm a_2275_1150# a_24050_1126# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4881 vcm a_2275_5166# a_23046_5142# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4882 a_11302_17230# rowon_n[15] a_10906_17190# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X4883 a_35398_13214# VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4884 a_33086_5142# a_2475_5166# a_32994_5142# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X4885 a_29070_17190# a_2475_17214# a_28978_17190# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X4886 VSS row_n[11] a_12306_13214# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4887 a_30074_12170# a_2475_12194# a_29982_12170# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X4888 a_16018_2130# a_2475_2154# a_15926_2130# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X4889 a_34490_15544# col_n[31] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X4890 a_30986_12170# row_n[10] a_31478_12532# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4891 a_12002_11166# a_2475_11190# a_11910_11166# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X4892 a_34090_11166# a_2475_11190# a_33998_11166# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X4893 a_9902_7150# row_n[5] a_10394_7512# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4894 VDD rowon_n[5] a_21950_7150# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4895 VSS row_n[1] a_34394_3174# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4896 VDD rowon_n[13] a_10906_15182# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4897 a_35002_11166# row_n[9] a_35494_11528# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4898 a_26362_9198# rowon_n[7] a_25966_9158# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X4899 a_8990_8154# a_2475_8178# a_8898_8154# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X4900 a_9994_4138# a_2475_4162# a_9902_4138# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X4901 a_12402_11528# col_n[9] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X4902 a_19334_11206# rowon_n[9] a_18938_11166# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X4903 VDD rowon_n[0] a_19942_2130# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4904 vcm a_2275_3158# a_28066_3134# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4905 vcm a_2275_6170# a_5978_6146# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4906 a_10298_18234# col_n[7] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4907 vcm a_2275_9182# a_18026_9158# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4908 a_2475_5166# a_1957_5166# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.342 pd=2.97 as=0.249 ps=1.62 w=1.2 l=0.15
X4909 a_25358_2170# rowon_n[0] a_24962_2130# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X4910 a_13310_2170# col_n[10] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4911 a_32994_8154# a_2275_8178# a_33086_8154# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4912 a_29070_2130# a_2475_2154# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4913 a_33998_4138# a_2275_4162# a_34090_4138# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4914 a_15318_8194# rowon_n[6] a_14922_8154# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X4915 vcm a_2275_17214# a_18026_17190# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4916 VDD rowon_n[7] a_25966_9158# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4917 a_14922_5142# row_n[3] a_15414_5504# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4918 vcm a_2275_2154# a_17022_2130# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4919 VDD rowon_n[3] a_26970_5142# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4920 vcm a_2275_17214# a_7986_17190# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4921 VDD rowon_n[6] a_4882_8154# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4922 a_9902_16186# row_n[14] a_10394_16548# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4923 a_21342_14218# rowon_n[12] a_20946_14178# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X4924 a_34394_13214# rowon_n[11] a_33998_13174# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X4925 a_27366_12210# col_n[24] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4926 VSS row_n[8] a_31382_10202# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4927 a_22042_17190# a_2475_17214# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4928 a_31990_11166# a_2275_11190# a_32082_11166# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4929 a_24354_6186# col_n[21] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4930 a_22954_13174# a_2275_13198# a_23046_13174# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4931 VDD rowon_n[15] a_28978_17190# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4932 a_17022_15182# a_2475_15206# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4933 a_26458_14540# col_n[23] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X4934 VDD rowon_n[10] a_29982_12170# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4935 a_26058_10162# a_2475_10186# a_25966_10162# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X4936 a_7286_7190# rowon_n[5] a_6890_7150# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X4937 a_6982_15182# a_2475_15206# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4938 VDD rowon_n[9] a_33998_11166# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4939 a_26970_10162# row_n[8] a_27462_10524# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4940 VSS VDD a_32386_18234# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4941 VDD rowon_n[0] a_28978_2130# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4942 a_19430_2492# col_n[16] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X4943 a_33390_14218# col_n[30] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4944 a_29374_4178# col_n[26] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4945 a_27062_18194# a_2475_18218# a_26970_18194# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X4946 vcm a_2275_15206# a_24050_15182# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4947 VSS row_n[12] a_10298_14218# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4948 a_12002_9158# a_2475_9182# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4949 a_28370_8194# col_n[25] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4950 a_18026_17190# a_2475_17214# a_17934_17190# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X4951 a_9294_15222# col_n[6] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4952 a_19334_15222# col_n[16] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4953 a_27974_18194# VDD a_28466_18556# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4954 a_7986_17190# a_2475_17214# a_7894_17190# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X4955 a_10906_17190# a_2275_17214# a_10998_17190# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4956 vcm a_2275_14202# a_28066_14178# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4957 a_14922_16186# a_2275_16210# a_15014_16186# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4958 a_32482_16548# col_n[29] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X4959 a_33390_2170# rowon_n[0] a_32994_2130# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X4960 a_10998_2130# a_2475_2154# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4961 a_4882_16186# a_2275_16210# a_4974_16186# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4962 a_27062_2130# a_2475_2154# a_26970_2130# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X4963 VSS row_n[2] a_14314_4178# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4964 a_8386_17552# col_n[5] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X4965 a_18426_17552# col_n[15] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X4966 vcm a_2275_8178# a_31078_8154# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4967 a_17326_7190# col_n[14] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4968 vcm a_2275_4162# a_32082_4138# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4969 a_18938_13174# row_n[11] a_19430_13536# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4970 a_28978_4138# row_n[2] a_29470_4500# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4971 a_8898_13174# row_n[11] a_9390_13536# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4972 a_3970_8154# a_2475_8178# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4973 a_6890_7150# row_n[5] a_7382_7512# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4974 a_4974_4138# a_2475_4162# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4975 a_33086_3134# a_2475_3158# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4976 a_22954_3134# a_2275_3158# a_23046_3134# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4977 a_2161_16210# sample VSS VSS sky130_fd_pr__nfet_01v8 ad=0.171 pd=1.77 as=0.171 ps=1.77 w=0.6 l=0.15
X4978 a_32082_7150# a_2475_7174# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4979 a_12914_9158# a_2275_9182# a_13006_9158# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4980 a_21438_6508# col_n[18] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X4981 a_30074_10162# a_2475_10186# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4982 VSS row_n[8] a_29374_10202# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4983 a_14410_4500# col_n[11] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X4984 vcm a_2275_18218# a_5978_18194# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4985 vcm a_2275_18218# a_16018_18194# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4986 a_11910_2130# a_2275_2154# a_12002_2130# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4987 VSS row_n[14] a_28370_16226# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4988 a_32386_14218# rowon_n[12] a_31990_14178# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X4989 a_20034_18194# a_2475_18218# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4990 VDD rowon_n[10] a_27974_12170# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4991 a_8990_6146# a_2475_6170# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4992 VSS row_n[3] a_23350_5182# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4993 a_10998_17190# a_2475_17214# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4994 a_33086_17190# a_2475_17214# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4995 a_27974_1126# a_2275_1150# a_28066_1126# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4996 a_20946_14178# a_2275_14202# a_21038_14178# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4997 a_33998_13174# a_2275_13198# a_34090_13174# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4998 a_4882_8154# a_2275_8178# a_4974_8154# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4999 a_5886_4138# a_2275_4162# a_5978_4138# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5000 VDD VDD a_26970_18194# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5001 a_4974_16186# a_2475_16210# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5002 a_15014_16186# a_2475_16210# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5003 a_25454_8516# col_n[22] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X5004 VDD rowon_n[6] a_35002_8154# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5005 a_2161_17214# sample VDD VDD sky130_fd_pr__pfet_01v8 ad=0.342 pd=2.97 as=0.342 ps=2.97 w=1.2 l=0.15
X5006 a_23446_3496# col_n[20] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X5007 a_22954_14178# row_n[12] a_23446_14540# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5008 a_8290_10202# col_n[5] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5009 a_18330_10202# col_n[15] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5010 vcm a_2275_10186# a_23046_10162# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5011 a_32386_9198# col_n[29] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5012 VSS row_n[5] a_27366_7190# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5013 VSS row_n[1] a_28370_3174# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5014 a_6982_12170# a_2475_12194# a_6890_12170# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X5015 a_9902_12170# a_2275_12194# a_9994_12170# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5016 a_17022_12170# a_2475_12194# a_16930_12170# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X5017 VSS row_n[4] a_6282_6186# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5018 a_1957_3158# VSS sample VDD sky130_fd_pr__pfet_01v8 ad=0.342 pd=2.97 as=0.342 ps=2.97 w=1.2 l=0.15
X5019 a_17326_16226# col_n[14] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5020 vcm a_2275_16210# a_22042_16186# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5021 VSS row_n[7] a_18330_9198# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5022 a_16018_18194# a_2475_18218# a_15926_18194# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X5023 a_7286_16226# col_n[4] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5024 a_2161_1150# sample VSS VSS sky130_fd_pr__nfet_01v8 ad=0.171 pd=1.77 as=0.171 ps=1.77 w=0.6 l=0.15
X5025 a_2966_4138# a_2475_4162# a_2874_4138# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X5026 a_5978_18194# a_2475_18218# a_5886_18194# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X5027 a_7382_12532# col_n[4] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X5028 a_17422_12532# col_n[14] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X5029 VDD VSS VSS sky130_fd_pr__cap_var_lvt w=16.4 l=16
X5030 a_13310_3174# rowon_n[1] a_12914_3134# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X5031 vcm a_2275_7174# a_20034_7150# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5032 a_28466_1488# col_n[25] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X5033 a_31078_3134# a_2475_3158# a_30986_3134# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X5034 vcm a_2275_3158# a_21038_3134# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5035 a_16418_18556# col_n[13] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X5036 a_26970_8154# a_2275_8178# a_27062_8154# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5037 a_30074_7150# a_2475_7174# a_29982_7150# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X5038 VDD VSS VSS sky130_fd_pr__cap_var_lvt w=16.4 l=16
X5039 a_6378_18556# col_n[3] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X5040 vcm a_2275_9182# a_10998_9158# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5041 a_31990_9158# row_n[7] a_32482_9520# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5042 a_22042_2130# a_2475_2154# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5043 a_18426_9520# col_n[15] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X5044 VDD VSS a_12914_1126# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5045 VDD rowon_n[3] a_19942_5142# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5046 a_14922_17190# row_n[15] a_15414_17552# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5047 a_26362_15222# rowon_n[13] a_25966_15182# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X5048 vcm a_2275_13198# a_15014_13174# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5049 VSS row_n[10] a_23350_12210# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5050 VSS VDD a_32386_1166# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5051 a_4882_17190# row_n[15] a_5374_17552# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5052 vcm a_2275_13198# a_4974_13174# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5053 a_6982_6146# a_2475_6170# a_6890_6146# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X5054 vcm a_2275_1150# a_26058_1126# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5055 VSS row_n[9] a_27366_11206# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5056 vcm a_2275_5166# a_25054_5142# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5057 vcm a_2275_8178# a_2966_8154# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5058 vcm a_2275_4162# a_3970_4138# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5059 a_35094_5142# a_2475_5166# a_35002_5142# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X5060 VDD VSS VSS sky130_fd_pr__cap_var_lvt w=16.4 l=16
X5061 VDD rowon_n[12] a_21950_14178# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5062 a_32082_12170# a_2475_12194# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5063 a_17326_10202# rowon_n[8] a_16930_10162# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X5064 VDD VSS sky130_fd_pr__cap_mim_m3_1 l=17.2 w=17.2
X5065 a_7286_10202# rowon_n[8] a_6890_10162# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X5066 a_18026_2130# a_2475_2154# a_17934_2130# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X5067 a_31078_18194# a_2475_18218# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5068 VDD rowon_n[11] a_25966_13174# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5069 a_23446_10524# col_n[20] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X5070 a_30986_6146# a_2275_6170# a_31078_6146# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5071 VDD rowon_n[5] a_23958_7150# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5072 a_21342_17230# col_n[18] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5073 a_31990_14178# a_2275_14202# a_32082_14178# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5074 a_25358_16226# col_n[22] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5075 a_28370_9198# rowon_n[7] a_27974_9158# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X5076 VDD rowon_n[0] a_21950_2130# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5077 a_29982_17190# a_2275_17214# a_30074_17190# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5078 vcm a_2275_6170# a_7986_6146# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5079 a_9902_2130# row_n[0] a_10394_2492# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5080 a_8290_18234# VDD a_7894_18194# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X5081 VSS row_n[13] a_5278_15222# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5082 VSS row_n[13] a_15318_15222# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5083 a_20034_15182# a_2475_15206# a_19942_15182# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X5084 a_12306_12210# col_n[9] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5085 a_21342_8194# col_n[18] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5086 a_27366_2170# rowon_n[0] a_26970_2130# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X5087 a_22346_4178# col_n[19] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5088 a_24450_18556# col_n[21] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X5089 a_24050_14178# a_2475_14202# a_23958_14178# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X5090 a_16322_11206# col_n[13] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5091 vcm a_2275_11190# a_21038_11166# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5092 VSS row_n[6] a_31382_8194# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5093 a_5278_5182# rowon_n[3] a_4882_5142# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X5094 a_15318_2170# col_n[12] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5095 a_20946_15182# row_n[13] a_21438_15544# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5096 VSS row_n[12] a_9294_14218# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5097 a_33998_14178# row_n[12] a_34490_14540# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5098 a_15014_13174# a_2475_13198# a_14922_13174# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X5099 a_6282_11206# col_n[3] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5100 vcm a_2275_10186# a_34090_10162# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5101 a_17326_8194# rowon_n[6] a_16930_8154# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X5102 a_35002_8154# a_2275_8178# a_35094_8154# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5103 a_19430_5504# col_n[16] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X5104 a_4974_13174# a_2475_13198# a_4882_13174# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X5105 VDD rowon_n[7] a_27974_9158# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5106 vcm a_2275_2154# a_19030_2130# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5107 VDD rowon_n[3] a_28978_5142# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5108 VDD rowon_n[15] a_3878_17190# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5109 VDD rowon_n[15] a_13918_17190# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5110 a_11398_14540# col_n[8] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X5111 VDD rowon_n[6] a_6890_8154# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5112 a_15414_13536# col_n[12] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X5113 a_11910_10162# row_n[8] a_12402_10524# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5114 a_20034_2130# a_2475_2154# a_19942_2130# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X5115 VDD rowon_n[14] a_7894_16186# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5116 a_5374_13536# col_n[2] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X5117 a_26058_7150# a_2475_7174# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5118 a_21950_4138# row_n[2] a_22442_4500# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5119 VDD rowon_n[1] a_4882_3134# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5120 a_26362_6186# col_n[23] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5121 vcm a_2275_18218# a_35094_18194# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5122 a_4274_9198# col_n[1] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5123 a_9294_7190# rowon_n[5] a_8898_7150# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X5124 a_20338_17230# rowon_n[15] a_19942_17190# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X5125 a_17022_10162# a_2475_10186# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5126 a_2874_18194# VDD a_3366_18556# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5127 a_12914_18194# VDD a_13406_18556# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5128 a_24354_16226# rowon_n[14] a_23958_16186# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X5129 vcm a_2275_14202# a_2966_14178# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5130 vcm a_2275_14202# a_13006_14178# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5131 VSS row_n[11] a_21342_13214# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5132 a_6982_10162# a_2475_10186# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5133 a_29070_18194# a_2475_18218# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5134 a_25966_15182# a_2275_15206# a_26058_15182# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5135 a_30074_13174# a_2475_13198# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5136 a_3878_9158# row_n[7] a_4370_9520# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5137 a_14010_9158# a_2475_9182# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5138 a_20946_1126# a_2275_1150# a_21038_1126# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5139 a_19942_5142# a_2275_5166# a_20034_5142# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5140 VDD rowon_n[13] a_19942_15182# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5141 a_5278_11206# rowon_n[9] a_4882_11166# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X5142 a_15318_11206# rowon_n[9] a_14922_11166# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X5143 a_16930_8154# row_n[6] a_17422_8516# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5144 a_31078_1126# a_2475_1150# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5145 a_30074_5142# a_2475_5166# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5146 a_9994_17190# a_2475_17214# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5147 a_20338_12210# col_n[17] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5148 a_21438_11528# col_n[18] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X5149 VSS en_C0_n a_4274_1166# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5150 a_30378_4178# col_n[27] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5151 a_18330_4178# rowon_n[2] a_17934_4138# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X5152 a_13006_2130# a_2475_2154# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5153 a_32386_17230# col_n[29] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5154 a_29070_2130# a_2475_2154# a_28978_2130# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X5155 VSS row_n[8] a_14314_10202# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5156 vcm a_2275_8178# a_33086_8154# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5157 a_19334_7190# col_n[16] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5158 vcm a_2275_4162# a_34090_4138# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5159 a_4882_11166# a_2275_11190# a_4974_11166# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5160 a_14922_11166# a_2275_11190# a_15014_11166# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5161 VSS row_n[8] a_4274_10202# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5162 VSS row_n[5] a_20338_7190# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5163 VSS row_n[1] a_21342_3174# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5164 a_6982_4138# a_2475_4162# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5165 VSS row_n[14] a_13310_16226# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5166 a_19942_10162# row_n[8] a_20434_10524# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5167 a_8898_7150# row_n[5] a_9390_7512# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5168 a_30378_7190# rowon_n[5] a_29982_7150# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X5169 a_24962_3134# a_2275_3158# a_25054_3134# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5170 vcm a_2275_17214# a_27062_17190# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5171 VSS row_n[14] a_3270_16226# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5172 a_31078_15182# a_2475_15206# a_30986_15182# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X5173 VSS row_n[7] a_11302_9198# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5174 a_34090_7150# a_2475_7174# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5175 a_2874_6146# a_2275_6170# a_2966_6146# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5176 a_35094_3134# a_2475_3158# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5177 VDD rowon_n[10] a_12914_12170# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5178 a_23446_6508# col_n[20] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X5179 a_6890_2130# row_n[0] a_7382_2492# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5180 a_29982_4138# row_n[2] a_30474_4500# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5181 VDD rowon_n[2] a_17934_4138# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5182 a_35494_18556# VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X5183 a_31990_15182# row_n[13] a_32482_15544# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5184 a_13006_14178# a_2475_14202# a_12914_14178# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X5185 a_35094_14178# a_2475_14202# a_35002_14178# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X5186 VDD rowon_n[10] a_2874_12170# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5187 vcm a_2275_11190# a_32082_11166# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5188 a_14922_9158# a_2275_9182# a_15014_9158# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5189 a_7894_18194# a_2275_18218# a_7986_18194# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5190 VDD VDD a_11910_18194# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5191 a_17934_18194# a_2275_18218# a_18026_18194# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5192 a_2966_14178# a_2475_14202# a_2874_14178# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X5193 a_2161_11190# sample VSS VSS sky130_fd_pr__nfet_01v8 ad=0.171 pd=1.77 as=0.171 ps=1.77 w=0.6 l=0.15
X5194 VDD a_2161_2154# a_2275_2154# VDD sky130_fd_pr__pfet_01v8 ad=0.249 pd=1.62 as=0.342 ps=2.97 w=1.2 l=0.15
X5195 a_21438_1488# col_n[18] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X5196 a_13918_2130# a_2275_2154# a_14010_2130# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5197 VSS VDD a_26362_1166# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5198 VSS row_n[3] a_25358_5182# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5199 a_11398_9520# col_n[8] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X5200 VSS row_n[6] a_3270_8194# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5201 a_35398_5182# rowon_n[3] a_35002_5142# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X5202 a_18330_17230# rowon_n[15] a_17934_17190# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X5203 a_7894_4138# a_2275_4162# a_7986_4138# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5204 a_27462_8516# col_n[24] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X5205 VSS row_n[11] a_19334_13214# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5206 a_23350_11206# rowon_n[9] a_22954_11166# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X5207 a_12002_9158# a_2475_9182# a_11910_9158# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X5208 a_11302_1166# VSS a_10906_1126# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X5209 a_4974_11166# a_2475_11190# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5210 a_15014_11166# a_2475_11190# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5211 a_25454_3496# col_n[22] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X5212 a_35398_16226# rowon_n[14] a_35002_16186# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X5213 VDD rowon_n[1] a_35002_3134# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5214 VDD rowon_n[13] a_17934_15182# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5215 a_10998_2130# a_2475_2154# a_10906_2130# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X5216 a_8990_12170# a_2475_12194# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5217 a_34394_9198# col_n[31] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5218 a_16418_7512# col_n[13] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X5219 VSS row_n[5] a_29374_7190# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5220 VSS row_n[4] a_8290_6186# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5221 a_23958_16186# a_2275_16210# a_24050_16186# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5222 a_19430_11528# col_n[16] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X5223 a_7986_18194# a_2475_18218# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5224 a_18026_18194# a_2475_18218# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5225 VSS row_n[13] a_34394_15222# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5226 a_31382_12210# col_n[28] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5227 a_21342_9198# rowon_n[7] a_20946_9158# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X5228 a_3970_8154# a_2475_8178# a_3878_8154# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X5229 a_2161_5166# sample VDD VDD sky130_fd_pr__pfet_01v8 ad=0.342 pd=2.97 as=0.342 ps=2.97 w=1.2 l=0.15
X5230 a_4974_4138# a_2475_4162# a_4882_4138# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X5231 vcm a_2275_3158# a_23046_3134# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5232 a_11302_15222# rowon_n[13] a_10906_15182# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X5233 a_35398_11206# VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5234 a_28978_8154# a_2275_8178# a_29070_8154# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5235 a_32082_7150# a_2475_7174# a_31990_7150# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X5236 a_33086_3134# a_2475_3158# a_32994_3134# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X5237 vcm a_2275_9182# a_13006_9158# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5238 a_20338_2170# rowon_n[0] a_19942_2130# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X5239 VDD rowon_n[15] a_32994_17190# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5240 a_29070_15182# a_2475_15206# a_28978_15182# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X5241 a_30474_14540# col_n[27] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X5242 vcm a_2275_12194# a_26058_12170# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5243 VSS row_n[9] a_12306_11206# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5244 a_30074_10162# a_2475_10186# a_29982_10162# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X5245 a_33998_9158# row_n[7] a_34490_9520# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5246 a_24050_2130# a_2475_2154# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5247 a_34490_13536# col_n[31] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X5248 a_30986_10162# row_n[8] a_31478_10524# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5249 a_10298_8194# rowon_n[6] a_9902_8154# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X5250 VDD rowon_n[3] a_21950_5142# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5251 VDD rowon_n[7] a_20946_9158# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5252 a_9902_5142# row_n[3] a_10394_5504# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5253 vcm a_2275_2154# a_12002_2130# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5254 VDD rowon_n[11] a_10906_13174# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5255 a_8990_6146# a_2475_6170# a_8898_6146# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X5256 vcm a_2275_1150# a_28066_1126# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5257 vcm a_2275_8178# a_4974_8154# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5258 vcm a_2275_4162# a_5978_4138# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5259 a_10298_16226# col_n[7] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5260 a_2475_3158# a_1957_3158# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.342 pd=2.97 as=0.249 ps=1.62 w=1.2 l=0.15
X5261 a_32994_6146# a_2275_6170# a_33086_6146# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5262 a_15318_6186# rowon_n[4] a_14922_6146# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X5263 a_29374_17230# rowon_n[15] a_28978_17190# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X5264 vcm a_2275_15206# a_18026_15182# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5265 VDD rowon_n[5] a_25966_7150# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5266 vcm a_2275_15206# a_7986_15182# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5267 a_30378_12210# rowon_n[10] a_29982_12170# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X5268 VDD rowon_n[4] a_4882_6146# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5269 a_34394_11206# rowon_n[9] a_33998_11166# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X5270 a_27366_10202# col_n[24] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5271 VDD rowon_n[0] a_23958_2130# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5272 a_22042_15182# a_2475_15206# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5273 VSS row_n[0] a_19334_2170# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5274 a_24354_4178# col_n[21] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5275 a_23350_8194# col_n[20] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5276 VSS row_n[6] a_33390_8194# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5277 a_29374_2170# rowon_n[0] a_28978_2130# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X5278 VDD rowon_n[13] a_28978_15182# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5279 a_17022_13174# a_2475_13198# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5280 a_26458_12532# col_n[23] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X5281 VDD rowon_n[8] a_29982_10162# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5282 a_7286_5182# rowon_n[3] a_6890_5142# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X5283 a_6982_13174# a_2475_13198# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5284 vcm a_2275_8178# a_27062_8154# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5285 VDD rowon_n[6] a_8898_8154# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5286 a_22042_2130# a_2475_2154# a_21950_2130# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X5287 a_28370_18234# col_n[25] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5288 VSS row_n[14] a_32386_16226# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5289 a_12306_7190# col_n[9] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5290 a_28066_7150# a_2475_7174# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5291 VDD VSS sky130_fd_pr__cap_mim_m3_1 l=17.2 w=17.2
X5292 VDD rowon_n[1] a_6890_3134# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5293 a_23958_4138# row_n[2] a_24450_4500# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5294 VSS row_n[15] a_8290_17230# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5295 VSS row_n[15] a_18330_17230# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5296 a_23046_17190# a_2475_17214# a_22954_17190# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X5297 a_27062_16186# a_2475_16210# a_26970_16186# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X5298 vcm a_2275_13198# a_24050_13174# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5299 a_28370_6186# col_n[25] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5300 VDD VDD a_30986_18194# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5301 a_23958_17190# row_n[15] a_24450_17552# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5302 a_18026_15182# a_2475_15206# a_17934_15182# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X5303 a_9294_13214# col_n[6] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5304 a_19334_13214# col_n[16] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5305 a_6282_9198# col_n[3] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5306 a_27974_16186# row_n[14] a_28466_16548# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5307 a_7986_15182# a_2475_15206# a_7894_15182# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X5308 a_10906_15182# a_2275_15206# a_10998_15182# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5309 a_14922_14178# a_2275_14202# a_15014_14178# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5310 a_4882_14178# a_2275_14202# a_4974_14178# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5311 a_8386_15544# col_n[5] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X5312 a_18426_15544# col_n[15] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X5313 vcm a_2275_6170# a_31078_6146# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5314 a_17326_5182# col_n[14] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5315 a_18938_11166# row_n[9] a_19430_11528# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5316 a_8898_11166# row_n[9] a_9390_11528# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5317 a_5886_9158# row_n[7] a_6378_9520# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5318 a_3970_6146# a_2475_6170# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5319 a_6890_5142# row_n[3] a_7382_5504# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5320 a_18938_8154# row_n[6] a_19430_8516# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5321 a_22954_1126# a_2275_1150# a_23046_1126# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5322 a_33086_1126# a_2475_1150# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5323 a_2161_14202# sample VSS VSS sky130_fd_pr__nfet_01v8 ad=0.171 pd=1.77 as=0.171 ps=1.77 w=0.6 l=0.15
X5324 a_32082_5142# a_2475_5166# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5325 vcm a_2275_17214# a_12002_17190# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5326 a_28370_12210# rowon_n[10] a_27974_12170# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X5327 a_25966_10162# a_2275_10186# a_26058_10162# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5328 a_20434_8516# col_n[17] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X5329 VDD rowon_n[6] a_29982_8154# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5330 a_15014_2130# a_2475_2154# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5331 a_16930_3134# row_n[1] a_17422_3496# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5332 a_27366_18234# VDD a_26970_18194# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X5333 vcm a_2275_16210# a_5978_16186# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5334 vcm a_2275_16210# a_16018_16186# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5335 vcm a_2275_8178# a_35094_8154# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5336 VSS row_n[12] a_28370_14218# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5337 a_28978_17190# a_2275_17214# a_29070_17190# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5338 a_20034_16186# a_2475_16210# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5339 VDD rowon_n[8] a_27974_10162# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5340 VSS row_n[5] a_22346_7190# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5341 VSS row_n[1] a_23350_3174# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5342 a_8990_4138# a_2475_4162# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5343 a_10998_15182# a_2475_15206# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5344 a_33086_15182# a_2475_15206# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5345 a_32386_7190# rowon_n[5] a_31990_7150# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X5346 VSS row_n[7] a_13310_9198# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5347 a_19030_9158# a_2475_9182# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5348 a_26058_7150# a_2475_7174# a_25966_7150# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X5349 a_4882_6146# a_2275_6170# a_4974_6146# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5350 VDD rowon_n[14] a_26970_16186# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5351 a_4974_14178# a_2475_14202# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5352 a_15014_14178# a_2475_14202# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5353 a_25454_6508# col_n[22] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X5354 a_8898_2130# row_n[0] a_9390_2492# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5355 VDD rowon_n[4] a_35002_6146# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5356 a_2161_15206# sample VDD VDD sky130_fd_pr__pfet_01v8 ad=0.342 pd=2.97 as=0.342 ps=2.97 w=1.2 l=0.15
X5357 a_23446_1488# col_n[20] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X5358 VSS row_n[10] a_17326_12210# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5359 a_22042_12170# a_2475_12194# a_21950_12170# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X5360 a_21950_8154# a_2275_8178# a_22042_8154# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5361 a_15926_2130# a_2275_2154# a_16018_2130# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5362 VSS row_n[10] a_7286_12210# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5363 VSS VDD a_16322_18234# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5364 a_21038_18194# a_2475_18218# a_20946_18194# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X5365 a_22954_12170# row_n[10] a_23446_12532# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5366 VSS VDD a_28370_1166# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5367 VSS row_n[3] a_27366_5182# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5368 VSS VDD a_6282_18234# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5369 a_6982_10162# a_2475_10186# a_6890_10162# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X5370 a_17022_10162# a_2475_10186# a_16930_10162# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X5371 a_13406_9520# col_n[10] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X5372 VSS row_n[6] a_5278_8194# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5373 a_1957_1150# VSS sample VDD sky130_fd_pr__pfet_01v8 ad=0.342 pd=2.97 as=0.342 ps=2.97 w=1.2 l=0.15
X5374 VSS row_n[2] a_6282_4178# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5375 a_21950_18194# VDD a_22442_18556# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5376 VDD rowon_n[12] a_15926_14178# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5377 a_17326_14218# col_n[14] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5378 vcm a_2275_14202# a_22042_14178# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5379 a_1957_17214# VDD sample VSS sky130_fd_pr__nfet_01v8 ad=0.171 pd=1.77 as=0.171 ps=1.77 w=0.6 l=0.15
X5380 a_16018_16186# a_2475_16210# a_15926_16186# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X5381 VDD rowon_n[12] a_5886_14178# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5382 a_7286_14218# col_n[4] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5383 a_29470_8516# col_n[26] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X5384 a_5978_16186# a_2475_16210# a_5886_16186# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X5385 a_7382_10524# col_n[4] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X5386 a_17422_10524# col_n[14] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X5387 a_13310_1166# VSS a_12914_1126# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X5388 vcm a_2275_1150# a_21038_1126# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5389 a_15318_17230# col_n[12] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5390 vcm a_2275_17214# a_20034_17190# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5391 a_14010_9158# a_2475_9182# a_13918_9158# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X5392 a_31078_1126# a_2475_1150# a_30986_1126# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X5393 vcm a_2275_5166# a_20034_5142# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5394 a_5278_17230# col_n[2] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5395 a_16418_16548# col_n[13] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X5396 a_26970_6146# a_2275_6170# a_27062_6146# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5397 a_27462_3496# col_n[24] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X5398 a_30074_5142# a_2475_5166# a_29982_5142# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X5399 a_6378_16548# col_n[3] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X5400 a_31990_7150# row_n[5] a_32482_7512# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5401 a_6378_4500# col_n[3] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X5402 a_13006_2130# a_2475_2154# a_12914_2130# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X5403 vcm a_2275_12194# a_10998_12170# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5404 a_18426_7512# col_n[15] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X5405 a_14922_15182# row_n[13] a_15414_15544# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5406 a_26362_13214# rowon_n[11] a_25966_13174# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X5407 vcm a_2275_11190# a_15014_11166# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5408 VSS row_n[8] a_23350_10202# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5409 a_16418_2492# col_n[13] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X5410 a_4882_15182# row_n[13] a_5374_15544# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5411 vcm a_2275_11190# a_4974_11166# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5412 a_23958_11166# a_2275_11190# a_24050_11166# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5413 a_23350_9198# rowon_n[7] a_22954_9158# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X5414 a_6982_4138# a_2475_4162# a_6890_4138# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X5415 a_35094_3134# a_2475_3158# a_35002_3134# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X5416 vcm a_2275_3158# a_25054_3134# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5417 a_1957_18218# VSS sample VDD sky130_fd_pr__pfet_01v8 ad=0.342 pd=2.97 as=0.342 ps=2.97 w=1.2 l=0.15
X5418 a_34090_7150# a_2475_7174# a_33998_7150# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X5419 vcm a_2275_6170# a_2966_6146# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5420 VDD rowon_n[10] a_21950_12170# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5421 a_27974_12170# a_2275_12194# a_28066_12170# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5422 vcm a_2275_9182# a_15014_9158# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5423 a_22346_2170# rowon_n[0] a_21950_2130# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X5424 a_10298_2170# col_n[7] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5425 a_26970_18194# a_2275_18218# a_27062_18194# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5426 a_31078_16186# a_2475_16210# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5427 VDD rowon_n[9] a_25966_11166# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5428 a_12306_8194# rowon_n[6] a_11910_8154# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X5429 a_29982_8154# a_2275_8178# a_30074_8154# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5430 a_30986_4138# a_2275_4162# a_31078_4138# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5431 VDD rowon_n[7] a_22954_9158# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5432 vcm a_2275_2154# a_14010_2130# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5433 VDD rowon_n[3] a_23958_5142# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5434 VSS VDD a_24354_18234# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5435 a_21342_15222# col_n[18] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5436 a_25358_14218# col_n[22] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5437 a_14314_17230# rowon_n[15] a_13918_17190# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X5438 a_21038_7150# a_2475_7174# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5439 a_19030_18194# a_2475_18218# a_18938_18194# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X5440 a_4274_17230# rowon_n[15] a_3878_17190# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X5441 a_29982_15182# a_2275_15206# a_30074_15182# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5442 vcm a_2275_4162# a_7986_4138# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5443 a_20434_17552# col_n[17] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X5444 a_8290_16226# rowon_n[14] a_7894_16186# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X5445 VSS row_n[11] a_5278_13214# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5446 VSS row_n[11] a_15318_13214# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5447 a_20034_13174# a_2475_13198# a_19942_13174# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X5448 a_33086_12170# a_2475_12194# a_32994_12170# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X5449 a_12306_10202# col_n[9] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5450 a_21342_6186# col_n[18] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5451 a_24450_16548# col_n[21] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X5452 a_20946_13174# row_n[11] a_21438_13536# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5453 a_10998_12170# a_2475_12194# a_10906_12170# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X5454 a_4274_7190# rowon_n[5] a_3878_7150# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X5455 VSS row_n[4] a_31382_6186# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5456 a_5278_3174# rowon_n[1] a_4882_3134# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X5457 a_33998_12170# row_n[10] a_34490_12532# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5458 a_15014_11166# a_2475_11190# a_14922_11166# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X5459 a_17326_6186# rowon_n[4] a_16930_6146# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X5460 a_35002_6146# a_2275_6170# a_35094_6146# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5461 a_4974_11166# a_2475_11190# a_4882_11166# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X5462 VDD rowon_n[5] a_27974_7150# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5463 VDD rowon_n[13] a_3878_15182# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5464 VDD rowon_n[13] a_13918_15182# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5465 a_11398_12532# col_n[8] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X5466 VDD rowon_n[4] a_6890_6146# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5467 a_15414_11528# col_n[12] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X5468 a_5374_11528# col_n[2] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X5469 VDD rowon_n[0] a_25966_2130# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5470 a_26058_5142# a_2475_5166# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5471 a_13310_18234# col_n[10] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5472 VDD VSS a_4882_1126# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5473 a_3270_18234# col_n[0] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5474 vcm a_2275_17214# a_31078_17190# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5475 a_25358_8194# col_n[22] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5476 a_26362_4178# col_n[23] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5477 vcm a_2275_16210# a_35094_16186# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5478 a_11910_8154# row_n[6] a_12402_8516# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5479 VSS row_n[6] a_35398_8194# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5480 a_9294_5182# rowon_n[3] a_8898_5142# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X5481 a_22042_10162# a_2475_10186# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5482 a_20338_15222# rowon_n[13] a_19942_15182# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X5483 vcm a_2275_8178# a_29070_8154# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5484 a_2874_16186# row_n[14] a_3366_16548# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5485 a_12914_16186# row_n[14] a_13406_16548# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5486 a_24354_14218# rowon_n[12] a_23958_14178# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X5487 VSS row_n[9] a_21342_11206# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5488 a_24050_2130# a_2475_2154# a_23958_2130# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X5489 a_25054_17190# a_2475_17214# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5490 a_14314_7190# col_n[11] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5491 VDD rowon_n[1] a_8898_3134# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5492 a_25966_4138# row_n[2] a_26458_4500# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5493 a_29070_16186# a_2475_16210# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5494 a_25966_13174# a_2275_13198# a_26058_13174# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5495 a_3878_7150# row_n[5] a_4370_7512# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5496 a_19942_3134# a_2275_3158# a_20034_3134# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5497 VDD VDD a_18938_18194# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5498 VDD rowon_n[11] a_19942_13174# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5499 a_8290_9198# col_n[5] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5500 a_16930_6146# row_n[4] a_17422_6508# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5501 a_30074_3134# a_2475_3158# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5502 a_9994_15182# a_2475_15206# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5503 a_20338_10202# col_n[17] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5504 a_2475_12194# a_1957_12194# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.342 pd=2.97 as=0.249 ps=1.62 w=1.2 l=0.15
X5505 a_9902_9158# a_2275_9182# a_9994_9158# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5506 a_13310_12210# rowon_n[10] a_12914_12170# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X5507 VSS VDD a_35398_18234# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5508 a_32386_15222# col_n[29] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5509 a_3270_12210# rowon_n[10] a_2874_12170# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X5510 a_10906_10162# a_2275_10186# a_10998_10162# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5511 a_7286_2170# col_n[4] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5512 vcm a_2275_6170# a_33086_6146# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5513 a_19334_5182# col_n[16] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5514 a_12306_18234# VDD a_11910_18194# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X5515 VSS VDD a_21342_1166# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5516 VSS row_n[3] a_20338_5182# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5517 VSS row_n[12] a_13310_14218# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5518 a_7894_9158# row_n[7] a_8386_9520# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5519 a_8898_5142# row_n[3] a_9390_5504# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5520 a_24962_1126# a_2275_1150# a_25054_1126# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5521 a_30378_5182# rowon_n[3] a_29982_5142# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X5522 a_31478_17552# col_n[28] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X5523 vcm a_2275_15206# a_27062_15182# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5524 VSS row_n[12] a_3270_14218# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5525 a_31078_13174# a_2475_13198# a_30986_13174# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X5526 a_35094_1126# a_2475_1150# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5527 a_2874_4138# a_2275_4162# a_2966_4138# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5528 a_34090_5142# a_2475_5166# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5529 a_3878_17190# a_2275_17214# a_3970_17190# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5530 a_13918_17190# a_2275_17214# a_14010_17190# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5531 VDD rowon_n[8] a_12914_10162# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5532 a_22442_8516# col_n[19] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X5533 a_35494_16548# VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X5534 a_31990_13174# row_n[11] a_32482_13536# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5535 VDD rowon_n[8] a_2874_10162# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5536 VDD rowon_n[6] a_31990_8154# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5537 a_18938_3134# row_n[1] a_19430_3496# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5538 a_7894_16186# a_2275_16210# a_7986_16186# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5539 VDD rowon_n[14] a_11910_16186# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5540 a_17934_16186# a_2275_16210# a_18026_16186# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5541 a_17022_2130# a_2475_2154# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5542 a_20434_3496# col_n[17] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X5543 vcm a_2275_12194# a_30074_12170# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5544 VDD rowon_n[1] a_29982_3134# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5545 VSS row_n[1] a_25358_3174# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5546 a_11398_7512# col_n[8] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X5547 VSS row_n[5] a_24354_7190# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5548 a_34394_7190# rowon_n[5] a_33998_7150# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X5549 VSS row_n[4] a_3270_6186# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5550 a_35398_3174# rowon_n[1] a_35002_3134# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X5551 a_18330_15222# rowon_n[13] a_17934_15182# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X5552 a_20034_11166# a_2475_11190# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5553 VSS row_n[7] a_15318_9198# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5554 a_28066_7150# a_2475_7174# a_27974_7150# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X5555 a_27462_6508# col_n[24] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X5556 VSS row_n[9] a_19334_11206# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5557 a_10998_10162# a_2475_10186# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5558 a_33086_10162# a_2475_10186# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5559 vcm a_2275_18218# a_19030_18194# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5560 a_5978_9158# a_2475_9182# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5561 vcm a_2275_18218# a_8990_18194# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5562 a_24050_12170# a_2475_12194# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5563 a_23958_8154# a_2275_8178# a_24050_8154# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5564 a_25454_1488# col_n[22] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X5565 a_35398_14218# rowon_n[12] a_35002_14178# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X5566 VDD VSS a_35002_1126# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5567 analog_in sw_n ctop VDD sky130_fd_pr__pfet_01v8 ad=0.275 pd=2.19 as=0.275 ps=2.19 w=1.9 l=0.22
X5568 a_17934_2130# a_2275_2154# a_18026_2130# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5569 a_23046_18194# a_2475_18218# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5570 VDD rowon_n[11] a_17934_13174# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5571 VSS row_n[3] a_29374_5182# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5572 a_15414_9520# col_n[12] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X5573 a_16418_5504# col_n[13] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X5574 VSS row_n[2] a_8290_4178# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5575 a_33390_17230# rowon_n[15] a_32994_17190# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X5576 a_23958_14178# a_2275_14202# a_24050_14178# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5577 VSS row_n[6] a_7286_8194# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5578 a_7986_16186# a_2475_16210# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5579 a_18026_16186# a_2475_16210# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5580 VSS row_n[11] a_34394_13214# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5581 a_31382_10202# col_n[28] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5582 a_3970_6146# a_2475_6170# a_3878_6146# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X5583 a_2161_3158# sample VDD VDD sky130_fd_pr__pfet_01v8 ad=0.342 pd=2.97 as=0.342 ps=2.97 w=1.2 l=0.15
X5584 vcm a_2275_1150# a_23046_1126# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5585 a_11302_13214# rowon_n[11] a_10906_13174# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X5586 a_1957_12194# VDD sample VSS sky130_fd_pr__nfet_01v8 ad=0.171 pd=1.77 as=0.171 ps=1.77 w=0.6 l=0.15
X5587 a_28978_6146# a_2275_6170# a_29070_6146# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5588 a_33086_1126# a_2475_1150# a_32994_1126# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X5589 a_29470_3496# col_n[26] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X5590 a_32082_5142# a_2475_5166# a_31990_5142# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X5591 a_6890_9158# a_2275_9182# a_6982_9158# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5592 a_29470_17552# col_n[26] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X5593 VDD rowon_n[13] a_32994_15182# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5594 a_25966_14178# row_n[12] a_26458_14540# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5595 a_29070_13174# a_2475_13198# a_28978_13174# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X5596 a_30474_12532# col_n[27] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X5597 vcm a_2275_10186# a_26058_10162# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5598 a_33998_7150# row_n[5] a_34490_7512# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5599 a_8386_4500# col_n[5] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X5600 a_9994_12170# a_2475_12194# a_9902_12170# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X5601 a_12914_12170# a_2275_12194# a_13006_12170# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5602 a_15014_2130# a_2475_2154# a_14922_2130# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X5603 a_2874_12170# a_2275_12194# a_2966_12170# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5604 a_34490_11528# col_n[31] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X5605 a_10298_6186# rowon_n[4] a_9902_6146# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X5606 a_31990_2130# row_n[0] a_32482_2492# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5607 VDD VSS VSS sky130_fd_pr__cap_var_lvt w=16.4 l=16
X5608 a_11910_18194# a_2275_18218# a_12002_18194# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5609 VDD rowon_n[9] a_10906_11166# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5610 VDD rowon_n[5] a_20946_7150# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5611 a_18426_2492# col_n[15] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X5612 a_8990_4138# a_2475_4162# a_8898_4138# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X5613 a_19030_9158# a_2475_9182# a_18938_9158# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X5614 vcm a_2275_6170# a_4974_6146# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5615 a_10298_14218# col_n[7] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5616 a_2475_1150# a_1957_1150# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.342 pd=2.97 as=0.249 ps=1.62 w=1.2 l=0.15
X5617 a_24354_2170# rowon_n[0] a_23958_2130# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X5618 a_32994_4138# a_2275_4162# a_33086_4138# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5619 a_14314_8194# rowon_n[6] a_13918_8154# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X5620 vcm a_2275_8178# a_22042_8154# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5621 a_15318_4178# rowon_n[2] a_14922_4138# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X5622 a_17934_17190# row_n[15] a_18426_17552# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5623 a_29374_15222# rowon_n[13] a_28978_15182# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X5624 vcm a_2275_13198# a_18026_13174# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5625 VSS row_n[10] a_26362_12210# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5626 vcm a_2275_2154# a_16018_2130# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5627 VDD rowon_n[3] a_25966_5142# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5628 a_7894_17190# row_n[15] a_8386_17552# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5629 vcm a_2275_13198# a_7986_13174# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5630 a_31078_11166# a_2475_11190# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5631 a_30378_10202# rowon_n[8] a_29982_10162# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X5632 VDD rowon_n[6] a_3878_8154# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5633 a_22042_13174# a_2475_13198# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5634 a_23046_7150# a_2475_7174# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5635 VDD rowon_n[12] a_24962_14178# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5636 a_13006_12170# a_2475_12194# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5637 a_35094_12170# a_2475_12194# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5638 a_2966_12170# a_2475_12194# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5639 a_23350_6186# col_n[20] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5640 VSS row_n[4] a_33390_6186# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5641 VDD rowon_n[2] a_14922_4138# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5642 VDD rowon_n[11] a_28978_13174# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5643 a_26458_10524# col_n[23] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X5644 a_29982_10162# a_2275_10186# a_30074_10162# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5645 a_6282_7190# rowon_n[5] a_5886_7150# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X5646 a_7286_3174# rowon_n[1] a_6890_3134# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X5647 vcm a_2275_6170# a_27062_6146# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5648 a_31382_18234# VDD a_30986_18194# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X5649 a_24354_17230# col_n[21] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5650 VDD rowon_n[4] a_8898_6146# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5651 a_28370_16226# col_n[25] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5652 VSS row_n[12] a_32386_14218# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5653 a_12306_5182# col_n[9] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5654 VDD rowon_n[0] a_27974_2130# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5655 a_28066_5142# a_2475_5166# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5656 a_19942_18194# a_2275_18218# a_20034_18194# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5657 a_32994_17190# a_2275_17214# a_33086_17190# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5658 VDD VSS a_6890_1126# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5659 VSS row_n[13] a_8290_15222# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5660 VSS row_n[13] a_18330_15222# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5661 a_23046_15182# a_2475_15206# a_22954_15182# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X5662 a_27062_14178# a_2475_14202# a_26970_14178# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X5663 a_19334_11206# col_n[16] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5664 vcm a_2275_11190# a_24050_11166# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5665 a_13918_8154# row_n[6] a_14410_8516# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5666 VDD VSS sky130_fd_pr__cap_mim_m3_1 l=17.2 w=17.2
X5667 a_28370_4178# col_n[25] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5668 a_27462_18556# col_n[24] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X5669 VDD rowon_n[14] a_30986_16186# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5670 a_23958_15182# row_n[13] a_24450_15544# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5671 a_18026_13174# a_2475_13198# a_17934_13174# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X5672 a_9294_11206# col_n[6] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5673 a_7986_13174# a_2475_13198# a_7894_13174# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X5674 a_10906_13174# a_2275_13198# a_10998_13174# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5675 VDD rowon_n[15] a_6890_17190# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5676 VDD rowon_n[15] a_16930_17190# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5677 a_11910_3134# row_n[1] a_12402_3496# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5678 a_18426_13536# col_n[15] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X5679 a_8386_13536# col_n[5] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X5680 vcm a_2275_8178# a_30074_8154# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5681 a_16322_7190# col_n[13] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5682 a_17326_3174# col_n[14] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5683 vcm a_2275_4162# a_31078_4138# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5684 ctop sw ctop VDD sky130_fd_pr__pfet_01v8 ad=0.503 pd=4.33 as=0 ps=0 w=1.9 l=0.22
X5685 a_27974_4138# row_n[2] a_28466_4500# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5686 a_5886_7150# row_n[5] a_6378_7512# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5687 a_3970_4138# a_2475_4162# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5688 a_18938_6146# row_n[4] a_19430_6508# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5689 a_21038_7150# a_2475_7174# a_20946_7150# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X5690 a_32082_3134# a_2475_3158# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5691 vcm a_2275_15206# a_12002_15182# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5692 a_29070_11166# a_2475_11190# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5693 a_28370_10202# rowon_n[8] a_27974_10162# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X5694 a_20434_6508# col_n[17] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X5695 a_3878_2130# row_n[0] a_4370_2492# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5696 VDD rowon_n[4] a_29982_6146# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5697 a_16930_1126# VDD a_17422_1488# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5698 a_15926_18194# VDD a_16418_18556# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5699 a_27366_16226# rowon_n[14] a_26970_16186# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X5700 vcm a_2275_14202# a_5978_14178# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5701 vcm a_2275_14202# a_16018_14178# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5702 a_9994_10162# a_2475_10186# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5703 a_9294_2170# col_n[6] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5704 a_5886_18194# VDD a_6378_18556# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5705 vcm a_2275_6170# a_35094_6146# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5706 a_10906_2130# a_2275_2154# a_10998_2130# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5707 a_28978_15182# a_2275_15206# a_29070_15182# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5708 a_20034_14178# a_2475_14202# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5709 VSS VDD a_23350_1166# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5710 VSS row_n[3] a_22346_5182# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5711 a_10998_13174# a_2475_13198# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5712 a_33086_13174# a_2475_13198# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5713 a_32386_5182# rowon_n[3] a_31990_5142# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X5714 a_23350_12210# col_n[20] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5715 a_4882_4138# a_2275_4162# a_4974_4138# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5716 a_26058_5142# a_2475_5166# a_25966_5142# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X5717 a_24450_8516# col_n[21] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X5718 a_22346_18234# col_n[19] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5719 VDD rowon_n[6] a_33998_8154# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5720 a_2161_13198# sample VDD VDD sky130_fd_pr__pfet_01v8 ad=0.342 pd=2.97 as=0.342 ps=2.97 w=1.2 l=0.15
X5721 a_22442_14540# col_n[19] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X5722 VSS row_n[8] a_17326_10202# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5723 a_22042_10162# a_2475_10186# a_21950_10162# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X5724 VSS a_2161_8178# a_2275_8178# VSS sky130_fd_pr__nfet_01v8 ad=0.124 pd=1.01 as=0.171 ps=1.77 w=0.6 l=0.15
X5725 a_21950_6146# a_2275_6170# a_22042_6146# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5726 VDD rowon_n[1] a_31990_3134# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5727 a_22442_3496# col_n[19] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X5728 a_7894_11166# a_2275_11190# a_7986_11166# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5729 a_17934_11166# a_2275_11190# a_18026_11166# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5730 VSS row_n[8] a_7286_10202# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5731 a_30986_18194# a_2275_18218# a_31078_18194# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5732 VSS row_n[14] a_16322_16226# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5733 a_21038_16186# a_2475_16210# a_20946_16186# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X5734 a_22954_10162# row_n[8] a_23446_10524# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5735 VSS row_n[1] a_27366_3174# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5736 VSS row_n[14] a_6282_16226# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5737 a_19334_9198# rowon_n[7] a_18938_9158# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X5738 a_31382_9198# col_n[28] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5739 a_13406_7512# col_n[10] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X5740 VSS row_n[4] a_5278_6186# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5741 a_21950_16186# row_n[14] a_22442_16548# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5742 VDD rowon_n[10] a_15926_12170# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5743 VSS row_n[7] a_17326_9198# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5744 a_1957_15206# VDD sample VSS sky130_fd_pr__nfet_01v8 ad=0.171 pd=1.77 as=0.171 ps=1.77 w=0.6 l=0.15
X5745 a_16018_14178# a_2475_14202# a_15926_14178# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X5746 VDD rowon_n[10] a_5886_12170# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5747 a_29470_6508# col_n[26] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X5748 a_11398_2492# col_n[8] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X5749 VDD VDD a_14922_18194# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5750 a_5978_14178# a_2475_14202# a_5886_14178# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X5751 VDD VDD a_4882_18194# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5752 a_15318_15222# col_n[12] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5753 vcm a_2275_15206# a_20034_15182# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5754 a_7986_9158# a_2475_9182# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5755 VSS row_n[0] a_16322_2170# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5756 a_30074_3134# a_2475_3158# a_29982_3134# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X5757 vcm a_2275_3158# a_20034_3134# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5758 a_14010_17190# a_2475_17214# a_13918_17190# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X5759 a_5278_15222# col_n[2] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5760 a_25966_8154# a_2275_8178# a_26058_8154# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5761 a_27462_1488# col_n[24] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X5762 a_26970_4138# a_2275_4162# a_27062_4138# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5763 a_3970_17190# a_2475_17214# a_3878_17190# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X5764 vcm a_2275_9182# a_9994_9158# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5765 VDD rowon_n[7] a_18938_9158# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5766 a_30986_9158# row_n[7] a_31478_9520# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5767 a_31990_5142# row_n[3] a_32482_5504# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5768 a_14410_17552# col_n[11] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X5769 a_10906_14178# row_n[12] a_11398_14540# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5770 vcm a_2275_10186# a_10998_10162# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5771 a_17422_9520# col_n[14] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X5772 VSS row_n[6] a_9294_8194# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5773 a_18426_5504# col_n[15] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X5774 a_4370_17552# col_n[1] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X5775 a_22346_12210# rowon_n[10] a_21950_12170# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X5776 a_14922_13174# row_n[11] a_15414_13536# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5777 a_26362_11206# rowon_n[9] a_25966_11166# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X5778 a_4882_13174# row_n[11] a_5374_13536# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5779 a_18026_11166# a_2475_11190# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5780 vcm a_2275_1150# a_25054_1126# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5781 a_35094_1126# a_2475_1150# a_35002_1126# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X5782 a_1957_16210# VSS sample VDD sky130_fd_pr__pfet_01v8 ad=0.342 pd=2.97 as=0.342 ps=2.97 w=1.2 l=0.15
X5783 a_7986_11166# a_2475_11190# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5784 a_1957_6170# VDD sample VSS sky130_fd_pr__nfet_01v8 ad=0.171 pd=1.77 as=0.171 ps=1.77 w=0.6 l=0.15
X5785 vcm a_2275_4162# a_2966_4138# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5786 a_34090_5142# a_2475_5166# a_33998_5142# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X5787 VDD rowon_n[8] a_21950_10162# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5788 a_8898_9158# a_2275_9182# a_8990_9158# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5789 a_17022_2130# a_2475_2154# a_16930_2130# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X5790 VSS row_n[15] a_20338_17230# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5791 a_26970_16186# a_2275_16210# a_27062_16186# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5792 a_31078_14178# a_2475_14202# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5793 a_12306_6186# rowon_n[4] a_11910_6146# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X5794 a_29982_6146# a_2275_6170# a_30074_6146# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5795 VDD rowon_n[5] a_22954_7150# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5796 a_33998_2130# row_n[0] a_34490_2492# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5797 VSS row_n[14] a_24354_16226# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5798 a_21342_13214# col_n[18] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5799 a_34394_12210# col_n[31] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5800 a_14314_15222# rowon_n[13] a_13918_15182# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X5801 VSS row_n[10] a_11302_12210# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5802 VDD rowon_n[0] a_20946_2130# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5803 a_21038_5142# a_2475_5166# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5804 a_19030_16186# a_2475_16210# a_18938_16186# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X5805 a_4274_15222# rowon_n[13] a_3878_15182# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X5806 a_29982_13174# a_2275_13198# a_30074_13174# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5807 VDD VDD a_22954_18194# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5808 a_20434_15544# col_n[17] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X5809 a_8290_14218# rowon_n[12] a_7894_14178# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X5810 a_33486_14540# col_n[30] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X5811 vcm a_2275_12194# a_29070_12170# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5812 VSS row_n[9] a_5278_11206# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5813 VSS row_n[9] a_15318_11206# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5814 a_20034_11166# a_2475_11190# a_19942_11166# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X5815 a_33086_10162# a_2475_10186# a_32994_10162# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X5816 a_20338_8194# col_n[17] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5817 a_26362_2170# rowon_n[0] a_25966_2130# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X5818 a_21342_4178# col_n[18] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5819 a_20946_11166# row_n[9] a_21438_11528# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5820 a_10998_10162# a_2475_10186# a_10906_10162# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X5821 a_5978_9158# a_2475_9182# a_5886_9158# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X5822 VSS row_n[6] a_30378_8194# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5823 a_4274_5182# rowon_n[3] a_3878_5142# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X5824 a_5278_1166# VSS a_4882_1126# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X5825 VSS row_n[2] a_31382_4178# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5826 VDD rowon_n[12] a_9902_14178# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5827 a_33998_10162# row_n[8] a_34490_10524# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5828 a_35002_4138# a_2275_4162# a_35094_4138# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5829 a_17326_4178# rowon_n[2] a_16930_4138# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X5830 a_16322_8194# rowon_n[6] a_15926_8154# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X5831 vcm a_2275_8178# a_24050_8154# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5832 vcm a_2275_2154# a_18026_2130# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5833 VDD rowon_n[3] a_27974_5142# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5834 VDD rowon_n[11] a_3878_13174# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5835 VDD rowon_n[11] a_13918_13174# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5836 a_11398_10524# col_n[8] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X5837 VDD rowon_n[6] a_5886_8154# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5838 a_25054_7150# a_2475_7174# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5839 a_26058_3134# a_2475_3158# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5840 a_13310_16226# col_n[10] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5841 VDD rowon_n[1] a_3878_3134# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5842 a_31478_4500# col_n[28] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X5843 a_20946_4138# row_n[2] a_21438_4500# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5844 a_12002_18194# a_2475_18218# a_11910_18194# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X5845 a_34090_18194# a_2475_18218# a_33998_18194# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X5846 a_3270_16226# col_n[0] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5847 vcm a_2275_15206# a_31078_15182# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5848 a_25358_6186# col_n[22] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5849 a_35002_18194# VDD a_35494_18556# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5850 vcm a_2275_14202# a_35094_14178# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5851 a_3270_9198# col_n[0] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5852 a_11910_6146# row_n[4] a_12402_6508# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5853 VSS row_n[4] a_35398_6186# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5854 a_9294_3174# rowon_n[1] a_8898_3134# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X5855 VDD rowon_n[2] a_16930_4138# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5856 a_8290_7190# rowon_n[5] a_7894_7150# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X5857 a_12402_18556# col_n[9] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X5858 a_19334_18234# VDD a_18938_18194# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X5859 a_20338_13214# rowon_n[11] a_19942_13174# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X5860 vcm a_2275_6170# a_29070_6146# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5861 vcm a_2275_9182# a_6982_9158# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5862 a_25054_15182# a_2475_15206# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5863 a_21950_12170# a_2275_12194# a_22042_12170# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5864 a_14314_5182# col_n[11] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5865 VDD VSS a_8898_1126# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5866 a_29070_14178# a_2475_14202# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5867 a_2874_9158# row_n[7] a_3366_9520# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5868 a_3878_5142# row_n[3] a_4370_5504# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5869 a_19942_1126# a_2275_1150# a_20034_1126# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5870 VDD rowon_n[14] a_18938_16186# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5871 VDD rowon_n[9] a_19942_11166# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5872 a_15926_8154# row_n[6] a_16418_8516# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5873 a_30074_1126# a_2475_1150# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5874 a_9994_13174# a_2475_13198# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5875 VSS row_n[15] a_31382_17230# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5876 a_2475_10186# a_1957_10186# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.342 pd=2.97 as=0.249 ps=1.62 w=1.2 l=0.15
X5877 a_13918_3134# row_n[1] a_14410_3496# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5878 a_13310_10202# rowon_n[8] a_12914_10162# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X5879 a_12002_2130# a_2475_2154# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5880 VSS row_n[14] a_35398_16226# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5881 a_32386_13214# col_n[29] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5882 a_3270_10202# rowon_n[8] a_2874_10162# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X5883 a_18330_7190# col_n[15] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5884 a_19334_3174# col_n[16] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5885 vcm a_2275_4162# a_33086_4138# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5886 a_26058_17190# a_2475_17214# a_25966_17190# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X5887 a_12306_16226# rowon_n[14] a_11910_16186# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X5888 VSS row_n[1] a_20338_3174# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5889 a_7894_7150# row_n[5] a_8386_7512# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5890 a_30378_3174# rowon_n[1] a_29982_3134# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X5891 VDD VDD a_33998_18194# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5892 a_26970_17190# row_n[15] a_27462_17552# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5893 a_31478_15544# col_n[28] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X5894 vcm a_2275_13198# a_27062_13174# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5895 a_31078_11166# a_2475_11190# a_30986_11166# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X5896 a_34090_3134# a_2475_3158# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5897 a_3878_15182# a_2275_15206# a_3970_15182# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5898 a_13918_15182# a_2275_15206# a_14010_15182# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5899 VSS row_n[7] a_10298_9198# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5900 a_23046_7150# a_2475_7174# a_22954_7150# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X5901 a_22442_6508# col_n[19] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X5902 a_5886_2130# row_n[0] a_6378_2492# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5903 a_17934_14178# a_2275_14202# a_18026_14178# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5904 a_31990_11166# row_n[9] a_32482_11528# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5905 VDD rowon_n[4] a_31990_6146# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5906 a_18938_1126# en_bit_n[2] a_19430_1488# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5907 a_7894_14178# a_2275_14202# a_7986_14178# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5908 a_20434_1488# en_bit_n[0] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X5909 a_29982_14178# row_n[12] a_30474_14540# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5910 vcm a_2275_10186# a_30074_10162# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5911 VDD VSS a_29982_1126# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5912 a_12914_2130# a_2275_2154# a_13006_2130# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5913 VSS VDD a_25358_1166# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5914 VSS row_n[3] a_24354_5182# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5915 a_10394_9520# col_n[7] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X5916 a_11398_5504# col_n[8] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X5917 a_35398_1166# VSS a_35002_1126# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X5918 VSS row_n[2] a_3270_4178# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5919 a_34394_5182# rowon_n[3] a_33998_5142# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X5920 a_18330_13214# rowon_n[11] a_17934_13174# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X5921 a_28978_10162# a_2275_10186# a_29070_10162# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5922 a_28066_5142# a_2475_5166# a_27974_5142# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X5923 vcm a_2275_16210# a_8990_16186# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5924 vcm a_2275_16210# a_19030_16186# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5925 a_23958_6146# a_2275_6170# a_24050_6146# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5926 a_24450_3496# col_n[21] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X5927 VDD rowon_n[1] a_33998_3134# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5928 a_23046_16186# a_2475_16210# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5929 VDD rowon_n[9] a_17934_11166# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5930 VSS row_n[1] a_29374_3174# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5931 a_3366_4500# col_n[0] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X5932 a_33390_9198# col_n[30] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5933 a_15414_7512# col_n[12] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X5934 VSS row_n[15] a_29374_17230# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5935 a_33390_15222# rowon_n[13] a_32994_15182# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X5936 VSS row_n[10] a_30378_12210# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5937 a_16018_7150# a_2475_7174# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5938 VSS row_n[4] a_7286_6186# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5939 a_7986_14178# a_2475_14202# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5940 a_18026_14178# a_2475_14202# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5941 VSS row_n[9] a_34394_11206# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5942 a_32386_2170# col_n[29] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5943 a_2161_1150# sample VDD VDD sky130_fd_pr__pfet_01v8 ad=0.342 pd=2.97 as=0.342 ps=2.97 w=1.2 l=0.15
X5944 a_13406_2492# col_n[10] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X5945 a_3970_4138# a_2475_4162# a_3878_4138# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X5946 a_9994_9158# a_2475_9182# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5947 a_25054_12170# a_2475_12194# a_24962_12170# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X5948 a_11302_11206# rowon_n[9] a_10906_11166# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X5949 a_1957_10186# VDD sample VSS sky130_fd_pr__nfet_01v8 ad=0.171 pd=1.77 as=0.171 ps=1.77 w=0.6 l=0.15
X5950 a_27974_8154# a_2275_8178# a_28066_8154# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5951 a_29470_1488# col_n[26] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X5952 VSS row_n[0] a_18330_2170# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5953 a_32082_3134# a_2475_3158# a_31990_3134# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X5954 a_28978_4138# a_2275_4162# a_29070_4138# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5955 a_29470_15544# col_n[26] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X5956 VDD rowon_n[11] a_32994_13174# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5957 a_25966_12170# row_n[10] a_26458_12532# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5958 a_29070_11166# a_2475_11190# a_28978_11166# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X5959 a_30474_10524# col_n[27] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X5960 a_32994_9158# row_n[7] a_33486_9520# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5961 a_33998_5142# row_n[3] a_34490_5504# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5962 a_9994_10162# a_2475_10186# a_9902_10162# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X5963 a_10298_4178# rowon_n[2] a_9902_4138# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X5964 a_11910_16186# a_2275_16210# a_12002_16186# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5965 VDD rowon_n[12] a_8898_14178# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5966 vcm a_2275_2154# a_10998_2130# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5967 VDD rowon_n[3] a_20946_5142# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5968 a_16930_7150# a_2275_7174# a_17022_7150# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5969 vcm a_2275_17214# a_23046_17190# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5970 a_8290_17230# col_n[5] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5971 a_18330_17230# col_n[15] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5972 vcm a_2275_4162# a_4974_4138# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5973 VDD rowon_n[2] a_9902_4138# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5974 vcm a_2275_12194# a_14010_12170# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5975 vcm a_2275_12194# a_3970_12170# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5976 a_14314_6186# rowon_n[4] a_13918_6146# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X5977 vcm a_2275_6170# a_22042_6146# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5978 a_17934_15182# row_n[13] a_18426_15544# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5979 a_29374_13214# rowon_n[11] a_28978_13174# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X5980 vcm a_2275_11190# a_18026_11166# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5981 VSS row_n[8] a_26362_10202# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5982 a_7894_15182# row_n[13] a_8386_15544# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5983 vcm a_2275_11190# a_7986_11166# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5984 a_26970_11166# a_2275_11190# a_27062_11166# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X5985 VDD rowon_n[4] a_3878_6146# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5986 VDD rowon_n[0] a_22954_2130# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5987 a_23046_5142# a_2475_5166# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5988 VDD rowon_n[10] a_24962_12170# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5989 a_28370_2170# rowon_n[0] a_27974_2130# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X5990 VSS row_n[2] a_33390_4178# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5991 a_23350_4178# col_n[20] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5992 VDD rowon_n[9] a_28978_11166# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X5993 a_7986_9158# a_2475_9182# a_7894_9158# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X5994 VSS row_n[6] a_32386_8194# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5995 a_6282_5182# rowon_n[3] a_5886_5142# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X5996 a_7286_1166# VSS a_6890_1126# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X5997 VSS a_2161_18218# a_2275_18218# VSS sky130_fd_pr__nfet_01v8 ad=0.124 pd=1.01 as=0.171 ps=1.77 w=0.6 l=0.15
X5998 vcm a_2275_8178# a_26058_8154# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5999 vcm a_2275_4162# a_27062_4138# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X6000 VSS VDD a_27366_18234# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X6001 a_31382_16226# rowon_n[14] a_30986_16186# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X6002 a_24354_15222# col_n[21] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X6003 VDD rowon_n[6] a_7894_8154# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X6004 a_2475_6170# a_1957_6170# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.171 pd=1.77 as=0.124 ps=1.01 w=0.6 l=0.15
X6005 a_17326_17230# rowon_n[15] a_16930_17190# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X6006 a_28370_14218# col_n[25] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X6007 a_11302_7190# col_n[8] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X6008 a_28066_3134# a_2475_3158# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X6009 a_12306_3174# col_n[9] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X6010 a_7286_17230# rowon_n[15] a_6890_17190# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X6011 a_19942_16186# a_2275_16210# a_20034_16186# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X6012 a_32994_15182# a_2275_15206# a_33086_15182# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X6013 a_31990_9158# a_2275_9182# a_32082_9158# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X6014 a_27062_7150# a_2475_7174# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X6015 a_22954_4138# row_n[2] a_23446_4500# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X6016 a_3970_18194# a_2475_18218# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X6017 a_14010_18194# a_2475_18218# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X6018 a_23446_17552# col_n[20] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X6019 VSS row_n[11] a_8290_13214# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X6020 VSS row_n[11] a_18330_13214# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X6021 a_23046_13174# a_2475_13198# a_22954_13174# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X6022 VDD rowon_n[1] a_5886_3134# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X6023 a_33486_4500# col_n[30] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X6024 a_13918_6146# row_n[4] a_14410_6508# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X6025 a_27462_16548# col_n[24] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X6026 a_23958_13174# row_n[11] a_24450_13536# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X6027 a_18026_11166# a_2475_11190# a_17934_11166# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X6028 a_5278_9198# col_n[2] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X6029 a_7986_11166# a_2475_11190# a_7894_11166# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X6030 VDD rowon_n[13] a_6890_15182# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X6031 VDD rowon_n[13] a_16930_15182# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X6032 vcm a_2275_9182# a_8990_9158# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X6033 a_11910_1126# VDD a_12402_1488# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X6034 a_18426_11528# col_n[15] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X6035 a_4274_2170# col_n[1] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X6036 a_8386_11528# col_n[5] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X6037 vcm a_2275_6170# a_30074_6146# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X6038 a_16322_5182# col_n[13] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X6039 a_17326_1166# col_n[14] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X6040 a_16322_18234# col_n[13] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X6041 vcm a_2275_18218# a_21038_18194# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X6042 a_6282_18234# col_n[3] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X6043 vcm a_2275_17214# a_34090_17190# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X6044 a_5886_5142# row_n[3] a_6378_5504# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X6045 a_4882_9158# row_n[7] a_5374_9520# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X6046 a_17934_8154# row_n[6] a_18426_8516# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X6047 a_25054_10162# a_2475_10186# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X6048 a_32082_1126# a_2475_1150# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X6049 a_21038_5142# a_2475_5166# a_20946_5142# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X6050 a_11910_17190# row_n[15] a_12402_17552# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X6051 vcm a_2275_13198# a_12002_13174# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X6052 a_14010_2130# a_2475_2154# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X6053 a_15926_3134# row_n[1] a_16418_3496# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X6054 a_5886_16186# row_n[14] a_6378_16548# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X6055 a_15926_16186# row_n[14] a_16418_16548# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X6056 a_27366_14218# rowon_n[12] a_26970_14178# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X6057 a_27366_9198# col_n[24] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X6058 vcm a_2275_4162# a_35094_4138# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X6059 a_28066_17190# a_2475_17214# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X6060 a_28978_13174# a_2275_13198# a_29070_13174# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X6061 VSS row_n[1] a_22346_3174# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X6062 a_31382_7190# rowon_n[5] a_30986_7150# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X6063 a_32386_3174# rowon_n[1] a_31990_3134# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X6064 a_23350_10202# col_n[20] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X6065 VSS row_n[7] a_12306_9198# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X6066 a_26058_3134# a_2475_3158# a_25966_3134# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X6067 a_25054_7150# a_2475_7174# a_24962_7150# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X6068 a_24450_6508# col_n[21] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X6069 a_7894_2130# row_n[0] a_8386_2492# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X6070 a_22346_16226# col_n[19] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X6071 a_16322_12210# rowon_n[10] a_15926_12170# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X6072 a_26970_9158# row_n[7] a_27462_9520# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X6073 VDD rowon_n[4] a_33998_6146# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X6074 a_6282_12210# rowon_n[10] a_5886_12170# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X6075 a_2161_11190# sample VDD VDD sky130_fd_pr__pfet_01v8 ad=0.342 pd=2.97 as=0.342 ps=2.97 w=1.2 l=0.15
X6076 a_13918_10162# a_2275_10186# a_14010_10162# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X6077 a_2966_9158# a_2475_9182# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X6078 VSS row_n[0] a_11302_2170# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X6079 a_22442_12532# col_n[19] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X6080 a_3878_10162# a_2275_10186# a_3970_10162# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X6081 a_20946_8154# a_2275_8178# a_21038_8154# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X6082 a_22442_1488# col_n[19] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X6083 VDD VSS a_31990_1126# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X6084 a_21950_4138# a_2275_4162# a_22042_4138# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X6085 a_5278_18234# VDD a_4882_18194# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X6086 a_15318_18234# VDD a_14922_18194# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X6087 a_31078_8154# a_2475_8178# vcm VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X6088 a_14922_2130# a_2275_2154# a_15014_2130# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X6089 a_21438_18556# col_n[18] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X6090 a_30986_16186# a_2275_16210# a_31078_16186# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X6091 VSS row_n[12] a_16322_14218# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X6092 a_21038_14178# a_2475_14202# a_20946_14178# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X6093 VSS VDD a_27366_1166# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X6094 VSS row_n[12] a_6282_14218# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X6095 a_12402_9520# col_n[9] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X6096 VSS row_n[6] a_4274_8194# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X6097 a_13406_5504# col_n[10] VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X6098 VSS row_n[2] a_5278_4178# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X6099 a_16930_17190# a_2275_17214# a_17022_17190# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X6100 VDD rowon_n[8] a_15926_10162# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X6101 a_6890_17190# a_2275_17214# a_6982_17190# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X6102 VDD rowon_n[8] a_5886_10162# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X6103 VSS row_n[15] a_4274_17230# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X6104 VSS row_n[15] a_14314_17230# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X6105 VDD rowon_n[14] a_14922_16186# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X6106 VDD rowon_n[14] a_4882_16186# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X6107 a_15318_13214# col_n[12] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X6108 vcm a_2275_13198# a_20034_13174# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X6109 vcm a_2275_1150# a_20034_1126# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X6110 a_30074_1126# a_2475_1150# a_29982_1126# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X6111 a_19942_17190# row_n[15] a_20434_17552# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X6112 a_14010_15182# a_2475_15206# a_13918_15182# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X6113 a_5278_13214# col_n[2] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X6114 vcm a_2275_12194# a_33086_12170# VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X6115 a_25966_6146# a_2275_6170# a_26058_6146# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
C0 row_n[14] a_20338_16226# 0.0117f
C1 a_3970_15182# a_3970_14178# 0.843f
C2 VDD a_24050_10162# 0.483f
C3 col_n[4] a_7382_2492# 0.0283f
C4 col_n[14] a_17422_14540# 0.0283f
C5 col[28] a_2475_13198# 0.136f
C6 row_n[4] a_30378_6186# 0.0117f
C7 a_26970_3134# a_27366_3174# 0.0313f
C8 vcm a_30074_5142# 0.56f
C9 a_2275_7174# a_6282_7190# 0.144f
C10 a_2475_7174# a_8898_7150# 0.264f
C11 rowoff_n[10] a_24050_12170# 0.294f
C12 rowoff_n[2] a_6982_4138# 0.294f
C13 row_n[6] a_20946_8154# 0.0437f
C14 a_2275_12194# a_31078_12170# 0.399f
C15 a_16930_12170# a_17422_12532# 0.0658f
C16 a_16018_12170# a_16322_12210# 0.0931f
C17 rowon_n[10] a_20034_12170# 0.248f
C18 rowon_n[15] col[6] 0.0323f
C19 rowon_n[4] rowon_n[3] 0.0632f
C20 rowon_n[12] col[0] 0.0318f
C21 row_n[14] col[3] 0.0342f
C22 rowon_n[14] col[4] 0.0323f
C23 rowon_n[9] ctop 0.203f
C24 row_n[13] col[1] 0.0342f
C25 rowon_n[13] col[2] 0.0323f
C26 row_n[15] col[5] 0.0342f
C27 col_n[5] rowoff_n[15] 0.0471f
C28 col_n[19] col[19] 0.489f
C29 row_n[0] m2_34288_2378# 0.0128f
C30 a_28066_17190# a_29070_17190# 0.843f
C31 VDD a_4974_13174# 0.483f
C32 col_n[28] a_31382_3174# 0.084f
C33 col_n[2] a_4974_2130# 0.251f
C34 col[8] rowoff_n[11] 0.0901f
C35 rowon_n[0] a_30074_2130# 0.248f
C36 rowoff_n[0] a_16018_2130# 0.294f
C37 col_n[12] a_15014_14178# 0.251f
C38 a_35002_5142# a_35398_5182# 0.0313f
C39 col_n[9] a_11910_4138# 0.0765f
C40 vcm a_10998_8154# 0.56f
C41 col[25] a_2275_16210# 0.0899f
C42 col_n[19] a_21950_16186# 0.0765f
C43 a_2275_9182# a_21342_9198# 0.144f
C44 a_2475_9182# a_23958_9158# 0.264f
C45 a_12914_9158# a_13006_9158# 0.326f
C46 col[30] a_2275_5166# 0.0899f
C47 row_n[0] a_7986_2130# 0.282f
C48 VDD a_20034_17190# 0.484f
C49 rowon_n[4] a_7894_6146# 0.118f
C50 col_n[3] a_6378_12532# 0.0283f
C51 vcm a_2275_2154# 6.51f
C52 a_7894_6146# a_8290_6186# 0.0313f
C53 a_2275_6170# a_14922_6146# 0.136f
C54 vcm a_26058_12170# 0.56f
C55 a_2966_11166# a_2966_10162# 0.843f
C56 col[29] a_31990_3134# 0.0682f
C57 VDD a_22954_2130# 0.181f
C58 m2_6176_9406# row_n[7] 0.0128f
C59 m2_12200_5390# row_n[3] 0.0128f
C60 ctop a_2966_6146# 4.06f
C61 col_n[15] a_2475_12194# 0.0531f
C62 a_31078_16186# a_31382_16226# 0.0931f
C63 row_n[11] a_28370_13214# 0.0117f
C64 a_31990_16186# a_32482_16548# 0.0658f
C65 col_n[20] a_2475_1150# 0.0531f
C66 a_3970_3134# a_4974_3134# 0.843f
C67 a_2475_3158# a_6982_3134# 0.316f
C68 rowoff_n[8] a_8898_10162# 0.202f
C69 col_n[17] a_20338_1166# 0.0572f
C70 row_n[13] a_18938_15182# 0.0437f
C71 vcm a_16322_6186# 0.155f
C72 col_n[1] a_3970_12170# 0.251f
C73 rowoff_n[11] a_12002_13174# 0.294f
C74 a_2275_8178# a_29982_8154# 0.136f
C75 col_n[27] a_30378_13214# 0.084f
C76 col[5] a_2475_9182# 0.136f
C77 vcm a_6982_15182# 0.56f
C78 col_n[8] a_10906_14178# 0.0765f
C79 a_27974_13174# a_28066_13174# 0.326f
C80 VDD a_3366_5504# 0.0779f
C81 row_n[3] a_28978_5142# 0.0437f
C82 rowon_n[7] a_28066_9158# 0.248f
C83 a_2275_17214# a_7986_17190# 0.399f
C84 m2_27260_14426# row_n[12] 0.0128f
C85 rowoff_n[6] a_17934_8154# 0.202f
C86 m2_33284_10410# row_n[8] 0.0128f
C87 col_n[12] a_2275_15206# 0.113f
C88 a_29070_6146# a_29070_5142# 0.843f
C89 a_2475_5166# a_22042_5142# 0.316f
C90 col_n[17] a_2275_4162# 0.113f
C91 vcm a_31382_10202# 0.155f
C92 rowoff_n[15] a_28066_17190# 0.294f
C93 a_22954_10162# a_23350_10202# 0.0313f
C94 m2_27260_16434# a_27062_16186# 0.165f
C95 rowoff_n[4] a_26970_6146# 0.202f
C96 ctop a_9994_4138# 4.11f
C97 m3_5880_1078# a_5978_2130# 0.0302f
C98 m2_9764_946# a_2475_1150# 0.286f
C99 col[21] a_24050_11166# 0.367f
C100 m2_4744_946# a_4882_1126# 0.225f
C101 row_n[7] a_5978_9158# 0.282f
C102 VDD a_18938_9158# 0.181f
C103 col[18] a_20946_1126# 0.0682f
C104 rowon_n[11] a_5886_13174# 0.118f
C105 col[28] a_30986_13174# 0.0682f
C106 col[2] a_2275_12194# 0.0899f
C107 VDD a_6282_18234# 0.019f
C108 col[7] a_2275_1150# 0.0899f
C109 a_2275_2154# a_13006_2130# 0.399f
C110 a_6982_2130# a_7286_2170# 0.0931f
C111 a_7894_2130# a_8386_2492# 0.0658f
C112 vcm a_24962_4138# 0.1f
C113 rowoff_n[9] a_18426_11528# 0.0133f
C114 rowon_n[1] a_15926_3134# 0.118f
C115 a_19030_7150# a_20034_7150# 0.843f
C116 col[28] a_2475_18218# 0.136f
C117 vcm a_12306_13214# 0.155f
C118 VDD a_10394_3496# 0.0779f
C119 col[22] a_2475_11190# 0.136f
C120 col_n[16] a_19334_11206# 0.084f
C121 m2_4744_18014# a_4974_18194# 0.0249f
C122 ctop a_25054_8154# 4.11f
C123 a_2275_16210# a_13310_16226# 0.144f
C124 a_2475_16210# a_15926_16186# 0.264f
C125 a_8898_16186# a_8990_16186# 0.326f
C126 VDD a_33998_13174# 0.181f
C127 a_23350_1166# m2_22816_946# 0.087f
C128 rowoff_n[7] a_27462_9520# 0.0133f
C129 col_n[27] a_30474_5504# 0.0283f
C130 a_2275_4162# a_28066_4138# 0.399f
C131 m3_33992_1078# ctop 0.355f
C132 col_n[29] a_2275_17214# 0.113f
C133 vcm a_5886_7150# 0.1f
C134 a_9994_9158# a_9994_8154# 0.843f
C135 rowoff_n[13] a_34490_15544# 0.0133f
C136 m2_18224_14426# a_18026_14178# 0.165f
C137 row_n[10] a_26970_12170# 0.0437f
C138 vcm a_27366_17230# 0.155f
C139 a_2275_13198# a_6890_13174# 0.136f
C140 rowon_n[14] a_26058_16186# 0.248f
C141 VDD a_25454_7512# 0.0779f
C142 ctop a_5978_11166# 4.11f
C143 a_2275_18218# a_28370_18234# 0.145f
C144 col[10] a_13006_9158# 0.367f
C145 VDD a_14922_16186# 0.181f
C146 col[19] a_2275_14202# 0.0899f
C147 a_2475_1150# a_20946_1126# 0.264f
C148 a_2275_1150# a_18330_1166# 0.126f
C149 m2_15212_2378# a_15014_2130# 0.165f
C150 col[24] a_2275_3158# 0.0899f
C151 col[17] a_19942_11166# 0.0682f
C152 a_22954_6146# a_23446_6508# 0.0658f
C153 a_22042_6146# a_22346_6186# 0.0931f
C154 m2_20808_946# m2_21812_946# 0.843f
C155 col_n[25] a_28066_5142# 0.251f
C156 vcm a_20946_11166# 0.1f
C157 a_33998_11166# a_34394_11206# 0.0313f
C158 row_n[14] a_3970_16186# 0.282f
C159 VDD a_17022_1126# 0.035f
C160 a_2275_15206# a_21950_15182# 0.136f
C161 VDD a_6378_10524# 0.0779f
C162 col_n[5] a_8290_9198# 0.084f
C163 ctop a_21038_15182# 4.11f
C164 row_n[4] a_14010_6146# 0.282f
C165 a_2275_3158# a_33390_3174# 0.144f
C166 a_18938_3134# a_19030_3134# 0.326f
C167 rowon_n[8] a_13918_10162# 0.118f
C168 rowoff_n[10] a_6378_12532# 0.0133f
C169 row_n[12] col[10] 0.0342f
C170 row_n[9] col[4] 0.0342f
C171 rowon_n[9] col[5] 0.0323f
C172 row_n[7] col[0] 0.0322f
C173 col_n[16] a_19430_3496# 0.0283f
C174 row_n[13] col[12] 0.0342f
C175 rowon_n[1] row_n[1] 18.9f
C176 rowon_n[15] col[17] 0.0323f
C177 col_n[16] rowoff_n[15] 0.0471f
C178 row_n[14] col[14] 0.0342f
C179 rowon_n[14] col[15] 0.0323f
C180 a_24354_1166# vcm 0.16f
C181 rowon_n[12] col[11] 0.0323f
C182 rowon_n[13] col[13] 0.0323f
C183 row_n[8] col[2] 0.0342f
C184 rowon_n[8] col[3] 0.0323f
C185 rowon_n[7] col[1] 0.0323f
C186 row_n[15] col[16] 0.0342f
C187 col_n[9] a_2475_10186# 0.0531f
C188 rowon_n[10] col[7] 0.0323f
C189 col_n[24] col[25] 7.13f
C190 rowon_n[11] col[9] 0.0323f
C191 row_n[10] col[6] 0.0342f
C192 row_n[4] ctop 0.186f
C193 row_n[11] col[8] 0.0342f
C194 m2_9188_12418# a_8990_12170# 0.165f
C195 row_n[6] a_2275_8178# 19.2f
C196 vcm a_34394_15222# 0.155f
C197 col_n[26] a_29470_15544# 0.0283f
C198 a_25054_13174# a_25054_12170# 0.843f
C199 m2_2160_4386# rowon_n[2] 0.0219f
C200 a_2475_12194# a_14010_12170# 0.316f
C201 VDD a_32082_5142# 0.483f
C202 rowon_n[10] a_1957_12194# 0.0172f
C203 col[19] rowoff_n[11] 0.0901f
C204 m2_22240_18442# VDD 0.0456f
C205 row_n[15] a_35398_17230# 0.0117f
C206 a_18938_17190# a_19334_17230# 0.0313f
C207 VDD a_21438_14540# 0.0779f
C208 m2_28264_8402# a_28066_8154# 0.165f
C209 col[6] a_8898_9158# 0.0682f
C210 a_3878_9158# a_3970_9158# 0.326f
C211 a_2874_9158# a_3270_9198# 0.0313f
C212 a_2275_9182# a_4974_9158# 0.399f
C213 rowoff_n[14] a_22442_16548# 0.0133f
C214 col_n[14] a_17022_3134# 0.251f
C215 vcm a_16930_18194# 0.101f
C216 a_2475_14202# a_29070_14178# 0.316f
C217 m2_11196_17438# rowon_n[15] 0.0322f
C218 a_15014_14178# a_16018_14178# 0.843f
C219 m2_17220_13422# rowon_n[11] 0.0322f
C220 row_n[7] a_35002_9158# 0.0437f
C221 VDD a_13006_8154# 0.483f
C222 m2_23244_9406# rowon_n[7] 0.0322f
C223 col_n[24] a_27062_15182# 0.251f
C224 m2_29268_5390# rowon_n[3] 0.0322f
C225 col_n[6] a_2275_13198# 0.113f
C226 col_n[21] a_23958_5142# 0.0765f
C227 m2_21812_946# vcm 0.353f
C228 rowon_n[11] a_34090_13174# 0.248f
C229 col_n[11] a_2275_2154# 0.113f
C230 VDD a_1957_17214# 0.196f
C231 col_n[31] a_33998_17190# 0.0765f
C232 vcm a_19030_3134# 0.56f
C233 a_33998_7150# a_34090_7150# 0.326f
C234 col[0] a_2966_17190# 0.367f
C235 col_n[26] a_2475_12194# 0.0531f
C236 a_2275_11190# a_20034_11166# 0.399f
C237 col[3] rowoff_n[12] 0.0901f
C238 col_n[5] a_8386_1488# 0.0283f
C239 col_n[31] a_2475_1150# 0.0971f
C240 m2_23820_18014# a_24050_18194# 0.0249f
C241 row_n[11] a_12002_13174# 0.282f
C242 col_n[15] a_18426_13536# 0.0283f
C243 a_5978_16186# a_5978_15182# 0.843f
C244 VDD a_28066_12170# 0.483f
C245 m2_16792_18014# m3_17928_18146# 0.0341f
C246 rowon_n[15] a_11910_17190# 0.118f
C247 a_28978_4138# a_29374_4178# 0.0313f
C248 row_n[1] a_22042_3134# 0.282f
C249 rowoff_n[1] a_7986_3134# 0.294f
C250 col[16] a_2475_9182# 0.136f
C251 m2_19228_6394# a_19030_6146# 0.165f
C252 vcm a_34090_7150# 0.56f
C253 rowon_n[5] a_21950_7150# 0.118f
C254 a_2475_8178# a_12914_8154# 0.264f
C255 a_2275_8178# a_10298_8194# 0.144f
C256 rowoff_n[12] a_28978_14178# 0.202f
C257 col_n[0] a_2874_9158# 0.0765f
C258 a_18026_13174# a_18330_13214# 0.0931f
C259 a_18938_13174# a_19430_13536# 0.0658f
C260 a_2275_13198# a_35094_13174# 0.0924f
C261 row_n[3] a_9294_5182# 0.0117f
C262 col_n[29] a_32386_2170# 0.084f
C263 VDD a_8990_15182# 0.483f
C264 col_n[23] a_2275_15206# 0.113f
C265 col_n[13] a_16018_13174# 0.251f
C266 col_n[28] a_2275_4162# 0.113f
C267 col_n[10] a_12914_3134# 0.0765f
C268 m3_2868_18146# a_2966_17190# 0.0303f
C269 col_n[20] a_22954_15182# 0.0765f
C270 a_2874_5142# a_2966_5142# 0.326f
C271 m2_20808_946# m3_20940_1078# 3.79f
C272 vcm a_15014_10162# 0.56f
C273 rowoff_n[15] a_10394_17552# 0.0133f
C274 m2_33860_18014# col[31] 0.347f
C275 a_2475_10186# a_27974_10162# 0.264f
C276 a_2275_10186# a_25358_10202# 0.144f
C277 a_14922_10162# a_15014_10162# 0.326f
C278 row_n[14] a_32994_16186# 0.0437f
C279 col[13] a_2275_12194# 0.0899f
C280 m2_10768_18014# ctop 0.0422f
C281 col[18] a_2275_1150# 0.0896f
C282 col_n[4] a_7382_11528# 0.0283f
C283 col_n[1] a_3878_1126# 0.0801f
C284 a_16018_3134# a_16018_2130# 0.843f
C285 m2_10192_4386# a_9994_4138# 0.165f
C286 m2_1732_2954# row_n[1] 0.292f
C287 vcm a_5278_4178# 0.155f
C288 a_9902_7150# a_10298_7190# 0.0313f
C289 a_2275_7174# a_18938_7150# 0.136f
C290 col[30] a_32994_2130# 0.0682f
C291 vcm a_30074_14178# 0.56f
C292 VDD a_26970_4138# 0.181f
C293 a_33086_17190# a_33390_17230# 0.0931f
C294 a_33998_17190# a_34490_17552# 0.0658f
C295 row_n[8] a_20034_10162# 0.282f
C296 rowoff_n[7] a_9902_9158# 0.202f
C297 col_n[3] a_2475_8178# 0.0531f
C298 rowon_n[12] a_19942_14178# 0.118f
C299 a_2475_4162# a_10998_4138# 0.316f
C300 a_5978_4138# a_6982_4138# 0.843f
C301 col_n[28] a_31382_12210# 0.084f
C302 m3_29976_18146# ctop 0.209f
C303 col_n[2] a_4974_11166# 0.251f
C304 m2_10192_16434# row_n[14] 0.0128f
C305 vcm a_20338_8194# 0.155f
C306 m2_16216_12418# row_n[10] 0.0128f
C307 rowoff_n[13] a_16930_15182# 0.202f
C308 m2_22240_8402# row_n[6] 0.0128f
C309 a_2275_9182# a_33998_9158# 0.136f
C310 col_n[9] a_11910_13174# 0.0765f
C311 m2_28264_4386# row_n[2] 0.0128f
C312 row_n[10] a_7286_12210# 0.0117f
C313 rowon_n[2] a_29982_4138# 0.118f
C314 ctop a_33086_3134# 4.11f
C315 vcm a_10998_17190# 0.56f
C316 a_29982_14178# a_30074_14178# 0.326f
C317 VDD a_7894_7150# 0.181f
C318 col[30] a_2275_14202# 0.0899f
C319 rowoff_n[5] a_18938_7150# 0.202f
C320 a_2275_18218# a_12002_18194# 0.0924f
C321 row_n[0] a_17326_2170# 0.0117f
C322 a_2475_1150# a_2275_1150# 2.68f
C323 a_1957_1150# a_2161_1150# 0.115f
C324 vcm a_13918_2130# 0.1f
C325 a_2475_6170# a_26058_6146# 0.316f
C326 a_31078_7150# a_31078_6146# 0.843f
C327 rowoff_n[3] a_27974_5142# 0.202f
C328 vcm a_2275_11190# 6.49f
C329 row_n[2] a_7894_4138# 0.0437f
C330 a_24962_11166# a_25358_11206# 0.0313f
C331 VDD a_33486_2492# 0.0779f
C332 col[22] a_25054_10162# 0.367f
C333 rowon_n[6] a_6982_8154# 0.248f
C334 ctop a_14010_6146# 4.11f
C335 a_2874_15182# a_3366_15544# 0.0658f
C336 a_2475_15206# a_4882_15182# 0.264f
C337 a_2275_15206# a_3878_15182# 0.136f
C338 VDD a_22954_11166# 0.181f
C339 col[29] a_31990_12170# 0.0682f
C340 ctop a_2966_15182# 4.06f
C341 row_n[7] col[11] 0.0342f
C342 row_n[13] col[23] 0.0342f
C343 rowon_n[12] col[22] 0.0323f
C344 row_n[9] col[15] 0.0342f
C345 row_n[5] col[7] 0.0342f
C346 col_n[27] rowoff_n[15] 0.0471f
C347 row_n[15] col[27] 0.0342f
C348 rowon_n[11] col[20] 0.0323f
C349 rowon_n[10] col[18] 0.0323f
C350 rowon_n[5] col[8] 0.0323f
C351 row_n[10] col[17] 0.0342f
C352 a_2275_3158# a_17022_3134# 0.399f
C353 rowon_n[13] col[24] 0.0323f
C354 row_n[4] col[5] 0.0342f
C355 rowon_n[7] col[12] 0.0323f
C356 rowon_n[4] col[6] 0.0323f
C357 row_n[8] col[13] 0.0342f
C358 rowon_n[3] col[4] 0.0323f
C359 col_n[30] col[30] 0.621f
C360 row_n[12] col[21] 0.0342f
C361 rowon_n[8] col[14] 0.0323f
C362 row_n[3] col[3] 0.0342f
C363 col_n[20] a_2475_10186# 0.0531f
C364 row_n[11] col[19] 0.0342f
C365 a_9902_3134# a_10394_3496# 0.0658f
C366 row_n[6] col[9] 0.0342f
C367 rowon_n[6] col[10] 0.0323f
C368 rowon_n[15] col[28] 0.0323f
C369 row_n[14] col[25] 0.0342f
C370 row_n[2] col[1] 0.0342f
C371 a_8990_3134# a_9294_3174# 0.0931f
C372 rowon_n[2] col[2] 0.0323f
C373 rowon_n[14] col[26] 0.0323f
C374 rowon_n[9] col[16] 0.0323f
C375 rowon_n[1] col[0] 0.0318f
C376 a_2475_18218# a_9994_18194# 0.0299f
C377 rowoff_n[8] a_19430_10524# 0.0133f
C378 a_30986_1126# a_2275_1150# 0.136f
C379 vcm a_28978_6146# 0.1f
C380 a_21038_8154# a_22042_8154# 0.843f
C381 col_n[17] a_20338_10202# 0.084f
C382 col[30] rowoff_n[11] 0.0901f
C383 vcm a_16322_15222# 0.155f
C384 VDD a_14410_5504# 0.0779f
C385 a_26362_1166# VDD 0.0149f
C386 ctop a_29070_10162# 4.11f
C387 row_n[15] a_18026_17190# 0.282f
C388 a_2475_17214# a_19942_17190# 0.264f
C389 a_10906_17190# a_10998_17190# 0.326f
C390 a_2275_17214# a_17326_17230# 0.144f
C391 col[10] a_2475_7174# 0.136f
C392 rowoff_n[6] a_28466_8516# 0.0133f
C393 VDD a_3366_14540# 0.0779f
C394 col_n[28] a_31478_4500# 0.0283f
C395 m3_25960_18146# a_26058_17190# 0.0303f
C396 row_n[5] a_28066_7150# 0.282f
C397 a_2275_5166# a_32082_5142# 0.399f
C398 rowon_n[9] a_27974_11166# 0.118f
C399 vcm a_9902_9158# 0.1f
C400 a_30986_1126# a_31478_1488# 0.0658f
C401 a_12002_10162# a_12002_9158# 0.843f
C402 rowoff_n[14] a_4882_16186# 0.202f
C403 col_n[17] a_2275_13198# 0.113f
C404 m2_34864_16006# a_35398_16226# 0.087f
C405 a_5886_14178# a_6282_14218# 0.0313f
C406 a_2275_14202# a_10906_14178# 0.136f
C407 col_n[22] a_2275_2154# 0.113f
C408 m2_32856_946# a_2475_1150# 0.284f
C409 VDD a_29470_9520# 0.0779f
C410 row_n[7] a_15318_9198# 0.0117f
C411 col[11] a_14010_8154# 0.367f
C412 ctop a_9994_13174# 4.11f
C413 VDD a_18938_18194# 0.343f
C414 col[18] a_20946_10162# 0.0682f
C415 a_2275_2154# a_22346_2170# 0.144f
C416 a_2475_2154# a_24962_2130# 0.264f
C417 m2_25828_946# VDD 1f
C418 row_n[9] a_5886_11166# 0.0437f
C419 col_n[26] a_29070_4138# 0.251f
C420 m2_1732_8978# m2_1732_7974# 0.843f
C421 col[14] rowoff_n[12] 0.0901f
C422 col[7] a_2275_10186# 0.0899f
C423 a_24050_7150# a_24354_7190# 0.0931f
C424 a_24962_7150# a_25454_7512# 0.0658f
C425 rowoff_n[9] a_29070_11166# 0.294f
C426 rowon_n[13] a_4974_15182# 0.248f
C427 vcm a_24962_13174# 0.1f
C428 a_2475_11190# a_2874_11166# 0.264f
C429 a_1957_11190# a_2275_11190# 0.158f
C430 VDD a_21038_3134# 0.483f
C431 m2_10768_18014# a_11302_18234# 0.087f
C432 m2_30848_18014# a_2275_18218# 0.28f
C433 col_n[6] a_9294_8194# 0.084f
C434 a_2275_16210# a_25966_16186# 0.136f
C435 rowon_n[3] a_15014_5142# 0.248f
C436 VDD a_10394_12532# 0.0779f
C437 ctop a_25054_17190# 4.06f
C438 col[27] a_2475_9182# 0.136f
C439 a_20946_4138# a_21038_4138# 0.326f
C440 col_n[17] a_20434_2492# 0.0283f
C441 rowon_n[5] a_3878_7150# 0.118f
C442 col_n[27] a_30474_14540# 0.0283f
C443 vcm a_5886_16186# 0.1f
C444 a_27062_14178# a_27062_13174# 0.843f
C445 a_2475_13198# a_18026_13174# 0.316f
C446 VDD a_2475_6170# 26.1f
C447 a_20946_18194# a_21342_18234# 0.0313f
C448 m2_26832_18014# a_2475_18218# 0.286f
C449 VDD a_25454_16548# 0.0779f
C450 a_15926_1126# a_16322_1166# 0.0313f
C451 col[0] a_2874_6146# 0.0682f
C452 row_n[12] a_26058_14178# 0.282f
C453 vcm a_7986_1126# 0.165f
C454 m2_6176_11414# rowon_n[9] 0.0322f
C455 col[7] a_9902_8154# 0.0682f
C456 m2_12200_7398# rowon_n[5] 0.0322f
C457 m2_31852_946# m2_32280_1374# 0.165f
C458 m2_18224_3382# rowon_n[1] 0.0322f
C459 col[24] a_2275_12194# 0.0899f
C460 a_4974_10162# a_5278_10202# 0.0931f
C461 a_2275_10186# a_8990_10162# 0.399f
C462 a_5886_10162# a_6378_10524# 0.0658f
C463 col_n[15] a_18026_2130# 0.25f
C464 col[29] a_2275_1150# 0.0899f
C465 row_n[14] a_13310_16226# 0.0117f
C466 m2_33284_17438# a_33086_17190# 0.165f
C467 col_n[25] a_28066_14178# 0.251f
C468 col_n[22] a_24962_4138# 0.0765f
C469 a_17022_15182# a_18026_15182# 0.843f
C470 a_2475_15206# a_33086_15182# 0.316f
C471 VDD a_17022_10162# 0.483f
C472 row_n[4] a_23350_6186# 0.0117f
C473 m2_1732_2954# col[0] 0.0137f
C474 col_n[5] a_8290_18234# 0.084f
C475 vcm a_23046_5142# 0.56f
C476 rowoff_n[10] a_17022_12170# 0.294f
C477 m2_27260_16434# rowon_n[14] 0.0322f
C478 m2_33284_12418# rowon_n[10] 0.0322f
C479 row_n[6] a_13918_8154# 0.0437f
C480 a_2275_12194# a_24050_12170# 0.399f
C481 rowon_n[10] a_13006_12170# 0.248f
C482 col_n[16] a_19430_12532# 0.0283f
C483 col_n[14] a_2475_8178# 0.0531f
C484 a_7986_17190# a_7986_16186# 0.843f
C485 VDD a_32082_14178# 0.483f
C486 row_n[8] a_1957_10186# 0.187f
C487 rowoff_n[0] a_8990_2130# 0.294f
C488 rowon_n[0] a_23046_2130# 0.248f
C489 a_30986_5142# a_31382_5182# 0.0313f
C490 m2_12776_946# ctop 0.0428f
C491 m2_1732_6970# a_2161_7174# 0.0454f
C492 vcm a_3970_8154# 0.56f
C493 a_2475_9182# a_16930_9158# 0.264f
C494 rowoff_n[14] a_33086_16186# 0.294f
C495 a_2275_9182# a_14314_9198# 0.144f
C496 col[4] a_2475_5166# 0.136f
C497 m2_24248_15430# a_24050_15182# 0.165f
C498 col[6] a_8898_18194# 0.0682f
C499 a_20034_14178# a_20338_14218# 0.0931f
C500 a_20946_14178# a_21438_14540# 0.0658f
C501 m2_34864_12994# ctop 0.0422f
C502 col_n[14] a_17022_12170# 0.251f
C503 VDD a_13006_17190# 0.484f
C504 col_n[11] a_13918_2130# 0.0765f
C505 a_27062_2130# a_28066_2130# 0.843f
C506 col_n[21] a_23958_14178# 0.0765f
C507 m3_28972_1078# VDD 0.0157f
C508 col_n[11] a_2275_11190# 0.113f
C509 vcm a_28370_3174# 0.155f
C510 row_n[9] a_34090_11166# 0.282f
C511 a_2275_6170# a_7894_6146# 0.136f
C512 rowon_n[13] a_33998_15182# 0.118f
C513 m2_34864_9982# a_2475_10186# 0.282f
C514 vcm a_19030_12170# 0.56f
C515 a_2475_11190# a_31990_11166# 0.264f
C516 a_2275_11190# a_29374_11206# 0.144f
C517 a_16930_11166# a_17022_11166# 0.326f
C518 VDD a_15926_2130# 0.181f
C519 m2_29844_18014# a_30378_18234# 0.087f
C520 row_n[11] a_21342_13214# 0.0117f
C521 rowon_n[1] col[11] 0.0323f
C522 col_n[31] a_2475_10186# 0.0531f
C523 col_n[5] a_8386_10524# 0.0283f
C524 rowon_n[5] col[19] 0.0323f
C525 row_n[8] col[24] 0.0342f
C526 rowon_n[9] col[27] 0.0323f
C527 rowon_n[7] col[23] 0.0323f
C528 row_n[6] col[20] 0.0342f
C529 rowon_n[6] col[21] 0.0323f
C530 row_n[11] col[30] 0.0342f
C531 row_n[4] col[16] 0.0342f
C532 rowon_n[10] col[29] 0.0323f
C533 rowon_n[3] col[15] 0.0323f
C534 ctop col[5] 0.123f
C535 row_n[0] col[8] 0.0342f
C536 row_n[9] col[26] 0.0342f
C537 row_n[12] sample_n 0.0596f
C538 row_n[5] col[18] 0.0342f
C539 rowon_n[11] col[31] 0.0323f
C540 row_n[10] col[28] 0.0342f
C541 row_n[2] col[12] 0.0342f
C542 row_n[3] col[14] 0.0342f
C543 rowon_n[0] col[9] 0.0323f
C544 row_n[1] col[10] 0.0342f
C545 row_n[7] col[22] 0.0342f
C546 rowon_n[4] col[17] 0.0323f
C547 m2_31852_18014# m3_30980_18146# 0.0341f
C548 rowon_n[2] col[13] 0.0323f
C549 rowon_n[8] col[25] 0.0323f
C550 col[1] a_2275_8178# 0.0899f
C551 a_18026_4138# a_18026_3134# 0.843f
C552 row_n[1] a_31382_3174# 0.0117f
C553 row_n[13] a_11910_15182# 0.0437f
C554 vcm a_9294_6186# 0.155f
C555 a_2275_8178# a_22954_8154# 0.136f
C556 a_11910_8154# a_12306_8194# 0.0313f
C557 rowoff_n[11] a_4974_13174# 0.294f
C558 m2_15212_13422# a_15014_13174# 0.165f
C559 vcm a_34090_16186# 0.56f
C560 col[21] a_2475_7174# 0.136f
C561 VDD a_30986_6146# 0.181f
C562 row_n[3] a_21950_5142# 0.0437f
C563 col_n[0] a_2874_18194# 0.0762f
C564 rowon_n[7] a_21038_9158# 0.248f
C565 rowoff_n[6] a_10906_8154# 0.202f
C566 m2_5172_10410# row_n[8] 0.0128f
C567 m2_11196_6394# row_n[4] 0.0128f
C568 m2_16216_2378# row_n[0] 0.0128f
C569 col_n[3] a_5978_10162# 0.251f
C570 col_n[29] a_32386_11206# 0.084f
C571 a_7986_5142# a_8990_5142# 0.843f
C572 a_2475_5166# a_15014_5142# 0.316f
C573 col_n[28] a_2275_13198# 0.113f
C574 m2_34288_9406# a_34090_9158# 0.165f
C575 col_n[10] a_12914_12170# 0.0765f
C576 vcm a_24354_10202# 0.155f
C577 rowoff_n[15] a_21038_17190# 0.294f
C578 rowoff_n[4] a_19942_6146# 0.202f
C579 a_31990_15182# a_32082_15182# 0.326f
C580 VDD a_11910_9158# 0.181f
C581 col[25] rowoff_n[12] 0.0901f
C582 col[18] a_2275_10186# 0.0899f
C583 m2_26256_15430# row_n[13] 0.0128f
C584 a_2275_2154# a_5978_2130# 0.399f
C585 m2_32280_11414# row_n[9] 0.0128f
C586 vcm a_17934_4138# 0.1f
C587 col_n[1] a_3878_10162# 0.0765f
C588 rowon_n[1] a_8898_3134# 0.118f
C589 rowoff_n[9] a_11398_11528# 0.0133f
C590 rowoff_n[2] a_28978_4138# 0.202f
C591 a_33086_8154# a_33086_7150# 0.843f
C592 a_2475_7174# a_30074_7150# 0.316f
C593 m2_6176_11414# a_5978_11166# 0.165f
C594 col[23] a_26058_9158# 0.367f
C595 vcm a_5278_13214# 0.155f
C596 a_26970_12170# a_27366_12210# 0.0313f
C597 VDD a_2966_3134# 0.485f
C598 col[30] a_32994_11166# 0.0682f
C599 ctop a_18026_8154# 4.11f
C600 a_2475_16210# a_8898_16186# 0.264f
C601 a_2275_16210# a_6282_16226# 0.144f
C602 VDD a_26970_13174# 0.181f
C603 row_n[8] a_29374_10202# 0.0117f
C604 rowoff_n[7] a_20434_9520# 0.0133f
C605 a_11910_4138# a_12402_4500# 0.0658f
C606 a_2275_4162# a_21038_4138# 0.399f
C607 a_10998_4138# a_11302_4178# 0.0931f
C608 m3_5880_1078# ctop 0.21f
C609 m2_25252_7398# a_25054_7150# 0.165f
C610 col_n[3] a_2475_17214# 0.0531f
C611 col_n[18] a_21342_9198# 0.084f
C612 vcm a_32994_8154# 0.1f
C613 rowoff_n[13] a_27462_15544# 0.0133f
C614 a_23046_9158# a_24050_9158# 0.843f
C615 col_n[8] a_2475_6170# 0.0531f
C616 row_n[10] a_19942_12170# 0.0437f
C617 vcm a_20338_17230# 0.155f
C618 rowon_n[14] a_19030_16186# 0.248f
C619 a_35002_14178# a_35398_14218# 0.0313f
C620 VDD a_18426_7512# 0.0779f
C621 rowoff_n[5] a_29470_7512# 0.0133f
C622 ctop a_33086_12170# 4.11f
C623 col_n[29] a_32482_3496# 0.0283f
C624 col[9] rowoff_n[13] 0.0901f
C625 a_2275_18218# a_21342_18234# 0.145f
C626 a_12914_18194# a_13006_18194# 0.0991f
C627 VDD a_7894_16186# 0.181f
C628 row_n[0] a_29982_2130# 0.0437f
C629 a_7894_1126# a_7986_1126# 0.0991f
C630 a_2275_1150# a_11302_1166# 0.145f
C631 a_2475_1150# a_13918_1126# 0.264f
C632 rowon_n[4] a_29070_6146# 0.248f
C633 vcm a_13918_11166# 0.1f
C634 a_14010_11166# a_14010_10162# 0.843f
C635 VDD a_9994_1126# 0.035f
C636 col[12] a_15014_7150# 0.367f
C637 a_7894_15182# a_8290_15222# 0.0313f
C638 a_2275_15206# a_14922_15182# 0.136f
C639 VDD a_33486_11528# 0.0779f
C640 col_n[5] a_2275_9182# 0.113f
C641 col[19] a_21950_9158# 0.0682f
C642 ctop a_14010_15182# 4.11f
C643 rowon_n[0] m2_23244_2378# 0.0322f
C644 row_n[4] a_6982_6146# 0.282f
C645 a_2275_3158# a_26362_3174# 0.144f
C646 a_2475_3158# a_28978_3134# 0.264f
C647 rowon_n[8] a_6890_10162# 0.118f
C648 col_n[27] a_30074_3134# 0.251f
C649 rowoff_n[8] a_30074_10162# 0.294f
C650 m2_16216_5390# a_16018_5142# 0.165f
C651 rowoff_n[11] a_33998_13174# 0.202f
C652 a_26970_8154# a_27462_8516# 0.0658f
C653 a_26058_8154# a_26362_8194# 0.0931f
C654 col_n[25] a_2475_8178# 0.0531f
C655 vcm a_28978_15182# 0.1f
C656 col_n[7] a_10298_7190# 0.084f
C657 a_3970_12170# a_4974_12170# 0.843f
C658 a_2475_12194# a_6982_12170# 0.316f
C659 VDD a_25054_5142# 0.483f
C660 m2_8184_18442# VDD 0.0456f
C661 row_n[15] a_27366_17230# 0.0117f
C662 a_2275_17214# a_29982_17190# 0.136f
C663 VDD a_14410_14540# 0.0779f
C664 m3_34996_17142# a_34090_17190# 0.0303f
C665 col_n[18] a_21438_1488# 0.0283f
C666 col[10] a_2475_16210# 0.136f
C667 a_22954_5142# a_23046_5142# 0.326f
C668 col_n[28] a_31478_13536# 0.0283f
C669 col[15] a_2475_5166# 0.136f
C670 rowoff_n[14] a_15414_16548# 0.0133f
C671 vcm a_9902_18194# 0.101f
C672 a_29070_15182# a_29070_14178# 0.843f
C673 a_2475_14202# a_22042_14178# 0.316f
C674 row_n[7] a_27974_9158# 0.0437f
C675 VDD a_5978_8154# 0.483f
C676 m2_1732_4962# rowon_n[3] 0.236f
C677 rowon_n[11] a_27062_13174# 0.248f
C678 col[1] a_3970_5142# 0.367f
C679 col_n[22] a_2275_11190# 0.113f
C680 VDD a_29470_18556# 0.0858f
C681 col[11] a_14010_17190# 0.367f
C682 a_17934_2130# a_18330_2170# 0.0313f
C683 a_2275_2154# a_35002_2130# 0.136f
C684 col[8] a_10906_7150# 0.0682f
C685 m2_7180_3382# a_6982_3134# 0.165f
C686 m3_24956_18146# VDD 0.0277f
C687 vcm a_12002_3134# 0.56f
C688 col_n[16] a_19030_1126# 0.303f
C689 col_n[26] a_29070_13174# 0.251f
C690 a_7894_11166# a_8386_11528# 0.0658f
C691 a_2275_11190# a_13006_11166# 0.399f
C692 a_6982_11166# a_7286_11206# 0.0931f
C693 col_n[23] a_25966_3134# 0.0765f
C694 row_n[1] col[21] 0.0342f
C695 rowon_n[6] sample_n 0.0692f
C696 rowon_n[0] col[20] 0.0323f
C697 rowon_n[4] col[28] 0.0323f
C698 row_n[0] col[19] 0.0342f
C699 row_n[2] col[23] 0.0342f
C700 ctop col[16] 0.129f
C701 row_n[6] col[31] 0.0342f
C702 rowon_n[5] col[30] 0.0323f
C703 row_n[5] col[29] 0.0342f
C704 rowon_n[1] col[22] 0.0323f
C705 row_n[4] col[27] 0.0342f
C706 rowon_n[2] col[24] 0.0323f
C707 row_n[3] col[25] 0.0342f
C708 rowon_n[3] col[26] 0.0323f
C709 col[12] a_2275_8178# 0.0899f
C710 row_n[11] a_4974_13174# 0.282f
C711 a_19030_16186# a_20034_16186# 0.843f
C712 VDD a_21038_12170# 0.483f
C713 m2_7756_18014# m3_7888_18146# 3.79f
C714 rowon_n[15] a_4882_17190# 0.118f
C715 col_n[6] a_9294_17230# 0.084f
C716 m2_16216_14426# rowon_n[12] 0.0322f
C717 m2_22240_10410# rowon_n[8] 0.0322f
C718 m2_28264_6394# rowon_n[4] 0.0322f
C719 row_n[1] a_15014_3134# 0.282f
C720 rowon_n[5] a_14922_7150# 0.118f
C721 vcm a_27062_7150# 0.56f
C722 a_2275_8178# a_3270_8194# 0.144f
C723 rowoff_n[12] a_21950_14178# 0.202f
C724 a_2475_8178# a_5886_8154# 0.264f
C725 col_n[17] a_20434_11528# 0.0283f
C726 a_2275_13198# a_28066_13174# 0.399f
C727 row_n[3] a_3878_5142# 0.0437f
C728 rowon_n[7] a_2966_9158# 0.248f
C729 VDD a_2475_15206# 26.1f
C730 col_n[2] a_2475_4162# 0.0531f
C731 vcm a_17326_1166# 0.16f
C732 a_32994_6146# a_33390_6186# 0.0313f
C733 col[0] a_2874_15182# 0.0682f
C734 m2_10768_946# m3_9896_1078# 0.0341f
C735 vcm a_7986_10162# 0.56f
C736 col[7] a_9902_17190# 0.0682f
C737 a_2275_10186# a_18330_10202# 0.144f
C738 rowoff_n[15] a_2966_17190# 0.294f
C739 a_2475_10186# a_20946_10162# 0.264f
C740 row_n[14] a_25966_16186# 0.0437f
C741 col_n[15] a_18026_11166# 0.251f
C742 a_22042_15182# a_22346_15222# 0.0931f
C743 a_22954_15182# a_23446_15544# 0.0658f
C744 col[29] a_2275_10186# 0.0899f
C745 col_n[12] a_14922_1126# 0.0765f
C746 row_n[4] a_34394_6186# 0.0117f
C747 col_n[22] a_24962_13174# 0.0765f
C748 a_29070_3134# a_30074_3134# 0.843f
C749 rowon_n[8] a_35094_10162# 0.0141f
C750 vcm a_32386_5182# 0.155f
C751 a_2275_7174# a_11910_7150# 0.136f
C752 m2_25828_18014# vcm 0.353f
C753 col_n[0] a_2275_7174# 0.113f
C754 vcm a_23046_14178# 0.56f
C755 a_2275_12194# a_33390_12210# 0.144f
C756 a_18938_12170# a_19030_12170# 0.326f
C757 VDD a_19942_4138# 0.181f
C758 col_n[6] a_9390_9520# 0.0283f
C759 col_n[14] a_2475_17214# 0.0531f
C760 row_n[8] a_13006_10162# 0.282f
C761 rowoff_n[7] a_2161_9182# 0.0226f
C762 col_n[19] a_2475_6170# 0.0531f
C763 rowon_n[12] a_12914_14178# 0.118f
C764 a_2475_4162# a_3970_4138# 0.316f
C765 a_2275_4162# a_2966_4138# 0.399f
C766 a_20034_5142# a_20034_4138# 0.843f
C767 m2_31852_18014# m2_32856_18014# 0.843f
C768 vcm a_13310_8194# 0.155f
C769 rowoff_n[13] a_9902_15182# 0.202f
C770 a_13918_9158# a_14314_9198# 0.0313f
C771 a_2275_9182# a_26970_9158# 0.136f
C772 rowon_n[2] a_22954_4138# 0.118f
C773 vcm a_3970_17190# 0.56f
C774 ctop a_26058_3134# 4.11f
C775 col[20] rowoff_n[13] 0.0901f
C776 m3_17928_1078# a_19030_1126# 0.0228f
C777 VDD a_35002_8154# 0.258f
C778 rowoff_n[5] a_11910_7150# 0.202f
C779 col[4] a_2475_14202# 0.136f
C780 a_2874_18194# a_3270_18234# 0.0313f
C781 col_n[1] rowoff_n[7] 0.0471f
C782 a_3878_18194# a_3970_18194# 0.0991f
C783 col_n[3] rowoff_n[9] 0.0471f
C784 VDD rowoff_n[3] 1.51f
C785 sample rowoff_n[4] 0.0775f
C786 col_n[0] rowoff_n[5] 0.0471f
C787 col_n[2] rowoff_n[8] 0.0471f
C788 a_2275_18218# a_4974_18194# 0.0924f
C789 vcm rowoff_n[6] 0.533f
C790 col[9] a_2475_3158# 0.136f
C791 col_n[30] a_33390_10202# 0.084f
C792 row_n[0] a_10298_2170# 0.0117f
C793 col_n[4] a_6982_9158# 0.251f
C794 a_32082_2130# a_32386_2170# 0.0931f
C795 a_32994_2130# a_33486_2492# 0.0658f
C796 col_n[11] a_13918_11166# 0.0765f
C797 m2_12776_18014# col_n[10] 0.243f
C798 vcm a_6890_2130# 0.1f
C799 a_2475_6170# a_19030_6146# 0.316f
C800 a_9994_6146# a_10998_6146# 0.843f
C801 rowoff_n[3] a_20946_5142# 0.202f
C802 vcm a_28370_12210# 0.155f
C803 VDD a_26458_2492# 0.0779f
C804 col_n[16] a_2275_9182# 0.113f
C805 m2_9188_17438# row_n[15] 0.0128f
C806 m2_15212_13422# row_n[11] 0.0128f
C807 m2_34864_7974# VDD 0.766f
C808 m2_21236_9406# row_n[7] 0.0128f
C809 m2_27260_5390# row_n[3] 0.0128f
C810 ctop a_6982_6146# 4.11f
C811 a_33998_16186# a_34090_16186# 0.326f
C812 row_n[11] a_33998_13174# 0.0437f
C813 VDD a_15926_11166# 0.181f
C814 rowon_n[15] a_33086_17190# 0.248f
C815 a_2275_3158# a_9994_3134# 0.399f
C816 a_2475_18218# a_2874_18194# 0.264f
C817 rowoff_n[8] a_12402_10524# 0.0133f
C818 rowoff_n[1] a_29982_3134# 0.202f
C819 col[1] a_2275_17214# 0.0899f
C820 m2_1732_4962# a_2475_5166# 0.139f
C821 col[24] a_27062_8154# 0.367f
C822 vcm a_21950_6146# 0.1f
C823 col[6] a_2275_6170# 0.0899f
C824 m2_34864_13998# m2_35292_14426# 0.165f
C825 a_2475_8178# a_34090_8154# 0.316f
C826 col[4] rowoff_n[14] 0.0901f
C827 col[31] a_33998_10162# 0.0682f
C828 vcm a_9294_15222# 0.155f
C829 a_28978_13174# a_29374_13214# 0.0313f
C830 VDD a_7382_5504# 0.0779f
C831 ctop a_22042_10162# 4.11f
C832 row_n[15] a_10998_17190# 0.282f
C833 a_2475_17214# a_12914_17190# 0.264f
C834 col[21] a_2475_16210# 0.136f
C835 a_2275_17214# a_10298_17230# 0.144f
C836 VDD a_30986_15182# 0.181f
C837 rowoff_n[6] a_21438_8516# 0.0133f
C838 col[26] a_2475_5166# 0.136f
C839 col_n[19] a_22346_8194# 0.084f
C840 a_2275_5166# a_25054_5142# 0.399f
C841 a_13918_5142# a_14410_5504# 0.0658f
C842 row_n[5] a_21038_7150# 0.282f
C843 a_13006_5142# a_13310_5182# 0.0931f
C844 rowon_n[9] a_20946_11166# 0.118f
C845 vcm a_2161_9182# 0.0169f
C846 a_25054_10162# a_26058_10162# 0.843f
C847 m2_30272_16434# a_30074_16186# 0.165f
C848 rowoff_n[4] a_30474_6508# 0.0133f
C849 m2_5748_946# a_6282_1166# 0.087f
C850 m2_15788_946# a_2275_1150# 0.28f
C851 m3_8892_1078# a_8990_2130# 0.0302f
C852 a_2874_14178# a_2966_14178# 0.326f
C853 row_n[7] a_8290_9198# 0.0117f
C854 VDD a_22442_9520# 0.0779f
C855 col_n[30] a_33486_2492# 0.0283f
C856 m2_1732_16006# ctop 0.0428f
C857 VDD a_11910_18194# 0.343f
C858 a_2475_2154# a_17934_2130# 0.264f
C859 a_9902_2130# a_9994_2130# 0.326f
C860 a_2275_2154# a_15318_2170# 0.144f
C861 m2_10192_1374# VDD 0.0194f
C862 vcm col_n[1] 1.93f
C863 VDD col_n[4] 5.17f
C864 row_n[1] sample_n 0.0596f
C865 rowon_n[0] col[31] 0.0323f
C866 rowoff_n[9] a_22042_11166# 0.294f
C867 col[10] col[11] 0.0355f
C868 ctop col[27] 0.123f
C869 row_n[0] col[30] 0.0342f
C870 col[23] a_2275_8178# 0.0899f
C871 vcm a_17934_13174# 0.1f
C872 col[13] a_16018_6146# 0.367f
C873 a_16018_12170# a_16018_11166# 0.843f
C874 VDD a_14010_3134# 0.483f
C875 m2_16792_18014# a_2275_18218# 0.28f
C876 col[20] a_22954_8154# 0.0682f
C877 a_9902_16186# a_10298_16226# 0.0313f
C878 a_2275_16210# a_18938_16186# 0.136f
C879 rowon_n[3] a_7986_5142# 0.248f
C880 VDD a_2966_12170# 0.485f
C881 a_26970_1126# m2_26832_946# 0.225f
C882 col_n[28] a_31078_2130# 0.251f
C883 ctop a_18026_17190# 4.06f
C884 rowoff_n[7] a_31078_9158# 0.294f
C885 a_2275_4162# a_30378_4178# 0.144f
C886 a_2475_4162# a_32994_4138# 0.264f
C887 rowoff_n[12] a_3878_14178# 0.202f
C888 a_28066_9158# a_28370_9198# 0.0931f
C889 col_n[8] a_11302_6186# 0.084f
C890 a_28978_9158# a_29470_9520# 0.0658f
C891 m2_21236_14426# a_21038_14178# 0.165f
C892 col_n[18] a_21342_18234# 0.084f
C893 vcm a_32994_17190# 0.1f
C894 col_n[8] a_2475_15206# 0.0531f
C895 a_5978_13174# a_6982_13174# 0.843f
C896 a_2475_13198# a_10998_13174# 0.316f
C897 VDD a_29070_7150# 0.483f
C898 col_n[13] a_2475_4162# 0.0531f
C899 a_2275_18218# a_33998_18194# 0.136f
C900 m2_12776_18014# a_2475_18218# 0.286f
C901 VDD a_18426_16548# 0.0779f
C902 a_2275_1150# a_23958_1126# 0.136f
C903 row_n[12] a_19030_14178# 0.282f
C904 m2_18224_2378# a_18026_2130# 0.165f
C905 col_n[29] a_32482_12532# 0.0283f
C906 vcm a_35094_2130# 0.165f
C907 a_24962_6146# a_25054_6146# 0.326f
C908 m2_24824_946# m2_25252_1374# 0.165f
C909 row_n[2] a_29070_4138# 0.282f
C910 a_1957_10186# a_2161_10186# 0.115f
C911 a_2475_10186# a_2275_10186# 2.76f
C912 col[3] a_2475_1150# 0.136f
C913 row_n[14] a_6282_16226# 0.0117f
C914 rowon_n[6] a_28978_8154# 0.118f
C915 m3_34996_4090# a_34090_4138# 0.0303f
C916 col[2] a_4974_4138# 0.367f
C917 a_31078_16186# a_31078_15182# 0.843f
C918 a_2475_15206# a_26058_15182# 0.316f
C919 VDD a_9994_10162# 0.483f
C920 col[12] a_15014_16186# 0.367f
C921 row_n[4] a_16322_6186# 0.0117f
C922 col[9] a_11910_6146# 0.0682f
C923 col_n[5] a_2275_18218# 0.113f
C924 a_19942_3134# a_20338_3174# 0.0313f
C925 col[19] a_21950_18194# 0.0682f
C926 a_2475_18218# a_31990_18194# 0.264f
C927 col_n[10] a_2275_7174# 0.113f
C928 vcm a_16018_5142# 0.56f
C929 rowoff_n[10] a_9994_12170# 0.294f
C930 col_n[27] a_30074_12170# 0.251f
C931 a_29982_1126# vcm 0.0989f
C932 col_n[24] a_26970_2130# 0.0765f
C933 m2_12200_12418# a_12002_12170# 0.165f
C934 m2_5172_12418# rowon_n[10] 0.0322f
C935 row_n[6] a_6890_8154# 0.0437f
C936 m2_11196_8402# rowon_n[6] 0.0322f
C937 m2_17220_4386# rowon_n[2] 0.0322f
C938 a_8990_12170# a_9294_12210# 0.0931f
C939 a_9902_12170# a_10394_12532# 0.0658f
C940 a_2275_12194# a_17022_12170# 0.399f
C941 VDD a_35398_5182# 0.0882f
C942 rowon_n[10] a_5978_12170# 0.248f
C943 col_n[25] a_2475_17214# 0.0531f
C944 m2_29844_18014# VDD 1f
C945 col_n[7] a_10298_16226# 0.084f
C946 a_21038_17190# a_22042_17190# 0.843f
C947 VDD a_25054_14178# 0.483f
C948 col_n[30] a_2475_6170# 0.0531f
C949 a_3270_1166# m2_2736_946# 0.087f
C950 col[0] a_2275_4162# 0.099f
C951 rowon_n[0] a_16018_2130# 0.248f
C952 rowoff_n[0] a_2475_2154# 3.9f
C953 en_bit_n[0] a_19942_1126# 0.0802f
C954 m2_31276_8402# a_31078_8154# 0.165f
C955 col_n[18] a_21438_10524# 0.0283f
C956 col[31] rowoff_n[13] 0.0901f
C957 vcm a_31078_9158# 0.56f
C958 a_2275_9182# a_7286_9198# 0.144f
C959 a_2475_9182# a_9902_9158# 0.264f
C960 rowoff_n[14] a_26058_16186# 0.294f
C961 a_5886_9158# a_5978_9158# 0.326f
C962 col[15] a_2475_14202# 0.136f
C963 col_n[6] rowoff_n[1] 0.0471f
C964 col[20] a_2475_3158# 0.136f
C965 col_n[8] rowoff_n[3] 0.0471f
C966 col_n[13] rowoff_n[8] 0.0471f
C967 col_n[11] rowoff_n[6] 0.0471f
C968 col_n[7] rowoff_n[2] 0.0471f
C969 col_n[10] rowoff_n[5] 0.0471f
C970 col_n[9] rowoff_n[4] 0.0471f
C971 col_n[14] rowoff_n[9] 0.0471f
C972 col_n[12] rowoff_n[7] 0.0471f
C973 col_n[5] rowoff_n[0] 0.0471f
C974 m2_26256_17438# rowon_n[15] 0.0322f
C975 a_2275_14202# a_32082_14178# 0.399f
C976 m2_32280_13422# rowon_n[11] 0.0322f
C977 VDD a_5978_17190# 0.484f
C978 col[1] a_3970_14178# 0.367f
C979 vcm a_21342_3174# 0.155f
C980 row_n[9] a_27062_11166# 0.282f
C981 col_n[27] a_2275_9182# 0.113f
C982 m2_1732_13998# sample_n 0.0522f
C983 col[8] a_10906_16186# 0.0682f
C984 rowon_n[13] a_26970_15182# 0.118f
C985 rowoff_n[3] a_2275_5166# 0.151f
C986 vcm a_12002_12170# 0.56f
C987 a_2275_11190# a_22346_11206# 0.144f
C988 a_2475_11190# a_24962_11166# 0.264f
C989 VDD a_8898_2130# 0.181f
C990 col_n[16] a_19030_10162# 0.251f
C991 a_24962_16186# a_25454_16548# 0.0658f
C992 a_24050_16186# a_24354_16226# 0.0931f
C993 row_n[11] a_14314_13214# 0.0117f
C994 col_n[23] a_25966_12170# 0.0765f
C995 m2_21812_18014# m3_22948_18146# 0.0341f
C996 col[12] a_2275_17214# 0.0899f
C997 col[17] a_2275_6170# 0.0899f
C998 a_31078_4138# a_32082_4138# 0.843f
C999 row_n[1] a_24354_3174# 0.0117f
C1000 col[15] rowoff_n[14] 0.0901f
C1001 m2_22240_6394# a_22042_6146# 0.165f
C1002 row_n[13] a_4882_15182# 0.0437f
C1003 vcm a_3878_6146# 0.1f
C1004 a_2275_8178# a_15926_8154# 0.136f
C1005 rowoff_n[12] a_32482_14540# 0.0133f
C1006 sample rowoff_n[10] 0.0775f
C1007 col_n[7] a_10394_8516# 0.0283f
C1008 vcm a_27062_16186# 0.56f
C1009 a_20946_13174# a_21038_13174# 0.326f
C1010 VDD a_23958_6146# 0.181f
C1011 row_n[3] a_14922_5142# 0.0437f
C1012 rowon_n[7] a_14010_9158# 0.248f
C1013 rowoff_n[6] a_3366_8516# 0.0133f
C1014 m2_34864_8978# rowoff_n[7] 0.278f
C1015 a_2475_5166# a_7986_5142# 0.316f
C1016 row_n[5] a_2966_7150# 0.281f
C1017 a_22042_6146# a_22042_5142# 0.843f
C1018 col_n[2] a_2475_13198# 0.0531f
C1019 m2_25828_946# m3_25960_1078# 3.79f
C1020 rowon_n[9] a_2275_11190# 1.79f
C1021 vcm a_17326_10202# 0.155f
C1022 col_n[7] a_2475_2154# 0.0531f
C1023 rowoff_n[15] a_14010_17190# 0.294f
C1024 a_15926_10162# a_16322_10202# 0.0313f
C1025 a_2275_10186# a_30986_10162# 0.136f
C1026 rowoff_n[4] a_12914_6146# 0.202f
C1027 ctop a_30074_5142# 4.11f
C1028 VDD a_4882_9158# 0.181f
C1029 col_n[5] a_7986_8154# 0.251f
C1030 VDD col_n[15] 4.83f
C1031 vcm col_n[12] 1.94f
C1032 col_n[12] a_14922_10162# 0.0765f
C1033 a_35002_3134# a_35494_3496# 0.0658f
C1034 m2_4168_11414# row_n[9] 0.0128f
C1035 m2_13204_4386# a_13006_4138# 0.165f
C1036 m2_10192_7398# row_n[5] 0.0128f
C1037 m2_16216_3382# row_n[1] 0.0128f
C1038 vcm a_10906_4138# 0.1f
C1039 rowoff_n[2] a_21950_4138# 0.202f
C1040 a_2475_7174# a_23046_7150# 0.316f
C1041 rowoff_n[9] a_4370_11528# 0.0133f
C1042 a_12002_7150# a_13006_7150# 0.843f
C1043 row_n[6] a_35094_8154# 0.0123f
C1044 vcm a_32386_14218# 0.155f
C1045 VDD a_30474_4500# 0.0779f
C1046 rowon_n[10] a_35002_12170# 0.118f
C1047 col_n[0] a_2275_16210# 0.113f
C1048 ctop a_10998_8154# 4.11f
C1049 VDD a_19942_13174# 0.181f
C1050 col_n[4] a_2275_5166# 0.113f
C1051 col_n[6] a_9390_18556# 0.0283f
C1052 row_n[8] a_22346_10202# 0.0117f
C1053 rowoff_n[0] a_30986_2130# 0.202f
C1054 rowoff_n[7] a_13406_9520# 0.0133f
C1055 col[25] a_28066_7150# 0.367f
C1056 a_2275_4162# a_14010_4138# 0.399f
C1057 m3_34996_13126# ctop 0.209f
C1058 m2_25252_16434# row_n[14] 0.0128f
C1059 col_n[19] a_2475_15206# 0.0531f
C1060 m2_31276_12418# row_n[10] 0.0128f
C1061 vcm a_25966_8154# 0.1f
C1062 rowoff_n[13] a_20434_15544# 0.0133f
C1063 col_n[24] a_2475_4162# 0.0531f
C1064 row_n[10] a_12914_12170# 0.0437f
C1065 ctop a_2275_2154# 0.0668f
C1066 vcm a_13310_17230# 0.155f
C1067 rowon_n[14] a_12002_16186# 0.248f
C1068 a_30986_14178# a_31382_14218# 0.0313f
C1069 VDD a_11398_7512# 0.0779f
C1070 rowoff_n[5] a_22442_7512# 0.0133f
C1071 ctop a_26058_12170# 4.11f
C1072 a_2275_18218# a_14314_18234# 0.145f
C1073 VDD a_35002_17190# 0.258f
C1074 row_n[0] a_22954_2130# 0.0437f
C1075 col_n[20] a_23350_7190# 0.084f
C1076 a_2475_1150# a_6890_1126# 0.264f
C1077 a_2275_1150# a_4274_1166# 0.126f
C1078 rowon_n[4] a_22042_6146# 0.248f
C1079 col[9] a_2475_12194# 0.136f
C1080 a_15926_6146# a_16418_6508# 0.0658f
C1081 a_15014_6146# a_15318_6186# 0.0931f
C1082 col[14] a_2475_1150# 0.136f
C1083 a_2275_6170# a_29070_6146# 0.399f
C1084 m2_34864_8978# vcm 0.408f
C1085 vcm a_6890_11166# 0.1f
C1086 rowoff_n[3] a_31478_5504# 0.0133f
C1087 a_27974_1126# col_n[25] 0.0786f
C1088 a_27062_11166# a_28066_11166# 0.843f
C1089 VDD a_2874_1126# 0.405f
C1090 a_2275_15206# a_7894_15182# 0.136f
C1091 m2_29844_946# col_n[27] 0.354f
C1092 VDD a_26458_11528# 0.0779f
C1093 col_n[16] a_2275_18218# 0.113f
C1094 m2_34864_16006# m3_34996_16138# 3.79f
C1095 col_n[21] a_2275_7174# 0.113f
C1096 ctop a_6982_15182# 4.11f
C1097 a_11910_3134# a_12002_3134# 0.326f
C1098 a_2475_3158# a_21950_3134# 0.264f
C1099 a_2275_3158# a_19334_3174# 0.144f
C1100 rowoff_n[8] a_23046_10162# 0.294f
C1101 m2_27836_18014# col[25] 0.347f
C1102 row_n[13] a_33086_15182# 0.282f
C1103 rowoff_n[11] a_26970_13174# 0.202f
C1104 col[14] a_17022_5142# 0.367f
C1105 col[24] a_27062_17190# 0.367f
C1106 vcm a_21950_15182# 0.1f
C1107 col[6] a_2275_15206# 0.0899f
C1108 a_18026_13174# a_18026_12170# 0.843f
C1109 col[21] a_23958_7150# 0.0682f
C1110 VDD a_18026_5142# 0.483f
C1111 col[11] a_2275_4162# 0.0899f
C1112 a_31990_1126# VDD 0.405f
C1113 row_n[15] a_20338_17230# 0.0117f
C1114 a_2275_17214# a_22954_17190# 0.136f
C1115 a_11910_17190# a_12306_17230# 0.0313f
C1116 rowoff_n[6] a_32082_8154# 0.294f
C1117 VDD a_7382_14540# 0.0779f
C1118 m3_28972_18146# a_29070_17190# 0.0303f
C1119 row_n[5] a_30378_7190# 0.0117f
C1120 col[26] a_2475_14202# 0.136f
C1121 a_2275_5166# a_35398_5182# 0.145f
C1122 col_n[9] a_12306_5182# 0.084f
C1123 m3_26964_1078# m3_27968_1078# 0.202f
C1124 col_n[17] rowoff_n[1] 0.0471f
C1125 col_n[19] rowoff_n[3] 0.0471f
C1126 col_n[23] rowoff_n[7] 0.0471f
C1127 col_n[24] rowoff_n[8] 0.0471f
C1128 col_n[16] rowoff_n[0] 0.0471f
C1129 col_n[18] rowoff_n[2] 0.0471f
C1130 col_n[21] rowoff_n[5] 0.0471f
C1131 col[31] a_2475_3158# 0.136f
C1132 col_n[25] rowoff_n[9] 0.0471f
C1133 col_n[20] rowoff_n[4] 0.0471f
C1134 col_n[22] rowoff_n[6] 0.0471f
C1135 a_32994_1126# a_33086_1126# 0.0991f
C1136 col_n[19] a_22346_17230# 0.084f
C1137 a_30074_10162# a_30378_10202# 0.0931f
C1138 rowoff_n[14] a_8386_16548# 0.0133f
C1139 a_30986_10162# a_31478_10524# 0.0658f
C1140 vcm a_2161_18218# 0.0168f
C1141 col_n[2] a_2475_18218# 0.0529f
C1142 a_7986_14178# a_8990_14178# 0.843f
C1143 a_2475_14202# a_15014_14178# 0.316f
C1144 VDD a_33086_9158# 0.483f
C1145 row_n[7] a_20946_9158# 0.0437f
C1146 rowon_n[11] a_20034_13174# 0.248f
C1147 col_n[30] a_33486_11528# 0.0283f
C1148 VDD a_22442_18556# 0.0858f
C1149 a_2275_2154# a_27974_2130# 0.136f
C1150 m2_33284_1374# VDD 0.0194f
C1151 vcm a_4974_3134# 0.56f
C1152 a_26970_7150# a_27062_7150# 0.326f
C1153 rowon_n[1] a_30074_3134# 0.248f
C1154 a_2275_11190# a_5978_11166# 0.399f
C1155 col[3] a_5978_3134# 0.367f
C1156 col[23] a_2275_17214# 0.0899f
C1157 m2_14784_18014# a_14922_18194# 0.225f
C1158 m2_1732_10986# VDD 0.856f
C1159 col[13] a_16018_15182# 0.367f
C1160 a_33086_17190# a_33086_16186# 0.843f
C1161 col[28] a_2275_6170# 0.0899f
C1162 a_2475_16210# a_30074_16186# 0.316f
C1163 col[10] a_12914_5142# 0.0682f
C1164 VDD a_14010_12170# 0.483f
C1165 a_35002_1126# m2_34864_946# 0.225f
C1166 col[26] rowoff_n[14] 0.0901f
C1167 col[20] a_22954_17190# 0.0682f
C1168 m2_5172_2378# rowon_n[0] 0.0322f
C1169 a_21950_4138# a_22346_4178# 0.0313f
C1170 row_n[1] a_7986_3134# 0.282f
C1171 col_n[28] a_31078_11166# 0.251f
C1172 col_n[9] rowoff_n[10] 0.0471f
C1173 rowon_n[5] a_7894_7150# 0.118f
C1174 vcm a_20034_7150# 0.56f
C1175 rowoff_n[12] a_14922_14178# 0.202f
C1176 a_11910_13174# a_12402_13536# 0.0658f
C1177 col_n[8] a_11302_15222# 0.084f
C1178 a_10998_13174# a_11302_13214# 0.0931f
C1179 a_2275_13198# a_21038_13174# 0.399f
C1180 col[1] a_3878_3134# 0.0682f
C1181 VDD a_29070_16186# 0.483f
C1182 a_18026_1126# a_19030_1126# 0.843f
C1183 col_n[13] a_2475_13198# 0.0531f
C1184 row_n[12] a_28370_14218# 0.0117f
C1185 col_n[18] a_2475_2154# 0.0531f
C1186 vcm a_10298_1166# 0.16f
C1187 col_n[19] a_22442_9520# 0.0283f
C1188 m2_15212_15430# rowon_n[13] 0.0322f
C1189 m2_21236_11414# rowon_n[9] 0.0322f
C1190 m2_27260_7398# rowon_n[5] 0.0322f
C1191 m2_33284_3382# rowon_n[1] 0.0322f
C1192 vcm a_35094_11166# 0.165f
C1193 a_2475_10186# a_13918_10162# 0.264f
C1194 a_2275_10186# a_11302_10202# 0.144f
C1195 a_7894_10162# a_7986_10162# 0.326f
C1196 row_n[14] a_18938_16186# 0.0437f
C1197 vcm col_n[23] 1.94f
C1198 VDD col_n[26] 5.17f
C1199 col_n[11] col_n[12] 0.0101f
C1200 col[10] rowoff_n[15] 0.0901f
C1201 col[21] col[22] 0.0355f
C1202 col[3] a_2475_10186# 0.136f
C1203 m2_34864_12994# m3_34996_13126# 3.79f
C1204 col[2] a_4974_13174# 0.367f
C1205 row_n[4] a_28978_6146# 0.0437f
C1206 rowon_n[8] a_28066_10162# 0.248f
C1207 a_8990_3134# a_8990_2130# 0.843f
C1208 col[9] a_11910_15182# 0.0682f
C1209 vcm a_25358_5182# 0.155f
C1210 rowoff_n[2] a_3878_4138# 0.202f
C1211 a_2966_7150# a_3970_7150# 0.843f
C1212 a_2275_7174# a_4882_7150# 0.136f
C1213 m2_11772_18014# vcm 0.353f
C1214 col_n[10] a_2275_16210# 0.113f
C1215 col_n[17] a_20034_9158# 0.251f
C1216 vcm a_16018_14178# 0.56f
C1217 col_n[15] a_2275_5166# 0.113f
C1218 a_2475_12194# a_28978_12170# 0.264f
C1219 a_2275_12194# a_26362_12210# 0.144f
C1220 VDD a_12914_4138# 0.181f
C1221 col_n[24] a_26970_11166# 0.0765f
C1222 a_26058_17190# a_26362_17230# 0.0931f
C1223 a_26970_17190# a_27462_17552# 0.0658f
C1224 row_n[0] m2_21236_2378# 0.0128f
C1225 VDD a_35398_14218# 0.0882f
C1226 row_n[8] a_5978_10162# 0.282f
C1227 col_n[30] a_2475_15206# 0.0531f
C1228 rowon_n[12] a_5886_14178# 0.118f
C1229 a_33086_5142# a_34090_5142# 0.843f
C1230 col[0] a_2275_13198# 0.099f
C1231 m2_21812_946# ctop 0.0428f
C1232 col[5] a_2275_2154# 0.0899f
C1233 vcm a_6282_8194# 0.155f
C1234 m2_24824_18014# m2_25828_18014# 0.843f
C1235 rowoff_n[13] a_2161_15206# 0.0226f
C1236 a_2275_9182# a_19942_9158# 0.136f
C1237 col_n[8] a_11398_7512# 0.0283f
C1238 m2_27260_15430# a_27062_15182# 0.165f
C1239 rowon_n[2] a_15926_4138# 0.118f
C1240 ctop a_19030_3134# 4.11f
C1241 vcm a_31078_18194# 0.165f
C1242 a_22954_14178# a_23046_14178# 0.326f
C1243 VDD a_27974_8154# 0.181f
C1244 rowoff_n[5] a_4882_7150# 0.202f
C1245 col[20] a_2475_12194# 0.136f
C1246 row_n[0] a_3270_2170# 0.0117f
C1247 col[25] a_2475_1150# 0.136f
C1248 vcm a_33998_3134# 0.1f
C1249 a_2475_6170# a_12002_6146# 0.316f
C1250 a_24050_7150# a_24050_6146# 0.843f
C1251 vcm a_21342_12210# 0.155f
C1252 rowoff_n[3] a_13918_5142# 0.202f
C1253 a_2275_11190# a_35002_11166# 0.136f
C1254 a_17934_11166# a_18330_11206# 0.0313f
C1255 col_n[27] a_2275_18218# 0.113f
C1256 VDD a_19430_2492# 0.0779f
C1257 m2_33860_18014# a_33998_18194# 0.225f
C1258 m2_10768_18014# a_10998_17190# 0.843f
C1259 col_n[6] a_8990_7150# 0.251f
C1260 ctop a_34090_7150# 4.06f
C1261 row_n[11] a_26970_13174# 0.0437f
C1262 VDD a_8898_11166# 0.181f
C1263 m2_1732_17010# m3_1864_16138# 0.0341f
C1264 rowon_n[15] a_26058_17190# 0.248f
C1265 col_n[13] a_15926_9158# 0.0765f
C1266 a_2275_3158# a_2874_3134# 0.136f
C1267 a_2475_3158# a_3878_3134# 0.264f
C1268 rowoff_n[1] a_22954_3134# 0.202f
C1269 rowoff_n[8] a_5374_10524# 0.0133f
C1270 col[17] a_2275_15206# 0.0899f
C1271 vcm a_14922_6146# 0.1f
C1272 a_2475_8178# a_27062_8154# 0.316f
C1273 a_14010_8154# a_15014_8154# 0.843f
C1274 col[22] a_2275_4162# 0.0899f
C1275 m2_18224_13422# a_18026_13174# 0.165f
C1276 vcm a_3878_15182# 0.1f
C1277 VDD a_34490_6508# 0.0779f
C1278 ctop a_15014_10162# 4.11f
C1279 col_n[7] a_10394_17552# 0.0283f
C1280 row_n[15] a_3970_17190# 0.282f
C1281 m2_14208_14426# row_n[12] 0.0128f
C1282 a_2275_17214# a_3270_17230# 0.144f
C1283 a_2475_17214# a_5886_17190# 0.264f
C1284 m2_20232_10410# row_n[8] 0.0128f
C1285 rowoff_n[6] a_14410_8516# 0.0133f
C1286 VDD a_23958_15182# 0.181f
C1287 m2_26256_6394# row_n[4] 0.0128f
C1288 col[26] a_29070_6146# 0.367f
C1289 col_n[29] rowoff_n[2] 0.0471f
C1290 col_n[31] rowoff_n[4] 0.0471f
C1291 col_n[27] rowoff_n[0] 0.0471f
C1292 col_n[30] rowoff_n[3] 0.0471f
C1293 col_n[28] rowoff_n[1] 0.0471f
C1294 m2_34864_3958# m2_34864_2954# 0.843f
C1295 a_2275_5166# a_18026_5142# 0.399f
C1296 row_n[5] a_14010_7150# 0.282f
C1297 m3_1864_6098# m3_1864_5094# 0.202f
C1298 col_n[13] a_2475_18218# 0.0529f
C1299 rowon_n[9] a_13918_11166# 0.118f
C1300 vcm a_29982_10162# 0.1f
C1301 en_C0_n a_3878_1126# 0.0802f
C1302 a_4974_10162# a_4974_9158# 0.843f
C1303 rowoff_n[4] a_23446_6508# 0.0133f
C1304 col_n[7] a_2475_11190# 0.0531f
C1305 a_32994_15182# a_33390_15222# 0.0313f
C1306 VDD a_15414_9520# 0.0779f
C1307 row_n[7] a_2275_9182# 19.2f
C1308 m2_34864_9982# m3_34996_10114# 3.79f
C1309 rowon_n[11] a_1957_13198# 0.0172f
C1310 ctop a_30074_14178# 4.11f
C1311 col_n[21] a_24354_6186# 0.084f
C1312 VDD a_4882_18194# 0.343f
C1313 col_n[5] a_7986_17190# 0.251f
C1314 a_2475_2154# a_10906_2130# 0.264f
C1315 a_2275_2154# a_8290_2170# 0.144f
C1316 col_n[2] a_4882_7150# 0.0765f
C1317 rowoff_n[9] a_15014_11166# 0.294f
C1318 a_17934_7150# a_18426_7512# 0.0658f
C1319 a_2275_7174# a_33086_7150# 0.399f
C1320 rowoff_n[2] a_32482_4500# 0.0133f
C1321 a_17022_7150# a_17326_7190# 0.0931f
C1322 m2_9188_11414# a_8990_11166# 0.165f
C1323 vcm a_10906_13174# 0.1f
C1324 a_29070_12170# a_30074_12170# 0.843f
C1325 VDD a_6982_3134# 0.483f
C1326 m2_2736_18014# a_2275_18218# 0.281f
C1327 a_2275_16210# a_11910_16186# 0.136f
C1328 VDD a_30474_13536# 0.0779f
C1329 col_n[20] rowoff_n[10] 0.0471f
C1330 row_n[8] a_35002_10162# 0.0437f
C1331 ctop a_10998_17190# 4.06f
C1332 rowoff_n[7] a_24050_9158# 0.294f
C1333 col_n[4] a_2275_14202# 0.113f
C1334 rowon_n[12] a_34090_14178# 0.248f
C1335 a_2275_4162# a_23350_4178# 0.144f
C1336 a_2475_4162# a_25966_4138# 0.264f
C1337 a_13918_4138# a_14010_4138# 0.326f
C1338 m3_20940_1078# ctop 0.21f
C1339 col_n[9] a_2275_3158# 0.113f
C1340 col[15] a_18026_4138# 0.367f
C1341 m2_28264_7398# a_28066_7150# 0.165f
C1342 col[25] a_28066_16186# 0.367f
C1343 vcm a_1957_7174# 0.139f
C1344 rowoff_n[13] a_31078_15182# 0.294f
C1345 col[22] a_24962_6146# 0.0682f
C1346 vcm a_25966_17190# 0.1f
C1347 a_20034_14178# a_20034_13174# 0.843f
C1348 a_2475_13198# a_3970_13174# 0.316f
C1349 a_2275_13198# a_2966_13174# 0.399f
C1350 VDD a_22042_7150# 0.483f
C1351 rowoff_n[5] a_33086_7150# 0.294f
C1352 col_n[24] a_2475_13198# 0.0531f
C1353 ctop a_2275_11190# 0.0683f
C1354 a_2275_18218# a_26970_18194# 0.136f
C1355 col_n[29] a_2475_2154# 0.0531f
C1356 a_13918_18194# a_14314_18234# 0.0313f
C1357 VDD a_11398_16548# 0.0779f
C1358 row_n[12] a_12002_14178# 0.282f
C1359 a_8898_1126# a_9294_1166# 0.0313f
C1360 a_2275_1150# a_16930_1126# 0.136f
C1361 col_n[10] a_13310_4178# 0.084f
C1362 vcm a_28066_2130# 0.56f
C1363 col_n[20] a_23350_16226# 0.084f
C1364 col_n[0] row_n[14] 0.298f
C1365 sample rowon_n[13] 0.0935f
C1366 row_n[2] a_22042_4138# 0.282f
C1367 vcm rowon_n[14] 0.65f
C1368 VDD row_n[13] 3.29f
C1369 col_n[2] rowon_n[15] 0.111f
C1370 col_n[1] row_n[15] 0.298f
C1371 col[21] rowoff_n[15] 0.0901f
C1372 a_32994_11166# a_33486_11528# 0.0658f
C1373 col[14] a_2475_10186# 0.136f
C1374 a_32082_11166# a_32386_11206# 0.0931f
C1375 VDD a_12306_1166# 0.0149f
C1376 m2_29844_18014# a_30074_17190# 0.843f
C1377 rowon_n[6] a_21950_8154# 0.118f
C1378 a_9994_15182# a_10998_15182# 0.843f
C1379 a_2475_15206# a_19030_15182# 0.316f
C1380 col_n[4] rowoff_n[11] 0.0471f
C1381 VDD a_2874_10162# 0.182f
C1382 col_n[31] a_34490_10524# 0.0283f
C1383 m2_1732_13998# m3_1864_13126# 0.0341f
C1384 row_n[4] a_9294_6186# 0.0117f
C1385 a_2275_3158# a_31990_3134# 0.136f
C1386 a_2475_18218# a_24962_18194# 0.264f
C1387 col_n[21] a_2275_16210# 0.113f
C1388 m2_19228_5390# a_19030_5142# 0.165f
C1389 a_24450_1488# a_23958_1126# 0.0658f
C1390 col_n[26] a_2275_5166# 0.113f
C1391 vcm a_8990_5142# 0.56f
C1392 a_28978_8154# a_29070_8154# 0.326f
C1393 rowoff_n[10] a_2874_12170# 0.202f
C1394 col[4] a_6982_2130# 0.367f
C1395 a_2275_12194# a_9994_12170# 0.399f
C1396 col[14] a_17022_14178# 0.367f
C1397 col[11] a_13918_4138# 0.0682f
C1398 m2_15788_18014# VDD 1.06f
C1399 row_n[15] a_32994_17190# 0.0437f
C1400 col[21] a_23958_16186# 0.0682f
C1401 a_2475_17214# a_34090_17190# 0.316f
C1402 VDD a_18026_14178# 0.483f
C1403 col[11] a_2275_13198# 0.0899f
C1404 col[16] a_2275_2154# 0.0899f
C1405 rowon_n[0] a_8990_2130# 0.248f
C1406 col_n[29] a_32082_10162# 0.251f
C1407 a_23958_5142# a_24354_5182# 0.0313f
C1408 vcm a_24050_9158# 0.56f
C1409 rowoff_n[14] a_19030_16186# 0.294f
C1410 col_n[9] a_12306_14218# 0.084f
C1411 col[31] a_2475_12194# 0.136f
C1412 m2_21812_946# a_22042_1126# 0.0249f
C1413 a_13918_14178# a_14410_14540# 0.0658f
C1414 a_13006_14178# a_13310_14218# 0.0931f
C1415 a_2275_14202# a_25054_14178# 0.399f
C1416 m2_4168_13422# rowon_n[11] 0.0322f
C1417 m2_34864_6970# m3_34996_7102# 3.79f
C1418 m2_10192_9406# rowon_n[7] 0.0322f
C1419 m2_16216_5390# rowon_n[3] 0.0322f
C1420 m2_13780_946# vcm 0.353f
C1421 VDD a_33086_18194# 0.0356f
C1422 a_20034_2130# a_21038_2130# 0.843f
C1423 col_n[20] a_23446_8516# 0.0283f
C1424 m2_10192_3382# a_9994_3134# 0.165f
C1425 vcm a_14314_3174# 0.155f
C1426 row_n[9] a_20034_11166# 0.282f
C1427 col_n[1] a_2475_9182# 0.0531f
C1428 m2_1732_11990# vcm 0.316f
C1429 rowon_n[13] a_19942_15182# 0.118f
C1430 vcm a_4974_12170# 0.56f
C1431 a_9902_11166# a_9994_11166# 0.326f
C1432 a_2275_11190# a_15318_11206# 0.144f
C1433 a_2475_11190# a_17934_11166# 0.264f
C1434 row_n[11] a_7286_13214# 0.0117f
C1435 rowon_n[3] a_29982_5142# 0.118f
C1436 col[3] a_5978_12170# 0.367f
C1437 m2_12776_18014# m3_12908_18146# 3.79f
C1438 m2_31276_14426# rowon_n[12] 0.0322f
C1439 col[28] a_2275_15206# 0.0899f
C1440 col[10] a_12914_14178# 0.0682f
C1441 a_10998_4138# a_10998_3134# 0.843f
C1442 row_n[1] a_17326_3174# 0.0117f
C1443 col_n[18] a_21038_8154# 0.251f
C1444 vcm a_29374_7190# 0.155f
C1445 rowoff_n[12] a_25454_14540# 0.0133f
C1446 a_2275_8178# a_8898_8154# 0.136f
C1447 a_4882_8154# a_5278_8194# 0.0313f
C1448 col_n[25] a_27974_10162# 0.0765f
C1449 vcm a_20034_16186# 0.56f
C1450 a_2275_13198# a_30378_13214# 0.144f
C1451 a_2475_13198# a_32994_13174# 0.264f
C1452 VDD a_16930_6146# 0.181f
C1453 row_n[3] a_7894_5142# 0.0437f
C1454 rowon_n[8] rowoff_n[8] 20.2f
C1455 col_n[3] a_2275_1150# 0.113f
C1456 rowon_n[7] a_6982_9158# 0.248f
C1457 a_28978_18194# a_29470_18556# 0.0658f
C1458 col[1] a_3878_12170# 0.0682f
C1459 col_n[24] a_2475_18218# 0.0529f
C1460 vcm a_22954_1126# 0.0989f
C1461 col_n[9] a_12402_6508# 0.0283f
C1462 m2_15788_946# m3_14916_1078# 0.0341f
C1463 m3_22948_18146# m3_23952_18146# 0.202f
C1464 col_n[18] a_2475_11190# 0.0531f
C1465 col_n[19] a_22442_18556# 0.0283f
C1466 vcm a_10298_10202# 0.155f
C1467 rowoff_n[15] a_6982_17190# 0.294f
C1468 a_2275_10186# a_23958_10162# 0.136f
C1469 rowoff_n[4] a_5886_6146# 0.202f
C1470 ctop a_23046_5142# 4.11f
C1471 a_24962_15182# a_25054_15182# 0.326f
C1472 VDD a_31990_10162# 0.181f
C1473 m2_1732_10986# m3_1864_10114# 0.0341f
C1474 col[8] a_2475_8178# 0.136f
C1475 rowoff_n[10] a_31990_12170# 0.202f
C1476 rowoff_n[2] a_14922_4138# 0.202f
C1477 a_2475_7174# a_16018_7150# 0.316f
C1478 a_26058_8154# a_26058_7150# 0.843f
C1479 row_n[6] a_28066_8154# 0.282f
C1480 vcm a_25358_14218# 0.155f
C1481 col_n[7] a_9994_6146# 0.251f
C1482 a_19942_12170# a_20338_12210# 0.0313f
C1483 VDD a_23446_4500# 0.0779f
C1484 rowon_n[10] a_27974_12170# 0.118f
C1485 col_n[31] rowoff_n[10] 0.0471f
C1486 ctop a_3970_8154# 4.11f
C1487 col_n[14] a_16930_8154# 0.0765f
C1488 col_n[15] a_2275_14202# 0.113f
C1489 VDD a_12914_13174# 0.181f
C1490 col_n[20] a_2275_3158# 0.113f
C1491 row_n[8] a_15318_10202# 0.0117f
C1492 rowoff_n[0] a_23958_2130# 0.202f
C1493 rowoff_n[7] a_6378_9520# 0.0133f
C1494 a_4882_4138# a_5374_4500# 0.0658f
C1495 a_3970_4138# a_4274_4178# 0.0931f
C1496 a_2275_4162# a_6982_4138# 0.399f
C1497 m3_16924_18146# ctop 0.209f
C1498 vcm a_18938_8154# 0.1f
C1499 m2_3164_12418# row_n[10] 0.0128f
C1500 m2_1732_17010# m2_2160_17438# 0.165f
C1501 a_16018_9158# a_17022_9158# 0.843f
C1502 m2_9188_8402# row_n[6] 0.0128f
C1503 a_2475_9182# a_31078_9158# 0.316f
C1504 rowoff_n[13] a_13406_15544# 0.0133f
C1505 m2_15212_4386# row_n[2] 0.0128f
C1506 row_n[10] a_5886_12170# 0.0437f
C1507 m2_34864_15002# a_35398_15222# 0.087f
C1508 col[5] a_2275_11190# 0.0899f
C1509 vcm a_6282_17230# 0.155f
C1510 col_n[8] a_11398_16548# 0.0283f
C1511 rowon_n[14] a_4974_16186# 0.248f
C1512 VDD a_4370_7512# 0.0779f
C1513 m2_34864_3958# m3_34996_4090# 3.79f
C1514 col_n[31] a_34394_7190# 0.084f
C1515 rowoff_n[5] a_15414_7512# 0.0133f
C1516 col[27] a_30074_5142# 0.367f
C1517 ctop a_19030_12170# 4.11f
C1518 a_5886_18194# a_5978_18194# 0.0991f
C1519 a_2275_18218# a_7286_18234# 0.145f
C1520 VDD a_27974_17190# 0.181f
C1521 row_n[0] a_15926_2130# 0.0437f
C1522 a_35002_2130# a_35094_2130# 0.0991f
C1523 a_34090_2130# a_34394_2170# 0.0931f
C1524 rowon_n[4] a_15014_6146# 0.248f
C1525 col_n[10] row_n[14] 0.298f
C1526 vcm row_n[9] 0.616f
C1527 sample row_n[8] 0.423f
C1528 col_n[22] col_n[23] 0.0101f
C1529 col_n[0] rowon_n[8] 0.111f
C1530 col_n[11] rowon_n[14] 0.111f
C1531 col_n[9] rowon_n[13] 0.111f
C1532 col_n[12] row_n[15] 0.298f
C1533 col_n[2] row_n[10] 0.298f
C1534 col_n[6] row_n[12] 0.298f
C1535 col_n[13] rowon_n[15] 0.111f
C1536 col_n[5] rowon_n[11] 0.111f
C1537 col_n[8] row_n[13] 0.298f
C1538 VDD rowon_n[7] 3.04f
C1539 col_n[3] rowon_n[10] 0.111f
C1540 col_n[7] rowon_n[12] 0.111f
C1541 col_n[4] row_n[11] 0.298f
C1542 col_n[1] rowon_n[9] 0.111f
C1543 sample_n rowoff_n[15] 0.142f
C1544 col[25] a_2475_10186# 0.136f
C1545 a_2275_6170# a_22042_6146# 0.399f
C1546 rowoff_n[3] a_24450_5504# 0.0133f
C1547 vcm a_33998_12170# 0.1f
C1548 a_6982_11166# a_6982_10162# 0.843f
C1549 col_n[15] rowoff_n[11] 0.0471f
C1550 VDD a_30074_2130# 0.483f
C1551 m2_24248_17438# row_n[15] 0.0128f
C1552 rowon_n[6] a_3878_8154# 0.118f
C1553 m2_30272_13422# row_n[11] 0.0128f
C1554 m2_35292_9406# row_n[7] 0.0128f
C1555 col_n[22] a_25358_5182# 0.084f
C1556 VDD a_19430_11528# 0.0779f
C1557 col_n[6] a_8990_16186# 0.251f
C1558 ctop a_34090_16186# 4.06f
C1559 col_n[3] a_5886_6146# 0.0765f
C1560 m3_1864_13126# a_2966_13174# 0.0302f
C1561 col_n[13] a_15926_18194# 0.0762f
C1562 a_2275_3158# a_12306_3174# 0.144f
C1563 a_2475_3158# a_14922_3134# 0.264f
C1564 rowoff_n[1] a_33486_3496# 0.0133f
C1565 rowoff_n[8] a_16018_10162# 0.294f
C1566 a_28066_1126# a_2475_1150# 0.0299f
C1567 row_n[13] a_26058_15182# 0.282f
C1568 rowoff_n[11] a_19942_13174# 0.202f
C1569 a_19030_8154# a_19334_8194# 0.0931f
C1570 a_19942_8154# a_20434_8516# 0.0658f
C1571 vcm a_14922_15182# 0.1f
C1572 a_31078_13174# a_32082_13174# 0.843f
C1573 col[22] a_2275_13198# 0.0899f
C1574 VDD a_10998_5142# 0.483f
C1575 a_24962_1126# VDD 0.405f
C1576 col[27] a_2275_2154# 0.0899f
C1577 row_n[15] a_13310_17230# 0.0117f
C1578 a_2275_17214# a_15926_17190# 0.136f
C1579 VDD a_34490_15544# 0.0779f
C1580 rowoff_n[6] a_25054_8154# 0.294f
C1581 col[16] a_19030_3134# 0.367f
C1582 a_2475_5166# a_29982_5142# 0.264f
C1583 row_n[5] a_23350_7190# 0.0117f
C1584 a_15926_5142# a_16018_5142# 0.326f
C1585 a_2275_5166# a_27366_5182# 0.144f
C1586 col[26] a_29070_15182# 0.367f
C1587 col[23] a_25966_5142# 0.0682f
C1588 m3_12908_1078# m3_13912_1078# 0.202f
C1589 col_n[0] rowoff_n[12] 0.0471f
C1590 m2_33284_16434# a_33086_16186# 0.165f
C1591 m2_13780_946# col_n[11] 0.331f
C1592 rowoff_n[4] a_34090_6146# 0.294f
C1593 a_22042_15182# a_22042_14178# 0.843f
C1594 m2_24824_946# a_2275_1150# 0.28f
C1595 m3_11904_1078# a_12002_2130# 0.0302f
C1596 a_2475_14202# a_7986_14178# 0.316f
C1597 m2_9764_946# a_9902_1126# 0.225f
C1598 row_n[7] a_13918_9158# 0.0437f
C1599 VDD a_26058_9158# 0.483f
C1600 m2_1732_7974# m3_1864_7102# 0.0341f
C1601 rowon_n[11] a_13006_13174# 0.248f
C1602 VDD a_15414_18556# 0.0858f
C1603 col_n[11] a_14314_3174# 0.084f
C1604 col_n[12] a_2475_9182# 0.0531f
C1605 a_2275_2154# a_20946_2130# 0.136f
C1606 a_10906_2130# a_11302_2170# 0.0313f
C1607 col_n[21] a_24354_15222# 0.084f
C1608 m2_18224_1374# VDD 0.0209f
C1609 vcm a_32082_4138# 0.56f
C1610 row_n[9] a_1957_11190# 0.187f
C1611 rowon_n[1] a_23046_3134# 0.248f
C1612 col_n[2] a_4882_16186# 0.0765f
C1613 a_35002_12170# a_35494_12532# 0.0658f
C1614 m2_9764_18014# a_9994_18194# 0.0249f
C1615 col[2] a_2475_6170# 0.136f
C1616 a_12002_16186# a_13006_16186# 0.843f
C1617 a_2475_16210# a_23046_16186# 0.316f
C1618 VDD a_6982_12170# 0.483f
C1619 a_28370_1166# m2_27836_946# 0.087f
C1620 m2_6752_18014# col_n[4] 0.243f
C1621 a_2275_4162# a_34394_4178# 0.144f
C1622 m2_1732_5966# a_2161_6170# 0.0454f
C1623 vcm a_13006_7150# 0.56f
C1624 rowoff_n[12] a_7894_14178# 0.202f
C1625 a_30986_9158# a_31078_9158# 0.326f
C1626 col_n[9] a_2275_12194# 0.113f
C1627 col[15] a_18026_13174# 0.367f
C1628 row_n[10] a_34090_12170# 0.282f
C1629 m2_24248_14426# a_24050_14178# 0.165f
C1630 row_n[5] rowoff_n[4] 0.085f
C1631 col[12] a_14922_3134# 0.0682f
C1632 col_n[14] a_2275_1150# 0.113f
C1633 vcm a_1957_16210# 0.139f
C1634 a_2275_13198# a_14010_13174# 0.399f
C1635 rowon_n[14] a_33998_16186# 0.118f
C1636 col[22] a_24962_15182# 0.0682f
C1637 col_n[30] a_33086_9158# 0.251f
C1638 VDD a_22042_16186# 0.483f
C1639 row_n[12] a_21342_14218# 0.0117f
C1640 col_n[29] a_2475_11190# 0.0531f
C1641 vcm a_3270_1166# 0.16f
C1642 a_25966_6146# a_26362_6186# 0.0313f
C1643 m2_34864_8978# a_2475_9182# 0.282f
C1644 m2_5172_3382# rowon_n[1] 0.0322f
C1645 col_n[10] a_13310_13214# 0.084f
C1646 vcm a_28066_11166# 0.56f
C1647 row_n[2] a_31382_4178# 0.0117f
C1648 a_2275_10186# a_4274_10202# 0.144f
C1649 a_2475_10186# a_6890_10162# 0.264f
C1650 row_n[14] a_11910_16186# 0.0437f
C1651 a_15014_15182# a_15318_15222# 0.0931f
C1652 a_15926_15182# a_16418_15544# 0.0658f
C1653 a_2275_15206# a_29070_15182# 0.399f
C1654 col[19] a_2475_8178# 0.136f
C1655 col_n[21] a_24450_7512# 0.0283f
C1656 row_n[4] a_21950_6146# 0.0437f
C1657 a_22042_3134# a_23046_3134# 0.843f
C1658 rowon_n[8] a_21038_10162# 0.248f
C1659 vcm a_18330_5182# 0.155f
C1660 rowon_n[10] rowoff_n[10] 20.2f
C1661 m2_14208_16434# rowon_n[14] 0.0322f
C1662 sample a_2161_1150# 0.0858f
C1663 m2_15212_12418# a_15014_12170# 0.165f
C1664 m2_20232_12418# rowon_n[10] 0.0322f
C1665 col_n[26] a_2275_14202# 0.113f
C1666 vcm a_8990_14178# 0.56f
C1667 m2_26256_8402# rowon_n[6] 0.0322f
C1668 a_11910_12170# a_12002_12170# 0.326f
C1669 m2_32280_4386# rowon_n[2] 0.0322f
C1670 a_2475_12194# a_21950_12170# 0.264f
C1671 a_2275_12194# a_19334_12210# 0.144f
C1672 VDD a_5886_4138# 0.181f
C1673 col_n[31] a_2275_3158# 0.113f
C1674 col[4] a_6982_11166# 0.367f
C1675 col[11] a_13918_13174# 0.0682f
C1676 col_n[19] a_22042_7150# 0.251f
C1677 a_13006_5142# a_13006_4138# 0.843f
C1678 col[16] a_2275_11190# 0.0899f
C1679 m2_34288_8402# a_34090_8154# 0.165f
C1680 col_n[26] a_28978_9158# 0.0765f
C1681 vcm a_33390_9198# 0.155f
C1682 m2_17796_18014# m2_18800_18014# 0.843f
C1683 a_6890_9158# a_7286_9198# 0.0313f
C1684 a_2275_9182# a_12914_9158# 0.136f
C1685 rowon_n[2] a_8898_4138# 0.118f
C1686 ctop a_12002_3134# 4.11f
C1687 vcm a_24050_18194# 0.165f
C1688 a_2275_14202# a_35398_14218# 0.145f
C1689 VDD a_20946_8154# 0.181f
C1690 m2_1732_4962# m3_1864_4090# 0.0341f
C1691 col_n[16] rowon_n[11] 0.111f
C1692 col_n[3] row_n[5] 0.298f
C1693 col_n[21] row_n[14] 0.298f
C1694 col_n[6] rowon_n[6] 0.111f
C1695 col_n[2] rowon_n[4] 0.111f
C1696 col_n[20] rowon_n[13] 0.111f
C1697 col_n[0] row_n[3] 0.298f
C1698 col_n[9] row_n[8] 0.298f
C1699 col_n[10] rowon_n[8] 0.111f
C1700 col_n[15] row_n[11] 0.298f
C1701 col_n[4] rowon_n[5] 0.111f
C1702 col_n[24] rowon_n[15] 0.111f
C1703 col_n[19] row_n[13] 0.298f
C1704 sample rowon_n[2] 0.0935f
C1705 col_n[1] row_n[4] 0.298f
C1706 col_n[5] row_n[6] 0.298f
C1707 col_n[13] row_n[10] 0.298f
C1708 col_n[7] row_n[7] 0.298f
C1709 vcm rowon_n[3] 0.65f
C1710 col_n[22] rowon_n[14] 0.111f
C1711 col_n[14] rowon_n[10] 0.111f
C1712 col_n[17] row_n[12] 0.298f
C1713 col_n[12] rowon_n[9] 0.111f
C1714 col_n[11] row_n[9] 0.298f
C1715 col_n[8] rowon_n[7] 0.111f
C1716 col_n[18] rowon_n[12] 0.111f
C1717 VDD row_n[2] 3.29f
C1718 col_n[23] row_n[15] 0.298f
C1719 a_25966_2130# a_26458_2492# 0.0658f
C1720 a_25054_2130# a_25358_2170# 0.0931f
C1721 col_n[10] a_13406_5504# 0.0283f
C1722 m3_15920_1078# VDD 0.0157f
C1723 row_n[9] a_29374_11206# 0.0117f
C1724 vcm a_26970_3134# 0.1f
C1725 col_n[26] rowoff_n[11] 0.0471f
C1726 a_2475_6170# a_4974_6146# 0.316f
C1727 col_n[20] a_23446_17552# 0.0283f
C1728 m2_6176_10410# a_5978_10162# 0.165f
C1729 rowoff_n[3] a_6890_5142# 0.202f
C1730 vcm a_14314_12210# 0.155f
C1731 a_2275_11190# a_27974_11166# 0.136f
C1732 VDD a_12402_2492# 0.0779f
C1733 m2_28840_18014# a_29070_18194# 0.0249f
C1734 col_n[6] a_2475_7174# 0.0531f
C1735 ctop a_27062_7150# 4.11f
C1736 a_26970_16186# a_27062_16186# 0.326f
C1737 row_n[11] a_19942_13174# 0.0437f
C1738 m2_26832_18014# m3_27968_18146# 0.0341f
C1739 rowon_n[15] a_19030_17190# 0.248f
C1740 row_n[1] a_29982_3134# 0.0437f
C1741 rowoff_n[1] a_15926_3134# 0.202f
C1742 m2_25252_6394# a_25054_6146# 0.165f
C1743 rowon_n[5] a_29070_7150# 0.248f
C1744 vcm a_7894_6146# 0.1f
C1745 a_28066_9158# a_28066_8154# 0.843f
C1746 a_2475_8178# a_20034_8154# 0.316f
C1747 col_n[8] a_10998_5142# 0.251f
C1748 col_n[18] a_21038_17190# 0.251f
C1749 vcm a_29374_16226# 0.155f
C1750 col_n[15] a_17934_7150# 0.0765f
C1751 a_21950_13174# a_22346_13214# 0.0313f
C1752 VDD a_27462_6508# 0.0779f
C1753 ctop a_7986_10162# 4.11f
C1754 VDD a_16930_15182# 0.181f
C1755 rowoff_n[6] a_7382_8516# 0.0133f
C1756 m2_3164_2378# row_n[0] 0.0128f
C1757 col_n[3] a_2275_10186# 0.113f
C1758 col_n[10] rowoff_n[12] 0.0471f
C1759 row_n[5] a_6982_7150# 0.282f
C1760 a_5978_5142# a_6282_5182# 0.0931f
C1761 a_6890_5142# a_7382_5504# 0.0658f
C1762 a_2275_5166# a_10998_5142# 0.399f
C1763 m2_30848_946# m3_30980_1078# 3.79f
C1764 m3_1864_13126# m3_1864_12122# 0.202f
C1765 rowon_n[9] a_6890_11166# 0.118f
C1766 vcm a_22954_10162# 0.1f
C1767 a_18026_10162# a_19030_10162# 0.843f
C1768 a_2475_10186# a_35094_10162# 0.0299f
C1769 col_n[9] a_12402_15544# 0.0283f
C1770 rowoff_n[4] a_16418_6508# 0.0133f
C1771 m2_20808_946# a_21038_2130# 0.843f
C1772 col[28] a_31078_4138# 0.367f
C1773 VDD a_8386_9520# 0.0779f
C1774 m2_25828_18014# ctop 0.0422f
C1775 col_n[23] a_2475_9182# 0.0531f
C1776 ctop a_23046_14178# 4.11f
C1777 m2_13204_15430# row_n[13] 0.0128f
C1778 m2_19228_11414# row_n[9] 0.0128f
C1779 m2_16216_4386# a_16018_4138# 0.165f
C1780 m2_25252_7398# row_n[5] 0.0128f
C1781 m2_31276_3382# row_n[1] 0.0128f
C1782 rowoff_n[9] a_7986_11166# 0.294f
C1783 a_2275_7174# a_26058_7150# 0.399f
C1784 rowoff_n[2] a_25454_4500# 0.0133f
C1785 col[8] a_2475_17214# 0.136f
C1786 col[13] a_2475_6170# 0.136f
C1787 a_8990_12170# a_8990_11166# 0.843f
C1788 col_n[23] a_26362_4178# 0.084f
C1789 VDD a_34090_4138# 0.483f
C1790 col_n[7] a_9994_15182# 0.251f
C1791 a_2966_16186# a_3970_16186# 0.843f
C1792 a_2275_16210# a_4882_16186# 0.136f
C1793 col_n[4] a_6890_5142# 0.0765f
C1794 VDD a_23446_13536# 0.0779f
C1795 row_n[8] a_27974_10162# 0.0437f
C1796 col_n[14] a_16930_17190# 0.0765f
C1797 ctop a_3970_17190# 4.06f
C1798 rowoff_n[0] a_34490_2492# 0.0133f
C1799 rowoff_n[7] a_17022_9158# 0.294f
C1800 rowon_n[12] a_27062_14178# 0.248f
C1801 a_2475_4162# a_18938_4138# 0.264f
C1802 a_2275_4162# a_16322_4178# 0.144f
C1803 col_n[20] a_2275_12194# 0.113f
C1804 m3_1864_5094# ctop 0.21f
C1805 ctop rowoff_n[6] 0.177f
C1806 row_n[1] rowoff_n[1] 0.209f
C1807 col_n[25] a_2275_1150# 0.113f
C1808 rowoff_n[13] a_24050_15182# 0.294f
C1809 a_21038_9158# a_21342_9198# 0.0931f
C1810 a_21950_9158# a_22442_9520# 0.0658f
C1811 vcm a_18938_17190# 0.1f
C1812 a_33086_14178# a_34090_14178# 0.843f
C1813 VDD a_15014_7150# 0.483f
C1814 rowoff_n[5] a_26058_7150# 0.294f
C1815 m2_2736_1950# m3_1864_2082# 0.0341f
C1816 a_2275_18218# a_19942_18194# 0.136f
C1817 VDD a_4370_16548# 0.0779f
C1818 col[17] a_20034_2130# 0.367f
C1819 col[10] a_2275_9182# 0.0899f
C1820 col_n[31] a_34394_16226# 0.084f
C1821 a_2275_1150# a_9902_1126# 0.136f
C1822 row_n[12] a_4974_14178# 0.282f
C1823 col[27] a_30074_14178# 0.367f
C1824 col[24] a_26970_4138# 0.0682f
C1825 vcm a_21038_2130# 0.56f
C1826 a_2475_6170# a_33998_6146# 0.264f
C1827 a_2275_6170# a_31382_6186# 0.144f
C1828 a_17934_6146# a_18026_6146# 0.326f
C1829 rowoff_n[3] a_35094_5142# 0.0135f
C1830 row_n[2] a_15014_4138# 0.282f
C1831 VDD a_5278_1166# 0.0149f
C1832 col[30] a_2475_8178# 0.136f
C1833 rowon_n[6] a_14922_8154# 0.118f
C1834 a_24050_16186# a_24050_15182# 0.843f
C1835 a_2475_15206# a_12002_15182# 0.316f
C1836 VDD a_30074_11166# 0.483f
C1837 col_n[12] a_15318_2170# 0.084f
C1838 col_n[22] a_25358_14218# 0.084f
C1839 row_n[4] a_3878_6146# 0.0437f
C1840 a_2275_3158# a_24962_3134# 0.136f
C1841 a_12914_3134# a_13310_3174# 0.0313f
C1842 rowon_n[8] a_2966_10162# 0.248f
C1843 a_2475_18218# a_17934_18194# 0.264f
C1844 col_n[3] a_5886_15182# 0.0765f
C1845 vcm a_2475_5166# 1.08f
C1846 rowoff_n[11] a_30474_13536# 0.0133f
C1847 a_2275_12194# a_2874_12170# 0.136f
C1848 a_2475_12194# a_3878_12170# 0.264f
C1849 m2_1732_18014# VDD 1.32f
C1850 row_n[15] a_25966_17190# 0.0437f
C1851 a_14010_17190# a_15014_17190# 0.843f
C1852 a_2475_17214# a_27062_17190# 0.316f
C1853 VDD a_10998_14178# 0.483f
C1854 col[27] a_2275_11190# 0.0899f
C1855 rowon_n[0] a_2475_2154# 0.31f
C1856 m3_31984_18146# a_32082_17190# 0.0303f
C1857 row_n[5] a_34394_7190# 0.0117f
C1858 col[16] a_19030_12170# 0.367f
C1859 rowon_n[9] a_35094_11166# 0.0141f
C1860 col[13] a_15926_2130# 0.0682f
C1861 vcm a_17022_9158# 0.56f
C1862 a_32994_10162# a_33086_10162# 0.326f
C1863 rowoff_n[14] a_12002_16186# 0.294f
C1864 col[23] a_25966_14178# 0.0682f
C1865 col_n[17] rowon_n[6] 0.111f
C1866 col_n[28] row_n[12] 0.298f
C1867 col_n[23] rowon_n[9] 0.111f
C1868 col_n[12] row_n[4] 0.298f
C1869 col_n[22] row_n[9] 0.298f
C1870 col_n[24] row_n[10] 0.298f
C1871 col_n[6] row_n[1] 0.298f
C1872 col_n[25] rowon_n[10] 0.111f
C1873 col_n[19] rowon_n[7] 0.111f
C1874 col_n[5] rowon_n[0] 0.111f
C1875 col_n[10] row_n[3] 0.298f
C1876 col_n[30] row_n[13] 0.298f
C1877 col_n[20] row_n[8] 0.298f
C1878 col_n[21] rowon_n[8] 0.111f
C1879 col_n[11] rowon_n[3] 0.111f
C1880 col_n[1] ctop 0.06f
C1881 col_n[29] rowon_n[12] 0.111f
C1882 col_n[4] row_n[0] 0.298f
C1883 col_n[18] row_n[7] 0.298f
C1884 col_n[7] rowon_n[1] 0.111f
C1885 col_n[15] rowon_n[5] 0.111f
C1886 vcm en_C0_n 0.0192f
C1887 col_n[9] rowon_n[2] 0.111f
C1888 col_n[26] row_n[11] 0.298f
C1889 col_n[31] rowon_n[13] 0.111f
C1890 col_n[14] row_n[5] 0.298f
C1891 col_n[27] rowon_n[11] 0.111f
C1892 col_n[13] rowon_n[4] 0.111f
C1893 VDD en_bit_n[0] 0.206f
C1894 col_n[16] row_n[6] 0.298f
C1895 col_n[8] row_n[2] 0.298f
C1896 a_2275_14202# a_18026_14178# 0.399f
C1897 VDD a_2275_8178# 1.95f
C1898 col_n[31] a_34090_8154# 0.251f
C1899 VDD a_26058_18194# 0.0356f
C1900 a_2475_2154# a_32082_2130# 0.316f
C1901 a_34090_3134# a_34090_2130# 0.843f
C1902 m3_11904_18146# VDD 0.0671f
C1903 col_n[11] a_14314_12210# 0.084f
C1904 vcm a_7286_3174# 0.155f
C1905 row_n[9] a_13006_11166# 0.282f
C1906 a_27974_7150# a_28370_7190# 0.0313f
C1907 rowon_n[13] a_12914_15182# 0.118f
C1908 col_n[17] a_2475_7174# 0.0531f
C1909 vcm a_32082_13174# 0.56f
C1910 a_2475_11190# a_10906_11166# 0.264f
C1911 a_2275_11190# a_8290_11206# 0.144f
C1912 VDD a_28978_3134# 0.181f
C1913 m2_15788_18014# a_16322_18234# 0.087f
C1914 col_n[22] a_25454_6508# 0.0283f
C1915 a_17022_16186# a_17326_16226# 0.0931f
C1916 a_2275_16210# a_33086_16186# 0.399f
C1917 a_17934_16186# a_18426_16548# 0.0658f
C1918 rowon_n[3] a_22954_5142# 0.118f
C1919 m2_3740_18014# m3_2868_18146# 0.0341f
C1920 m2_3164_14426# rowon_n[12] 0.0322f
C1921 col[2] a_2475_15206# 0.136f
C1922 m2_9188_10410# rowon_n[8] 0.0322f
C1923 m2_15212_6394# rowon_n[4] 0.0322f
C1924 col[7] a_2475_4162# 0.136f
C1925 a_24050_4138# a_25054_4138# 0.843f
C1926 row_n[1] a_10298_3174# 0.0117f
C1927 vcm a_22346_7190# 0.155f
C1928 a_2475_8178# a_1957_8178# 0.0734f
C1929 rowoff_n[12] a_18426_14540# 0.0133f
C1930 m2_23820_946# col_n[21] 0.331f
C1931 col[5] a_7986_10162# 0.367f
C1932 vcm a_13006_16186# 0.56f
C1933 a_2275_13198# a_23350_13214# 0.144f
C1934 a_13918_13174# a_14010_13174# 0.326f
C1935 a_2475_13198# a_25966_13174# 0.264f
C1936 VDD a_9902_6146# 0.181f
C1937 col[12] a_14922_12170# 0.0682f
C1938 col_n[21] rowoff_n[12] 0.0471f
C1939 col_n[14] a_2275_10186# 0.113f
C1940 m2_21812_18014# col[19] 0.347f
C1941 row_n[12] a_33998_14178# 0.0437f
C1942 col_n[20] a_23046_6146# 0.251f
C1943 vcm a_15926_1126# 0.0989f
C1944 m2_30272_15430# rowon_n[13] 0.0322f
C1945 col_n[27] a_29982_8154# 0.0765f
C1946 m2_35292_11414# rowon_n[9] 0.0322f
C1947 a_15014_6146# a_15014_5142# 0.843f
C1948 m3_8892_18146# m3_9896_18146# 0.202f
C1949 m2_5748_946# m3_6884_1078# 0.0341f
C1950 vcm a_3270_10202# 0.155f
C1951 a_8898_10162# a_9294_10202# 0.0313f
C1952 a_2275_10186# a_16930_10162# 0.136f
C1953 col[4] a_2275_7174# 0.0899f
C1954 ctop a_16018_5142# 4.11f
C1955 VDD a_24962_10162# 0.181f
C1956 col_n[11] a_14410_4500# 0.0283f
C1957 a_27062_3134# a_27366_3174# 0.0931f
C1958 a_27974_3134# a_28466_3496# 0.0658f
C1959 col[19] a_2475_17214# 0.136f
C1960 col_n[21] a_24450_16548# 0.0283f
C1961 m2_1732_3958# a_2475_4162# 0.139f
C1962 col[24] a_2475_6170# 0.136f
C1963 vcm a_30986_5142# 0.1f
C1964 a_2475_7174# a_8990_7150# 0.316f
C1965 rowoff_n[2] a_7894_4138# 0.202f
C1966 a_4974_7150# a_5978_7150# 0.843f
C1967 rowoff_n[10] a_24962_12170# 0.202f
C1968 row_n[6] a_21038_8154# 0.282f
C1969 vcm a_18330_14218# 0.155f
C1970 a_2275_12194# a_31990_12170# 0.136f
C1971 VDD a_16418_4500# 0.0779f
C1972 rowon_n[10] a_20946_12170# 0.118f
C1973 col_n[5] rowoff_n[13] 0.0471f
C1974 sample a_2161_10186# 0.0858f
C1975 ctop a_31078_9158# 4.11f
C1976 row_n[0] m2_35292_2378# 0.0128f
C1977 a_28978_17190# a_29070_17190# 0.326f
C1978 VDD a_5886_13174# 0.181f
C1979 col_n[31] a_2275_12194# 0.113f
C1980 col[2] rowoff_n[3] 0.0901f
C1981 col[8] rowoff_n[9] 0.0901f
C1982 row_n[8] a_8290_10202# 0.0117f
C1983 col[4] rowoff_n[5] 0.0901f
C1984 col[1] rowoff_n[2] 0.0901f
C1985 col[7] rowoff_n[8] 0.0901f
C1986 col[0] rowoff_n[1] 0.0901f
C1987 col[5] rowoff_n[6] 0.0901f
C1988 col[6] rowoff_n[7] 0.0901f
C1989 col[3] rowoff_n[4] 0.0901f
C1990 rowon_n[0] a_30986_2130# 0.118f
C1991 rowoff_n[0] a_16930_2130# 0.202f
C1992 col_n[9] a_12002_4138# 0.251f
C1993 col_n[19] a_22042_16186# 0.251f
C1994 vcm a_11910_8154# 0.1f
C1995 m2_28840_18014# m2_29268_18442# 0.165f
C1996 a_2475_9182# a_24050_9158# 0.316f
C1997 rowoff_n[13] a_6378_15544# 0.0133f
C1998 a_30074_10162# a_30074_9158# 0.843f
C1999 col_n[16] a_18938_6146# 0.0765f
C2000 m2_30272_15430# a_30074_15182# 0.165f
C2001 vcm a_33390_18234# 0.16f
C2002 col_n[26] a_28978_18194# 0.0762f
C2003 col[21] a_2275_9182# 0.0899f
C2004 a_23958_14178# a_24354_14218# 0.0313f
C2005 VDD a_31478_8516# 0.0779f
C2006 rowoff_n[5] a_8386_7512# 0.0133f
C2007 ctop a_12002_12170# 4.11f
C2008 row_n[0] a_8898_2130# 0.0437f
C2009 VDD a_20946_17190# 0.181f
C2010 rowon_n[4] a_7986_6146# 0.248f
C2011 m2_1732_6970# m2_1732_5966# 0.843f
C2012 vcm a_2966_2130# 0.165f
C2013 a_8898_6146# a_9390_6508# 0.0658f
C2014 a_2275_6170# a_15014_6146# 0.399f
C2015 a_7986_6146# a_8290_6186# 0.0931f
C2016 col_n[10] a_13406_14540# 0.0283f
C2017 rowoff_n[3] a_17422_5504# 0.0133f
C2018 vcm a_26970_12170# 0.1f
C2019 a_20034_11166# a_21038_11166# 0.843f
C2020 col[29] a_32082_3134# 0.367f
C2021 VDD a_23046_2130# 0.483f
C2022 m2_2160_13422# row_n[11] 0.0194f
C2023 m2_1732_17010# a_1957_17214# 0.245f
C2024 m2_8184_9406# row_n[7] 0.0128f
C2025 m2_14208_5390# row_n[3] 0.0128f
C2026 VDD a_12402_11528# 0.0779f
C2027 col_n[6] a_2475_16210# 0.0531f
C2028 ctop a_27062_16186# 4.11f
C2029 col_n[11] a_2475_5166# 0.0531f
C2030 a_2275_3158# a_5278_3174# 0.144f
C2031 a_3878_3134# a_4274_3174# 0.0313f
C2032 a_2475_3158# a_7894_3134# 0.264f
C2033 a_4882_3134# a_4974_3134# 0.326f
C2034 rowoff_n[1] a_26458_3496# 0.0133f
C2035 rowoff_n[8] a_8990_10162# 0.294f
C2036 row_n[13] a_19030_15182# 0.282f
C2037 rowoff_n[11] a_12914_13174# 0.202f
C2038 a_2275_8178# a_30074_8154# 0.399f
C2039 col_n[24] a_27366_3174# 0.084f
C2040 m2_21236_13422# a_21038_13174# 0.165f
C2041 vcm a_7894_15182# 0.1f
C2042 a_10998_13174# a_10998_12170# 0.843f
C2043 col_n[8] a_10998_14178# 0.251f
C2044 VDD a_3970_5142# 0.483f
C2045 row_n[3] a_29070_5142# 0.282f
C2046 col_n[5] a_7894_4138# 0.0765f
C2047 row_n[15] a_6282_17230# 0.0117f
C2048 col[1] a_2475_2154# 0.136f
C2049 m2_29268_14426# row_n[12] 0.0128f
C2050 rowon_n[7] a_28978_9158# 0.118f
C2051 col_n[15] a_17934_16186# 0.0765f
C2052 a_4882_17190# a_5278_17230# 0.0313f
C2053 a_2275_17214# a_8898_17190# 0.136f
C2054 rowoff_n[6] a_18026_8154# 0.294f
C2055 VDD a_27462_15544# 0.0779f
C2056 m2_34864_9982# row_n[8] 0.267f
C2057 a_2275_5166# a_20338_5182# 0.144f
C2058 a_2475_5166# a_22954_5142# 0.264f
C2059 row_n[5] a_16322_7190# 0.0117f
C2060 m3_1864_2082# m3_2868_2082# 0.202f
C2061 m3_34996_3086# m3_34996_2082# 0.202f
C2062 col_n[12] ctop 0.0594f
C2063 col_n[17] row_n[1] 0.298f
C2064 col_n[29] row_n[7] 0.298f
C2065 col_n[26] rowon_n[5] 0.111f
C2066 VDD col[9] 3.83f
C2067 rowon_n[12] rowon_n[11] 0.0632f
C2068 col_n[21] row_n[3] 0.298f
C2069 col_n[30] rowon_n[7] 0.111f
C2070 col_n[18] rowon_n[1] 0.111f
C2071 col_n[22] rowon_n[3] 0.111f
C2072 col_n[19] row_n[2] 0.298f
C2073 col_n[23] row_n[4] 0.298f
C2074 col_n[27] row_n[6] 0.298f
C2075 col_n[24] rowon_n[4] 0.111f
C2076 col_n[25] row_n[5] 0.298f
C2077 col_n[20] rowon_n[2] 0.111f
C2078 col_n[31] row_n[8] 0.298f
C2079 vcm col[6] 5.46f
C2080 col_n[28] rowon_n[6] 0.111f
C2081 col_n[15] row_n[0] 0.297f
C2082 col_n[3] col[3] 0.489f
C2083 col_n[16] rowon_n[0] 0.111f
C2084 a_25966_1126# a_26058_1126# 0.0991f
C2085 a_23958_10162# a_24450_10524# 0.0658f
C2086 rowoff_n[15] a_28978_17190# 0.202f
C2087 col_n[8] a_2275_8178# 0.113f
C2088 a_23046_10162# a_23350_10202# 0.0931f
C2089 rowoff_n[4] a_27062_6146# 0.294f
C2090 m2_4744_946# a_4974_1126# 0.0249f
C2091 m2_10768_946# a_2475_1150# 0.286f
C2092 row_n[7] a_6890_9158# 0.0437f
C2093 VDD a_19030_9158# 0.483f
C2094 rowon_n[11] a_5978_13174# 0.248f
C2095 col[28] a_31078_13174# 0.367f
C2096 VDD a_8386_18556# 0.0858f
C2097 col[25] a_27974_3134# 0.0682f
C2098 a_2275_2154# a_13918_2130# 0.136f
C2099 col_n[28] a_2475_7174# 0.0531f
C2100 vcm a_25054_4138# 0.56f
C2101 a_2275_7174# a_2275_6170# 0.0715f
C2102 rowon_n[1] a_16018_3134# 0.248f
C2103 a_19942_7150# a_20034_7150# 0.326f
C2104 m2_12200_11414# a_12002_11166# 0.165f
C2105 col_n[13] a_16322_1166# 0.0839f
C2106 col[13] a_2475_15206# 0.136f
C2107 a_26058_17190# a_26058_16186# 0.843f
C2108 a_2475_16210# a_16018_16186# 0.316f
C2109 VDD a_34090_13174# 0.483f
C2110 col_n[23] a_26362_13214# 0.084f
C2111 col[18] a_2475_4162# 0.136f
C2112 col_n[4] a_6890_14178# 0.0765f
C2113 a_2275_4162# a_28978_4138# 0.136f
C2114 a_14922_4138# a_15318_4178# 0.0313f
C2115 m2_31276_7398# a_31078_7150# 0.165f
C2116 vcm a_5978_7150# 0.56f
C2117 row_n[10] a_27062_12170# 0.282f
C2118 col_n[25] a_2275_10186# 0.113f
C2119 m2_1732_15002# sample 0.2f
C2120 rowon_n[14] a_26970_16186# 0.118f
C2121 a_3970_13174# a_4274_13214# 0.0931f
C2122 a_4882_13174# a_5374_13536# 0.0658f
C2123 a_2275_13198# a_6982_13174# 0.399f
C2124 m2_34864_8978# ctop 0.0422f
C2125 VDD a_15014_16186# 0.483f
C2126 a_2475_1150# a_21038_1126# 0.0299f
C2127 row_n[12] a_14314_14218# 0.0117f
C2128 col[10] a_2275_18218# 0.0899f
C2129 col[17] a_20034_11166# 0.367f
C2130 vcm a_30378_2170# 0.155f
C2131 col[14] a_16930_1126# 0.0682f
C2132 col[15] a_2275_7174# 0.0899f
C2133 col[24] a_26970_13174# 0.0682f
C2134 row_n[2] a_24354_4178# 0.0117f
C2135 vcm a_21038_11166# 0.56f
C2136 a_34090_11166# a_34394_11206# 0.0931f
C2137 a_35002_11166# a_35094_11166# 0.0991f
C2138 VDD a_17934_1126# 0.403f
C2139 row_n[14] a_4882_16186# 0.0437f
C2140 a_2275_15206# a_22042_15182# 0.399f
C2141 col[30] a_2475_17214# 0.136f
C2142 row_n[4] a_14922_6146# 0.0437f
C2143 col_n[12] a_15318_11206# 0.084f
C2144 rowon_n[8] a_14010_10162# 0.248f
C2145 a_2475_3158# a_2475_2154# 0.0666f
C2146 m2_22240_5390# a_22042_5142# 0.165f
C2147 vcm a_11302_5182# 0.155f
C2148 a_29982_8154# a_30378_8194# 0.0313f
C2149 col_n[16] rowoff_n[13] 0.0471f
C2150 row_n[6] a_2966_8154# 0.281f
C2151 vcm a_2475_14202# 1.08f
C2152 a_2475_12194# a_14922_12170# 0.264f
C2153 m2_4168_4386# rowon_n[2] 0.0322f
C2154 a_2275_12194# a_12306_12210# 0.144f
C2155 VDD a_32994_5142# 0.181f
C2156 rowon_n[10] a_2275_12194# 1.79f
C2157 col_n[23] a_26458_5504# 0.0283f
C2158 col_n[5] a_2475_3158# 0.0531f
C2159 col[19] rowoff_n[9] 0.0901f
C2160 col[13] rowoff_n[3] 0.0901f
C2161 col[18] rowoff_n[8] 0.0901f
C2162 col[17] rowoff_n[7] 0.0901f
C2163 col[15] rowoff_n[5] 0.0901f
C2164 col[12] rowoff_n[2] 0.0901f
C2165 m2_23244_18442# VDD 0.0456f
C2166 col[16] rowoff_n[6] 0.0901f
C2167 col[10] rowoff_n[0] 0.0901f
C2168 col[11] rowoff_n[1] 0.0901f
C2169 col[14] rowoff_n[4] 0.0901f
C2170 a_19942_17190# a_20434_17552# 0.0658f
C2171 a_19030_17190# a_19334_17230# 0.0931f
C2172 a_2475_1150# m2_1732_946# 0.139f
C2173 a_26058_5142# a_27062_5142# 0.843f
C2174 col[6] a_8990_9158# 0.367f
C2175 vcm a_26362_9198# 0.155f
C2176 m2_10768_18014# m2_11772_18014# 0.843f
C2177 a_2275_9182# a_5886_9158# 0.136f
C2178 ctop a_4974_3134# 4.11f
C2179 vcm a_17022_18194# 0.165f
C2180 col[13] a_15926_11166# 0.0682f
C2181 m2_13204_17438# rowon_n[15] 0.0322f
C2182 a_15926_14178# a_16018_14178# 0.326f
C2183 a_2475_14202# a_29982_14178# 0.264f
C2184 a_2275_14202# a_27366_14218# 0.144f
C2185 VDD a_13918_8154# 0.181f
C2186 row_n[7] a_35094_9158# 0.0123f
C2187 m2_19228_13422# rowon_n[11] 0.0322f
C2188 m2_25252_9406# rowon_n[7] 0.0322f
C2189 m2_31276_5390# rowon_n[3] 0.0322f
C2190 rowon_n[11] a_35002_13174# 0.118f
C2191 m2_22816_946# vcm 0.353f
C2192 col_n[21] a_24050_5142# 0.251f
C2193 VDD a_2275_17214# 1.96f
C2194 col_n[31] a_34090_17190# 0.251f
C2195 col_n[2] a_2275_6170# 0.113f
C2196 col_n[28] a_30986_7150# 0.0765f
C2197 m2_13204_3382# a_13006_3134# 0.165f
C2198 vcm a_19942_3134# 0.1f
C2199 vcm rowoff_n[14] 0.533f
C2200 row_n[9] a_22346_11206# 0.0117f
C2201 col_n[1] a_4274_9198# 0.084f
C2202 a_17022_7150# a_17022_6146# 0.843f
C2203 vcm a_7286_12210# 0.155f
C2204 a_2275_11190# a_20946_11166# 0.136f
C2205 a_10906_11166# a_11302_11206# 0.0313f
C2206 VDD a_5374_2492# 0.0779f
C2207 col[3] rowoff_n[10] 0.0901f
C2208 col_n[17] a_2475_16210# 0.0531f
C2209 ctop a_20034_7150# 4.11f
C2210 col_n[22] a_2475_5166# 0.0531f
C2211 row_n[11] a_12914_13174# 0.0437f
C2212 VDD a_28978_12170# 0.181f
C2213 col_n[12] a_15414_3496# 0.0283f
C2214 m2_17796_18014# m3_17928_18146# 3.79f
C2215 rowon_n[15] a_12002_17190# 0.248f
C2216 col_n[22] a_25454_15544# 0.0283f
C2217 a_29070_4138# a_29374_4178# 0.0931f
C2218 a_29982_4138# a_30474_4500# 0.0658f
C2219 row_n[1] a_22954_3134# 0.0437f
C2220 rowoff_n[1] a_8898_3134# 0.202f
C2221 rowon_n[5] a_22042_7150# 0.248f
C2222 vcm a_35002_7150# 0.101f
C2223 col[7] a_2475_13198# 0.136f
C2224 a_6982_8154# a_7986_8154# 0.843f
C2225 a_2475_8178# a_13006_8154# 0.316f
C2226 rowoff_n[12] a_29070_14178# 0.294f
C2227 col_n[0] a_3366_9520# 0.0283f
C2228 col[12] a_2475_2154# 0.136f
C2229 vcm a_22346_16226# 0.155f
C2230 a_2275_13198# a_34394_13214# 0.144f
C2231 VDD a_20434_6508# 0.0779f
C2232 col[2] a_4882_9158# 0.0682f
C2233 a_30986_18194# a_31078_18194# 0.0991f
C2234 VDD a_9902_15182# 0.181f
C2235 vcm col[17] 5.46f
C2236 col_n[31] rowon_n[2] 0.111f
C2237 col_n[29] rowon_n[1] 0.111f
C2238 col_n[26] row_n[0] 0.298f
C2239 col_n[8] col[9] 7.13f
C2240 col_n[27] rowon_n[0] 0.111f
C2241 col_n[23] ctop 0.0594f
C2242 col_n[30] row_n[2] 0.298f
C2243 col_n[28] row_n[1] 0.298f
C2244 col_n[10] a_13006_3134# 0.251f
C2245 VDD col[20] 3.83f
C2246 rowon_n[9] row_n[9] 18.9f
C2247 col_n[19] a_2275_8178# 0.113f
C2248 a_2275_5166# a_3970_5142# 0.399f
C2249 col_n[20] a_23046_15182# 0.251f
C2250 m2_21812_946# m3_20940_1078# 0.0341f
C2251 col_n[17] a_19942_5142# 0.0765f
C2252 vcm a_15926_10162# 0.1f
C2253 a_32082_11166# a_32082_10162# 0.843f
C2254 a_2475_10186# a_28066_10162# 0.316f
C2255 col_n[27] a_29982_17190# 0.0765f
C2256 row_n[14] a_33086_16186# 0.282f
C2257 rowoff_n[4] a_9390_6508# 0.0133f
C2258 a_25966_15182# a_26362_15222# 0.0313f
C2259 VDD a_35494_10524# 0.106f
C2260 m2_11772_18014# ctop 0.0422f
C2261 col[4] a_2275_16210# 0.0899f
C2262 ctop a_16018_14178# 4.11f
C2263 col[9] a_2275_5166# 0.0899f
C2264 col_n[11] a_14410_13536# 0.0283f
C2265 m2_3164_3382# row_n[1] 0.0128f
C2266 a_2275_7174# a_19030_7150# 0.399f
C2267 a_10906_7150# a_11398_7512# 0.0658f
C2268 rowoff_n[2] a_18426_4500# 0.0133f
C2269 a_9994_7150# a_10298_7190# 0.0931f
C2270 rowoff_n[10] a_35494_12532# 0.0133f
C2271 col[30] a_33086_2130# 0.367f
C2272 row_n[6] a_30378_8194# 0.0117f
C2273 col[24] a_2475_15206# 0.136f
C2274 vcm a_30986_14178# 0.1f
C2275 a_22042_12170# a_23046_12170# 0.843f
C2276 VDD a_27062_4138# 0.483f
C2277 col[29] a_2475_4162# 0.136f
C2278 VDD a_16418_13536# 0.0779f
C2279 row_n[8] a_20946_10162# 0.0437f
C2280 rowoff_n[0] a_27462_2492# 0.0133f
C2281 rowoff_n[7] a_9994_9158# 0.294f
C2282 rowon_n[12] a_20034_14178# 0.248f
C2283 a_2475_4162# a_11910_4138# 0.264f
C2284 a_2275_4162# a_9294_4178# 0.144f
C2285 a_6890_4138# a_6982_4138# 0.326f
C2286 m3_31984_18146# ctop 0.209f
C2287 col_n[25] a_28370_2170# 0.084f
C2288 col_n[0] a_2475_1150# 0.0532f
C2289 m2_12200_16434# row_n[14] 0.0128f
C2290 m2_18224_12418# row_n[10] 0.0128f
C2291 rowoff_n[13] a_17022_15182# 0.294f
C2292 m2_24248_8402# row_n[6] 0.0128f
C2293 a_2275_9182# a_34090_9158# 0.399f
C2294 col_n[9] a_12002_13174# 0.251f
C2295 m2_30272_4386# row_n[2] 0.0128f
C2296 col_n[6] a_8898_3134# 0.0765f
C2297 rowon_n[2] a_30074_4138# 0.248f
C2298 vcm a_11910_17190# 0.1f
C2299 a_13006_14178# a_13006_13174# 0.843f
C2300 col_n[16] a_18938_15182# 0.0765f
C2301 VDD a_7986_7150# 0.483f
C2302 rowoff_n[5] a_19030_7150# 0.294f
C2303 a_2275_18218# a_12914_18194# 0.136f
C2304 a_6890_18194# a_7286_18234# 0.0313f
C2305 col[21] a_2275_18218# 0.0899f
C2306 VDD a_31478_17552# 0.0779f
C2307 a_2161_1150# a_2275_1150# 0.183f
C2308 col[26] a_2275_7174# 0.0899f
C2309 a_2475_1150# a_2966_1126# 0.0299f
C2310 vcm a_14010_2130# 0.56f
C2311 a_2475_6170# a_26970_6146# 0.264f
C2312 a_2275_6170# a_24354_6186# 0.144f
C2313 vcm a_2966_11166# 0.56f
C2314 row_n[2] a_7986_4138# 0.282f
C2315 rowoff_n[3] a_28066_5142# 0.294f
C2316 a_25966_11166# a_26458_11528# 0.0658f
C2317 a_25054_11166# a_25358_11206# 0.0931f
C2318 rowon_n[6] a_7894_8154# 0.118f
C2319 a_2475_15206# a_4974_15182# 0.316f
C2320 VDD a_23046_11166# 0.483f
C2321 col[29] a_32082_12170# 0.367f
C2322 col[26] a_28978_2130# 0.0682f
C2323 a_2275_3158# a_17934_3134# 0.136f
C2324 a_2475_18218# a_10906_18194# 0.264f
C2325 col_n[27] rowoff_n[13] 0.0471f
C2326 a_31078_1126# a_2275_1150# 0.0924f
C2327 row_n[13] a_28370_15222# 0.0117f
C2328 col_n[11] a_2475_14202# 0.0531f
C2329 vcm a_29070_6146# 0.56f
C2330 rowoff_n[11] a_23446_13536# 0.0133f
C2331 a_21950_8154# a_22042_8154# 0.326f
C2332 col_n[16] a_2475_3158# 0.0531f
C2333 col[29] rowoff_n[8] 0.0901f
C2334 col[21] rowoff_n[0] 0.0901f
C2335 col[25] rowoff_n[4] 0.0901f
C2336 col[23] rowoff_n[2] 0.0901f
C2337 col[28] rowoff_n[7] 0.0901f
C2338 col[22] rowoff_n[1] 0.0901f
C2339 col[30] rowoff_n[9] 0.0901f
C2340 col[26] rowoff_n[5] 0.0901f
C2341 col[27] rowoff_n[6] 0.0901f
C2342 col[24] rowoff_n[3] 0.0901f
C2343 col_n[24] a_27366_12210# 0.084f
C2344 a_28466_1488# VDD 0.0977f
C2345 col[7] a_2475_18218# 0.136f
C2346 row_n[15] a_18938_17190# 0.0437f
C2347 a_2475_17214# a_20034_17190# 0.316f
C2348 VDD a_3970_14178# 0.483f
C2349 col_n[5] a_7894_13174# 0.0765f
C2350 a_22042_2130# m2_22240_2378# 0.165f
C2351 col[1] a_2475_11190# 0.136f
C2352 a_16930_5142# a_17326_5182# 0.0313f
C2353 row_n[5] a_28978_7150# 0.0437f
C2354 a_2275_5166# a_32994_5142# 0.136f
C2355 rowon_n[9] a_28066_11166# 0.248f
C2356 vcm a_9994_9158# 0.56f
C2357 rowoff_n[14] a_4974_16186# 0.294f
C2358 m2_33860_946# a_2475_1150# 0.18f
C2359 m2_10768_946# a_11302_1166# 0.087f
C2360 m3_14916_1078# a_15014_2130# 0.0302f
C2361 a_2275_14202# a_10998_14178# 0.399f
C2362 col_n[8] a_2275_17214# 0.113f
C2363 a_5978_14178# a_6282_14218# 0.0931f
C2364 a_6890_14178# a_7382_14540# 0.0658f
C2365 col_n[13] a_2275_6170# 0.113f
C2366 col_n[11] rowoff_n[14] 0.0471f
C2367 VDD a_19030_18194# 0.0356f
C2368 col[18] a_21038_10162# 0.367f
C2369 a_2475_2154# a_25054_2130# 0.316f
C2370 a_13006_2130# a_14010_2130# 0.843f
C2371 m2_26832_946# VDD 1f
C2372 vcm a_35398_4178# 0.161f
C2373 col[25] a_27974_12170# 0.0682f
C2374 row_n[9] a_5978_11166# 0.282f
C2375 col[14] rowoff_n[10] 0.0901f
C2376 rowoff_n[9] a_29982_11166# 0.202f
C2377 col_n[28] a_2475_16210# 0.0531f
C2378 rowon_n[13] a_5886_15182# 0.118f
C2379 col_n[0] a_3270_6186# 0.084f
C2380 vcm a_25054_13174# 0.56f
C2381 VDD a_21950_3134# 0.181f
C2382 col[3] a_2275_3158# 0.0899f
C2383 m2_31852_18014# a_2275_18218# 0.28f
C2384 a_2275_16210# a_26058_16186# 0.399f
C2385 rowon_n[3] a_15926_5142# 0.118f
C2386 a_31990_1126# m2_31852_946# 0.225f
C2387 col_n[13] a_16322_10202# 0.084f
C2388 col[18] a_2475_13198# 0.136f
C2389 a_3970_4138# a_3970_3134# 0.843f
C2390 row_n[1] a_3270_3174# 0.0117f
C2391 col[23] a_2475_2154# 0.136f
C2392 vcm a_15318_7190# 0.155f
C2393 rowoff_n[12] a_11398_14540# 0.0133f
C2394 a_31990_9158# a_32386_9198# 0.0313f
C2395 col_n[24] a_27462_4500# 0.0283f
C2396 m2_27260_14426# a_27062_14178# 0.165f
C2397 ctop a_28066_2130# 4.06f
C2398 vcm a_5978_16186# 0.56f
C2399 a_2475_13198# a_18938_13174# 0.264f
C2400 a_2275_13198# a_16322_13214# 0.144f
C2401 VDD a_2161_6170# 0.187f
C2402 VDD col[31] 3.79f
C2403 vcm col[28] 5.46f
C2404 col_n[14] col[14] 0.489f
C2405 rowon_n[14] ctop 0.203f
C2406 m2_27836_18014# a_2475_18218# 0.286f
C2407 a_21950_18194# a_22442_18556# 0.0658f
C2408 col_n[30] a_2275_8178# 0.113f
C2409 a_16930_1126# a_17422_1488# 0.0658f
C2410 row_n[12] a_26970_14178# 0.0437f
C2411 vcm a_8898_1126# 0.0989f
C2412 m2_2160_15430# rowon_n[13] 0.0219f
C2413 m2_8184_11414# rowon_n[9] 0.0322f
C2414 col[7] a_9994_8154# 0.367f
C2415 a_28066_6146# a_29070_6146# 0.843f
C2416 m2_14208_7398# rowon_n[5] 0.0322f
C2417 m2_20232_3382# rowon_n[1] 0.0322f
C2418 vcm a_30378_11206# 0.155f
C2419 col[14] a_16930_10162# 0.0682f
C2420 a_2275_10186# a_9902_10162# 0.136f
C2421 col[15] a_2275_16210# 0.0899f
C2422 m2_34864_3958# VDD 0.772f
C2423 ctop a_8990_5142# 4.11f
C2424 col[20] a_2275_5166# 0.0899f
C2425 col_n[22] a_25054_4138# 0.251f
C2426 a_17934_15182# a_18026_15182# 0.326f
C2427 a_2475_15206# a_33998_15182# 0.264f
C2428 a_2275_15206# a_31382_15222# 0.144f
C2429 VDD a_17934_10162# 0.181f
C2430 col_n[29] a_31990_6146# 0.0765f
C2431 col_n[2] a_5278_8194# 0.084f
C2432 m2_34864_11990# m2_35292_12418# 0.165f
C2433 vcm a_23958_5142# 0.1f
C2434 m2_7756_946# col_n[5] 0.331f
C2435 a_19030_8154# a_19030_7150# 0.843f
C2436 rowoff_n[10] a_17934_12170# 0.202f
C2437 a_29374_1166# col_n[26] 0.084f
C2438 m2_29268_16434# rowon_n[14] 0.0322f
C2439 m2_18224_12418# a_18026_12170# 0.165f
C2440 row_n[6] a_14010_8154# 0.282f
C2441 m2_34864_11990# rowon_n[10] 0.231f
C2442 vcm a_11302_14218# 0.155f
C2443 a_2275_12194# a_24962_12170# 0.136f
C2444 a_12914_12170# a_13310_12210# 0.0313f
C2445 VDD a_9390_4500# 0.0779f
C2446 rowon_n[10] a_13918_12170# 0.118f
C2447 col_n[13] a_16418_2492# 0.0283f
C2448 ctop a_24050_9158# 4.11f
C2449 VDD a_32994_14178# 0.181f
C2450 col_n[23] a_26458_14540# 0.0283f
C2451 col_n[5] a_2475_12194# 0.0531f
C2452 row_n[8] a_2275_10186# 19.2f
C2453 col_n[10] a_2475_1150# 0.0531f
C2454 rowoff_n[0] a_9902_2130# 0.202f
C2455 rowon_n[0] a_23958_2130# 0.118f
C2456 rowon_n[12] a_1957_14202# 0.0172f
C2457 a_31990_5142# a_32482_5504# 0.0658f
C2458 a_31078_5142# a_31382_5182# 0.0931f
C2459 m2_13780_946# ctop 0.0428f
C2460 vcm a_4882_8154# 0.1f
C2461 m2_21812_18014# m2_22240_18442# 0.165f
C2462 a_2475_9182# a_17022_9158# 0.316f
C2463 a_8990_9158# a_9994_9158# 0.843f
C2464 rowoff_n[14] a_33998_16186# 0.202f
C2465 vcm a_26362_18234# 0.16f
C2466 VDD a_24450_8516# 0.0779f
C2467 col[3] a_5886_8154# 0.0682f
C2468 m2_1732_11990# ctop 0.0428f
C2469 ctop a_4974_12170# 4.11f
C2470 VDD a_13918_17190# 0.181f
C2471 a_29982_1126# col[27] 0.0682f
C2472 col_n[11] a_14010_2130# 0.251f
C2473 a_27974_2130# a_28066_2130# 0.326f
C2474 col_n[21] a_24050_14178# 0.251f
C2475 m3_30980_1078# VDD 0.0157f
C2476 col_n[18] a_20946_4138# 0.0765f
C2477 row_n[9] a_35002_11166# 0.0437f
C2478 a_2275_6170# a_7986_6146# 0.399f
C2479 col_n[28] a_30986_16186# 0.0765f
C2480 col_n[2] a_2275_15206# 0.113f
C2481 rowon_n[13] a_34090_15182# 0.248f
C2482 m2_9188_10410# a_8990_10162# 0.165f
C2483 rowoff_n[3] a_10394_5504# 0.0133f
C2484 col_n[7] a_2275_4162# 0.113f
C2485 vcm a_19942_12170# 0.1f
C2486 a_34090_12170# a_34090_11166# 0.843f
C2487 col_n[1] a_4274_18234# 0.084f
C2488 a_2475_11190# a_32082_11166# 0.316f
C2489 VDD a_16018_2130# 0.483f
C2490 sample a_1957_8178# 0.345f
C2491 a_27974_16186# a_28370_16226# 0.0313f
C2492 VDD a_5374_11528# 0.0779f
C2493 m2_31852_18014# m3_32988_18146# 0.0341f
C2494 ctop a_20034_16186# 4.11f
C2495 col_n[22] a_2475_14202# 0.0531f
C2496 col_n[12] a_15414_12532# 0.0283f
C2497 col_n[27] a_2475_3158# 0.0531f
C2498 sample_n rowoff_n[0] 0.14f
C2499 rowoff_n[1] a_19430_3496# 0.0133f
C2500 rowoff_n[8] a_2475_10186# 3.9f
C2501 en_bit_n[2] a_2275_1150# 0.0364f
C2502 m2_28264_6394# a_28066_6146# 0.165f
C2503 row_n[13] a_12002_15182# 0.282f
C2504 a_12914_8154# a_13406_8516# 0.0658f
C2505 rowoff_n[11] a_5886_13174# 0.202f
C2506 a_2275_8178# a_23046_8154# 0.399f
C2507 a_12002_8154# a_12306_8194# 0.0931f
C2508 col[18] a_2475_18218# 0.136f
C2509 vcm a_35002_16186# 0.101f
C2510 a_24050_13174# a_25054_13174# 0.843f
C2511 VDD a_31078_6146# 0.483f
C2512 row_n[3] a_22042_5142# 0.282f
C2513 col_n[0] a_3366_18556# 0.0283f
C2514 col[12] a_2475_11190# 0.136f
C2515 m2_1732_13998# row_n[12] 0.292f
C2516 rowon_n[7] a_21950_9158# 0.118f
C2517 a_2475_17214# a_1957_17214# 0.0734f
C2518 m2_7180_10410# row_n[8] 0.0128f
C2519 VDD a_20434_15544# 0.0779f
C2520 rowoff_n[6] a_10998_8154# 0.294f
C2521 m2_13204_6394# row_n[4] 0.0128f
C2522 m2_18224_2378# row_n[0] 0.0128f
C2523 col[2] a_4882_18194# 0.0682f
C2524 a_2475_5166# a_15926_5142# 0.264f
C2525 a_8898_5142# a_8990_5142# 0.326f
C2526 a_2275_5166# a_13310_5182# 0.144f
C2527 row_n[5] a_9294_7190# 0.0117f
C2528 col_n[10] a_13006_12170# 0.251f
C2529 col_n[7] a_9902_2130# 0.0765f
C2530 col_n[19] a_2275_17214# 0.113f
C2531 rowoff_n[15] a_21950_17190# 0.202f
C2532 col_n[17] a_19942_14178# 0.0765f
C2533 col_n[24] a_2275_6170# 0.113f
C2534 rowoff_n[4] a_20034_6146# 0.294f
C2535 a_15014_15182# a_15014_14178# 0.843f
C2536 col_n[22] rowoff_n[14] 0.0471f
C2537 VDD a_12002_9158# 0.483f
C2538 col[25] rowoff_n[10] 0.0901f
C2539 a_2275_2154# a_6890_2130# 0.136f
C2540 m2_28264_15430# row_n[13] 0.0128f
C2541 m2_34288_11414# row_n[9] 0.0128f
C2542 m2_19228_4386# a_19030_4138# 0.165f
C2543 col[9] a_2275_14202# 0.0899f
C2544 vcm a_18026_4138# 0.56f
C2545 rowoff_n[2] a_29070_4138# 0.294f
C2546 a_2475_7174# a_30986_7150# 0.264f
C2547 a_2275_7174# a_28370_7190# 0.144f
C2548 col_n[1] a_4370_10524# 0.0283f
C2549 col[14] a_2275_3158# 0.0899f
C2550 rowon_n[1] a_8990_3134# 0.248f
C2551 a_27974_12170# a_28466_12532# 0.0658f
C2552 a_27062_12170# a_27366_12210# 0.0931f
C2553 VDD a_3878_3134# 0.181f
C2554 col[30] a_33086_11166# 0.367f
C2555 a_2475_16210# a_8990_16186# 0.316f
C2556 a_4974_16186# a_5978_16186# 0.843f
C2557 col[29] a_2475_13198# 0.136f
C2558 VDD a_27062_13174# 0.483f
C2559 a_2275_4162# a_21950_4138# 0.136f
C2560 m3_7888_1078# ctop 0.21f
C2561 vcm a_33086_8154# 0.56f
C2562 a_23958_9158# a_24050_9158# 0.326f
C2563 row_n[10] a_20034_12170# 0.282f
C2564 rowon_n[13] col[3] 0.0323f
C2565 row_n[13] col[2] 0.0342f
C2566 row_n[9] ctop 0.186f
C2567 row_n[15] col[6] 0.0342f
C2568 rowon_n[14] col[5] 0.0323f
C2569 col_n[0] a_2475_10186# 0.0532f
C2570 col_n[19] col[20] 7.13f
C2571 rowon_n[15] col[7] 0.0323f
C2572 rowon_n[12] col[1] 0.0323f
C2573 row_n[14] col[4] 0.0342f
C2574 col_n[25] a_28370_11206# 0.084f
C2575 col_n[6] rowoff_n[15] 0.0471f
C2576 row_n[12] col[0] 0.0322f
C2577 rowon_n[14] a_19942_16186# 0.118f
C2578 col_n[6] a_8898_12170# 0.0765f
C2579 col[9] rowoff_n[11] 0.0901f
C2580 row_n[0] a_30074_2130# 0.282f
C2581 VDD a_7986_16186# 0.483f
C2582 a_2475_1150# a_14010_1126# 0.0299f
C2583 row_n[12] a_7286_14218# 0.0117f
C2584 rowon_n[4] a_29982_6146# 0.118f
C2585 vcm a_23350_2170# 0.155f
C2586 a_18938_6146# a_19334_6186# 0.0313f
C2587 col[26] a_2275_16210# 0.0899f
C2588 m2_1732_9982# sample_n 0.0522f
C2589 m2_12776_946# m2_13780_946# 0.843f
C2590 col[31] a_2275_5166# 0.0899f
C2591 row_n[2] a_17326_4178# 0.0117f
C2592 vcm a_14010_11166# 0.56f
C2593 VDD a_10906_1126# 0.405f
C2594 a_8898_15182# a_9390_15544# 0.0658f
C2595 a_7986_15182# a_8290_15222# 0.0931f
C2596 a_2275_15206# a_15014_15182# 0.399f
C2597 col[19] a_22042_9158# 0.367f
C2598 rowon_n[0] m2_25252_2378# 0.0322f
C2599 row_n[4] a_7894_6146# 0.0437f
C2600 a_15014_3134# a_16018_3134# 0.843f
C2601 col_n[1] a_2275_2154# 0.113f
C2602 a_2475_3158# a_29070_3134# 0.316f
C2603 rowon_n[8] a_6982_10162# 0.248f
C2604 col[26] a_28978_11166# 0.0682f
C2605 rowoff_n[8] a_30986_10162# 0.202f
C2606 vcm a_4274_5182# 0.155f
C2607 rowoff_n[11] a_34090_13174# 0.294f
C2608 vcm a_29070_15182# 0.56f
C2609 a_2475_12194# a_7894_12170# 0.264f
C2610 a_4882_12170# a_4974_12170# 0.326f
C2611 a_3878_12170# a_4274_12210# 0.0313f
C2612 a_2275_12194# a_5278_12210# 0.144f
C2613 VDD a_25966_5142# 0.181f
C2614 col_n[16] a_2475_12194# 0.0531f
C2615 m2_9188_18442# VDD 0.0456f
C2616 col_n[21] a_2475_1150# 0.0531f
C2617 col_n[14] a_17326_9198# 0.084f
C2618 a_2275_17214# a_30074_17190# 0.399f
C2619 a_5978_5142# a_5978_4138# 0.843f
C2620 col_n[25] a_28466_3496# 0.0283f
C2621 vcm a_19334_9198# 0.155f
C2622 col[6] a_2475_9182# 0.136f
C2623 m2_3740_18014# m2_4744_18014# 0.843f
C2624 ctop a_32082_4138# 4.11f
C2625 vcm a_9994_18194# 0.165f
C2626 a_2275_14202# a_20338_14218# 0.144f
C2627 a_2475_14202# a_22954_14178# 0.264f
C2628 VDD a_6890_8154# 0.181f
C2629 row_n[7] a_28066_9158# 0.282f
C2630 m2_3164_5390# rowon_n[3] 0.0322f
C2631 rowon_n[11] a_27974_13174# 0.118f
C2632 VDD a_28370_18234# 0.019f
C2633 a_2275_2154# a_35094_2130# 0.0924f
C2634 a_18026_2130# a_18330_2170# 0.0931f
C2635 col_n[13] a_2275_15206# 0.113f
C2636 a_18938_2130# a_19430_2492# 0.0658f
C2637 col[8] a_10998_7150# 0.367f
C2638 col_n[18] a_2275_4162# 0.113f
C2639 m3_26964_18146# VDD 0.0898f
C2640 vcm a_12914_3134# 0.1f
C2641 row_n[9] a_15318_11206# 0.0117f
C2642 a_30074_7150# a_31078_7150# 0.843f
C2643 col[15] a_17934_9158# 0.0682f
C2644 vcm a_35398_13214# 0.161f
C2645 a_2275_11190# a_13918_11166# 0.136f
C2646 VDD a_32482_3496# 0.0779f
C2647 col_n[23] a_26058_3134# 0.251f
C2648 m2_19804_18014# a_19942_18194# 0.225f
C2649 col_n[0] a_3270_15222# 0.084f
C2650 ctop a_13006_7150# 4.11f
C2651 row_n[11] a_5886_13174# 0.0437f
C2652 a_2275_16210# a_2275_15206# 0.0715f
C2653 a_19942_16186# a_20034_16186# 0.326f
C2654 col_n[30] a_32994_5142# 0.0765f
C2655 col[3] a_2275_12194# 0.0899f
C2656 VDD a_21950_12170# 0.181f
C2657 m2_8760_18014# m3_7888_18146# 0.0341f
C2658 rowon_n[15] a_4974_17190# 0.248f
C2659 m2_18224_14426# rowon_n[12] 0.0322f
C2660 col[8] a_2275_1150# 0.0899f
C2661 col_n[3] a_6282_7190# 0.084f
C2662 m2_24248_10410# rowon_n[8] 0.0322f
C2663 m2_30272_6394# rowon_n[4] 0.0322f
C2664 row_n[1] a_15926_3134# 0.0437f
C2665 col[29] a_2475_18218# 0.136f
C2666 vcm a_27974_7150# 0.1f
C2667 rowon_n[5] a_15014_7150# 0.248f
C2668 a_21038_9158# a_21038_8154# 0.843f
C2669 a_2966_8154# a_3270_8194# 0.0931f
C2670 a_3878_8154# a_4370_8516# 0.0658f
C2671 a_2475_8178# a_5978_8154# 0.316f
C2672 rowoff_n[12] a_22042_14178# 0.294f
C2673 m2_34864_13998# a_35398_14218# 0.087f
C2674 col[23] a_2475_11190# 0.136f
C2675 col_n[14] a_17422_1488# 0.0283f
C2676 vcm a_15318_16226# 0.155f
C2677 a_2275_13198# a_28978_13174# 0.136f
C2678 a_14922_13174# a_15318_13214# 0.0313f
C2679 VDD a_13406_6508# 0.0779f
C2680 col_n[24] a_27462_13536# 0.0283f
C2681 ctop a_28066_11166# 4.11f
C2682 rowon_n[7] a_3878_9158# 0.118f
C2683 VDD a_2161_15206# 0.187f
C2684 col_n[30] a_2275_17214# 0.113f
C2685 a_33086_6146# a_33390_6186# 0.0931f
C2686 a_33998_6146# a_34490_6508# 0.0658f
C2687 m2_34864_4962# vcm 0.408f
C2688 m2_10768_946# m3_11904_1078# 0.0341f
C2689 row_n[15] rowoff_n[14] 0.085f
C2690 vcm a_8898_10162# 0.1f
C2691 a_10998_10162# a_12002_10162# 0.843f
C2692 a_2475_10186# a_21038_10162# 0.316f
C2693 rowoff_n[15] a_3878_17190# 0.202f
C2694 col[7] a_9994_17190# 0.367f
C2695 row_n[14] a_26058_16186# 0.282f
C2696 col[4] a_6890_7150# 0.0682f
C2697 rowoff_n[4] a_1957_6170# 0.0219f
C2698 VDD a_28466_10524# 0.0779f
C2699 col[20] a_2275_14202# 0.0899f
C2700 ctop a_8990_14178# 4.11f
C2701 col_n[22] a_25054_13174# 0.251f
C2702 col[25] a_2275_3158# 0.0899f
C2703 col_n[19] a_21950_3134# 0.0765f
C2704 a_29982_3134# a_30074_3134# 0.326f
C2705 col_n[29] a_31990_15182# 0.0765f
C2706 rowoff_n[2] a_11398_4500# 0.0133f
C2707 rowoff_n[10] a_28466_12532# 0.0133f
C2708 a_2275_7174# a_12002_7150# 0.399f
C2709 col_n[2] a_5278_17230# 0.084f
C2710 m2_26832_18014# vcm 0.353f
C2711 col_n[0] a_2966_7150# 0.251f
C2712 row_n[6] a_23350_8194# 0.0117f
C2713 vcm a_23958_14178# 0.1f
C2714 a_2475_12194# a_2475_11190# 0.0666f
C2715 VDD a_20034_4138# 0.483f
C2716 a_29982_17190# a_30378_17230# 0.0313f
C2717 VDD a_9390_13536# 0.0779f
C2718 col_n[13] a_16418_11528# 0.0283f
C2719 row_n[8] a_13918_10162# 0.0437f
C2720 rowoff_n[7] a_2874_9158# 0.202f
C2721 rowoff_n[0] a_20434_2492# 0.0133f
C2722 rowon_n[12] a_13006_14178# 0.248f
C2723 a_2275_4162# a_3878_4138# 0.136f
C2724 a_2874_4138# a_3366_4500# 0.0658f
C2725 a_2475_4162# a_4882_4138# 0.264f
C2726 m3_3872_18146# ctop 0.209f
C2727 rowon_n[14] col[16] 0.0323f
C2728 row_n[12] col[11] 0.0342f
C2729 rowon_n[10] col[8] 0.0323f
C2730 col_n[17] rowoff_n[15] 0.0471f
C2731 rowon_n[11] col[10] 0.0323f
C2732 row_n[10] col[7] 0.0342f
C2733 row_n[8] col[3] 0.0342f
C2734 row_n[7] col[1] 0.0342f
C2735 row_n[13] col[13] 0.0342f
C2736 rowon_n[13] col[14] 0.0323f
C2737 col_n[10] a_2475_10186# 0.0531f
C2738 rowon_n[7] col[2] 0.0323f
C2739 rowon_n[12] col[12] 0.0323f
C2740 rowon_n[9] col[6] 0.0323f
C2741 rowon_n[6] col[0] 0.0318f
C2742 row_n[15] col[17] 0.0342f
C2743 rowon_n[1] rowon_n[0] 0.0632f
C2744 rowon_n[3] ctop 0.203f
C2745 col_n[25] col[25] 0.541f
C2746 row_n[14] col[15] 0.0342f
C2747 row_n[11] col[9] 0.0342f
C2748 row_n[9] col[5] 0.0342f
C2749 rowon_n[8] col[4] 0.0323f
C2750 rowon_n[15] col[18] 0.0323f
C2751 a_14922_9158# a_15414_9520# 0.0658f
C2752 rowoff_n[13] a_9994_15182# 0.294f
C2753 a_14010_9158# a_14314_9198# 0.0931f
C2754 a_2275_9182# a_27062_9158# 0.399f
C2755 m2_2160_4386# row_n[2] 0.0194f
C2756 m2_33284_15430# a_33086_15182# 0.165f
C2757 row_n[10] a_1957_12194# 0.187f
C2758 rowon_n[2] a_23046_4138# 0.248f
C2759 col[20] rowoff_n[11] 0.0901f
C2760 vcm a_4882_17190# 0.1f
C2761 a_26058_14178# a_27062_14178# 0.843f
C2762 m3_19936_1078# a_19030_1126# 0.0206f
C2763 rowoff_n[5] a_12002_7150# 0.294f
C2764 a_2275_18218# a_5886_18194# 0.136f
C2765 VDD a_24450_17552# 0.0779f
C2766 col[3] a_5886_17190# 0.0682f
C2767 col[0] a_2475_7174# 0.148f
C2768 col_n[11] a_14010_11166# 0.251f
C2769 vcm a_6982_2130# 0.56f
C2770 a_2275_6170# a_17326_6186# 0.144f
C2771 a_2475_6170# a_19942_6146# 0.264f
C2772 col_n[8] a_10906_1126# 0.0765f
C2773 a_10906_6146# a_10998_6146# 0.326f
C2774 col_n[18] a_20946_13174# 0.0765f
C2775 rowoff_n[3] a_21038_5142# 0.294f
C2776 m2_11196_17438# row_n[15] 0.0128f
C2777 m2_15788_18014# col[13] 0.347f
C2778 m2_5172_17438# a_4974_17190# 0.165f
C2779 m2_17220_13422# row_n[11] 0.0128f
C2780 m2_15788_18014# a_16018_17190# 0.843f
C2781 m2_1732_6970# VDD 0.856f
C2782 m2_23244_9406# row_n[7] 0.0128f
C2783 col_n[7] a_2275_13198# 0.113f
C2784 m2_29268_5390# row_n[3] 0.0128f
C2785 row_n[11] a_34090_13174# 0.282f
C2786 a_17022_16186# a_17022_15182# 0.843f
C2787 VDD a_16018_11166# 0.483f
C2788 col_n[12] a_2275_2154# 0.113f
C2789 sample a_1957_17214# 0.345f
C2790 rowon_n[15] a_33998_17190# 0.118f
C2791 a_5886_3134# a_6282_3174# 0.0313f
C2792 a_2275_3158# a_10906_3134# 0.136f
C2793 rowoff_n[1] a_30074_3134# 0.294f
C2794 col_n[2] a_5374_9520# 0.0283f
C2795 m2_1732_4962# a_2161_5166# 0.0454f
C2796 a_24050_1126# a_2275_1150# 0.0924f
C2797 row_n[13] a_21342_15222# 0.0117f
C2798 vcm a_22042_6146# 0.56f
C2799 rowoff_n[11] a_16418_13536# 0.0133f
C2800 a_2275_8178# a_32386_8194# 0.144f
C2801 col_n[27] a_2475_12194# 0.0531f
C2802 a_2475_8178# a_35002_8154# 0.264f
C2803 col[4] rowoff_n[12] 0.0901f
C2804 m2_24248_13422# a_24050_13174# 0.165f
C2805 col[31] a_34090_10162# 0.367f
C2806 a_29982_13174# a_30474_13536# 0.0658f
C2807 a_29070_13174# a_29374_13214# 0.0931f
C2808 row_n[3] a_31382_5182# 0.0117f
C2809 row_n[15] a_11910_17190# 0.0437f
C2810 a_6982_17190# a_7986_17190# 0.843f
C2811 a_2475_17214# a_13006_17190# 0.316f
C2812 VDD a_31078_15182# 0.483f
C2813 col[17] a_2475_9182# 0.136f
C2814 row_n[5] a_21950_7150# 0.0437f
C2815 a_2275_5166# a_25966_5142# 0.136f
C2816 m2_34864_7974# a_2475_8178# 0.282f
C2817 rowon_n[9] a_21038_11166# 0.248f
C2818 col_n[26] a_29374_10202# 0.084f
C2819 vcm a_2874_9158# 0.1f
C2820 a_26970_1126# a_27366_1166# 0.0313f
C2821 rowoff_n[15] a_32482_17552# 0.0133f
C2822 a_25966_10162# a_26058_10162# 0.326f
C2823 col_n[7] a_9902_11166# 0.0765f
C2824 a_2275_14202# a_3970_14178# 0.399f
C2825 m2_16792_946# a_2275_1150# 0.28f
C2826 col_n[24] a_2275_15206# 0.113f
C2827 col_n[29] a_2275_4162# 0.113f
C2828 VDD a_12002_18194# 0.0356f
C2829 m2_31852_18014# col_n[29] 0.243f
C2830 a_2475_2154# a_18026_2130# 0.316f
C2831 a_27062_3134# a_27062_2130# 0.843f
C2832 m2_11196_1374# VDD 0.0194f
C2833 vcm a_27366_4178# 0.155f
C2834 a_20946_7150# a_21342_7190# 0.0313f
C2835 rowoff_n[9] a_22954_11166# 0.202f
C2836 m2_15212_11414# a_15014_11166# 0.165f
C2837 vcm a_18026_13174# 0.56f
C2838 col[14] a_2275_12194# 0.0899f
C2839 VDD a_14922_3134# 0.181f
C2840 m2_17796_18014# a_2275_18218# 0.28f
C2841 col[19] a_2275_1150# 0.0899f
C2842 col[20] a_23046_8154# 0.367f
C2843 a_2275_16210# a_19030_16186# 0.399f
C2844 a_10906_16186# a_11398_16548# 0.0658f
C2845 a_9994_16186# a_10298_16226# 0.0931f
C2846 VDD a_3878_12170# 0.181f
C2847 rowon_n[3] a_8898_5142# 0.118f
C2848 a_27062_1126# m2_26832_946# 0.0249f
C2849 col[27] a_29982_10162# 0.0682f
C2850 rowoff_n[7] a_31990_9158# 0.202f
C2851 a_2475_4162# a_33086_4138# 0.316f
C2852 a_17022_4138# a_18026_4138# 0.843f
C2853 m2_34288_7398# a_34090_7150# 0.165f
C2854 vcm a_8290_7190# 0.155f
C2855 rowoff_n[12] a_4370_14540# 0.0133f
C2856 row_n[10] a_29374_12210# 0.0117f
C2857 vcm a_33086_17190# 0.56f
C2858 ctop a_21038_2130# 4.06f
C2859 a_2475_13198# a_11910_13174# 0.264f
C2860 col_n[15] a_18330_8194# 0.084f
C2861 a_6890_13174# a_6982_13174# 0.326f
C2862 a_2275_13198# a_9294_13214# 0.144f
C2863 VDD a_29982_7150# 0.181f
C2864 m2_13780_18014# a_2475_18218# 0.286f
C2865 a_2275_18218# a_34090_18194# 0.0924f
C2866 col_n[4] a_2475_8178# 0.0531f
C2867 row_n[12] a_19942_14178# 0.0437f
C2868 col_n[26] a_29470_2492# 0.0283f
C2869 vcm a_34394_2170# 0.155f
C2870 a_7986_6146# a_7986_5142# 0.843f
C2871 m2_6176_9406# a_5978_9158# 0.165f
C2872 row_n[2] a_29982_4138# 0.0437f
C2873 vcm a_23350_11206# 0.155f
C2874 a_2161_10186# a_2275_10186# 0.183f
C2875 a_2475_10186# a_2966_10162# 0.317f
C2876 VDD a_21438_1488# 0.0977f
C2877 rowon_n[6] a_29070_8154# 0.248f
C2878 col[31] a_2275_14202# 0.0899f
C2879 ctop a_2475_5166# 0.0488f
C2880 a_2275_15206# a_24354_15222# 0.144f
C2881 a_2475_15206# a_26970_15182# 0.264f
C2882 VDD a_10906_10162# 0.181f
C2883 col[9] a_12002_6146# 0.367f
C2884 a_20034_3134# a_20338_3174# 0.0931f
C2885 a_20946_3134# a_21438_3496# 0.0658f
C2886 a_2475_18218# a_32082_18194# 0.0299f
C2887 m2_25252_5390# a_25054_5142# 0.165f
C2888 col[16] a_18938_8154# 0.0682f
C2889 vcm a_16930_5142# 0.1f
C2890 col_n[1] a_2275_11190# 0.113f
C2891 a_32082_8154# a_33086_8154# 0.843f
C2892 rowoff_n[10] a_10906_12170# 0.202f
C2893 a_30074_1126# vcm 0.165f
C2894 m2_1732_16006# rowon_n[14] 0.236f
C2895 col_n[24] a_27062_2130# 0.251f
C2896 m2_7180_12418# rowon_n[10] 0.0322f
C2897 row_n[6] a_6982_8154# 0.282f
C2898 m2_13204_8402# rowon_n[6] 0.0322f
C2899 vcm a_4274_14218# 0.155f
C2900 m2_19228_4386# rowon_n[2] 0.0322f
C2901 a_2275_12194# a_17934_12170# 0.136f
C2902 m2_34864_5966# rowoff_n[4] 0.278f
C2903 VDD a_1957_4162# 0.196f
C2904 rowon_n[10] a_6890_12170# 0.118f
C2905 col_n[31] a_33998_4138# 0.0765f
C2906 m2_30848_18014# VDD 1.11f
C2907 ctop a_17022_9158# 4.11f
C2908 a_21950_17190# a_22042_17190# 0.326f
C2909 VDD a_25966_14178# 0.181f
C2910 col_n[4] a_7286_6186# 0.084f
C2911 col[0] a_2966_4138# 0.367f
C2912 row_n[6] col[10] 0.0342f
C2913 row_n[13] col[24] 0.0342f
C2914 row_n[7] col[12] 0.0342f
C2915 rowon_n[5] col[9] 0.0323f
C2916 rowon_n[15] col[29] 0.0323f
C2917 col_n[21] a_2475_10186# 0.0531f
C2918 rowon_n[7] col[13] 0.0323f
C2919 row_n[8] col[14] 0.0342f
C2920 row_n[5] col[8] 0.0342f
C2921 rowon_n[1] col[1] 0.0323f
C2922 rowon_n[12] col[23] 0.0323f
C2923 row_n[14] col[26] 0.0342f
C2924 rowon_n[3] col[5] 0.0323f
C2925 row_n[11] col[20] 0.0342f
C2926 rowon_n[14] col[27] 0.0323f
C2927 row_n[1] col[0] 0.0322f
C2928 col_n[28] rowoff_n[15] 0.0471f
C2929 row_n[2] col[2] 0.0342f
C2930 rowon_n[6] col[11] 0.0323f
C2931 row_n[12] col[22] 0.0342f
C2932 rowon_n[13] col[25] 0.0323f
C2933 rowon_n[2] col[3] 0.0323f
C2934 row_n[9] col[16] 0.0342f
C2935 col_n[30] col[31] 7.27f
C2936 rowon_n[10] col[19] 0.0323f
C2937 rowon_n[11] col[21] 0.0323f
C2938 row_n[10] col[18] 0.0342f
C2939 rowon_n[9] col[17] 0.0323f
C2940 rowon_n[4] col[7] 0.0323f
C2941 rowon_n[8] col[15] 0.0323f
C2942 row_n[4] col[6] 0.0342f
C2943 row_n[3] col[4] 0.0342f
C2944 row_n[15] col[28] 0.0342f
C2945 col_n[14] a_17326_18234# 0.084f
C2946 rowon_n[0] a_16930_2130# 0.118f
C2947 rowoff_n[0] a_2161_2154# 0.0226f
C2948 en_bit_n[0] a_20034_1126# 0.208f
C2949 col[31] rowoff_n[11] 0.0901f
C2950 m2_14784_18014# m2_15212_18442# 0.165f
C2951 vcm a_31990_9158# 0.1f
C2952 rowoff_n[14] a_26970_16186# 0.202f
C2953 a_2475_9182# a_9994_9158# 0.316f
C2954 a_23046_10162# a_23046_9158# 0.843f
C2955 VDD m2_2160_1374# 0.0268f
C2956 col_n[25] a_28466_12532# 0.0283f
C2957 vcm a_19334_18234# 0.16f
C2958 m2_28264_17438# rowon_n[15] 0.0322f
C2959 a_2275_14202# a_32994_14178# 0.136f
C2960 a_16930_14178# a_17326_14218# 0.0313f
C2961 VDD a_17422_8516# 0.0779f
C2962 m2_34288_13422# rowon_n[11] 0.0322f
C2963 col[11] a_2475_7174# 0.136f
C2964 ctop a_32082_13174# 4.11f
C2965 m3_34996_11118# a_34090_11166# 0.0303f
C2966 VDD a_6890_17190# 0.181f
C2967 m2_16216_3382# a_16018_3134# 0.165f
C2968 m3_2868_1078# VDD 0.0166f
C2969 row_n[9] a_27974_11166# 0.0437f
C2970 col[8] a_10998_16186# 0.367f
C2971 rowon_n[13] a_27062_15182# 0.248f
C2972 col_n[18] a_2275_13198# 0.113f
C2973 col[5] a_7894_6146# 0.0682f
C2974 vcm a_12914_12170# 0.1f
C2975 rowoff_n[3] a_2966_5142# 0.294f
C2976 a_13006_11166# a_14010_11166# 0.843f
C2977 a_2475_11190# a_25054_11166# 0.316f
C2978 col_n[23] a_2275_2154# 0.113f
C2979 col[15] a_17934_18194# 0.0682f
C2980 VDD a_8990_2130# 0.483f
C2981 VDD a_32482_12532# 0.0779f
C2982 col_n[23] a_26058_12170# 0.251f
C2983 m2_22816_18014# m3_22948_18146# 3.79f
C2984 col_n[20] a_22954_2130# 0.0765f
C2985 ctop a_13006_16186# 4.11f
C2986 col_n[30] a_32994_14178# 0.0765f
C2987 a_31990_4138# a_32082_4138# 0.326f
C2988 rowoff_n[1] a_12402_3496# 0.0133f
C2989 col[15] rowoff_n[12] 0.0901f
C2990 col[8] a_2275_10186# 0.0899f
C2991 col_n[3] a_6282_16226# 0.084f
C2992 row_n[13] a_4974_15182# 0.282f
C2993 a_2275_8178# a_16018_8154# 0.399f
C2994 vcm a_27974_16186# 0.1f
C2995 a_3970_13174# a_3970_12170# 0.843f
C2996 VDD a_24050_6146# 0.483f
C2997 row_n[3] a_15014_5142# 0.282f
C2998 col_n[14] a_17422_10524# 0.0283f
C2999 col[28] a_2475_9182# 0.136f
C3000 rowon_n[7] a_14922_9158# 0.118f
C3001 a_31990_18194# a_32386_18234# 0.0313f
C3002 VDD a_13406_15544# 0.0779f
C3003 rowoff_n[6] a_3970_8154# 0.294f
C3004 a_2475_5166# a_8898_5142# 0.264f
C3005 a_2275_5166# a_6282_5182# 0.144f
C3006 row_n[5] a_3878_7150# 0.0437f
C3007 m2_26832_946# m3_25960_1078# 0.0341f
C3008 rowon_n[9] a_2966_11166# 0.248f
C3009 rowoff_n[15] a_14922_17190# 0.202f
C3010 a_2275_10186# a_31078_10162# 0.399f
C3011 a_16018_10162# a_16322_10202# 0.0931f
C3012 a_16930_10162# a_17422_10524# 0.0658f
C3013 rowoff_n[4] a_13006_6146# 0.294f
C3014 a_28066_15182# a_29070_15182# 0.843f
C3015 VDD a_4974_9158# 0.483f
C3016 col[4] a_6890_16186# 0.0682f
C3017 col_n[12] a_15014_10162# 0.251f
C3018 a_35002_3134# a_35398_3174# 0.0313f
C3019 m2_6176_11414# row_n[9] 0.0128f
C3020 m2_12200_7398# row_n[5] 0.0128f
C3021 m2_18224_3382# row_n[1] 0.0128f
C3022 vcm a_10998_4138# 0.56f
C3023 col_n[19] a_21950_12170# 0.0765f
C3024 col[25] a_2275_12194# 0.0899f
C3025 a_12914_7150# a_13006_7150# 0.326f
C3026 a_2275_7174# a_21342_7190# 0.144f
C3027 a_2475_7174# a_23958_7150# 0.264f
C3028 rowoff_n[2] a_22042_4138# 0.294f
C3029 rowon_n[1] a_2475_3158# 0.31f
C3030 col[30] a_2275_1150# 0.0899f
C3031 row_n[6] a_34394_8194# 0.0117f
C3032 rowon_n[10] a_35094_12170# 0.0141f
C3033 col_n[0] a_2966_16186# 0.251f
C3034 a_19030_17190# a_19030_16186# 0.843f
C3035 VDD a_20034_13174# 0.483f
C3036 rowoff_n[0] a_31078_2130# 0.294f
C3037 m2_1732_13998# col[0] 0.0137f
C3038 col_n[3] a_6378_8516# 0.0283f
C3039 a_7894_4138# a_8290_4178# 0.0313f
C3040 a_2275_4162# a_14922_4138# 0.136f
C3041 m3_34996_12122# ctop 0.209f
C3042 a_30474_1488# col_n[27] 0.0283f
C3043 m2_27260_16434# row_n[14] 0.0128f
C3044 m2_33284_12418# row_n[10] 0.0128f
C3045 vcm a_26058_8154# 0.56f
C3046 a_2966_9158# a_2966_8154# 0.843f
C3047 row_n[10] a_13006_12170# 0.282f
C3048 rowon_n[14] a_12914_16186# 0.118f
C3049 a_31990_14178# a_32482_14540# 0.0658f
C3050 col_n[15] a_2475_8178# 0.0531f
C3051 a_31078_14178# a_31382_14218# 0.0931f
C3052 row_n[0] a_23046_2130# 0.282f
C3053 a_2475_1150# a_6982_1126# 0.0299f
C3054 rowon_n[4] a_22954_6146# 0.118f
C3055 m2_2736_1950# a_3270_2170# 0.087f
C3056 vcm a_16322_2170# 0.155f
C3057 a_2275_6170# a_29982_6146# 0.136f
C3058 col[0] a_2475_16210# 0.148f
C3059 col_n[27] a_30378_9198# 0.084f
C3060 col_n[1] a_3970_8154# 0.251f
C3061 m2_1732_7974# vcm 0.316f
C3062 m2_5748_946# m2_6752_946# 0.843f
C3063 col[5] a_2475_5166# 0.136f
C3064 row_n[2] a_10298_4178# 0.0117f
C3065 vcm a_6982_11166# 0.56f
C3066 a_27974_11166# a_28066_11166# 0.326f
C3067 col_n[8] a_10906_10162# 0.0765f
C3068 VDD a_3366_1488# 0.0978f
C3069 a_2275_15206# a_7986_15182# 0.399f
C3070 m2_34864_16006# m3_34996_15134# 0.0341f
C3071 m2_32856_946# col[30] 0.425f
C3072 col_n[12] a_2275_11190# 0.113f
C3073 a_29070_4138# a_29070_3134# 0.843f
C3074 a_2475_3158# a_22042_3134# 0.316f
C3075 rowoff_n[8] a_23958_10162# 0.202f
C3076 a_35398_1166# a_2275_1150# 0.145f
C3077 row_n[13] a_33998_15182# 0.0437f
C3078 vcm a_31382_6186# 0.155f
C3079 rowoff_n[11] a_27062_13174# 0.294f
C3080 a_22954_8154# a_23350_8194# 0.0313f
C3081 col_n[2] a_5374_18556# 0.0283f
C3082 vcm a_22042_15182# 0.56f
C3083 col[21] a_24050_7150# 0.367f
C3084 VDD a_18938_5142# 0.181f
C3085 rowon_n[3] col[16] 0.0323f
C3086 rowon_n[1] col[12] 0.0323f
C3087 rowon_n[0] col[10] 0.0323f
C3088 row_n[9] col[27] 0.0342f
C3089 row_n[5] col[19] 0.0342f
C3090 rowon_n[10] col[30] 0.0323f
C3091 row_n[0] col[9] 0.0342f
C3092 row_n[4] col[17] 0.0342f
C3093 rowon_n[6] col[22] 0.0323f
C3094 rowon_n[7] col[24] 0.0323f
C3095 rowon_n[9] col[28] 0.0323f
C3096 rowon_n[8] col[26] 0.0323f
C3097 rowon_n[4] col[18] 0.0323f
C3098 row_n[11] col[31] 0.0342f
C3099 row_n[2] col[13] 0.0342f
C3100 rowon_n[5] col[20] 0.0323f
C3101 row_n[6] col[21] 0.0342f
C3102 row_n[8] col[25] 0.0342f
C3103 row_n[1] col[11] 0.0342f
C3104 rowon_n[2] col[14] 0.0323f
C3105 rowon_n[11] sample_n 0.0692f
C3106 a_32082_1126# VDD 0.035f
C3107 row_n[7] col[23] 0.0342f
C3108 row_n[3] col[15] 0.0342f
C3109 ctop col[6] 0.123f
C3110 row_n[10] col[29] 0.0342f
C3111 a_12914_17190# a_13406_17552# 0.0658f
C3112 a_2275_17214# a_23046_17190# 0.399f
C3113 col[2] a_2275_8178# 0.0899f
C3114 a_12002_17190# a_12306_17230# 0.0931f
C3115 col[28] a_30986_9158# 0.0682f
C3116 rowoff_n[6] a_32994_8154# 0.202f
C3117 a_25054_2130# m2_25252_2378# 0.165f
C3118 a_19030_5142# a_20034_5142# 0.843f
C3119 m3_27968_1078# m3_28972_1078# 0.202f
C3120 vcm a_12306_9198# 0.155f
C3121 col_n[16] a_19334_7190# 0.084f
C3122 col[22] a_2475_7174# 0.136f
C3123 ctop a_25054_4138# 4.11f
C3124 vcm a_2874_18194# 0.101f
C3125 a_8898_14178# a_8990_14178# 0.326f
C3126 a_2475_14202# a_15926_14178# 0.264f
C3127 a_2275_14202# a_13310_14218# 0.144f
C3128 m2_14784_946# a_14922_1126# 0.225f
C3129 VDD a_33998_9158# 0.181f
C3130 row_n[7] a_21038_9158# 0.282f
C3131 rowon_n[11] a_20946_13174# 0.118f
C3132 VDD a_21342_18234# 0.019f
C3133 a_2275_2154# a_28066_2130# 0.399f
C3134 m2_1732_2954# a_2475_3158# 0.139f
C3135 col_n[29] a_2275_13198# 0.113f
C3136 m2_34864_946# VDD 1.3f
C3137 vcm a_5886_3134# 0.1f
C3138 row_n[9] a_8290_11206# 0.0117f
C3139 rowon_n[1] a_30986_3134# 0.118f
C3140 rowoff_n[9] a_33486_11528# 0.0133f
C3141 a_9994_7150# a_9994_6146# 0.843f
C3142 vcm a_27366_13214# 0.155f
C3143 a_2275_11190# a_6890_11166# 0.136f
C3144 VDD a_25454_3496# 0.0779f
C3145 m2_14784_18014# a_15014_18194# 0.0249f
C3146 ctop a_5978_7150# 4.11f
C3147 a_2475_16210# a_30986_16186# 0.264f
C3148 a_2275_16210# a_28370_16226# 0.144f
C3149 col[10] a_13006_5142# 0.367f
C3150 VDD a_14922_12170# 0.181f
C3151 a_35094_1126# m2_34864_946# 0.0249f
C3152 col[19] a_2275_10186# 0.0899f
C3153 col[26] rowoff_n[12] 0.0901f
C3154 col[20] a_23046_17190# 0.367f
C3155 col[17] a_19942_7150# 0.0682f
C3156 m2_2160_6394# rowon_n[4] 0.0219f
C3157 m2_7180_2378# rowon_n[0] 0.0322f
C3158 a_22954_4138# a_23446_4500# 0.0658f
C3159 a_22042_4138# a_22346_4178# 0.0931f
C3160 row_n[1] a_8898_3134# 0.0437f
C3161 rowon_n[5] a_7986_7150# 0.248f
C3162 m2_1732_15002# m2_2160_15430# 0.165f
C3163 vcm a_20946_7150# 0.1f
C3164 rowoff_n[12] a_15014_14178# 0.294f
C3165 a_33998_9158# a_34394_9198# 0.0313f
C3166 m2_30272_14426# a_30074_14178# 0.165f
C3167 vcm a_8290_16226# 0.155f
C3168 a_2275_13198# a_21950_13174# 0.136f
C3169 VDD a_6378_6508# 0.0779f
C3170 col_n[5] a_8290_5182# 0.084f
C3171 ctop a_21038_11166# 4.11f
C3172 col_n[15] a_18330_17230# 0.084f
C3173 a_23958_18194# a_24050_18194# 0.0991f
C3174 VDD a_29982_16186# 0.181f
C3175 a_18938_1126# a_19030_1126# 0.361f
C3176 col_n[4] a_2475_17214# 0.0531f
C3177 m2_17220_15430# rowon_n[13] 0.0322f
C3178 m2_23244_11414# rowon_n[9] 0.0322f
C3179 col_n[9] a_2475_6170# 0.0531f
C3180 m2_29268_7398# rowon_n[5] 0.0322f
C3181 m2_34864_2954# rowon_n[1] 0.231f
C3182 col_n[26] a_29470_11528# 0.0283f
C3183 vcm a_34394_11206# 0.155f
C3184 a_2475_10186# a_14010_10162# 0.316f
C3185 a_25054_11166# a_25054_10162# 0.843f
C3186 row_n[14] a_19030_16186# 0.282f
C3187 m2_1732_16006# a_1957_16210# 0.245f
C3188 a_18938_15182# a_19334_15222# 0.0313f
C3189 VDD a_21438_10524# 0.0779f
C3190 col[10] rowoff_n[13] 0.0901f
C3191 m2_34864_12994# m3_34996_12122# 0.0341f
C3192 ctop a_2475_14202# 0.0488f
C3193 row_n[4] a_29070_6146# 0.282f
C3194 rowon_n[8] a_28978_10162# 0.118f
C3195 col[9] a_12002_15182# 0.367f
C3196 col[6] a_8898_5142# 0.0682f
C3197 a_3878_7150# a_3970_7150# 0.326f
C3198 a_2275_7174# a_4974_7150# 0.399f
C3199 rowoff_n[2] a_4370_4500# 0.0133f
C3200 rowoff_n[10] a_21438_12532# 0.0133f
C3201 a_2874_7150# a_3270_7190# 0.0313f
C3202 m2_12776_18014# vcm 0.353f
C3203 m2_21236_12418# a_21038_12170# 0.165f
C3204 col[16] a_18938_17190# 0.0682f
C3205 row_n[6] a_16322_8194# 0.0117f
C3206 vcm a_16930_14178# 0.1f
C3207 a_15014_12170# a_16018_12170# 0.843f
C3208 a_2475_12194# a_29070_12170# 0.316f
C3209 VDD a_13006_4138# 0.483f
C3210 col_n[24] a_27062_11166# 0.251f
C3211 col_n[6] a_2275_9182# 0.113f
C3212 col_n[21] a_23958_1126# 0.0765f
C3213 row_n[0] m2_23244_2378# 0.0128f
C3214 VDD a_1957_13198# 0.196f
C3215 col_n[31] a_33998_13174# 0.0765f
C3216 row_n[8] a_6890_10162# 0.0437f
C3217 rowoff_n[0] a_13406_2492# 0.0133f
C3218 col_n[4] a_7286_15222# 0.084f
C3219 rowon_n[12] a_5978_14178# 0.248f
C3220 col[0] a_2966_13174# 0.367f
C3221 a_33998_5142# a_34090_5142# 0.326f
C3222 m2_22816_946# ctop 0.0428f
C3223 col_n[26] a_2475_8178# 0.0531f
C3224 rowoff_n[13] a_2874_15182# 0.202f
C3225 a_2275_9182# a_20034_9158# 0.399f
C3226 rowon_n[2] a_16018_4138# 0.248f
C3227 vcm a_31990_18194# 0.101f
C3228 ctop rowoff_n[14] 0.177f
C3229 a_5978_14178# a_5978_13174# 0.843f
C3230 col_n[15] a_18426_9520# 0.0283f
C3231 VDD a_28066_8154# 0.483f
C3232 rowoff_n[5] a_4974_7150# 0.294f
C3233 VDD a_17422_17552# 0.0779f
C3234 col[11] a_2475_16210# 0.136f
C3235 a_28978_2130# a_29374_2170# 0.0313f
C3236 col[16] a_2475_5166# 0.136f
C3237 vcm a_34090_3134# 0.56f
C3238 a_2275_6170# a_10298_6186# 0.144f
C3239 a_2475_6170# a_12914_6146# 0.264f
C3240 m2_12200_10410# a_12002_10162# 0.165f
C3241 col_n[0] a_2874_5142# 0.0765f
C3242 rowoff_n[3] a_14010_5142# 0.294f
C3243 a_18938_11166# a_19430_11528# 0.0658f
C3244 a_2275_11190# a_35094_11166# 0.0924f
C3245 a_18026_11166# a_18330_11206# 0.0931f
C3246 m2_33860_18014# a_34090_18194# 0.0249f
C3247 col[5] a_7894_15182# 0.0682f
C3248 m2_1732_4962# row_n[3] 0.292f
C3249 row_n[11] a_27062_13174# 0.282f
C3250 a_30074_16186# a_31078_16186# 0.843f
C3251 col_n[23] a_2275_11190# 0.113f
C3252 VDD a_8990_11166# 0.483f
C3253 col_n[13] a_16018_9158# 0.251f
C3254 rowon_n[15] a_26970_17190# 0.118f
C3255 a_2874_3134# a_2966_3134# 0.326f
C3256 col_n[20] a_22954_11166# 0.0765f
C3257 rowoff_n[1] a_23046_3134# 0.294f
C3258 m2_31276_6394# a_31078_6146# 0.165f
C3259 row_n[13] a_14314_15222# 0.0117f
C3260 vcm a_15014_6146# 0.56f
C3261 rowoff_n[11] a_9390_13536# 0.0133f
C3262 a_2475_8178# a_27974_8154# 0.264f
C3263 a_2275_8178# a_25358_8194# 0.144f
C3264 a_14922_8154# a_15014_8154# 0.326f
C3265 en_bit_n[1] col[15] 0.142f
C3266 ctop col[17] 0.127f
C3267 row_n[1] col[22] 0.0342f
C3268 row_n[2] col[24] 0.0342f
C3269 row_n[3] col[26] 0.0342f
C3270 col[5] col[6] 0.0355f
C3271 rowon_n[3] col[27] 0.0323f
C3272 rowon_n[4] col[29] 0.0323f
C3273 rowon_n[0] col[21] 0.0323f
C3274 row_n[6] sample_n 0.0596f
C3275 row_n[5] col[30] 0.0342f
C3276 row_n[4] col[28] 0.0342f
C3277 row_n[0] col[20] 0.0342f
C3278 rowon_n[5] col[31] 0.0323f
C3279 rowon_n[1] col[23] 0.0323f
C3280 rowon_n[2] col[25] 0.0323f
C3281 col[13] a_2275_8178# 0.0899f
C3282 row_n[3] a_24354_5182# 0.0117f
C3283 row_n[15] a_4882_17190# 0.0437f
C3284 m2_16216_14426# row_n[12] 0.0128f
C3285 a_3878_17190# a_4370_17552# 0.0658f
C3286 a_2966_17190# a_3270_17230# 0.0931f
C3287 a_2475_17214# a_5978_17190# 0.316f
C3288 m2_22240_10410# row_n[8] 0.0128f
C3289 VDD a_24050_15182# 0.483f
C3290 col_n[4] a_7382_7512# 0.0283f
C3291 m2_28264_6394# row_n[4] 0.0128f
C3292 row_n[5] a_14922_7150# 0.0437f
C3293 a_9902_5142# a_10298_5182# 0.0313f
C3294 a_2275_5166# a_18938_5142# 0.136f
C3295 m3_34996_6098# m3_34996_5094# 0.202f
C3296 rowon_n[9] a_14010_11166# 0.248f
C3297 vcm a_30074_10162# 0.56f
C3298 en_C0_n a_4370_1488# 0.018f
C3299 rowoff_n[15] a_25454_17552# 0.0133f
C3300 m2_25828_946# a_26058_2130# 0.843f
C3301 a_33998_15182# a_34490_15544# 0.0658f
C3302 a_33086_15182# a_33390_15222# 0.0931f
C3303 row_n[7] a_2966_9158# 0.281f
C3304 m2_34864_9982# m3_34996_9110# 0.0341f
C3305 rowon_n[11] a_2275_13198# 1.79f
C3306 col_n[3] a_2475_4162# 0.0531f
C3307 VDD a_4974_18194# 0.0356f
C3308 a_5978_2130# a_6982_2130# 0.843f
C3309 a_2475_2154# a_10998_2130# 0.316f
C3310 col_n[2] a_4974_7150# 0.251f
C3311 col_n[28] a_31382_8194# 0.084f
C3312 m2_22240_4386# a_22042_4138# 0.165f
C3313 vcm a_20338_4178# 0.155f
C3314 a_2275_7174# a_33998_7150# 0.136f
C3315 rowoff_n[9] a_15926_11166# 0.202f
C3316 col_n[9] a_11910_9158# 0.0765f
C3317 vcm a_10998_13174# 0.56f
C3318 a_29982_12170# a_30074_12170# 0.326f
C3319 VDD a_7894_3134# 0.181f
C3320 m2_2736_18014# a_2966_18194# 0.0249f
C3321 m2_3740_18014# a_2275_18218# 0.28f
C3322 col[30] a_2275_10186# 0.0899f
C3323 sw_n a_2475_1150# 0.0185f
C3324 a_2275_16210# a_12002_16186# 0.399f
C3325 row_n[8] a_35094_10162# 0.0123f
C3326 rowoff_n[7] a_24962_9158# 0.202f
C3327 rowon_n[12] a_35002_14178# 0.118f
C3328 a_2475_4162# a_26058_4138# 0.316f
C3329 a_31078_5142# a_31078_4138# 0.843f
C3330 m3_22948_1078# ctop 0.21f
C3331 col_n[3] a_6378_17552# 0.0283f
C3332 vcm a_2275_7174# 6.49f
C3333 rowoff_n[13] a_31990_15182# 0.202f
C3334 a_24962_9158# a_25358_9198# 0.0313f
C3335 col[22] a_25054_6146# 0.367f
C3336 row_n[10] a_22346_12210# 0.0117f
C3337 ctop a_14010_2130# 4.06f
C3338 vcm a_26058_17190# 0.56f
C3339 a_2874_13174# a_3366_13536# 0.0658f
C3340 a_2475_13198# a_4882_13174# 0.264f
C3341 a_2275_13198# a_3878_13174# 0.136f
C3342 VDD a_22954_7150# 0.181f
C3343 col[29] a_31990_8154# 0.0682f
C3344 rowoff_n[5] a_33998_7150# 0.202f
C3345 ctop a_2966_11166# 4.06f
C3346 a_14922_18194# a_15414_18556# 0.0658f
C3347 col_n[15] a_2475_17214# 0.0531f
C3348 a_2275_18218# a_27062_18194# 0.0924f
C3349 row_n[0] a_32386_2170# 0.0117f
C3350 a_9902_1126# a_10394_1488# 0.0658f
C3351 a_2275_1150# a_17022_1126# 0.0924f
C3352 row_n[12] a_12914_14178# 0.0437f
C3353 col_n[20] a_2475_6170# 0.0531f
C3354 vcm a_28978_2130# 0.1f
C3355 a_21038_6146# a_22042_6146# 0.843f
C3356 m2_16792_946# m2_17220_1374# 0.165f
C3357 col_n[17] a_20338_6186# 0.084f
C3358 vcm a_16322_11206# 0.155f
C3359 row_n[2] a_22954_4138# 0.0437f
C3360 col_n[27] a_30378_18234# 0.084f
C3361 col[21] rowoff_n[13] 0.0901f
C3362 col_n[1] a_3970_17190# 0.251f
C3363 VDD a_14410_1488# 0.0977f
C3364 rowon_n[6] a_22042_8154# 0.248f
C3365 col[5] a_2475_14202# 0.136f
C3366 ctop a_29070_6146# 4.11f
C3367 a_10906_15182# a_10998_15182# 0.326f
C3368 a_2475_15206# a_19942_15182# 0.264f
C3369 a_2275_15206# a_17326_15222# 0.144f
C3370 col[10] a_2475_3158# 0.136f
C3371 col_n[4] rowoff_n[9] 0.0471f
C3372 vcm rowoff_n[5] 0.533f
C3373 col_n[2] rowoff_n[7] 0.0471f
C3374 col_n[0] rowoff_n[4] 0.0471f
C3375 VDD rowoff_n[2] 1.51f
C3376 col_n[1] rowoff_n[6] 0.0471f
C3377 sample rowoff_n[3] 0.0775f
C3378 col_n[3] rowoff_n[8] 0.0471f
C3379 VDD a_3366_10524# 0.0779f
C3380 a_2275_3158# a_32082_3134# 0.399f
C3381 a_2475_18218# a_25054_18194# 0.0299f
C3382 rowoff_n[8] a_34490_10524# 0.0133f
C3383 vcm a_9902_5142# 0.1f
C3384 rowoff_n[10] a_3366_12532# 0.0133f
C3385 a_12002_8154# a_12002_7150# 0.843f
C3386 col_n[17] a_2275_9182# 0.113f
C3387 vcm a_31382_15222# 0.155f
C3388 a_2275_12194# a_10906_12170# 0.136f
C3389 a_5886_12170# a_6282_12210# 0.0313f
C3390 VDD a_29470_5504# 0.0779f
C3391 col[11] a_14010_4138# 0.367f
C3392 m2_16792_18014# VDD 0.993f
C3393 ctop a_9994_9158# 4.11f
C3394 row_n[15] a_33086_17190# 0.282f
C3395 a_2275_17214# a_32386_17230# 0.144f
C3396 col[21] a_24050_16186# 0.367f
C3397 a_2475_17214# a_35002_17190# 0.264f
C3398 VDD a_18938_14178# 0.181f
C3399 col[18] a_20946_6146# 0.0682f
C3400 rowon_n[0] a_9902_2130# 0.118f
C3401 col[28] a_30986_18194# 0.0682f
C3402 col[2] a_2275_17214# 0.0899f
C3403 a_24050_5142# a_24354_5182# 0.0931f
C3404 col[7] a_2275_6170# 0.0899f
C3405 a_24962_5142# a_25454_5504# 0.0658f
C3406 col[5] rowoff_n[14] 0.0901f
C3407 vcm a_24962_9158# 0.1f
C3408 m2_7756_18014# m2_8184_18442# 0.165f
C3409 a_1957_9182# a_2275_9182# 0.158f
C3410 rowoff_n[14] a_19942_16186# 0.202f
C3411 a_2475_9182# a_2874_9158# 0.264f
C3412 col_n[6] a_9294_4178# 0.084f
C3413 vcm a_12306_18234# 0.16f
C3414 a_2275_14202# a_25966_14178# 0.136f
C3415 VDD a_10394_8516# 0.0779f
C3416 col_n[16] a_19334_16226# 0.084f
C3417 row_n[7] a_30378_9198# 0.0117f
C3418 m2_6176_13422# rowon_n[11] 0.0322f
C3419 col[22] a_2475_16210# 0.136f
C3420 m2_34864_6970# m3_34996_6098# 0.0341f
C3421 m2_12200_9406# rowon_n[7] 0.0322f
C3422 m2_18224_5390# rowon_n[3] 0.0322f
C3423 m2_14784_946# vcm 0.353f
C3424 ctop a_25054_13174# 4.11f
C3425 col[27] a_2475_5166# 0.136f
C3426 VDD a_33998_18194# 0.343f
C3427 a_20946_2130# a_21038_2130# 0.326f
C3428 m2_2736_1950# a_2966_3134# 0.843f
C3429 row_n[9] a_20946_11166# 0.0437f
C3430 col_n[27] a_30474_10524# 0.0283f
C3431 rowon_n[13] a_20034_15182# 0.248f
C3432 vcm a_5886_12170# 0.1f
C3433 a_27062_12170# a_27062_11166# 0.843f
C3434 a_2475_11190# a_18026_11166# 0.316f
C3435 VDD a_2475_2154# 26.1f
C3436 m2_20808_18014# a_21342_18234# 0.087f
C3437 a_20946_16186# a_21342_16226# 0.0313f
C3438 VDD a_25454_12532# 0.0779f
C3439 rowon_n[3] a_30074_5142# 0.248f
C3440 m2_13780_18014# m3_12908_18146# 0.0341f
C3441 col[0] a_2874_2130# 0.0682f
C3442 m2_33284_14426# rowon_n[12] 0.0322f
C3443 ctop a_5978_16186# 4.11f
C3444 col[10] a_13006_14178# 0.367f
C3445 VDD col_n[5] 5.17f
C3446 col[7] a_9902_4138# 0.0682f
C3447 vcm col_n[2] 1.94f
C3448 rowoff_n[1] a_5374_3496# 0.0133f
C3449 rowon_n[0] sample_n 0.0692f
C3450 ctop col[28] 0.123f
C3451 row_n[0] col[31] 0.0342f
C3452 col[24] a_2275_8178# 0.0899f
C3453 col[17] a_19942_16186# 0.0682f
C3454 a_4974_8154# a_5278_8194# 0.0931f
C3455 a_5886_8154# a_6378_8516# 0.0658f
C3456 a_2275_8178# a_8990_8154# 0.399f
C3457 col_n[25] a_28066_10162# 0.251f
C3458 vcm a_20946_16186# 0.1f
C3459 a_2475_13198# a_33086_13174# 0.316f
C3460 a_17022_13174# a_18026_13174# 0.843f
C3461 VDD a_17022_6146# 0.483f
C3462 row_n[3] a_7986_5142# 0.282f
C3463 rowon_n[7] a_7894_9158# 0.118f
C3464 VDD a_6378_15544# 0.0779f
C3465 col_n[5] a_8290_14218# 0.084f
C3466 vcm a_23046_1126# 0.165f
C3467 m2_15788_946# m3_16924_1078# 0.0341f
C3468 m3_23952_18146# m3_24956_18146# 0.202f
C3469 a_2275_10186# a_24050_10162# 0.399f
C3470 rowoff_n[15] a_7894_17190# 0.202f
C3471 row_n[14] a_28370_16226# 0.0117f
C3472 col_n[16] a_19430_8516# 0.0283f
C3473 col_n[9] a_2475_15206# 0.0531f
C3474 rowoff_n[4] a_5978_6146# 0.294f
C3475 col_n[14] a_2475_4162# 0.0531f
C3476 a_7986_15182# a_7986_14178# 0.843f
C3477 VDD a_32082_10162# 0.483f
C3478 a_30986_3134# a_31382_3174# 0.0313f
C3479 vcm a_3970_4138# 0.56f
C3480 rowoff_n[2] a_15014_4138# 0.294f
C3481 a_2475_7174# a_16930_7150# 0.264f
C3482 rowoff_n[10] a_32082_12170# 0.294f
C3483 a_2275_7174# a_14314_7190# 0.144f
C3484 col[4] a_2475_1150# 0.136f
C3485 row_n[6] a_28978_8154# 0.0437f
C3486 col[6] a_8898_14178# 0.0682f
C3487 a_20946_12170# a_21438_12532# 0.0658f
C3488 a_20034_12170# a_20338_12210# 0.0931f
C3489 rowon_n[10] a_28066_12170# 0.248f
C3490 col_n[14] a_17022_8154# 0.251f
C3491 a_32082_17190# a_33086_17190# 0.843f
C3492 VDD a_13006_13174# 0.483f
C3493 col_n[6] a_2275_18218# 0.113f
C3494 col_n[21] a_23958_10162# 0.0765f
C3495 rowoff_n[0] a_24050_2130# 0.294f
C3496 col_n[11] a_2275_7174# 0.113f
C3497 a_2275_4162# a_7894_4138# 0.136f
C3498 m3_18932_18146# ctop 0.209f
C3499 vcm a_19030_8154# 0.56f
C3500 m2_5172_12418# row_n[10] 0.0128f
C3501 a_2475_9182# a_31990_9158# 0.264f
C3502 a_16930_9158# a_17022_9158# 0.326f
C3503 a_2275_9182# a_29374_9198# 0.144f
C3504 m2_11196_8402# row_n[6] 0.0128f
C3505 m2_17220_4386# row_n[2] 0.0128f
C3506 row_n[10] a_5978_12170# 0.282f
C3507 col_n[26] a_2475_17214# 0.0531f
C3508 rowon_n[14] a_5886_16186# 0.118f
C3509 col_n[5] a_8386_6508# 0.0283f
C3510 m2_34864_3958# m3_34996_3086# 0.0341f
C3511 col_n[31] a_2475_6170# 0.0531f
C3512 col[1] a_2275_4162# 0.0899f
C3513 col_n[15] a_18426_18556# 0.0283f
C3514 VDD a_28066_17190# 0.484f
C3515 row_n[0] a_16018_2130# 0.282f
C3516 a_18026_2130# a_18026_1126# 0.843f
C3517 rowon_n[4] a_15926_6146# 0.118f
C3518 vcm a_9294_2170# 0.155f
C3519 sample_n rowoff_n[13] 0.14f
C3520 a_11910_6146# a_12306_6186# 0.0313f
C3521 a_2275_6170# a_22954_6146# 0.136f
C3522 col[16] a_2475_14202# 0.136f
C3523 vcm a_34090_12170# 0.56f
C3524 row_n[2] a_3270_4178# 0.0117f
C3525 col_n[13] rowoff_n[7] 0.0471f
C3526 col_n[7] rowoff_n[1] 0.0471f
C3527 col_n[12] rowoff_n[6] 0.0471f
C3528 col_n[14] rowoff_n[8] 0.0471f
C3529 col_n[10] rowoff_n[4] 0.0471f
C3530 col_n[8] rowoff_n[2] 0.0471f
C3531 col_n[15] rowoff_n[9] 0.0471f
C3532 col[21] a_2475_3158# 0.136f
C3533 col_n[9] rowoff_n[3] 0.0471f
C3534 col_n[11] rowoff_n[5] 0.0471f
C3535 col_n[6] rowoff_n[0] 0.0471f
C3536 VDD a_30986_2130# 0.181f
C3537 m2_26256_17438# row_n[15] 0.0128f
C3538 m2_8184_17438# a_7986_17190# 0.165f
C3539 m2_32280_13422# row_n[11] 0.0128f
C3540 col_n[0] a_2874_14178# 0.0765f
C3541 col_n[29] a_32386_7190# 0.084f
C3542 col_n[3] a_5978_6146# 0.251f
C3543 a_7986_3134# a_8990_3134# 0.843f
C3544 a_2475_3158# a_15014_3134# 0.316f
C3545 rowoff_n[8] a_16930_10162# 0.202f
C3546 col_n[28] a_2275_9182# 0.113f
C3547 a_28978_1126# a_2475_1150# 0.264f
C3548 m2_34864_15002# rowoff_n[13] 0.278f
C3549 col_n[10] a_12914_8154# 0.0765f
C3550 a_26362_1166# a_2275_1150# 0.145f
C3551 row_n[13] a_26970_15182# 0.0437f
C3552 vcm a_24354_6186# 0.155f
C3553 rowoff_n[11] a_20034_13174# 0.294f
C3554 m2_27260_13422# a_27062_13174# 0.165f
C3555 vcm a_15014_15182# 0.56f
C3556 a_31990_13174# a_32082_13174# 0.326f
C3557 VDD a_11910_5142# 0.181f
C3558 a_25054_1126# VDD 0.035f
C3559 col[13] a_2275_17214# 0.0899f
C3560 a_2275_17214# a_16018_17190# 0.399f
C3561 rowoff_n[6] a_25966_8154# 0.202f
C3562 col[18] a_2275_6170# 0.0899f
C3563 col[16] rowoff_n[14] 0.0901f
C3564 col_n[4] a_7382_16548# 0.0283f
C3565 m2_2736_1950# m2_3164_2378# 0.165f
C3566 col_n[1] a_3878_6146# 0.0765f
C3567 a_33086_6146# a_33086_5142# 0.843f
C3568 a_2475_5166# a_30074_5142# 0.316f
C3569 m3_13912_1078# m3_14916_1078# 0.202f
C3570 col[23] a_26058_5142# 0.367f
C3571 col_n[0] rowoff_n[10] 0.0471f
C3572 vcm a_5278_9198# 0.155f
C3573 a_26970_10162# a_27366_10202# 0.0313f
C3574 col[30] a_32994_7150# 0.0682f
C3575 rowoff_n[4] a_35002_6146# 0.202f
C3576 ctop a_18026_4138# 4.11f
C3577 m2_25828_946# a_2275_1150# 0.28f
C3578 m2_9764_946# a_9994_1126# 0.0249f
C3579 a_2475_14202# a_8898_14178# 0.264f
C3580 a_2275_14202# a_6282_14218# 0.144f
C3581 row_n[7] a_14010_9158# 0.282f
C3582 VDD a_26970_9158# 0.181f
C3583 rowon_n[11] a_13918_13174# 0.118f
C3584 m2_16792_946# col[14] 0.425f
C3585 VDD a_14314_18234# 0.019f
C3586 a_2275_2154# a_21038_2130# 0.399f
C3587 a_11910_2130# a_12402_2492# 0.0658f
C3588 a_10998_2130# a_11302_2170# 0.0931f
C3589 col_n[3] a_2475_13198# 0.0531f
C3590 col_n[18] a_21342_5182# 0.084f
C3591 m2_20232_1374# VDD 0.0208f
C3592 row_n[9] a_2275_11190# 19.2f
C3593 vcm a_32994_4138# 0.1f
C3594 rowon_n[1] a_23958_3134# 0.118f
C3595 rowoff_n[9] a_26458_11528# 0.0133f
C3596 col_n[8] a_2475_2154# 0.0531f
C3597 a_23046_7150# a_24050_7150# 0.843f
C3598 col_n[28] a_31382_17230# 0.084f
C3599 col_n[2] a_4974_16186# 0.251f
C3600 m2_18224_11414# a_18026_11166# 0.165f
C3601 rowon_n[13] a_1957_15206# 0.0172f
C3602 vcm a_20338_13214# 0.155f
C3603 a_35002_12170# a_35398_12210# 0.0313f
C3604 col_n[9] a_11910_18194# 0.0762f
C3605 VDD a_18426_3496# 0.0779f
C3606 ctop a_33086_8154# 4.11f
C3607 a_2275_16210# a_21342_16226# 0.144f
C3608 a_2475_16210# a_23958_16186# 0.264f
C3609 a_12914_16186# a_13006_16186# 0.326f
C3610 VDD a_7894_12170# 0.181f
C3611 col_n[6] col_n[7] 0.0101f
C3612 vcm col_n[13] 1.94f
C3613 VDD col_n[16] 4.83f
C3614 col[0] rowoff_n[15] 0.0901f
C3615 col[16] col[17] 0.0337f
C3616 rowoff_n[7] a_35494_9520# 0.0133f
C3617 m2_9764_18014# col[7] 0.347f
C3618 vcm a_13918_7150# 0.1f
C3619 a_14010_9158# a_14010_8154# 0.843f
C3620 rowoff_n[12] a_7986_14178# 0.294f
C3621 row_n[10] a_35002_12170# 0.0437f
C3622 col[12] a_15014_3134# 0.367f
C3623 vcm a_2275_16210# 6.49f
C3624 a_7894_13174# a_8290_13214# 0.0313f
C3625 a_2275_13198# a_14922_13174# 0.136f
C3626 rowon_n[14] a_34090_16186# 0.248f
C3627 col[22] a_25054_15182# 0.367f
C3628 VDD a_33486_7512# 0.0779f
C3629 col_n[5] a_2275_5166# 0.113f
C3630 col[19] a_21950_5142# 0.0682f
C3631 ctop a_14010_11166# 4.11f
C3632 col[29] a_31990_17190# 0.0682f
C3633 VDD a_22954_16186# 0.181f
C3634 m2_1732_4962# m2_1732_3958# 0.843f
C3635 a_26058_6146# a_26362_6186# 0.0931f
C3636 a_26970_6146# a_27462_6508# 0.0658f
C3637 col_n[20] a_2475_15206# 0.0531f
C3638 m2_1732_6970# rowon_n[5] 0.236f
C3639 m2_28840_946# m2_29844_946# 0.843f
C3640 m2_7180_3382# rowon_n[1] 0.0322f
C3641 m2_9188_9406# a_8990_9158# 0.165f
C3642 col_n[25] a_2475_4162# 0.0531f
C3643 vcm a_28978_11166# 0.1f
C3644 col_n[7] a_10298_3174# 0.084f
C3645 a_2475_10186# a_6982_10162# 0.316f
C3646 a_3970_10162# a_4974_10162# 0.843f
C3647 row_n[14] a_12002_16186# 0.282f
C3648 col_n[17] a_20338_15222# 0.084f
C3649 m3_2868_2082# a_2966_3134# 0.0303f
C3650 a_2275_15206# a_29982_15182# 0.136f
C3651 VDD a_14410_10524# 0.0779f
C3652 ctop a_29070_15182# 4.11f
C3653 row_n[4] a_22042_6146# 0.282f
C3654 col[10] a_2475_12194# 0.136f
C3655 rowon_n[8] a_21950_10162# 0.118f
C3656 a_22954_3134# a_23046_3134# 0.326f
C3657 col[15] a_2475_1150# 0.136f
C3658 col_n[28] a_31478_9520# 0.0283f
C3659 m2_1732_10986# rowoff_n[9] 0.415f
C3660 m2_28264_5390# a_28066_5142# 0.165f
C3661 rowoff_n[10] a_14410_12532# 0.0133f
C3662 a_32386_1166# vcm 0.16f
C3663 m2_16216_16434# rowon_n[14] 0.0322f
C3664 row_n[6] a_9294_8194# 0.0117f
C3665 m2_22240_12418# rowon_n[10] 0.0322f
C3666 vcm a_9902_14178# 0.1f
C3667 m2_28264_8402# rowon_n[6] 0.0322f
C3668 a_29070_13174# a_29070_12170# 0.843f
C3669 m2_34288_4386# rowon_n[2] 0.0322f
C3670 a_2475_12194# a_22042_12170# 0.316f
C3671 VDD a_5978_4138# 0.483f
C3672 col_n[17] a_2275_18218# 0.113f
C3673 m2_25828_18014# col_n[23] 0.243f
C3674 col[1] a_3970_1126# 0.428f
C3675 a_22954_17190# a_23350_17230# 0.0313f
C3676 col_n[22] a_2275_7174# 0.113f
C3677 VDD a_29470_14540# 0.0779f
C3678 col[11] a_14010_13174# 0.367f
C3679 col[8] a_10906_3134# 0.0682f
C3680 rowoff_n[0] a_6378_2492# 0.0133f
C3681 col[18] a_20946_15182# 0.0682f
C3682 col_n[26] a_29070_9158# 0.251f
C3683 m2_1732_18014# m2_1732_17010# 0.843f
C3684 a_2275_9182# a_13006_9158# 0.399f
C3685 a_7894_9158# a_8386_9520# 0.0658f
C3686 a_6982_9158# a_7286_9198# 0.0931f
C3687 rowoff_n[14] a_30474_16548# 0.0133f
C3688 col[7] a_2275_15206# 0.0899f
C3689 col[12] a_2275_4162# 0.0899f
C3690 rowon_n[2] a_8990_4138# 0.248f
C3691 vcm a_24962_18194# 0.101f
C3692 a_19030_14178# a_20034_14178# 0.843f
C3693 VDD a_21038_8154# 0.483f
C3694 col_n[6] a_9294_13214# 0.084f
C3695 VDD a_10394_17552# 0.0779f
C3696 col[27] a_2475_14202# 0.136f
C3697 m2_19228_3382# a_19030_3134# 0.165f
C3698 col_n[19] rowoff_n[2] 0.0471f
C3699 col_n[26] rowoff_n[9] 0.0471f
C3700 col_n[25] rowoff_n[8] 0.0471f
C3701 col_n[17] rowoff_n[0] 0.0471f
C3702 col_n[22] rowoff_n[5] 0.0471f
C3703 col_n[21] rowoff_n[4] 0.0471f
C3704 col_n[23] rowoff_n[6] 0.0471f
C3705 col_n[24] rowoff_n[7] 0.0471f
C3706 col_n[20] rowoff_n[3] 0.0471f
C3707 vcm a_27062_3134# 0.56f
C3708 col_n[18] rowoff_n[1] 0.0471f
C3709 a_2475_6170# a_5886_6146# 0.264f
C3710 a_2275_6170# a_3270_6186# 0.144f
C3711 col_n[17] a_20434_7512# 0.0283f
C3712 rowoff_n[3] a_6982_5142# 0.294f
C3713 col_n[3] a_2475_18218# 0.0529f
C3714 a_2275_11190# a_28066_11166# 0.399f
C3715 a_9994_16186# a_9994_15182# 0.843f
C3716 row_n[11] a_20034_13174# 0.282f
C3717 VDD a_2475_11190# 26.1f
C3718 m2_27836_18014# m3_27968_18146# 3.79f
C3719 rowon_n[15] a_19942_17190# 0.118f
C3720 a_32994_4138# a_33390_4178# 0.0313f
C3721 col[0] a_2874_11166# 0.0682f
C3722 rowoff_n[1] a_16018_3134# 0.294f
C3723 row_n[1] a_30074_3134# 0.282f
C3724 m2_1732_16006# rowoff_n[14] 0.415f
C3725 row_n[13] a_7286_15222# 0.0117f
C3726 vcm a_7986_6146# 0.56f
C3727 rowon_n[5] a_29982_7150# 0.118f
C3728 a_2475_8178# a_20946_8154# 0.264f
C3729 col[7] a_9902_13174# 0.0682f
C3730 rowoff_n[11] a_1957_13198# 0.0219f
C3731 a_2275_8178# a_18330_8194# 0.144f
C3732 col[24] a_2275_17214# 0.0899f
C3733 m2_1732_10986# sample 0.2f
C3734 col_n[15] a_18026_7150# 0.251f
C3735 a_22954_13174# a_23446_13536# 0.0658f
C3736 a_22042_13174# a_22346_13214# 0.0931f
C3737 col[29] a_2275_6170# 0.0899f
C3738 m2_34864_4962# ctop 0.0422f
C3739 row_n[3] a_17326_5182# 0.0117f
C3740 col[27] rowoff_n[14] 0.0901f
C3741 col_n[22] a_24962_9158# 0.0765f
C3742 a_33998_18194# a_34394_18234# 0.0313f
C3743 VDD a_17022_15182# 0.483f
C3744 m2_5172_2378# row_n[0] 0.0128f
C3745 col_n[10] rowoff_n[10] 0.0471f
C3746 row_n[5] a_7894_7150# 0.0437f
C3747 a_2275_5166# a_11910_5142# 0.136f
C3748 m3_34996_13126# m3_34996_12122# 0.202f
C3749 m2_31852_946# m3_30980_1078# 0.0341f
C3750 col_n[0] a_2275_3158# 0.113f
C3751 rowon_n[9] a_6982_11166# 0.248f
C3752 vcm a_23046_10162# 0.56f
C3753 a_18938_10162# a_19030_10162# 0.326f
C3754 a_2275_10186# a_33390_10202# 0.144f
C3755 rowoff_n[15] a_18426_17552# 0.0133f
C3756 col_n[6] a_9390_5504# 0.0283f
C3757 col_n[16] a_19430_17552# 0.0283f
C3758 m2_26832_18014# ctop 0.0422f
C3759 col_n[14] a_2475_13198# 0.0531f
C3760 col_n[19] a_2475_2154# 0.0531f
C3761 a_2475_2154# a_3970_2130# 0.316f
C3762 a_20034_3134# a_20034_2130# 0.843f
C3763 a_2275_2154# a_2966_2130# 0.0924f
C3764 m2_15212_15430# row_n[13] 0.0128f
C3765 m2_21236_11414# row_n[9] 0.0128f
C3766 m2_27260_7398# row_n[5] 0.0128f
C3767 m2_33284_3382# row_n[1] 0.0128f
C3768 vcm a_13310_4178# 0.155f
C3769 a_2275_7174# a_26970_7150# 0.136f
C3770 a_13918_7150# a_14314_7190# 0.0313f
C3771 rowoff_n[9] a_8898_11166# 0.202f
C3772 vcm a_3970_13174# 0.56f
C3773 VDD col_n[27] 5.17f
C3774 vcm col_n[24] 1.94f
C3775 VDD a_35002_4138# 0.258f
C3776 col[4] a_2475_10186# 0.136f
C3777 col[11] rowoff_n[15] 0.0901f
C3778 a_2275_16210# a_4974_16186# 0.399f
C3779 a_2874_16186# a_3270_16226# 0.0313f
C3780 a_3878_16186# a_3970_16186# 0.326f
C3781 col_n[4] a_6982_5142# 0.251f
C3782 col_n[30] a_33390_6186# 0.084f
C3783 col_n[14] a_17022_17190# 0.251f
C3784 row_n[8] a_28066_10162# 0.282f
C3785 rowoff_n[7] a_17934_9158# 0.202f
C3786 col_n[11] a_13918_7150# 0.0765f
C3787 rowon_n[12] a_27974_14178# 0.118f
C3788 a_9994_4138# a_10998_4138# 0.843f
C3789 a_2475_4162# a_19030_4138# 0.316f
C3790 m3_1864_4090# ctop 0.21f
C3791 col_n[11] a_2275_16210# 0.113f
C3792 vcm a_28370_8194# 0.155f
C3793 rowoff_n[13] a_24962_15182# 0.202f
C3794 col_n[16] a_2275_5166# 0.113f
C3795 row_n[10] a_15318_12210# 0.0117f
C3796 vcm a_19030_17190# 0.56f
C3797 ctop a_6982_2130# 4.06f
C3798 a_33998_14178# a_34090_14178# 0.326f
C3799 VDD a_15926_7150# 0.181f
C3800 rowoff_n[5] a_26970_7150# 0.202f
C3801 a_2275_18218# a_20034_18194# 0.0924f
C3802 row_n[0] a_25358_2170# 0.0117f
C3803 col_n[31] a_2475_15206# 0.0531f
C3804 col_n[5] a_8386_15544# 0.0283f
C3805 row_n[12] a_5886_14178# 0.0437f
C3806 a_2275_1150# a_9994_1126# 0.0924f
C3807 col[1] a_2275_13198# 0.0899f
C3808 col[24] a_27062_4138# 0.367f
C3809 vcm a_21950_2130# 0.1f
C3810 col[6] a_2275_2154# 0.0899f
C3811 a_2475_6170# a_34090_6146# 0.316f
C3812 m2_9764_946# m2_10192_1374# 0.165f
C3813 col[31] a_33998_6146# 0.0682f
C3814 row_n[2] a_15926_4138# 0.0437f
C3815 vcm a_9294_11206# 0.155f
C3816 a_28978_11166# a_29374_11206# 0.0313f
C3817 VDD a_7382_1488# 0.0977f
C3818 rowon_n[6] a_15014_8154# 0.248f
C3819 ctop a_22042_6146# 4.11f
C3820 col[21] a_2475_12194# 0.136f
C3821 a_2275_15206# a_10298_15222# 0.144f
C3822 a_2475_15206# a_12914_15182# 0.264f
C3823 VDD a_30986_11166# 0.181f
C3824 col[26] a_2475_1150# 0.136f
C3825 col_n[19] a_22346_4178# 0.084f
C3826 a_13918_3134# a_14410_3496# 0.0658f
C3827 a_13006_3134# a_13310_3174# 0.0931f
C3828 a_2275_3158# a_25054_3134# 0.399f
C3829 a_2475_18218# a_18026_18194# 0.0299f
C3830 rowon_n[8] a_3878_10162# 0.118f
C3831 rowoff_n[8] a_27462_10524# 0.0133f
C3832 col_n[29] a_32386_16226# 0.084f
C3833 col_n[3] a_5978_15182# 0.251f
C3834 vcm a_2161_5166# 0.0169f
C3835 a_25054_8154# a_26058_8154# 0.843f
C3836 col_n[28] a_2275_18218# 0.113f
C3837 col_n[10] a_12914_17190# 0.0765f
C3838 m2_34864_12994# a_35398_13214# 0.087f
C3839 vcm a_24354_15222# 0.155f
C3840 a_2874_12170# a_2966_12170# 0.326f
C3841 VDD a_22442_5504# 0.0779f
C3842 m2_2736_18014# VDD 1.09f
C3843 row_n[15] a_26058_17190# 0.282f
C3844 m3_1864_7102# a_2966_7150# 0.0302f
C3845 a_14922_17190# a_15014_17190# 0.326f
C3846 a_2275_17214# a_25358_17230# 0.144f
C3847 a_2475_17214# a_27974_17190# 0.264f
C3848 VDD a_11910_14178# 0.181f
C3849 a_28066_2130# m2_28264_2378# 0.165f
C3850 rowon_n[0] a_2161_2154# 0.0177f
C3851 col[18] a_2275_15206# 0.0899f
C3852 col[23] a_2275_4162# 0.0899f
C3853 vcm a_17934_9158# 0.1f
C3854 col[13] a_16018_2130# 0.367f
C3855 col_n[1] a_3878_15182# 0.0765f
C3856 rowoff_n[14] a_12914_16186# 0.202f
C3857 a_16018_10162# a_16018_9158# 0.843f
C3858 col[23] a_26058_14178# 0.367f
C3859 vcm a_5278_18234# 0.16f
C3860 col[20] a_22954_4138# 0.0682f
C3861 m3_20940_1078# a_21038_2130# 0.0302f
C3862 m2_15788_946# a_16322_1166# 0.087f
C3863 a_2275_14202# a_18938_14178# 0.136f
C3864 a_9902_14178# a_10298_14218# 0.0313f
C3865 row_n[7] a_23350_9198# 0.0117f
C3866 VDD a_2966_8154# 0.485f
C3867 col[30] a_32994_16186# 0.0682f
C3868 ctop a_18026_13174# 4.11f
C3869 VDD a_26970_18194# 0.343f
C3870 col_n[31] rowoff_n[3] 0.0471f
C3871 col_n[30] rowoff_n[2] 0.0471f
C3872 col_n[29] rowoff_n[1] 0.0471f
C3873 col_n[28] rowoff_n[0] 0.0471f
C3874 a_2475_2154# a_32994_2130# 0.264f
C3875 a_2275_2154# a_30378_2170# 0.144f
C3876 m3_13912_18146# VDD 0.0312f
C3877 col_n[14] a_2475_18218# 0.0529f
C3878 row_n[9] a_13918_11166# 0.0437f
C3879 col_n[8] a_11302_2170# 0.084f
C3880 a_28066_7150# a_28370_7190# 0.0931f
C3881 a_28978_7150# a_29470_7512# 0.0658f
C3882 rowon_n[13] a_13006_15182# 0.248f
C3883 col_n[18] a_21342_14218# 0.084f
C3884 vcm a_32994_13174# 0.1f
C3885 a_5978_11166# a_6982_11166# 0.843f
C3886 col_n[8] a_2475_11190# 0.0531f
C3887 a_2475_11190# a_10998_11166# 0.316f
C3888 VDD a_29070_3134# 0.483f
C3889 row_n[11] a_1957_13198# 0.187f
C3890 a_2275_16210# a_33998_16186# 0.136f
C3891 rowon_n[3] a_23046_5142# 0.248f
C3892 VDD a_18426_12532# 0.0779f
C3893 m2_3740_18014# m3_4876_18146# 0.0341f
C3894 m2_5172_14426# rowon_n[12] 0.0322f
C3895 ctop a_33086_17190# 4.06f
C3896 col_n[29] a_32482_8516# 0.0283f
C3897 m2_11196_10410# rowon_n[8] 0.0322f
C3898 m2_17220_6394# rowon_n[4] 0.0322f
C3899 a_24962_4138# a_25054_4138# 0.326f
C3900 a_1957_8178# a_2161_8178# 0.115f
C3901 a_2475_8178# a_2275_8178# 2.76f
C3902 m2_33284_14426# a_33086_14178# 0.165f
C3903 vcm a_13918_16186# 0.1f
C3904 a_2475_13198# a_26058_13174# 0.316f
C3905 a_31078_14178# a_31078_13174# 0.843f
C3906 VDD a_9994_6146# 0.483f
C3907 m2_26832_946# col[24] 0.425f
C3908 col[12] a_15014_12170# 0.367f
C3909 col_n[21] rowoff_n[10] 0.0471f
C3910 col[9] a_11910_2130# 0.0682f
C3911 a_24962_18194# a_25358_18234# 0.0313f
C3912 VDD a_33486_16548# 0.0779f
C3913 col_n[5] a_2275_14202# 0.113f
C3914 a_19942_1126# a_20338_1166# 0.0342f
C3915 col[19] a_21950_14178# 0.0682f
C3916 row_n[12] a_34090_14178# 0.282f
C3917 col_n[10] a_2275_3158# 0.113f
C3918 vcm a_16018_1126# 0.165f
C3919 m2_32280_15430# rowon_n[13] 0.0322f
C3920 col_n[27] a_30074_8154# 0.251f
C3921 m2_6752_946# m3_6884_1078# 3.79f
C3922 m3_9896_18146# m3_10900_18146# 0.202f
C3923 a_8990_10162# a_9294_10202# 0.0931f
C3924 a_9902_10162# a_10394_10524# 0.0658f
C3925 a_2275_10186# a_17022_10162# 0.399f
C3926 row_n[14] a_21342_16226# 0.0117f
C3927 m2_5172_16434# a_4974_16186# 0.165f
C3928 col_n[25] a_2475_13198# 0.0531f
C3929 col_n[7] a_10298_12210# 0.084f
C3930 m2_8760_946# a_8990_2130# 0.843f
C3931 a_21038_15182# a_22042_15182# 0.843f
C3932 col_n[30] a_2475_2154# 0.0531f
C3933 VDD a_25054_10162# 0.483f
C3934 row_n[4] a_31382_6186# 0.0117f
C3935 m2_1732_3958# a_2161_4162# 0.0454f
C3936 col_n[18] a_21438_6508# 0.0283f
C3937 vcm a_31078_5142# 0.56f
C3938 col_n[1] rowon_n[14] 0.111f
C3939 col_n[0] rowon_n[13] 0.111f
C3940 rowoff_n[10] a_25054_12170# 0.294f
C3941 col_n[3] rowon_n[15] 0.111f
C3942 VDD rowon_n[12] 3.04f
C3943 vcm row_n[14] 0.616f
C3944 sample row_n[13] 0.423f
C3945 col_n[2] row_n[15] 0.298f
C3946 a_2475_7174# a_9902_7150# 0.264f
C3947 rowoff_n[2] a_7986_4138# 0.294f
C3948 a_2275_7174# a_7286_7190# 0.144f
C3949 a_5886_7150# a_5978_7150# 0.326f
C3950 col[22] rowoff_n[15] 0.0901f
C3951 col_n[28] a_31478_18556# 0.0283f
C3952 col[15] a_2475_10186# 0.136f
C3953 col[27] col[28] 0.0355f
C3954 m2_24248_12418# a_24050_12170# 0.165f
C3955 row_n[6] a_21950_8154# 0.0437f
C3956 a_2275_12194# a_32082_12170# 0.399f
C3957 rowon_n[10] a_21038_12170# 0.248f
C3958 col_n[5] rowoff_n[11] 0.0471f
C3959 a_12002_17190# a_12002_16186# 0.843f
C3960 VDD a_5978_13174# 0.483f
C3961 col[1] a_3970_10162# 0.367f
C3962 rowon_n[0] a_31078_2130# 0.248f
C3963 rowoff_n[0] a_17022_2130# 0.294f
C3964 col_n[22] a_2275_16210# 0.113f
C3965 col_n[27] a_2275_5166# 0.113f
C3966 col[8] a_10906_12170# 0.0682f
C3967 m2_34864_6970# a_2475_7174# 0.282f
C3968 vcm a_12002_8154# 0.56f
C3969 a_2275_9182# a_22346_9198# 0.144f
C3970 a_2475_9182# a_24962_9158# 0.264f
C3971 col_n[16] a_19030_6146# 0.251f
C3972 a_24962_14178# a_25454_14540# 0.0658f
C3973 a_24050_14178# a_24354_14218# 0.0931f
C3974 col_n[23] a_25966_8154# 0.0765f
C3975 col[12] a_2275_13198# 0.0899f
C3976 a_1957_18218# a_2275_18218# 0.158f
C3977 VDD a_21038_17190# 0.484f
C3978 row_n[0] a_8990_2130# 0.282f
C3979 col[17] a_2275_2154# 0.0899f
C3980 a_31078_2130# a_32082_2130# 0.843f
C3981 rowon_n[4] a_8898_6146# 0.118f
C3982 vcm a_3878_2130# 0.1f
C3983 a_2275_6170# a_15926_6146# 0.136f
C3984 m2_15212_10410# a_15014_10162# 0.165f
C3985 vcm a_27062_12170# 0.56f
C3986 col_n[7] a_10394_4500# 0.0283f
C3987 a_20946_11166# a_21038_11166# 0.326f
C3988 VDD a_23958_2130# 0.181f
C3989 m2_4168_13422# row_n[11] 0.0128f
C3990 m2_1732_17010# a_2275_17214# 0.191f
C3991 col_n[17] a_20434_16548# 0.0283f
C3992 m2_10192_9406# row_n[7] 0.0128f
C3993 m2_16216_5390# row_n[3] 0.0128f
C3994 row_n[11] a_29374_13214# 0.0117f
C3995 m2_34864_1950# m2_35292_2378# 0.165f
C3996 a_2475_3158# a_7986_3134# 0.316f
C3997 a_22042_4138# a_22042_3134# 0.843f
C3998 col_n[2] a_2475_9182# 0.0531f
C3999 rowoff_n[8] a_9902_10162# 0.202f
C4000 m2_34288_6394# a_34090_6146# 0.165f
C4001 row_n[13] a_19942_15182# 0.0437f
C4002 vcm a_17326_6186# 0.155f
C4003 a_2275_8178# a_30986_8154# 0.136f
C4004 rowoff_n[11] a_13006_13174# 0.294f
C4005 a_15926_8154# a_16322_8194# 0.0313f
C4006 m3_34996_2082# m2_34864_1950# 3.79f
C4007 vcm a_7986_15182# 0.56f
C4008 m3_1864_2082# m2_1732_946# 0.0341f
C4009 VDD a_4882_5142# 0.181f
C4010 row_n[3] a_29982_5142# 0.0437f
C4011 col_n[5] a_7986_4138# 0.251f
C4012 a_5886_17190# a_6378_17552# 0.0658f
C4013 a_2275_17214# a_8990_17190# 0.399f
C4014 col_n[15] a_18026_16186# 0.251f
C4015 m2_31276_14426# row_n[12] 0.0128f
C4016 rowon_n[7] a_29070_9158# 0.248f
C4017 a_4974_17190# a_5278_17230# 0.0931f
C4018 col[29] a_2275_15206# 0.0899f
C4019 rowoff_n[6] a_18938_8154# 0.202f
C4020 col_n[12] a_14922_6146# 0.0765f
C4021 col_n[22] a_24962_18194# 0.0762f
C4022 a_12002_5142# a_13006_5142# 0.843f
C4023 a_2475_5166# a_23046_5142# 0.316f
C4024 m3_1864_2082# m3_1864_1078# 0.202f
C4025 m2_6176_8402# a_5978_8154# 0.165f
C4026 vcm a_32386_10202# 0.155f
C4027 rowoff_n[15] a_29070_17190# 0.294f
C4028 col_n[0] a_2275_12194# 0.113f
C4029 rowoff_n[4] a_27974_6146# 0.202f
C4030 ctop a_10998_4138# 4.11f
C4031 m2_11772_946# a_2475_1150# 0.286f
C4032 row_n[8] rowoff_n[8] 0.209f
C4033 col_n[4] a_2275_1150# 0.113f
C4034 VDD a_19942_9158# 0.181f
C4035 row_n[7] a_6982_9158# 0.282f
C4036 col_n[6] a_9390_14540# 0.0283f
C4037 rowon_n[11] a_6890_13174# 0.118f
C4038 VDD a_7286_18234# 0.019f
C4039 col_n[25] a_2475_18218# 0.0529f
C4040 col[25] a_28066_3134# 0.367f
C4041 a_2275_2154# a_14010_2130# 0.399f
C4042 m2_25252_4386# a_25054_4138# 0.165f
C4043 m2_4744_946# VDD 0.999f
C4044 vcm a_25966_4138# 0.1f
C4045 m2_34864_9982# m2_35292_10410# 0.165f
C4046 col_n[19] a_2475_11190# 0.0531f
C4047 rowon_n[1] a_16930_3134# 0.118f
C4048 rowoff_n[9] a_19430_11528# 0.0133f
C4049 vcm a_13310_13214# 0.155f
C4050 a_30986_12170# a_31382_12210# 0.0313f
C4051 VDD a_11398_3496# 0.0779f
C4052 m2_5748_18014# a_5886_18194# 0.225f
C4053 ctop a_26058_8154# 4.11f
C4054 a_2275_16210# a_14314_16226# 0.144f
C4055 a_2475_16210# a_16930_16186# 0.264f
C4056 VDD a_35002_13174# 0.258f
C4057 col_n[20] a_23350_3174# 0.084f
C4058 rowoff_n[7] a_28466_9520# 0.0133f
C4059 col[9] a_2475_8178# 0.136f
C4060 col_n[4] a_6982_14178# 0.251f
C4061 col_n[30] a_33390_15222# 0.084f
C4062 a_15926_4138# a_16418_4500# 0.0658f
C4063 a_2275_4162# a_29070_4138# 0.399f
C4064 a_15014_4138# a_15318_4178# 0.0931f
C4065 col_n[11] a_13918_16186# 0.0765f
C4066 vcm a_6890_7150# 0.1f
C4067 a_27062_9158# a_28066_9158# 0.843f
C4068 rowoff_n[13] a_35494_15544# 0.0133f
C4069 row_n[10] a_27974_12170# 0.0437f
C4070 vcm a_28370_17230# 0.155f
C4071 a_2275_13198# a_7894_13174# 0.136f
C4072 rowon_n[14] a_27062_16186# 0.248f
C4073 VDD a_26458_7512# 0.0779f
C4074 m2_1732_7974# ctop 0.0428f
C4075 col_n[16] a_2275_14202# 0.113f
C4076 ctop a_6982_11166# 4.11f
C4077 col_n[21] a_2275_3158# 0.113f
C4078 a_2275_18218# a_29374_18234# 0.145f
C4079 a_16930_18194# a_17022_18194# 0.0991f
C4080 VDD a_15926_16186# 0.181f
C4081 a_2275_1150# a_19334_1166# 0.126f
C4082 a_2475_1150# a_21950_1126# 0.264f
C4083 a_11910_1126# a_12002_1126# 0.0991f
C4084 m2_21812_946# m2_22816_946# 0.843f
C4085 col[24] a_27062_13174# 0.367f
C4086 vcm a_21950_11166# 0.1f
C4087 col[6] a_2275_11190# 0.0899f
C4088 a_18026_11166# a_18026_10162# 0.843f
C4089 col[21] a_23958_3134# 0.0682f
C4090 row_n[14] a_4974_16186# 0.282f
C4091 VDD a_18026_1126# 0.994f
C4092 col[31] a_33998_15182# 0.0682f
C4093 a_11910_15182# a_12306_15222# 0.0313f
C4094 a_2275_15206# a_22954_15182# 0.136f
C4095 VDD a_7382_10524# 0.0779f
C4096 ctop a_22042_15182# 4.11f
C4097 row_n[4] a_15014_6146# 0.282f
C4098 col_n[14] rowon_n[15] 0.111f
C4099 col_n[9] row_n[13] 0.298f
C4100 col_n[2] rowon_n[9] 0.111f
C4101 col_n[10] rowon_n[13] 0.111f
C4102 col_n[0] row_n[8] 0.298f
C4103 col_n[4] rowon_n[10] 0.111f
C4104 VDD row_n[7] 3.29f
C4105 col_n[3] row_n[10] 0.298f
C4106 col_n[5] row_n[11] 0.298f
C4107 col_n[11] row_n[14] 0.298f
C4108 col_n[7] row_n[12] 0.298f
C4109 col_n[6] rowon_n[11] 0.111f
C4110 col_n[13] row_n[15] 0.298f
C4111 col_n[1] row_n[9] 0.298f
C4112 col_n[8] rowon_n[12] 0.111f
C4113 col_n[12] rowon_n[14] 0.111f
C4114 sample rowon_n[7] 0.0935f
C4115 vcm rowon_n[8] 0.65f
C4116 a_2275_3158# a_35398_3174# 0.145f
C4117 col[26] a_2475_10186# 0.136f
C4118 rowon_n[8] a_14922_10162# 0.118f
C4119 col_n[9] a_12306_1166# 0.0839f
C4120 col_n[19] a_22346_13214# 0.084f
C4121 a_30074_8154# a_30378_8194# 0.0931f
C4122 a_30986_8154# a_31478_8516# 0.0658f
C4123 rowoff_n[10] a_7382_12532# 0.0133f
C4124 a_25358_1166# vcm 0.16f
C4125 col_n[16] rowoff_n[11] 0.0471f
C4126 row_n[6] a_3878_8154# 0.0437f
C4127 vcm a_2161_14202# 0.0169f
C4128 m2_6176_4386# rowon_n[2] 0.0322f
C4129 a_2475_12194# a_15014_12170# 0.316f
C4130 a_7986_12170# a_8990_12170# 0.843f
C4131 rowon_n[10] a_2966_12170# 0.248f
C4132 VDD a_33086_5142# 0.483f
C4133 m2_24248_18442# VDD 0.0456f
C4134 col_n[30] a_33486_7512# 0.0283f
C4135 VDD a_22442_14540# 0.0779f
C4136 a_2161_1150# m2_1732_946# 0.0454f
C4137 a_2475_1150# m2_2736_946# 0.287f
C4138 a_26970_5142# a_27062_5142# 0.326f
C4139 rowoff_n[14] a_23446_16548# 0.0133f
C4140 a_2275_9182# a_5978_9158# 0.399f
C4141 col[23] a_2275_13198# 0.0899f
C4142 rowon_n[2] a_2475_4162# 0.31f
C4143 col[13] a_16018_11166# 0.367f
C4144 vcm a_17934_18194# 0.101f
C4145 col[28] a_2275_2154# 0.0899f
C4146 a_33086_15182# a_33086_14178# 0.843f
C4147 m2_15212_17438# rowon_n[15] 0.0322f
C4148 a_2475_14202# a_30074_14178# 0.316f
C4149 col[10] a_12914_1126# 0.0682f
C4150 m2_21236_13422# rowon_n[11] 0.0322f
C4151 VDD a_14010_8154# 0.483f
C4152 row_n[7] a_34394_9198# 0.0117f
C4153 m2_27260_9406# rowon_n[7] 0.0322f
C4154 m2_33284_5390# rowon_n[3] 0.0322f
C4155 rowon_n[11] a_35094_13174# 0.0141f
C4156 col[20] a_22954_13174# 0.0682f
C4157 m2_23820_946# vcm 0.353f
C4158 VDD a_2966_17190# 0.486f
C4159 a_21950_2130# a_22346_2170# 0.0313f
C4160 col_n[28] a_31078_7150# 0.251f
C4161 vcm rowoff_n[12] 0.533f
C4162 vcm a_20034_3134# 0.56f
C4163 a_11910_11166# a_12402_11528# 0.0658f
C4164 a_2275_11190# a_21038_11166# 0.399f
C4165 a_10998_11166# a_11302_11206# 0.0931f
C4166 col_n[8] a_11302_11206# 0.084f
C4167 m2_24824_18014# a_24962_18194# 0.225f
C4168 a_23046_16186# a_24050_16186# 0.843f
C4169 row_n[11] a_13006_13174# 0.282f
C4170 VDD a_29070_12170# 0.483f
C4171 m2_18800_18014# m3_17928_18146# 0.0341f
C4172 col_n[13] a_2475_9182# 0.0531f
C4173 rowon_n[15] a_12914_17190# 0.118f
C4174 col_n[19] a_22442_5504# 0.0283f
C4175 row_n[1] a_23046_3134# 0.282f
C4176 rowoff_n[1] a_8990_3134# 0.294f
C4177 col_n[29] a_32482_17552# 0.0283f
C4178 rowon_n[5] a_22954_7150# 0.118f
C4179 vcm a_35094_7150# 0.165f
C4180 rowoff_n[12] a_29982_14178# 0.202f
C4181 a_2275_8178# a_11302_8194# 0.144f
C4182 a_2475_8178# a_13918_8154# 0.264f
C4183 a_7894_8154# a_7986_8154# 0.326f
C4184 col[3] a_2475_6170# 0.136f
C4185 row_n[3] a_10298_5182# 0.0117f
C4186 col[2] a_4974_9158# 0.367f
C4187 VDD a_9994_15182# 0.483f
C4188 m3_3872_18146# a_3970_17190# 0.0303f
C4189 col[9] a_11910_11166# 0.0682f
C4190 a_2275_5166# a_4882_5142# 0.136f
C4191 a_2966_5142# a_3970_5142# 0.843f
C4192 m2_1732_5966# sample_n 0.0522f
C4193 col_n[17] a_20034_5142# 0.251f
C4194 m2_21812_946# m3_22948_1078# 0.0341f
C4195 col_n[10] a_2275_12194# 0.113f
C4196 vcm a_16018_10162# 0.56f
C4197 rowon_n[4] rowoff_n[4] 20.2f
C4198 col_n[15] a_2275_1150# 0.0948f
C4199 a_2475_10186# a_28978_10162# 0.264f
C4200 col_n[27] a_30074_17190# 0.251f
C4201 a_2275_10186# a_26362_10202# 0.144f
C4202 rowoff_n[15] a_11398_17552# 0.0133f
C4203 row_n[14] a_33998_16186# 0.0437f
C4204 col_n[24] a_26970_7150# 0.0765f
C4205 a_26058_15182# a_26362_15222# 0.0931f
C4206 a_26970_15182# a_27462_15544# 0.0658f
C4207 VDD a_35398_10202# 0.0882f
C4208 m2_12776_18014# ctop 0.0422f
C4209 col_n[30] a_2475_11190# 0.0531f
C4210 col[0] a_2275_9182# 0.099f
C4211 a_33086_3134# a_34090_3134# 0.843f
C4212 m2_5172_3382# row_n[1] 0.0128f
C4213 vcm a_6282_4178# 0.155f
C4214 col_n[8] a_11398_3496# 0.0283f
C4215 a_2275_7174# a_19942_7150# 0.136f
C4216 col_n[18] a_21438_15544# 0.0283f
C4217 vcm a_31078_14178# 0.56f
C4218 a_22954_12170# a_23046_12170# 0.326f
C4219 VDD a_27974_4138# 0.181f
C4220 col[20] a_2475_8178# 0.136f
C4221 row_n[8] a_21038_10162# 0.282f
C4222 rowoff_n[7] a_10906_9158# 0.202f
C4223 rowon_n[12] a_20946_14178# 0.118f
C4224 a_2475_4162# a_12002_4138# 0.316f
C4225 a_24050_5142# a_24050_4138# 0.843f
C4226 m3_33992_18146# ctop 0.209f
C4227 row_n[10] rowoff_n[10] 0.209f
C4228 m2_14208_16434# row_n[14] 0.0128f
C4229 m2_20232_12418# row_n[10] 0.0128f
C4230 vcm a_21342_8194# 0.155f
C4231 m2_26256_8402# row_n[6] 0.0128f
C4232 a_2275_9182# a_35002_9158# 0.136f
C4233 col_n[27] a_2275_14202# 0.113f
C4234 rowoff_n[13] a_17934_15182# 0.202f
C4235 a_17934_9158# a_18330_9198# 0.0313f
C4236 m2_32280_4386# row_n[2] 0.0128f
C4237 row_n[10] a_8290_12210# 0.0117f
C4238 rowon_n[2] a_30986_4138# 0.118f
C4239 col_n[6] a_8990_3134# 0.251f
C4240 ctop a_34090_3134# 4.06f
C4241 vcm a_12002_17190# 0.56f
C4242 col_n[16] a_19030_15182# 0.251f
C4243 VDD a_8898_7150# 0.181f
C4244 rowoff_n[5] a_19942_7150# 0.202f
C4245 col_n[13] a_15926_5142# 0.0765f
C4246 a_7894_18194# a_8386_18556# 0.0658f
C4247 a_2275_18218# a_13006_18194# 0.0924f
C4248 row_n[0] a_18330_2170# 0.0117f
C4249 col_n[23] a_25966_17190# 0.0765f
C4250 a_2475_1150# a_3878_1126# 0.285f
C4251 a_2275_1150# a_2874_1126# 0.136f
C4252 m2_1732_1950# a_2475_2154# 0.139f
C4253 col[17] a_2275_11190# 0.0899f
C4254 vcm a_14922_2130# 0.1f
C4255 a_14010_6146# a_15014_6146# 0.843f
C4256 a_2475_6170# a_27062_6146# 0.316f
C4257 rowoff_n[3] a_28978_5142# 0.202f
C4258 row_n[2] a_8898_4138# 0.0437f
C4259 vcm a_3878_11166# 0.1f
C4260 VDD a_34490_2492# 0.0779f
C4261 rowon_n[6] a_7986_8154# 0.248f
C4262 m2_11196_17438# a_10998_17190# 0.165f
C4263 m2_20808_18014# a_21038_17190# 0.843f
C4264 col_n[7] a_10394_13536# 0.0283f
C4265 ctop a_15014_6146# 4.11f
C4266 a_2275_15206# a_3270_15222# 0.144f
C4267 a_2475_15206# a_5886_15182# 0.264f
C4268 col_n[1] rowon_n[3] 0.111f
C4269 sample row_n[2] 0.423f
C4270 col_n[20] row_n[13] 0.298f
C4271 col_n[25] rowon_n[15] 0.111f
C4272 col_n[7] rowon_n[6] 0.111f
C4273 col_n[16] row_n[11] 0.298f
C4274 col_n[14] row_n[10] 0.298f
C4275 col_n[21] rowon_n[13] 0.111f
C4276 col_n[10] row_n[8] 0.298f
C4277 col_n[19] rowon_n[12] 0.111f
C4278 VDD rowon_n[1] 3.04f
C4279 col_n[15] rowon_n[10] 0.111f
C4280 col_n[23] rowon_n[14] 0.111f
C4281 col_n[4] row_n[5] 0.298f
C4282 col_n[9] rowon_n[7] 0.111f
C4283 col_n[0] rowon_n[2] 0.111f
C4284 col_n[24] row_n[15] 0.298f
C4285 col_n[18] row_n[12] 0.298f
C4286 col_n[8] row_n[7] 0.298f
C4287 col_n[28] col_n[29] 0.0104f
C4288 col_n[6] row_n[6] 0.298f
C4289 col_n[12] row_n[9] 0.298f
C4290 col_n[2] row_n[4] 0.298f
C4291 VDD a_23958_11166# 0.181f
C4292 col_n[11] rowon_n[8] 0.111f
C4293 col_n[5] rowon_n[5] 0.111f
C4294 col_n[22] row_n[14] 0.298f
C4295 col_n[17] rowon_n[11] 0.111f
C4296 vcm row_n[3] 0.616f
C4297 col_n[3] rowon_n[4] 0.111f
C4298 col_n[13] rowon_n[9] 0.111f
C4299 col[26] a_29070_2130# 0.367f
C4300 a_2275_3158# a_18026_3134# 0.399f
C4301 col_n[27] rowoff_n[11] 0.0471f
C4302 a_2475_18218# a_10998_18194# 0.0299f
C4303 rowoff_n[8] a_20434_10524# 0.0133f
C4304 a_31990_1126# a_2275_1150# 0.136f
C4305 vcm a_29982_6146# 0.1f
C4306 a_4974_8154# a_4974_7150# 0.843f
C4307 m2_30272_13422# a_30074_13174# 0.165f
C4308 col_n[7] a_2475_7174# 0.0531f
C4309 vcm a_17326_15222# 0.155f
C4310 a_32994_13174# a_33390_13214# 0.0313f
C4311 VDD a_15414_5504# 0.0779f
C4312 a_27366_1166# VDD 0.0149f
C4313 col_n[21] a_24354_2170# 0.084f
C4314 ctop a_30074_10162# 4.11f
C4315 row_n[15] a_19030_17190# 0.282f
C4316 a_2275_17214# a_18330_17230# 0.144f
C4317 a_2475_17214# a_20946_17190# 0.264f
C4318 rowoff_n[6] a_29470_8516# 0.0133f
C4319 VDD a_4882_14178# 0.181f
C4320 col_n[5] a_7986_13174# 0.251f
C4321 col_n[2] a_4882_3134# 0.0765f
C4322 col_n[12] a_14922_15182# 0.0765f
C4323 a_17022_5142# a_17326_5182# 0.0931f
C4324 a_17934_5142# a_18426_5504# 0.0658f
C4325 row_n[5] a_29070_7150# 0.282f
C4326 a_2275_5166# a_33086_5142# 0.399f
C4327 rowon_n[9] a_28978_11166# 0.118f
C4328 vcm a_10906_9158# 0.1f
C4329 a_29070_10162# a_30074_10162# 0.843f
C4330 rowoff_n[14] a_5886_16186# 0.202f
C4331 m2_1732_15002# a_1957_15206# 0.245f
C4332 a_2275_14202# a_11910_14178# 0.136f
C4333 row_n[7] a_16322_9198# 0.0117f
C4334 VDD a_30474_9520# 0.0779f
C4335 ctop a_10998_13174# 4.11f
C4336 col_n[11] rowoff_n[12] 0.0471f
C4337 VDD a_19942_18194# 0.343f
C4338 col_n[4] a_2275_10186# 0.113f
C4339 a_2475_2154# a_25966_2130# 0.264f
C4340 a_2275_2154# a_23350_2170# 0.144f
C4341 a_13918_2130# a_14010_2130# 0.326f
C4342 m2_27836_946# VDD 1f
C4343 vcm a_1957_3158# 0.139f
C4344 row_n[9] a_6890_11166# 0.0437f
C4345 col[25] a_28066_12170# 0.367f
C4346 rowoff_n[9] a_30074_11166# 0.294f
C4347 col[22] a_24962_2130# 0.0682f
C4348 rowon_n[13] a_5978_15182# 0.248f
C4349 m2_21236_11414# a_21038_11166# 0.165f
C4350 vcm a_25966_13174# 0.1f
C4351 a_2275_11190# a_2966_11166# 0.399f
C4352 a_20034_12170# a_20034_11166# 0.843f
C4353 a_2475_11190# a_3970_11166# 0.316f
C4354 VDD a_22042_3134# 0.483f
C4355 col_n[24] a_2475_9182# 0.0531f
C4356 m2_32856_18014# a_2275_18218# 0.28f
C4357 ctop a_2275_7174# 0.0683f
C4358 a_13918_16186# a_14314_16226# 0.0313f
C4359 a_2275_16210# a_26970_16186# 0.136f
C4360 VDD a_11398_12532# 0.0779f
C4361 rowon_n[3] a_16018_5142# 0.248f
C4362 a_32082_1126# m2_31852_946# 0.0249f
C4363 ctop a_26058_17190# 4.06f
C4364 col_n[20] a_23350_12210# 0.084f
C4365 col[9] a_2475_17214# 0.136f
C4366 a_32082_9158# a_32386_9198# 0.0931f
C4367 a_32994_9158# a_33486_9520# 0.0658f
C4368 col[14] a_2475_6170# 0.136f
C4369 vcm a_6890_16186# 0.1f
C4370 a_2475_13198# a_19030_13174# 0.316f
C4371 a_9994_13174# a_10998_13174# 0.843f
C4372 VDD a_2874_6146# 0.182f
C4373 col_n[31] a_34490_6508# 0.0283f
C4374 m2_28840_18014# a_2475_18218# 0.286f
C4375 VDD a_26458_16548# 0.0779f
C4376 row_n[12] a_27062_14178# 0.282f
C4377 col_n[21] a_2275_12194# 0.113f
C4378 ctop rowoff_n[5] 0.177f
C4379 row_n[1] rowoff_n[0] 0.085f
C4380 vcm a_8990_1126# 0.165f
C4381 col_n[26] a_2275_1150# 0.113f
C4382 m2_4168_15430# rowon_n[13] 0.0322f
C4383 a_28978_6146# a_29070_6146# 0.326f
C4384 m2_10192_11414# rowon_n[9] 0.0322f
C4385 m2_16216_7398# rowon_n[5] 0.0322f
C4386 m2_32856_946# m2_33284_1374# 0.165f
C4387 m2_22240_3382# rowon_n[1] 0.0322f
C4388 m2_12200_9406# a_12002_9158# 0.165f
C4389 a_2275_10186# a_9994_10162# 0.399f
C4390 col[14] a_17022_10162# 0.367f
C4391 row_n[14] a_14314_16226# 0.0117f
C4392 m2_1732_2954# VDD 0.856f
C4393 col[21] a_23958_12170# 0.0682f
C4394 a_2475_15206# a_34090_15182# 0.316f
C4395 VDD a_18026_10162# 0.483f
C4396 col[11] a_2275_9182# 0.0899f
C4397 row_n[4] a_24354_6186# 0.0117f
C4398 col_n[29] a_32082_6146# 0.251f
C4399 a_23958_3134# a_24354_3174# 0.0313f
C4400 m2_31276_5390# a_31078_5142# 0.165f
C4401 vcm a_24050_5142# 0.56f
C4402 rowoff_n[10] a_18026_12170# 0.294f
C4403 col_n[9] a_12306_10202# 0.084f
C4404 m2_31276_16434# rowon_n[14] 0.0322f
C4405 row_n[6] a_14922_8154# 0.0437f
C4406 col[31] a_2475_8178# 0.136f
C4407 a_13918_12170# a_14410_12532# 0.0658f
C4408 a_2275_12194# a_25054_12170# 0.399f
C4409 a_13006_12170# a_13310_12210# 0.0931f
C4410 m2_10768_946# col[8] 0.425f
C4411 rowon_n[10] a_14010_12170# 0.248f
C4412 a_25054_17190# a_26058_17190# 0.843f
C4413 VDD a_33086_14178# 0.483f
C4414 col_n[20] a_23446_4500# 0.0283f
C4415 row_n[8] a_2966_10162# 0.281f
C4416 rowon_n[0] a_24050_2130# 0.248f
C4417 rowoff_n[0] a_9994_2130# 0.294f
C4418 col_n[30] a_33486_16548# 0.0283f
C4419 rowon_n[12] a_2275_14202# 1.79f
C4420 col_n[1] a_2475_5166# 0.0531f
C4421 m2_14784_946# ctop 0.0428f
C4422 vcm a_4974_8154# 0.56f
C4423 a_2275_9182# a_15318_9198# 0.144f
C4424 a_9902_9158# a_9994_9158# 0.326f
C4425 a_2475_9182# a_17934_9158# 0.264f
C4426 rowoff_n[14] a_34090_16186# 0.294f
C4427 m2_1732_18014# sample 0.2f
C4428 col[3] a_5978_8154# 0.367f
C4429 col[28] a_2275_11190# 0.0899f
C4430 m2_3740_18014# col[1] 0.347f
C4431 row_n[0] a_2475_2154# 0.405f
C4432 col[10] a_12914_10162# 0.0682f
C4433 VDD a_14010_17190# 0.484f
C4434 m2_22240_3382# a_22042_3134# 0.165f
C4435 col_n[18] a_21038_4138# 0.251f
C4436 m3_32988_1078# VDD 0.0157f
C4437 vcm a_29374_3174# 0.155f
C4438 row_n[9] a_35094_11166# 0.0123f
C4439 a_4882_6146# a_5278_6186# 0.0313f
C4440 a_2275_6170# a_8898_6146# 0.136f
C4441 col_n[28] a_31078_16186# 0.251f
C4442 rowon_n[13] a_35002_15182# 0.118f
C4443 col_n[25] a_27974_6146# 0.0765f
C4444 vcm a_20034_12170# 0.56f
C4445 col_n[20] rowon_n[7] 0.111f
C4446 vcm en_bit_n[1] 0.0193f
C4447 col_n[29] row_n[12] 0.298f
C4448 col_n[9] row_n[2] 0.298f
C4449 col_n[16] rowon_n[5] 0.111f
C4450 col_n[28] rowon_n[11] 0.111f
C4451 col_n[1] en_C0_n 0.186f
C4452 col_n[10] rowon_n[2] 0.111f
C4453 col_n[13] row_n[4] 0.298f
C4454 col_n[6] rowon_n[0] 0.111f
C4455 col_n[31] row_n[13] 0.298f
C4456 col_n[30] rowon_n[12] 0.111f
C4457 col_n[8] rowon_n[1] 0.111f
C4458 a_2475_11190# a_32994_11166# 0.264f
C4459 col_n[2] ctop 0.0594f
C4460 col_n[14] rowon_n[4] 0.111f
C4461 col_n[17] row_n[6] 0.298f
C4462 a_2275_11190# a_30378_11206# 0.144f
C4463 col_n[15] row_n[5] 0.298f
C4464 col_n[11] row_n[3] 0.298f
C4465 col_n[27] row_n[11] 0.298f
C4466 col_n[24] rowon_n[9] 0.111f
C4467 col_n[26] rowon_n[10] 0.111f
C4468 col_n[12] rowon_n[3] 0.111f
C4469 col_n[25] row_n[10] 0.298f
C4470 col_n[23] row_n[9] 0.298f
C4471 col_n[22] rowon_n[8] 0.111f
C4472 col_n[21] row_n[8] 0.298f
C4473 col_n[5] row_n[0] 0.298f
C4474 col_n[19] row_n[7] 0.298f
C4475 col_n[7] row_n[1] 0.298f
C4476 col_n[18] rowon_n[6] 0.111f
C4477 VDD analog_in 0.396f
C4478 VDD a_16930_2130# 0.181f
C4479 row_n[11] a_22346_13214# 0.0117f
C4480 a_28978_16186# a_29470_16548# 0.0658f
C4481 a_28066_16186# a_28370_16226# 0.0931f
C4482 a_25358_1166# col_n[22] 0.0839f
C4483 m2_32856_18014# m3_32988_18146# 3.79f
C4484 col[1] a_3878_8154# 0.0682f
C4485 row_n[1] a_32386_3174# 0.0117f
C4486 col_n[9] a_12402_2492# 0.0283f
C4487 rowoff_n[8] a_2161_10186# 0.0226f
C4488 col_n[18] a_2475_7174# 0.0531f
C4489 row_n[13] a_12914_15182# 0.0437f
C4490 vcm a_10298_6186# 0.155f
C4491 col_n[19] a_22442_14540# 0.0283f
C4492 rowoff_n[11] a_5978_13174# 0.294f
C4493 a_2275_8178# a_23958_8154# 0.136f
C4494 vcm a_35094_16186# 0.165f
C4495 a_24962_13174# a_25054_13174# 0.326f
C4496 VDD a_31990_6146# 0.181f
C4497 row_n[3] a_22954_5142# 0.0437f
C4498 m2_3164_14426# row_n[12] 0.0128f
C4499 rowon_n[7] a_22042_9158# 0.248f
C4500 a_2475_17214# a_2275_17214# 2.76f
C4501 a_1957_17214# a_2161_17214# 0.115f
C4502 rowoff_n[6] a_11910_8154# 0.202f
C4503 m2_9188_10410# row_n[8] 0.0128f
C4504 col[3] a_2475_15206# 0.136f
C4505 m2_15212_6394# row_n[4] 0.0128f
C4506 col[8] a_2475_4162# 0.136f
C4507 a_2475_5166# a_16018_5142# 0.316f
C4508 a_26058_6146# a_26058_5142# 0.843f
C4509 m2_19804_18014# col_n[17] 0.243f
C4510 vcm a_25358_10202# 0.155f
C4511 a_25966_1126# col[23] 0.0682f
C4512 col_n[7] a_9994_2130# 0.251f
C4513 a_19942_10162# a_20338_10202# 0.0313f
C4514 rowoff_n[15] a_22042_17190# 0.294f
C4515 col_n[17] a_20034_14178# 0.251f
C4516 rowoff_n[4] a_20946_6146# 0.202f
C4517 col_n[14] a_16930_4138# 0.0765f
C4518 ctop a_3970_4138# 4.11f
C4519 col_n[22] rowoff_n[12] 0.0471f
C4520 col_n[15] a_2275_10186# 0.113f
C4521 VDD a_12914_9158# 0.181f
C4522 col_n[24] a_26970_16186# 0.0765f
C4523 m2_30272_15430# row_n[13] 0.0128f
C4524 a_3970_2130# a_4274_2170# 0.0931f
C4525 a_4882_2130# a_5374_2492# 0.0658f
C4526 a_2275_2154# a_6982_2130# 0.399f
C4527 m2_35292_11414# row_n[9] 0.0128f
C4528 vcm a_18938_4138# 0.1f
C4529 rowoff_n[9] a_12402_11528# 0.0133f
C4530 rowon_n[1] a_9902_3134# 0.118f
C4531 a_2475_7174# a_31078_7150# 0.316f
C4532 rowoff_n[2] a_29982_4138# 0.202f
C4533 a_16018_7150# a_17022_7150# 0.843f
C4534 col[0] a_2275_18218# 0.099f
C4535 col[5] a_2275_7174# 0.0899f
C4536 vcm a_6282_13214# 0.155f
C4537 col_n[8] a_11398_12532# 0.0283f
C4538 VDD a_4370_3496# 0.0779f
C4539 col_n[31] a_34394_3174# 0.084f
C4540 ctop a_19030_8154# 4.11f
C4541 a_2475_16210# a_9902_16186# 0.264f
C4542 a_2275_16210# a_7286_16226# 0.144f
C4543 a_5886_16186# a_5978_16186# 0.326f
C4544 VDD a_27974_13174# 0.181f
C4545 col[20] a_2475_17214# 0.136f
C4546 row_n[8] a_30378_10202# 0.0117f
C4547 rowoff_n[7] a_21438_9520# 0.0133f
C4548 col[25] a_2475_6170# 0.136f
C4549 a_2275_4162# a_22042_4138# 0.399f
C4550 m3_9896_1078# ctop 0.21f
C4551 vcm a_33998_8154# 0.1f
C4552 rowoff_n[13] a_28466_15544# 0.0133f
C4553 a_6982_9158# a_6982_8154# 0.843f
C4554 row_n[10] a_20946_12170# 0.0437f
C4555 col_n[6] rowoff_n[13] 0.0471f
C4556 vcm a_21342_17230# 0.155f
C4557 rowon_n[14] a_20034_16186# 0.248f
C4558 VDD a_19430_7512# 0.0779f
C4559 rowoff_n[5] a_30474_7512# 0.0133f
C4560 col_n[6] a_8990_12170# 0.251f
C4561 ctop a_34090_12170# 4.06f
C4562 col[9] rowoff_n[9] 0.0901f
C4563 col[7] rowoff_n[7] 0.0901f
C4564 col[4] rowoff_n[4] 0.0901f
C4565 col[6] rowoff_n[6] 0.0901f
C4566 col[2] rowoff_n[2] 0.0901f
C4567 col[0] rowoff_n[0] 0.0901f
C4568 col_n[3] a_5886_2130# 0.0765f
C4569 col[8] rowoff_n[8] 0.0901f
C4570 col[1] rowoff_n[1] 0.0901f
C4571 col[3] rowoff_n[3] 0.0901f
C4572 col[5] rowoff_n[5] 0.0901f
C4573 a_2275_18218# a_22346_18234# 0.145f
C4574 row_n[0] a_30986_2130# 0.0437f
C4575 VDD a_8898_16186# 0.181f
C4576 a_2275_1150# a_12306_1166# 0.145f
C4577 a_2475_1150# a_14922_1126# 0.264f
C4578 col_n[13] a_15926_14178# 0.0765f
C4579 rowon_n[4] a_30074_6146# 0.248f
C4580 a_19942_6146# a_20434_6508# 0.0658f
C4581 a_19030_6146# a_19334_6186# 0.0931f
C4582 vcm a_14922_11166# 0.1f
C4583 a_31078_11166# a_32082_11166# 0.843f
C4584 col[22] a_2275_9182# 0.0899f
C4585 VDD a_10998_1126# 0.035f
C4586 a_2275_15206# a_15926_15182# 0.136f
C4587 VDD a_34490_11528# 0.0779f
C4588 ctop a_15014_15182# 4.11f
C4589 rowon_n[0] m2_27260_2378# 0.0322f
C4590 row_n[4] a_7986_6146# 0.282f
C4591 rowon_n[8] a_7894_10162# 0.118f
C4592 a_15926_3134# a_16018_3134# 0.326f
C4593 col[26] a_29070_11166# 0.367f
C4594 a_2275_3158# a_27366_3174# 0.144f
C4595 a_2475_3158# a_29982_3134# 0.264f
C4596 rowoff_n[8] a_31078_10162# 0.294f
C4597 rowoff_n[11] a_35002_13174# 0.202f
C4598 vcm a_29982_15182# 0.1f
C4599 a_22042_13174# a_22042_12170# 0.843f
C4600 a_2475_12194# a_7986_12170# 0.316f
C4601 VDD a_26058_5142# 0.483f
C4602 m2_10192_18442# VDD 0.0456f
C4603 row_n[15] a_28370_17230# 0.0117f
C4604 col_n[7] a_2475_16210# 0.0531f
C4605 a_2275_17214# a_30986_17190# 0.136f
C4606 a_15926_17190# a_16322_17230# 0.0313f
C4607 VDD a_15414_14540# 0.0779f
C4608 col_n[12] a_2475_5166# 0.0531f
C4609 a_31078_2130# m2_31276_2378# 0.165f
C4610 col_n[21] a_24354_11206# 0.084f
C4611 col_n[2] a_4882_12170# 0.0765f
C4612 a_35002_10162# a_35494_10524# 0.0658f
C4613 rowoff_n[14] a_16418_16548# 0.0133f
C4614 vcm a_10906_18194# 0.101f
C4615 m2_20232_1374# a_20034_1126# 0.165f
C4616 m3_23952_1078# a_24050_2130# 0.0302f
C4617 a_12002_14178# a_13006_14178# 0.843f
C4618 col[2] a_2475_2154# 0.136f
C4619 a_2475_14202# a_23046_14178# 0.316f
C4620 row_n[7] a_28978_9158# 0.0437f
C4621 VDD a_6982_8154# 0.483f
C4622 m2_5172_5390# rowon_n[3] 0.0322f
C4623 rowon_n[11] a_28066_13174# 0.248f
C4624 VDD a_30474_18556# 0.0858f
C4625 a_2275_2154# a_34394_2170# 0.144f
C4626 m3_28972_18146# VDD 0.0277f
C4627 col_n[28] row_n[6] 0.298f
C4628 vcm col[7] 5.46f
C4629 col_n[24] row_n[4] 0.298f
C4630 col_n[30] row_n[7] 0.298f
C4631 col_n[26] row_n[5] 0.298f
C4632 col_n[20] row_n[2] 0.298f
C4633 col_n[21] rowon_n[2] 0.111f
C4634 vcm a_13006_3134# 0.56f
C4635 col_n[23] rowon_n[3] 0.111f
C4636 col_n[3] col[4] 7.13f
C4637 col_n[13] ctop 0.0594f
C4638 col_n[25] rowon_n[4] 0.111f
C4639 col_n[17] rowon_n[0] 0.111f
C4640 col_n[16] row_n[0] 0.297f
C4641 col_n[31] rowon_n[7] 0.111f
C4642 col_n[29] rowon_n[6] 0.111f
C4643 VDD col[10] 3.83f
C4644 col_n[22] row_n[3] 0.298f
C4645 col_n[18] row_n[1] 0.298f
C4646 col_n[19] rowon_n[1] 0.111f
C4647 col_n[27] rowon_n[5] 0.111f
C4648 a_30986_7150# a_31078_7150# 0.326f
C4649 col_n[9] a_2275_8178# 0.113f
C4650 col[15] a_18026_9158# 0.367f
C4651 vcm a_1957_12194# 0.139f
C4652 a_2275_11190# a_14010_11166# 0.399f
C4653 col[22] a_24962_11166# 0.0682f
C4654 m2_19804_18014# a_20034_18194# 0.0249f
C4655 row_n[11] a_5978_13174# 0.282f
C4656 col_n[30] a_33086_5142# 0.251f
C4657 VDD a_22042_12170# 0.483f
C4658 m2_8760_18014# m3_9896_18146# 0.0341f
C4659 rowon_n[15] a_5886_17190# 0.118f
C4660 ctop a_2275_16210# 0.0683f
C4661 m2_20232_14426# rowon_n[12] 0.0322f
C4662 m2_1732_9982# col[0] 0.0137f
C4663 m2_26256_10410# rowon_n[8] 0.0322f
C4664 col_n[29] a_2475_7174# 0.0531f
C4665 m2_32280_6394# rowon_n[4] 0.0322f
C4666 a_25966_4138# a_26362_4178# 0.0313f
C4667 row_n[1] a_16018_3134# 0.282f
C4668 rowoff_n[1] a_2475_3158# 3.9f
C4669 col_n[10] a_13310_9198# 0.084f
C4670 rowon_n[5] a_15926_7150# 0.118f
C4671 vcm a_28066_7150# 0.56f
C4672 rowoff_n[12] a_22954_14178# 0.202f
C4673 a_2275_8178# a_4274_8194# 0.144f
C4674 a_2475_8178# a_6890_8154# 0.264f
C4675 a_2275_13198# a_29070_13174# 0.399f
C4676 a_15014_13174# a_15318_13214# 0.0931f
C4677 a_15926_13174# a_16418_13536# 0.0658f
C4678 col[14] a_2475_15206# 0.136f
C4679 row_n[3] a_3270_5182# 0.0117f
C4680 col[19] a_2475_4162# 0.136f
C4681 col_n[21] a_24450_3496# 0.0283f
C4682 VDD a_2874_15182# 0.182f
C4683 col_n[31] a_34490_15544# 0.0283f
C4684 vcm a_18330_1166# 0.155f
C4685 m2_1732_3958# vcm 0.316f
C4686 m2_11772_946# m3_11904_1078# 3.79f
C4687 col_n[26] a_2275_10186# 0.113f
C4688 vcm a_8990_10162# 0.56f
C4689 a_2275_10186# a_19334_10202# 0.144f
C4690 a_11910_10162# a_12002_10162# 0.326f
C4691 a_2475_10186# a_21950_10162# 0.264f
C4692 rowoff_n[15] a_4370_17552# 0.0133f
C4693 row_n[14] a_26970_16186# 0.0437f
C4694 col[4] a_6982_7150# 0.367f
C4695 m2_8184_16434# a_7986_16186# 0.165f
C4696 rowoff_n[4] a_2275_6170# 0.151f
C4697 col[11] a_13918_9158# 0.0682f
C4698 col[11] a_2275_18218# 0.0899f
C4699 col_n[19] a_22042_3134# 0.251f
C4700 a_13006_3134# a_13006_2130# 0.843f
C4701 col_n[29] a_32082_15182# 0.251f
C4702 col[16] a_2275_7174# 0.0899f
C4703 col_n[26] a_28978_5142# 0.0765f
C4704 vcm a_33390_5182# 0.155f
C4705 a_2275_7174# a_12914_7150# 0.136f
C4706 a_6890_7150# a_7286_7190# 0.0313f
C4707 m2_27836_18014# vcm 0.353f
C4708 m2_27260_12418# a_27062_12170# 0.165f
C4709 vcm a_24050_14178# 0.56f
C4710 a_2275_12194# a_35398_12210# 0.145f
C4711 VDD a_20946_4138# 0.181f
C4712 col[31] a_2475_17214# 0.136f
C4713 a_30986_17190# a_31478_17552# 0.0658f
C4714 a_30074_17190# a_30378_17230# 0.0931f
C4715 row_n[8] a_14010_10162# 0.282f
C4716 col_n[10] a_13406_1488# 0.0283f
C4717 rowoff_n[7] a_3366_9520# 0.0133f
C4718 rowon_n[12] a_13918_14178# 0.118f
C4719 col_n[20] a_23446_13536# 0.0283f
C4720 a_2475_4162# a_4974_4138# 0.316f
C4721 m3_5880_18146# ctop 0.209f
C4722 col_n[17] rowoff_n[13] 0.0471f
C4723 m2_32856_18014# m2_33860_18014# 0.843f
C4724 vcm a_14314_8194# 0.155f
C4725 a_2275_9182# a_27974_9158# 0.136f
C4726 rowoff_n[13] a_10906_15182# 0.202f
C4727 col_n[1] a_2475_14202# 0.0531f
C4728 m2_4168_4386# row_n[2] 0.0128f
C4729 row_n[10] a_2275_12194# 19.2f
C4730 rowon_n[2] a_23958_4138# 0.118f
C4731 col_n[6] a_2475_3158# 0.0531f
C4732 col[13] rowoff_n[2] 0.0901f
C4733 ctop a_27062_3134# 4.11f
C4734 col[15] rowoff_n[4] 0.0901f
C4735 col[17] rowoff_n[6] 0.0901f
C4736 col[19] rowoff_n[8] 0.0901f
C4737 col[11] rowoff_n[0] 0.0901f
C4738 vcm a_4974_17190# 0.56f
C4739 col[20] rowoff_n[9] 0.0901f
C4740 col[18] rowoff_n[7] 0.0901f
C4741 col[12] rowoff_n[1] 0.0901f
C4742 col[14] rowoff_n[3] 0.0901f
C4743 col[16] rowoff_n[5] 0.0901f
C4744 rowon_n[14] a_1957_16210# 0.0172f
C4745 a_26970_14178# a_27062_14178# 0.326f
C4746 rowoff_n[5] a_12914_7150# 0.202f
C4747 a_2275_18218# a_5978_18194# 0.0924f
C4748 row_n[0] a_11302_2170# 0.0117f
C4749 col[3] a_5978_17190# 0.367f
C4750 vcm a_7894_2130# 0.1f
C4751 a_28066_7150# a_28066_6146# 0.843f
C4752 a_2475_6170# a_20034_6146# 0.316f
C4753 m2_18224_10410# a_18026_10162# 0.165f
C4754 col_n[18] a_21038_13174# 0.251f
C4755 m2_20808_946# col[18] 0.425f
C4756 rowoff_n[3] a_21950_5142# 0.202f
C4757 vcm a_29374_12210# 0.155f
C4758 col_n[15] a_17934_3134# 0.0765f
C4759 a_21950_11166# a_22346_11206# 0.0313f
C4760 VDD a_27462_2492# 0.0779f
C4761 m2_13204_17438# row_n[15] 0.0128f
C4762 m2_19228_13422# row_n[11] 0.0128f
C4763 m2_25252_9406# row_n[7] 0.0128f
C4764 col_n[25] a_27974_15182# 0.0765f
C4765 ctop a_7986_6146# 4.11f
C4766 m2_31276_5390# row_n[3] 0.0128f
C4767 row_n[11] a_35002_13174# 0.0437f
C4768 VDD a_16930_11166# 0.181f
C4769 rowon_n[15] a_34090_17190# 0.248f
C4770 col_n[3] a_2275_6170# 0.113f
C4771 a_2275_3158# a_10998_3134# 0.399f
C4772 a_5978_3134# a_6282_3174# 0.0931f
C4773 a_6890_3134# a_7382_3496# 0.0658f
C4774 col_n[1] rowoff_n[14] 0.0471f
C4775 a_2475_18218# a_3970_18194# 0.0299f
C4776 rowoff_n[8] a_13406_10524# 0.0133f
C4777 rowoff_n[1] a_30986_3134# 0.202f
C4778 col[1] a_3878_17190# 0.0682f
C4779 a_24962_1126# a_2275_1150# 0.136f
C4780 vcm a_22954_6146# 0.1f
C4781 m2_1732_12994# m2_2160_13422# 0.165f
C4782 a_2475_8178# a_35094_8154# 0.0299f
C4783 a_18026_8154# a_19030_8154# 0.843f
C4784 col_n[9] a_12402_11528# 0.0283f
C4785 col[4] rowoff_n[10] 0.0901f
C4786 col_n[18] a_2475_16210# 0.0531f
C4787 vcm a_10298_15222# 0.155f
C4788 col_n[23] a_2475_5166# 0.0531f
C4789 VDD a_8386_5504# 0.0779f
C4790 ctop a_23046_10162# 4.11f
C4791 row_n[15] a_12002_17190# 0.282f
C4792 a_2275_17214# a_11302_17230# 0.144f
C4793 a_2475_17214# a_13918_17190# 0.264f
C4794 a_7894_17190# a_7986_17190# 0.326f
C4795 rowoff_n[6] a_22442_8516# 0.0133f
C4796 VDD a_31990_15182# 0.181f
C4797 a_2275_5166# a_26058_5142# 0.399f
C4798 row_n[5] a_22042_7150# 0.282f
C4799 col[8] a_2475_13198# 0.136f
C4800 m2_9188_8402# a_8990_8154# 0.165f
C4801 rowon_n[9] a_21950_11166# 0.118f
C4802 col[13] a_2475_2154# 0.136f
C4803 a_27974_1126# a_28466_1488# 0.0658f
C4804 a_8990_10162# a_8990_9158# 0.843f
C4805 rowoff_n[4] a_31478_6508# 0.0133f
C4806 col_n[7] a_9994_11166# 0.251f
C4807 m2_30848_946# a_31078_2130# 0.843f
C4808 m2_20808_946# a_2475_1150# 0.286f
C4809 a_2275_14202# a_4882_14178# 0.136f
C4810 a_2966_14178# a_3970_14178# 0.843f
C4811 col_n[4] a_6890_1126# 0.0765f
C4812 VDD a_23446_9520# 0.0779f
C4813 row_n[7] a_9294_9198# 0.0117f
C4814 ctop a_3970_13174# 4.11f
C4815 col_n[14] a_16930_13174# 0.0765f
C4816 col_n[27] row_n[0] 0.298f
C4817 col_n[24] ctop 0.0594f
C4818 col_n[28] rowon_n[0] 0.111f
C4819 col_n[30] rowon_n[1] 0.111f
C4820 VDD col[21] 3.83f
C4821 col_n[29] row_n[1] 0.298f
C4822 vcm col[18] 5.46f
C4823 rowon_n[9] rowon_n[8] 0.0632f
C4824 col_n[31] row_n[2] 0.298f
C4825 col_n[9] col[9] 0.489f
C4826 VDD a_12914_18194# 0.343f
C4827 col_n[20] a_2275_8178# 0.113f
C4828 a_2475_2154# a_18938_2130# 0.264f
C4829 a_2275_2154# a_16322_2170# 0.144f
C4830 m2_28264_4386# a_28066_4138# 0.165f
C4831 m2_34864_2954# rowoff_n[1] 0.278f
C4832 m2_12200_1374# VDD 0.0194f
C4833 a_21038_7150# a_21342_7190# 0.0931f
C4834 rowoff_n[9] a_23046_11166# 0.294f
C4835 a_21950_7150# a_22442_7512# 0.0658f
C4836 vcm a_18938_13174# 0.1f
C4837 a_33086_12170# a_34090_12170# 0.843f
C4838 VDD a_15014_3134# 0.483f
C4839 m2_18800_18014# a_2275_18218# 0.28f
C4840 m2_6752_18014# a_7286_18234# 0.087f
C4841 col[5] a_2275_16210# 0.0899f
C4842 a_2275_16210# a_19942_16186# 0.136f
C4843 rowon_n[3] a_8990_5142# 0.248f
C4844 col[10] a_2275_5166# 0.0899f
C4845 VDD a_4370_12532# 0.0779f
C4846 col_n[31] a_34394_12210# 0.084f
C4847 col[27] a_30074_10162# 0.367f
C4848 ctop a_19030_17190# 4.06f
C4849 rowoff_n[7] a_32082_9158# 0.294f
C4850 a_17934_4138# a_18026_4138# 0.326f
C4851 a_2275_4162# a_31382_4178# 0.144f
C4852 a_2475_4162# a_33998_4138# 0.264f
C4853 col[25] a_2475_15206# 0.136f
C4854 m2_34864_17010# m2_34864_16006# 0.843f
C4855 col[30] a_2475_4162# 0.136f
C4856 vcm a_33998_17190# 0.1f
C4857 a_2475_13198# a_12002_13174# 0.316f
C4858 a_24050_14178# a_24050_13174# 0.843f
C4859 VDD a_30074_7150# 0.483f
C4860 col_n[22] a_25358_10202# 0.084f
C4861 a_17934_18194# a_18330_18234# 0.0313f
C4862 a_2275_18218# a_35002_18194# 0.136f
C4863 m2_14784_18014# a_2475_18218# 0.286f
C4864 VDD a_19430_16548# 0.0779f
C4865 a_12914_1126# a_13310_1166# 0.0313f
C4866 row_n[12] a_20034_14178# 0.282f
C4867 col_n[3] a_5886_11166# 0.0765f
C4868 vcm a_2475_1150# 1.05f
C4869 m2_25828_946# m2_26256_1374# 0.165f
C4870 row_n[2] a_30074_4138# 0.282f
C4871 a_2275_10186# a_2874_10162# 0.136f
C4872 a_2475_10186# a_3878_10162# 0.264f
C4873 row_n[14] a_7286_16226# 0.0117f
C4874 rowon_n[6] a_29982_8154# 0.118f
C4875 a_2475_15206# a_27062_15182# 0.316f
C4876 a_14010_15182# a_15014_15182# 0.843f
C4877 VDD a_10998_10162# 0.483f
C4878 col[22] a_2275_18218# 0.0899f
C4879 col[27] a_2275_7174# 0.0899f
C4880 row_n[4] a_17326_6186# 0.0117f
C4881 a_2475_18218# a_32994_18194# 0.264f
C4882 col[16] a_19030_8154# 0.367f
C4883 vcm a_17022_5142# 0.56f
C4884 a_32994_8154# a_33086_8154# 0.326f
C4885 rowoff_n[10] a_10998_12170# 0.294f
C4886 a_30986_1126# vcm 0.0989f
C4887 col[23] a_25966_10162# 0.0682f
C4888 m2_3164_16434# rowon_n[14] 0.0322f
C4889 row_n[6] a_7894_8154# 0.0437f
C4890 m2_9188_12418# rowon_n[10] 0.0322f
C4891 m2_15212_8402# rowon_n[6] 0.0322f
C4892 a_2275_12194# a_18026_12170# 0.399f
C4893 m2_21236_4386# rowon_n[2] 0.0322f
C4894 rowon_n[10] a_6982_12170# 0.248f
C4895 VDD a_2275_4162# 1.96f
C4896 col_n[31] a_34090_4138# 0.251f
C4897 m2_31852_18014# VDD 1.06f
C4898 a_4974_17190# a_4974_16186# 0.843f
C4899 VDD a_26058_14178# 0.483f
C4900 col_n[28] rowoff_n[13] 0.0471f
C4901 rowon_n[0] a_17022_2130# 0.248f
C4902 rowoff_n[0] a_2874_2130# 0.202f
C4903 col_n[11] a_14314_8194# 0.084f
C4904 col_n[12] a_2475_14202# 0.0531f
C4905 a_27974_5142# a_28370_5182# 0.0313f
C4906 col_n[17] a_2475_3158# 0.0531f
C4907 col[22] rowoff_n[0] 0.0901f
C4908 col[24] rowoff_n[2] 0.0901f
C4909 col[27] rowoff_n[5] 0.0901f
C4910 col[25] rowoff_n[3] 0.0901f
C4911 col[23] rowoff_n[1] 0.0901f
C4912 col[26] rowoff_n[4] 0.0901f
C4913 col[29] rowoff_n[7] 0.0901f
C4914 col[28] rowoff_n[6] 0.0901f
C4915 col[31] rowoff_n[9] 0.0901f
C4916 col[30] rowoff_n[8] 0.0901f
C4917 vcm a_32082_9158# 0.56f
C4918 a_2475_9182# a_10906_9158# 0.264f
C4919 rowoff_n[14] a_27062_16186# 0.294f
C4920 a_2275_9182# a_8290_9198# 0.144f
C4921 col[8] a_2475_18218# 0.136f
C4922 a_2275_14202# a_33086_14178# 0.399f
C4923 a_17934_14178# a_18426_14540# 0.0658f
C4924 col_n[22] a_25454_2492# 0.0283f
C4925 a_17022_14178# a_17326_14218# 0.0931f
C4926 m2_30272_17438# rowon_n[15] 0.0322f
C4927 m2_35292_13422# rowon_n[11] 0.0322f
C4928 col[2] a_2475_11190# 0.136f
C4929 VDD a_6982_17190# 0.484f
C4930 a_24050_2130# a_25054_2130# 0.843f
C4931 m3_4876_1078# VDD 0.0157f
C4932 vcm a_22346_3174# 0.155f
C4933 row_n[9] a_28066_11166# 0.282f
C4934 a_2475_6170# a_1957_6170# 0.0734f
C4935 en_bit_n[1] a_18426_1488# 0.018f
C4936 rowon_n[13] a_27974_15182# 0.118f
C4937 col[5] a_7986_6146# 0.367f
C4938 rowoff_n[3] a_3878_5142# 0.202f
C4939 vcm a_13006_12170# 0.56f
C4940 a_13918_11166# a_14010_11166# 0.326f
C4941 a_2475_11190# a_25966_11166# 0.264f
C4942 a_2275_11190# a_23350_11206# 0.144f
C4943 col_n[9] a_2275_17214# 0.113f
C4944 VDD a_9902_2130# 0.181f
C4945 m2_25828_18014# a_26362_18234# 0.087f
C4946 col[12] a_14922_8154# 0.0682f
C4947 col_n[14] a_2275_6170# 0.113f
C4948 row_n[11] a_15318_13214# 0.0117f
C4949 m2_23820_18014# m3_22948_18146# 0.0341f
C4950 col_n[12] rowoff_n[14] 0.0471f
C4951 col_n[20] a_23046_2130# 0.251f
C4952 col_n[30] a_33086_14178# 0.251f
C4953 a_15014_4138# a_15014_3134# 0.843f
C4954 col_n[27] a_29982_4138# 0.0765f
C4955 col[15] rowoff_n[10] 0.0901f
C4956 row_n[1] a_25358_3174# 0.0117f
C4957 col_n[29] a_2475_16210# 0.0531f
C4958 row_n[13] a_5886_15182# 0.0437f
C4959 vcm a_3270_6186# 0.155f
C4960 rowoff_n[12] a_33486_14540# 0.0133f
C4961 a_2275_8178# a_16930_8154# 0.136f
C4962 a_8898_8154# a_9294_8194# 0.0313f
C4963 col[4] a_2275_3158# 0.0899f
C4964 col_n[10] a_13310_18234# 0.084f
C4965 vcm a_28066_16186# 0.56f
C4966 VDD a_24962_6146# 0.181f
C4967 row_n[3] a_15926_5142# 0.0437f
C4968 a_32994_18194# a_33486_18556# 0.0658f
C4969 rowon_n[7] a_15014_9158# 0.248f
C4970 rowoff_n[6] a_4882_8154# 0.202f
C4971 col[19] a_2475_13198# 0.136f
C4972 col_n[21] a_24450_12532# 0.0283f
C4973 m3_6884_18146# a_6982_17190# 0.0303f
C4974 col[24] a_2475_2154# 0.136f
C4975 a_2475_5166# a_8990_5142# 0.316f
C4976 a_4974_5142# a_5978_5142# 0.843f
C4977 m2_26832_946# m3_27968_1078# 0.0341f
C4978 m3_32988_1078# col_n[30] 0.0116f
C4979 rowon_n[9] a_3878_11166# 0.118f
C4980 vcm a_18330_10202# 0.155f
C4981 a_2275_10186# a_31990_10162# 0.136f
C4982 rowoff_n[15] a_15014_17190# 0.294f
C4983 sample a_2161_6170# 0.0858f
C4984 rowoff_n[4] a_13918_6146# 0.202f
C4985 ctop a_31078_5142# 4.11f
C4986 a_28978_15182# a_29070_15182# 0.326f
C4987 rowon_n[6] row_n[6] 18.9f
C4988 VDD sample_n 14.5f
C4989 vcm col[29] 5.46f
C4990 col_n[14] col[15] 7.13f
C4991 row_n[14] ctop 0.186f
C4992 VDD a_5886_9158# 0.181f
C4993 col_n[31] a_2275_8178# 0.113f
C4994 col[4] a_6982_16186# 0.367f
C4995 col[11] a_13918_18194# 0.0682f
C4996 m2_2160_15430# row_n[13] 0.0194f
C4997 m2_8184_11414# row_n[9] 0.0128f
C4998 m2_14208_7398# row_n[5] 0.0128f
C4999 m2_20232_3382# row_n[1] 0.0128f
C5000 vcm a_11910_4138# 0.1f
C5001 col_n[19] a_22042_12170# 0.251f
C5002 a_2475_7174# a_24050_7150# 0.316f
C5003 a_30074_8154# a_30074_7150# 0.843f
C5004 rowoff_n[9] a_5374_11528# 0.0133f
C5005 rowon_n[1] a_2161_3158# 0.0177f
C5006 rowoff_n[2] a_22954_4138# 0.202f
C5007 col_n[16] a_18938_2130# 0.0765f
C5008 m2_34864_11990# a_35398_12210# 0.087f
C5009 col[16] a_2275_16210# 0.0899f
C5010 col_n[26] a_28978_14178# 0.0765f
C5011 vcm a_33390_14218# 0.155f
C5012 col[21] a_2275_5166# 0.0899f
C5013 a_23958_12170# a_24354_12210# 0.0313f
C5014 VDD a_31478_4500# 0.0779f
C5015 m2_34864_15002# VDD 0.772f
C5016 ctop a_12002_8154# 4.11f
C5017 VDD a_20946_13174# 0.181f
C5018 row_n[8] a_23350_10202# 0.0117f
C5019 rowoff_n[7] a_14410_9520# 0.0133f
C5020 rowoff_n[0] a_31990_2130# 0.202f
C5021 a_8898_4138# a_9390_4500# 0.0658f
C5022 a_7986_4138# a_8290_4178# 0.0931f
C5023 a_2275_4162# a_15014_4138# 0.399f
C5024 m3_34996_11118# ctop 0.209f
C5025 col_n[10] a_13406_10524# 0.0283f
C5026 m2_29268_16434# row_n[14] 0.0128f
C5027 m2_34864_11990# row_n[10] 0.267f
C5028 vcm a_26970_8154# 0.1f
C5029 a_20034_9158# a_21038_9158# 0.843f
C5030 rowoff_n[13] a_21438_15544# 0.0133f
C5031 row_n[10] a_13918_12170# 0.0437f
C5032 vcm a_14314_17230# 0.155f
C5033 rowon_n[14] a_13006_16186# 0.248f
C5034 VDD a_12402_7512# 0.0779f
C5035 rowoff_n[5] a_23446_7512# 0.0133f
C5036 col_n[6] a_2475_12194# 0.0531f
C5037 ctop a_27062_12170# 4.11f
C5038 a_2275_18218# a_15318_18234# 0.145f
C5039 a_9902_18194# a_9994_18194# 0.0991f
C5040 row_n[0] a_23958_2130# 0.0437f
C5041 col_n[11] a_2475_1150# 0.0531f
C5042 a_2475_1150# a_7894_1126# 0.264f
C5043 a_3878_1126# a_4274_1166# 0.0342f
C5044 a_2275_1150# a_5278_1166# 0.145f
C5045 a_4882_1126# a_4974_1126# 0.0991f
C5046 row_n[12] a_1957_14202# 0.187f
C5047 rowon_n[4] a_23046_6146# 0.248f
C5048 a_2275_6170# a_30074_6146# 0.399f
C5049 rowoff_n[3] a_32482_5504# 0.0133f
C5050 vcm a_7894_11166# 0.1f
C5051 a_10998_11166# a_10998_10162# 0.843f
C5052 col_n[8] a_10998_10162# 0.251f
C5053 VDD a_3970_1126# 0.995f
C5054 m2_14208_17438# a_14010_17190# 0.165f
C5055 a_4882_15182# a_5278_15222# 0.0313f
C5056 col_n[15] a_17934_12170# 0.0765f
C5057 a_2275_15206# a_8898_15182# 0.136f
C5058 VDD a_27462_11528# 0.0779f
C5059 ctop a_7986_15182# 4.11f
C5060 a_2475_3158# a_22954_3134# 0.264f
C5061 a_2275_3158# a_20338_3174# 0.144f
C5062 rowoff_n[8] a_24050_10162# 0.294f
C5063 col_n[3] a_2275_15206# 0.113f
C5064 row_n[13] a_34090_15182# 0.282f
C5065 rowoff_n[11] a_27974_13174# 0.202f
C5066 a_23046_8154# a_23350_8194# 0.0931f
C5067 col_n[8] a_2275_4162# 0.113f
C5068 a_23958_8154# a_24450_8516# 0.0658f
C5069 m2_33284_13422# a_33086_13174# 0.165f
C5070 vcm a_22954_15182# 0.1f
C5071 VDD a_19030_5142# 0.483f
C5072 a_32994_1126# VDD 0.412f
C5073 a_26458_1488# col_n[23] 0.0283f
C5074 row_n[15] a_21342_17230# 0.0117f
C5075 col[28] a_31078_9158# 0.367f
C5076 a_2275_17214# a_23958_17190# 0.136f
C5077 rowoff_n[6] a_33086_8154# 0.294f
C5078 col_n[23] a_2475_14202# 0.0531f
C5079 VDD a_8386_14540# 0.0779f
C5080 col_n[28] a_2475_3158# 0.0531f
C5081 en_bit_n[0] a_2275_1150# 0.0363f
C5082 a_19942_5142# a_20034_5142# 0.326f
C5083 row_n[5] a_31382_7190# 0.0117f
C5084 a_2275_5166# a_2275_4162# 0.0715f
C5085 m3_28972_1078# m3_29976_1078# 0.202f
C5086 col[19] a_2475_18218# 0.136f
C5087 rowoff_n[14] a_9390_16548# 0.0133f
C5088 m2_5172_15430# a_4974_15182# 0.165f
C5089 col[13] a_2475_11190# 0.136f
C5090 m2_14784_946# a_15014_1126# 0.0249f
C5091 a_2475_14202# a_16018_14178# 0.316f
C5092 a_26058_15182# a_26058_14178# 0.843f
C5093 col_n[23] a_26362_9198# 0.084f
C5094 VDD a_34090_9158# 0.483f
C5095 row_n[7] a_21950_9158# 0.0437f
C5096 rowon_n[11] a_21038_13174# 0.248f
C5097 col_n[4] a_6890_10162# 0.0765f
C5098 VDD a_23446_18556# 0.0858f
C5099 a_2275_2154# a_28978_2130# 0.136f
C5100 a_14922_2130# a_15318_2170# 0.0313f
C5101 m2_1732_2954# a_2161_3158# 0.0454f
C5102 m3_1046_19620# VDD 0.204f
C5103 vcm a_5978_3134# 0.56f
C5104 rowon_n[1] a_31078_3134# 0.248f
C5105 col_n[20] a_2275_17214# 0.113f
C5106 m2_24248_11414# a_24050_11166# 0.165f
C5107 col_n[25] a_2275_6170# 0.113f
C5108 a_4882_11166# a_5374_11528# 0.0658f
C5109 a_2275_11190# a_6982_11166# 0.399f
C5110 a_3970_11166# a_4274_11206# 0.0931f
C5111 col_n[23] rowoff_n[14] 0.0471f
C5112 a_16018_16186# a_17022_16186# 0.843f
C5113 a_2475_16210# a_31078_16186# 0.316f
C5114 VDD a_15014_12170# 0.483f
C5115 col[26] rowoff_n[10] 0.0901f
C5116 col[10] a_2275_14202# 0.0899f
C5117 col[17] a_20034_7150# 0.367f
C5118 m2_4168_6394# rowon_n[4] 0.0322f
C5119 m2_9188_2378# rowon_n[0] 0.0322f
C5120 col[15] a_2275_3158# 0.0899f
C5121 row_n[1] a_8990_3134# 0.282f
C5122 m2_34864_5966# a_2475_6170# 0.282f
C5123 col[24] a_26970_9158# 0.0682f
C5124 vcm a_21038_7150# 0.56f
C5125 rowon_n[5] a_8898_7150# 0.118f
C5126 a_34090_9158# a_34394_9198# 0.0931f
C5127 rowoff_n[12] a_15926_14178# 0.202f
C5128 a_35002_9158# a_35094_9158# 0.0991f
C5129 a_2275_13198# a_22042_13174# 0.399f
C5130 col[30] a_2475_13198# 0.136f
C5131 VDD a_30074_16186# 0.483f
C5132 col_n[12] a_15318_7190# 0.084f
C5133 row_n[12] a_29374_14218# 0.0117f
C5134 vcm a_11302_1166# 0.16f
C5135 m2_19228_15430# rowon_n[13] 0.0322f
C5136 a_29982_6146# a_30378_6186# 0.0313f
C5137 m2_25252_11414# rowon_n[9] 0.0322f
C5138 m2_31276_7398# rowon_n[5] 0.0322f
C5139 m2_15212_9406# a_15014_9158# 0.165f
C5140 rowon_n[11] col[0] 0.0318f
C5141 rowon_n[8] ctop 0.203f
C5142 row_n[13] col[3] 0.0342f
C5143 vcm a_2475_10186# 1.08f
C5144 col_n[20] col[20] 0.489f
C5145 row_n[12] col[1] 0.0342f
C5146 row_n[14] col[5] 0.0342f
C5147 rowon_n[12] col[2] 0.0323f
C5148 row_n[15] col[7] 0.0342f
C5149 rowon_n[14] col[6] 0.0323f
C5150 rowon_n[13] col[4] 0.0323f
C5151 rowon_n[15] col[8] 0.0323f
C5152 col_n[7] rowoff_n[15] 0.0471f
C5153 a_2475_10186# a_14922_10162# 0.264f
C5154 a_2275_10186# a_12306_10202# 0.144f
C5155 row_n[14] a_19942_16186# 0.0437f
C5156 m2_1732_16006# a_2275_16210# 0.191f
C5157 a_19942_15182# a_20434_15544# 0.0658f
C5158 a_19030_15182# a_19334_15222# 0.0931f
C5159 col[10] rowoff_n[11] 0.0901f
C5160 row_n[4] a_29982_6146# 0.0437f
C5161 a_26058_3134# a_27062_3134# 0.843f
C5162 rowon_n[8] a_29070_10162# 0.248f
C5163 col[27] a_2275_16210# 0.0899f
C5164 m2_34288_5390# a_34090_5142# 0.165f
C5165 vcm a_26362_5182# 0.155f
C5166 col[6] a_8990_5142# 0.367f
C5167 a_2275_7174# a_5886_7150# 0.136f
C5168 m2_13780_18014# vcm 0.353f
C5169 col[16] a_19030_17190# 0.367f
C5170 vcm a_17022_14178# 0.56f
C5171 col[13] a_15926_7150# 0.0682f
C5172 a_15926_12170# a_16018_12170# 0.326f
C5173 a_2475_12194# a_29982_12170# 0.264f
C5174 a_2275_12194# a_27366_12210# 0.144f
C5175 VDD a_13918_4138# 0.181f
C5176 row_n[0] m2_25252_2378# 0.0128f
C5177 VDD a_2275_13198# 1.96f
C5178 col_n[31] a_34090_13174# 0.251f
C5179 row_n[8] a_6982_10162# 0.282f
C5180 col_n[2] a_2275_2154# 0.113f
C5181 col_n[28] a_30986_3134# 0.0765f
C5182 rowon_n[12] a_6890_14178# 0.118f
C5183 a_17022_5142# a_17022_4138# 0.843f
C5184 col_n[1] a_4274_5182# 0.084f
C5185 m2_23820_946# ctop 0.0428f
C5186 m2_6176_7398# a_5978_7150# 0.165f
C5187 col_n[11] a_14314_17230# 0.084f
C5188 vcm a_7286_8194# 0.155f
C5189 m2_25828_18014# m2_26832_18014# 0.843f
C5190 rowoff_n[13] a_3366_15544# 0.0133f
C5191 a_2275_9182# a_20946_9158# 0.136f
C5192 a_10906_9158# a_11302_9198# 0.0313f
C5193 col_n[17] a_2475_12194# 0.0531f
C5194 rowon_n[2] a_16930_4138# 0.118f
C5195 vcm a_32082_18194# 0.165f
C5196 ctop rowoff_n[12] 0.177f
C5197 ctop a_20034_3134# 4.11f
C5198 col_n[22] a_2475_1150# 0.0531f
C5199 VDD a_28978_8154# 0.181f
C5200 rowoff_n[5] a_5886_7150# 0.202f
C5201 col_n[22] a_25454_11528# 0.0283f
C5202 row_n[0] a_4274_2170# 0.0117f
C5203 a_29982_2130# a_30474_2492# 0.0658f
C5204 a_29070_2130# a_29374_2170# 0.0931f
C5205 m2_25252_3382# a_25054_3134# 0.165f
C5206 vcm a_35002_3134# 0.101f
C5207 a_2475_6170# a_13006_6146# 0.316f
C5208 col[7] a_2475_9182# 0.136f
C5209 a_6982_6146# a_7986_6146# 0.843f
C5210 col_n[0] a_3366_5504# 0.0283f
C5211 rowoff_n[3] a_14922_5142# 0.202f
C5212 vcm a_22346_12210# 0.155f
C5213 a_2275_11190# a_34394_11206# 0.144f
C5214 VDD a_20434_2492# 0.0779f
C5215 col[5] a_7986_15182# 0.367f
C5216 m2_3164_5390# row_n[3] 0.0128f
C5217 m3_34996_5094# a_34090_5142# 0.0303f
C5218 col[2] a_4882_5142# 0.0682f
C5219 a_30986_16186# a_31078_16186# 0.326f
C5220 row_n[11] a_27974_13174# 0.0437f
C5221 VDD a_9902_11166# 0.181f
C5222 rowon_n[15] a_27062_17190# 0.248f
C5223 col[12] a_14922_17190# 0.0682f
C5224 col_n[14] a_2275_15206# 0.113f
C5225 col_n[19] a_2275_4162# 0.113f
C5226 col_n[20] a_23046_11166# 0.251f
C5227 a_2275_3158# a_3970_3134# 0.399f
C5228 rowoff_n[1] a_23958_3134# 0.202f
C5229 rowoff_n[8] a_6378_10524# 0.0133f
C5230 col_n[17] a_19942_1126# 0.0801f
C5231 vcm a_15926_6146# 0.1f
C5232 a_2475_8178# a_28066_8154# 0.316f
C5233 col_n[27] a_29982_13174# 0.0765f
C5234 a_32082_9158# a_32082_8154# 0.843f
C5235 vcm a_3270_15222# 0.155f
C5236 a_25966_13174# a_26362_13214# 0.0313f
C5237 VDD a_35494_6508# 0.106f
C5238 col[4] a_2275_12194# 0.0899f
C5239 ctop a_16018_10162# 4.11f
C5240 row_n[15] a_4974_17190# 0.282f
C5241 a_2475_17214# a_6890_17190# 0.264f
C5242 m2_18224_14426# row_n[12] 0.0128f
C5243 col[9] a_2275_1150# 0.0899f
C5244 a_2275_17214# a_4274_17230# 0.144f
C5245 m2_24248_10410# row_n[8] 0.0128f
C5246 rowoff_n[6] a_15414_8516# 0.0133f
C5247 VDD a_24962_15182# 0.181f
C5248 m2_30272_6394# row_n[4] 0.0128f
C5249 col[30] a_2475_18218# 0.136f
C5250 col_n[11] a_14410_9520# 0.0283f
C5251 m2_1732_2954# m2_1732_1950# 0.843f
C5252 a_9994_5142# a_10298_5182# 0.0931f
C5253 a_10906_5142# a_11398_5504# 0.0658f
C5254 a_2275_5166# a_19030_5142# 0.399f
C5255 row_n[5] a_15014_7150# 0.282f
C5256 m2_4744_946# col[2] 0.425f
C5257 m3_1864_5094# m3_1864_4090# 0.202f
C5258 rowon_n[9] a_14922_11166# 0.118f
C5259 col[24] a_2475_11190# 0.136f
C5260 vcm a_30986_10162# 0.1f
C5261 a_22042_10162# a_23046_10162# 0.843f
C5262 rowoff_n[4] a_24450_6508# 0.0133f
C5263 VDD a_16418_9520# 0.0779f
C5264 row_n[7] a_3878_9158# 0.0437f
C5265 sample a_2161_15206# 0.0858f
C5266 rowon_n[11] a_2966_13174# 0.248f
C5267 ctop a_31078_14178# 4.11f
C5268 VDD a_5886_18194# 0.343f
C5269 col_n[31] a_2275_17214# 0.113f
C5270 a_2275_2154# a_9294_2170# 0.144f
C5271 a_6890_2130# a_6982_2130# 0.326f
C5272 a_2475_2154# a_11910_2130# 0.264f
C5273 a_2275_7174# a_34090_7150# 0.399f
C5274 rowon_n[14] rowoff_n[14] 20.2f
C5275 rowoff_n[9] a_16018_11166# 0.294f
C5276 rowoff_n[2] a_33486_4500# 0.0133f
C5277 col_n[9] a_12002_9158# 0.251f
C5278 m2_34864_16006# vcm 0.395f
C5279 vcm a_11910_13174# 0.1f
C5280 a_13006_12170# a_13006_11166# 0.843f
C5281 VDD a_7986_3134# 0.483f
C5282 col_n[16] a_18938_11166# 0.0765f
C5283 m2_4744_18014# a_2275_18218# 0.28f
C5284 a_2275_16210# a_12914_16186# 0.136f
C5285 col[21] a_2275_14202# 0.0899f
C5286 a_6890_16186# a_7286_16226# 0.0313f
C5287 VDD a_31478_13536# 0.0779f
C5288 rowon_n[3] a_2475_5166# 0.31f
C5289 col[26] a_2275_3158# 0.0899f
C5290 ctop a_12002_17190# 4.06f
C5291 row_n[8] a_34394_10202# 0.0117f
C5292 rowoff_n[7] a_25054_9158# 0.294f
C5293 rowon_n[12] a_35094_14178# 0.0141f
C5294 a_2475_4162# a_26970_4138# 0.264f
C5295 a_2275_4162# a_24354_4178# 0.144f
C5296 m3_24956_1078# ctop 0.21f
C5297 vcm a_2966_7150# 0.56f
C5298 a_25966_9158# a_26458_9520# 0.0658f
C5299 rowoff_n[13] a_32082_15182# 0.294f
C5300 a_25054_9158# a_25358_9198# 0.0931f
C5301 vcm a_26970_17190# 0.1f
C5302 a_2475_13198# a_4974_13174# 0.316f
C5303 VDD a_23046_7150# 0.483f
C5304 col[29] a_32082_8154# 0.367f
C5305 rowoff_n[5] a_34090_7150# 0.294f
C5306 a_2275_18218# a_27974_18194# 0.136f
C5307 VDD a_12402_16548# 0.0779f
C5308 row_n[12] a_13006_14178# 0.282f
C5309 a_2275_1150# a_17934_1126# 0.138f
C5310 col_n[25] col[26] 7.03f
C5311 row_n[3] ctop 0.186f
C5312 row_n[13] col[14] 0.0342f
C5313 row_n[7] col[2] 0.0342f
C5314 row_n[12] col[12] 0.0342f
C5315 rowon_n[14] col[17] 0.0323f
C5316 row_n[9] col[6] 0.0342f
C5317 rowon_n[11] col[11] 0.0323f
C5318 row_n[11] col[10] 0.0342f
C5319 row_n[15] col[18] 0.0342f
C5320 rowon_n[7] col[3] 0.0323f
C5321 rowon_n[12] col[13] 0.0323f
C5322 rowon_n[15] col[19] 0.0323f
C5323 row_n[14] col[16] 0.0342f
C5324 row_n[10] col[8] 0.0342f
C5325 row_n[8] col[4] 0.0342f
C5326 rowon_n[8] col[5] 0.0323f
C5327 rowon_n[13] col[15] 0.0323f
C5328 col_n[11] a_2475_10186# 0.0531f
C5329 col_n[18] rowoff_n[15] 0.0471f
C5330 rowon_n[6] col[1] 0.0323f
C5331 rowon_n[10] col[9] 0.0323f
C5332 rowon_n[9] col[7] 0.0323f
C5333 row_n[6] col[0] 0.0322f
C5334 vcm a_29070_2130# 0.56f
C5335 a_21950_6146# a_22042_6146# 0.326f
C5336 row_n[2] a_23046_4138# 0.282f
C5337 col[21] rowoff_n[11] 0.0901f
C5338 VDD a_13310_1166# 0.0149f
C5339 rowon_n[6] a_22954_8154# 0.118f
C5340 col_n[24] a_27366_8194# 0.084f
C5341 a_28066_16186# a_28066_15182# 0.843f
C5342 a_2475_15206# a_20034_15182# 0.316f
C5343 VDD a_3970_10162# 0.483f
C5344 col_n[5] a_7894_9158# 0.0765f
C5345 col[1] a_2475_7174# 0.136f
C5346 row_n[4] a_10298_6186# 0.0117f
C5347 a_2275_3158# a_32994_3134# 0.136f
C5348 a_16930_3134# a_17326_3174# 0.0313f
C5349 a_2475_18218# a_25966_18194# 0.264f
C5350 m2_13780_18014# col_n[11] 0.243f
C5351 vcm a_9994_5142# 0.56f
C5352 rowoff_n[10] a_3970_12170# 0.294f
C5353 m2_1732_6970# sample 0.2f
C5354 a_2275_12194# a_10998_12170# 0.399f
C5355 col_n[8] a_2275_13198# 0.113f
C5356 a_5978_12170# a_6282_12210# 0.0931f
C5357 a_6890_12170# a_7382_12532# 0.0658f
C5358 col_n[13] a_2275_2154# 0.113f
C5359 m2_17796_18014# VDD 1f
C5360 row_n[15] a_33998_17190# 0.0437f
C5361 a_2475_17214# a_35094_17190# 0.0299f
C5362 a_18026_17190# a_19030_17190# 0.843f
C5363 VDD a_19030_14178# 0.483f
C5364 col[18] a_21038_6146# 0.367f
C5365 a_34090_2130# m2_34288_2378# 0.165f
C5366 rowon_n[0] a_9994_2130# 0.248f
C5367 col[25] a_27974_8154# 0.0682f
C5368 col_n[28] a_2475_12194# 0.0531f
C5369 col[5] rowoff_n[12] 0.0901f
C5370 col_n[0] a_3270_2170# 0.084f
C5371 vcm a_25054_9158# 0.56f
C5372 rowoff_n[14] a_20034_16186# 0.294f
C5373 m2_22816_946# a_22954_1126# 0.225f
C5374 m3_26964_1078# a_27062_2130# 0.0302f
C5375 m2_2160_17438# rowon_n[15] 0.0219f
C5376 a_2275_14202# a_26058_14178# 0.399f
C5377 m2_8184_13422# rowon_n[11] 0.0322f
C5378 m2_14208_9406# rowon_n[7] 0.0322f
C5379 m2_20232_5390# rowon_n[3] 0.0322f
C5380 col_n[13] a_16322_6186# 0.084f
C5381 m2_15788_946# vcm 0.353f
C5382 col_n[23] a_26362_18234# 0.084f
C5383 VDD a_34090_18194# 0.0356f
C5384 col[18] a_2475_9182# 0.136f
C5385 a_3970_2130# a_3970_1126# 0.843f
C5386 vcm a_15318_3174# 0.155f
C5387 row_n[9] a_21038_11166# 0.282f
C5388 a_31990_7150# a_32386_7190# 0.0313f
C5389 rowon_n[13] a_20946_15182# 0.118f
C5390 vcm a_5978_12170# 0.56f
C5391 a_2475_11190# a_18938_11166# 0.264f
C5392 a_2275_11190# a_16322_11206# 0.144f
C5393 VDD a_2161_2154# 0.187f
C5394 col_n[25] a_2275_15206# 0.113f
C5395 a_21950_16186# a_22442_16548# 0.0658f
C5396 row_n[11] a_8290_13214# 0.0117f
C5397 a_21038_16186# a_21342_16226# 0.0931f
C5398 col_n[30] a_2275_4162# 0.113f
C5399 rowon_n[3] a_30986_5142# 0.118f
C5400 m2_13780_18014# m3_14916_18146# 0.0341f
C5401 m2_34864_13998# rowon_n[12] 0.231f
C5402 a_28066_4138# a_29070_4138# 0.843f
C5403 col[7] a_9994_4138# 0.367f
C5404 row_n[1] a_18330_3174# 0.0117f
C5405 col[17] a_20034_16186# 0.367f
C5406 vcm a_30378_7190# 0.155f
C5407 col[14] a_16930_6146# 0.0682f
C5408 a_2275_8178# a_9902_8154# 0.136f
C5409 rowoff_n[12] a_26458_14540# 0.0133f
C5410 col[15] a_2275_12194# 0.0899f
C5411 col[24] a_26970_18194# 0.0682f
C5412 col[20] a_2275_1150# 0.0899f
C5413 vcm a_21038_16186# 0.56f
C5414 a_2475_13198# a_33998_13174# 0.264f
C5415 a_2275_13198# a_31382_13214# 0.144f
C5416 a_17934_13174# a_18026_13174# 0.326f
C5417 VDD a_17934_6146# 0.181f
C5418 row_n[3] a_8898_5142# 0.0437f
C5419 rowon_n[7] a_7986_9158# 0.248f
C5420 col_n[29] a_31990_2130# 0.0765f
C5421 col_n[2] a_5278_4178# 0.084f
C5422 vcm a_23958_1126# 0.0989f
C5423 col_n[12] a_15318_16226# 0.084f
C5424 a_19030_6146# a_19030_5142# 0.843f
C5425 m3_24956_18146# m3_25960_18146# 0.202f
C5426 m2_16792_946# m3_16924_1078# 3.79f
C5427 vcm a_11302_10202# 0.155f
C5428 a_2275_10186# a_24962_10162# 0.136f
C5429 rowoff_n[15] a_7986_17190# 0.294f
C5430 a_12914_10162# a_13310_10202# 0.0313f
C5431 m2_11196_16434# a_10998_16186# 0.165f
C5432 rowoff_n[4] a_6890_6146# 0.202f
C5433 ctop a_24050_5142# 4.11f
C5434 m2_13780_946# a_14010_2130# 0.843f
C5435 VDD a_32994_10162# 0.181f
C5436 col_n[23] a_26458_10524# 0.0283f
C5437 col_n[5] a_2475_8178# 0.0531f
C5438 a_31990_3134# a_32482_3496# 0.0658f
C5439 a_31078_3134# a_31382_3174# 0.0931f
C5440 vcm a_4882_4138# 0.1f
C5441 a_8990_7150# a_9994_7150# 0.843f
C5442 rowoff_n[10] a_32994_12170# 0.202f
C5443 rowoff_n[2] a_15926_4138# 0.202f
C5444 a_2475_7174# a_17022_7150# 0.316f
C5445 m2_30272_12418# a_30074_12170# 0.165f
C5446 row_n[6] a_29070_8154# 0.282f
C5447 vcm a_26362_14218# 0.155f
C5448 col[6] a_8990_14178# 0.367f
C5449 VDD a_24450_4500# 0.0779f
C5450 col[3] a_5886_4138# 0.0682f
C5451 rowon_n[10] a_28978_12170# 0.118f
C5452 col[13] a_15926_16186# 0.0682f
C5453 ctop a_4974_8154# 4.11f
C5454 a_32994_17190# a_33086_17190# 0.326f
C5455 VDD a_13918_13174# 0.181f
C5456 col_n[21] a_24050_10162# 0.251f
C5457 row_n[8] a_16322_10202# 0.0117f
C5458 rowoff_n[7] a_7382_9520# 0.0133f
C5459 rowoff_n[0] a_24962_2130# 0.202f
C5460 a_2275_4162# a_7986_4138# 0.399f
C5461 col_n[28] a_30986_12170# 0.0765f
C5462 col_n[2] a_2275_11190# 0.113f
C5463 m3_20940_18146# ctop 0.209f
C5464 m2_1732_16006# row_n[14] 0.292f
C5465 vcm a_19942_8154# 0.1f
C5466 m2_7180_12418# row_n[10] 0.0128f
C5467 col_n[1] a_4274_14218# 0.084f
C5468 a_2475_9182# a_32082_9158# 0.316f
C5469 m2_13204_8402# row_n[6] 0.0128f
C5470 a_34090_10162# a_34090_9158# 0.843f
C5471 rowoff_n[13] a_14410_15544# 0.0133f
C5472 m2_19228_4386# row_n[2] 0.0128f
C5473 m2_1732_13998# a_1957_14202# 0.245f
C5474 sample a_1957_4162# 0.345f
C5475 row_n[10] a_6890_12170# 0.0437f
C5476 vcm a_7286_17230# 0.155f
C5477 a_27974_14178# a_28370_14218# 0.0313f
C5478 rowon_n[14] a_5978_16186# 0.248f
C5479 VDD a_5374_7512# 0.0779f
C5480 rowoff_n[5] a_16418_7512# 0.0133f
C5481 ctop a_20034_12170# 4.11f
C5482 rowon_n[13] col[26] 0.0323f
C5483 rowon_n[4] col[8] 0.0323f
C5484 row_n[5] col[9] 0.0342f
C5485 rowon_n[1] col[2] 0.0323f
C5486 row_n[6] col[11] 0.0342f
C5487 col_n[22] a_2475_10186# 0.0531f
C5488 rowon_n[14] col[28] 0.0323f
C5489 row_n[2] col[3] 0.0342f
C5490 row_n[4] col[7] 0.0342f
C5491 row_n[10] col[19] 0.0342f
C5492 rowon_n[10] col[20] 0.0323f
C5493 row_n[15] col[29] 0.0342f
C5494 rowon_n[12] col[24] 0.0323f
C5495 rowon_n[7] col[14] 0.0323f
C5496 row_n[13] col[25] 0.0342f
C5497 col_n[29] rowoff_n[15] 0.0471f
C5498 rowon_n[9] col[18] 0.0323f
C5499 rowon_n[5] col[10] 0.0323f
C5500 row_n[8] col[15] 0.0342f
C5501 rowon_n[8] col[16] 0.0323f
C5502 row_n[11] col[21] 0.0342f
C5503 row_n[9] col[17] 0.0342f
C5504 rowon_n[6] col[12] 0.0323f
C5505 row_n[3] col[5] 0.0342f
C5506 rowon_n[3] col[6] 0.0323f
C5507 row_n[14] col[27] 0.0342f
C5508 row_n[1] col[1] 0.0342f
C5509 rowon_n[11] col[22] 0.0323f
C5510 row_n[12] col[23] 0.0342f
C5511 rowon_n[0] col[0] 0.0318f
C5512 col_n[31] col[31] 0.665f
C5513 rowon_n[15] col[30] 0.0323f
C5514 rowon_n[2] col[4] 0.0323f
C5515 row_n[7] col[13] 0.0342f
C5516 a_2275_18218# a_8290_18234# 0.145f
C5517 row_n[0] a_16930_2130# 0.0437f
C5518 VDD a_28978_17190# 0.181f
C5519 col_n[12] a_15414_8516# 0.0283f
C5520 rowon_n[4] a_16018_6146# 0.248f
C5521 sample_n rowoff_n[11] 0.14f
C5522 a_2275_6170# a_23046_6146# 0.399f
C5523 a_12914_6146# a_13406_6508# 0.0658f
C5524 a_12002_6146# a_12306_6186# 0.0931f
C5525 m2_21236_10410# a_21038_10162# 0.165f
C5526 rowoff_n[3] a_25454_5504# 0.0133f
C5527 vcm a_35002_12170# 0.101f
C5528 a_24050_11166# a_25054_11166# 0.843f
C5529 m2_28264_17438# row_n[15] 0.0128f
C5530 VDD a_31078_2130# 0.483f
C5531 m2_34288_13422# row_n[11] 0.0128f
C5532 col[12] a_2475_7174# 0.136f
C5533 col_n[0] a_3366_14540# 0.0283f
C5534 a_2475_15206# a_1957_15206# 0.0734f
C5535 VDD a_20434_11528# 0.0779f
C5536 col[2] a_4882_14178# 0.0682f
C5537 a_2275_3158# a_13310_3174# 0.144f
C5538 a_8898_3134# a_8990_3134# 0.326f
C5539 a_2475_3158# a_15926_3134# 0.264f
C5540 rowoff_n[1] a_34490_3496# 0.0133f
C5541 rowoff_n[8] a_17022_10162# 0.294f
C5542 col_n[10] a_13006_8154# 0.251f
C5543 a_29070_1126# a_2475_1150# 0.0299f
C5544 row_n[13] a_27062_15182# 0.282f
C5545 col_n[19] a_2275_13198# 0.113f
C5546 rowoff_n[11] a_20946_13174# 0.202f
C5547 col_n[17] a_19942_10162# 0.0765f
C5548 col_n[24] a_2275_2154# 0.113f
C5549 vcm a_15926_15182# 0.1f
C5550 a_15014_13174# a_15014_12170# 0.843f
C5551 VDD a_12002_5142# 0.483f
C5552 a_25966_1126# VDD 0.405f
C5553 row_n[15] a_14314_17230# 0.0117f
C5554 a_2275_17214# a_16930_17190# 0.136f
C5555 a_8898_17190# a_9294_17230# 0.0313f
C5556 rowoff_n[6] a_26058_8154# 0.294f
C5557 VDD a_35494_15544# 0.106f
C5558 col[16] rowoff_n[12] 0.0901f
C5559 col[9] a_2275_10186# 0.0899f
C5560 a_2275_5166# a_28370_5182# 0.144f
C5561 a_2475_5166# a_30986_5142# 0.264f
C5562 row_n[5] a_24354_7190# 0.0117f
C5563 col_n[1] a_4370_6508# 0.0283f
C5564 m3_14916_1078# m3_15920_1078# 0.202f
C5565 m2_12200_8402# a_12002_8154# 0.165f
C5566 col_n[11] a_14410_18556# 0.0283f
C5567 a_29982_1126# a_30074_1126# 0.0991f
C5568 rowoff_n[14] a_1957_16210# 0.0219f
C5569 a_27974_10162# a_28466_10524# 0.0658f
C5570 a_27062_10162# a_27366_10202# 0.0931f
C5571 col[30] a_33086_7150# 0.367f
C5572 rowoff_n[4] a_35094_6146# 0.0135f
C5573 a_4974_14178# a_5978_14178# 0.843f
C5574 m2_26832_946# a_2275_1150# 0.28f
C5575 a_2475_14202# a_8990_14178# 0.316f
C5576 col[29] a_2475_9182# 0.136f
C5577 VDD a_27062_9158# 0.483f
C5578 row_n[7] a_14922_9158# 0.0437f
C5579 m2_1732_7974# rowoff_n[6] 0.415f
C5580 rowon_n[11] a_14010_13174# 0.248f
C5581 VDD a_16418_18556# 0.0858f
C5582 a_2275_2154# a_21950_2130# 0.136f
C5583 m2_31276_4386# a_31078_4138# 0.165f
C5584 m2_21236_1374# VDD 0.0193f
C5585 vcm a_33086_4138# 0.56f
C5586 row_n[9] a_2966_11166# 0.281f
C5587 a_23958_7150# a_24050_7150# 0.326f
C5588 rowon_n[1] a_24050_3134# 0.248f
C5589 rowon_n[13] a_2275_15206# 1.79f
C5590 col_n[0] a_2475_6170# 0.0532f
C5591 col_n[25] a_28370_7190# 0.084f
C5592 m2_10768_18014# a_10906_18194# 0.225f
C5593 col_n[6] a_8898_8154# 0.0765f
C5594 a_2475_16210# a_24050_16186# 0.316f
C5595 a_30074_17190# a_30074_16186# 0.843f
C5596 VDD a_7986_12170# 0.483f
C5597 col[0] rowoff_n[13] 0.0901f
C5598 a_32994_1126# col_n[30] 0.0784f
C5599 a_18938_4138# a_19334_4178# 0.0313f
C5600 col[26] a_2275_12194# 0.0899f
C5601 row_n[1] a_2475_3158# 0.405f
C5602 col[31] a_2275_1150# 0.0508f
C5603 vcm a_14010_7150# 0.56f
C5604 rowoff_n[12] a_8898_14178# 0.202f
C5605 row_n[10] a_35094_12170# 0.0123f
C5606 vcm a_2966_16186# 0.56f
C5607 a_2275_13198# a_15014_13174# 0.399f
C5608 rowon_n[14] a_35002_16186# 0.118f
C5609 a_8898_13174# a_9390_13536# 0.0658f
C5610 a_7986_13174# a_8290_13214# 0.0931f
C5611 col[19] a_22042_5142# 0.367f
C5612 VDD a_23046_16186# 0.483f
C5613 col[29] a_32082_17190# 0.367f
C5614 col[26] a_28978_7150# 0.0682f
C5615 row_n[12] a_22346_14218# 0.0117f
C5616 vcm a_4274_1166# 0.155f
C5617 m2_3164_7398# rowon_n[5] 0.0322f
C5618 m2_9188_3382# rowon_n[1] 0.0322f
C5619 row_n[2] a_32386_4178# 0.0117f
C5620 vcm a_29070_11166# 0.56f
C5621 a_2275_10186# a_5278_10202# 0.144f
C5622 a_3878_10162# a_4274_10202# 0.0313f
C5623 a_4882_10162# a_4974_10162# 0.326f
C5624 a_2475_10186# a_7894_10162# 0.264f
C5625 col_n[16] a_2475_8178# 0.0531f
C5626 row_n[14] a_12914_16186# 0.0437f
C5627 col_n[14] a_17326_5182# 0.084f
C5628 a_2275_15206# a_30074_15182# 0.399f
C5629 col_n[24] a_27366_17230# 0.084f
C5630 row_n[4] a_22954_6146# 0.0437f
C5631 col_n[5] a_7894_18194# 0.0762f
C5632 a_5978_3134# a_5978_2130# 0.843f
C5633 rowon_n[8] a_22042_10162# 0.248f
C5634 col[1] a_2475_16210# 0.136f
C5635 vcm a_19334_5182# 0.155f
C5636 col[6] a_2475_5166# 0.136f
C5637 m2_18224_16434# rowon_n[14] 0.0322f
C5638 m2_24248_12418# rowon_n[10] 0.0322f
C5639 vcm a_9994_14178# 0.56f
C5640 m2_30272_8402# rowon_n[6] 0.0322f
C5641 a_2275_12194# a_20338_12210# 0.144f
C5642 m2_35292_4386# rowon_n[2] 0.0322f
C5643 a_2475_12194# a_22954_12170# 0.264f
C5644 VDD a_6890_4138# 0.181f
C5645 m2_30848_946# col_n[28] 0.349f
C5646 a_23958_17190# a_24450_17552# 0.0658f
C5647 a_23046_17190# a_23350_17230# 0.0931f
C5648 col_n[13] a_2275_11190# 0.113f
C5649 m2_32856_946# col[31] 0.0132f
C5650 col[8] a_10998_3134# 0.367f
C5651 m2_28840_18014# col[26] 0.347f
C5652 col[18] a_21038_15182# 0.367f
C5653 a_30074_5142# a_31078_5142# 0.843f
C5654 col[15] a_17934_5142# 0.0682f
C5655 col[25] a_27974_17190# 0.0682f
C5656 m2_18800_18014# m2_19804_18014# 0.843f
C5657 vcm a_35398_9198# 0.161f
C5658 a_2275_9182# a_13918_9158# 0.136f
C5659 rowon_n[2] a_9902_4138# 0.118f
C5660 col_n[0] a_3270_11206# 0.084f
C5661 row_n[8] col[26] 0.0342f
C5662 rowon_n[3] col[17] 0.0323f
C5663 rowon_n[0] col[11] 0.0323f
C5664 row_n[2] col[14] 0.0342f
C5665 ctop col[7] 0.123f
C5666 rowon_n[6] col[23] 0.0323f
C5667 rowon_n[7] col[25] 0.0323f
C5668 rowon_n[9] col[29] 0.0323f
C5669 ctop a_13006_3134# 4.11f
C5670 rowon_n[10] col[31] 0.0323f
C5671 col[0] col[1] 0.0354f
C5672 row_n[5] col[20] 0.0342f
C5673 row_n[11] sample_n 0.0596f
C5674 row_n[1] col[12] 0.0342f
C5675 row_n[3] col[16] 0.0342f
C5676 row_n[6] col[22] 0.0342f
C5677 vcm a_25054_18194# 0.165f
C5678 row_n[0] col[10] 0.0342f
C5679 row_n[10] col[30] 0.0342f
C5680 rowon_n[4] col[19] 0.0323f
C5681 row_n[4] col[18] 0.0342f
C5682 row_n[7] col[24] 0.0342f
C5683 rowon_n[8] col[27] 0.0323f
C5684 rowon_n[5] col[21] 0.0323f
C5685 rowon_n[2] col[15] 0.0323f
C5686 row_n[9] col[28] 0.0342f
C5687 rowon_n[1] col[13] 0.0323f
C5688 a_19942_14178# a_20034_14178# 0.326f
C5689 a_2275_14202# a_2275_13198# 0.0715f
C5690 col[3] a_2275_8178# 0.0899f
C5691 VDD a_21950_8154# 0.181f
C5692 col_n[3] a_6282_3174# 0.084f
C5693 col_n[13] a_16322_15222# 0.084f
C5694 m3_19936_1078# VDD 0.0122f
C5695 row_n[9] a_30378_11206# 0.0117f
C5696 m2_34864_7974# m2_35292_8402# 0.165f
C5697 vcm a_27974_3134# 0.1f
C5698 a_2966_6146# a_3270_6186# 0.0931f
C5699 a_3878_6146# a_4370_6508# 0.0658f
C5700 a_21038_7150# a_21038_6146# 0.843f
C5701 a_2475_6170# a_5978_6146# 0.316f
C5702 col[23] a_2475_7174# 0.136f
C5703 rowoff_n[3] a_7894_5142# 0.202f
C5704 vcm a_15318_12210# 0.155f
C5705 a_2275_11190# a_28978_11166# 0.136f
C5706 a_14922_11166# a_15318_11206# 0.0313f
C5707 VDD a_13406_2492# 0.0779f
C5708 m2_6752_18014# a_6982_17190# 0.843f
C5709 m2_29844_18014# a_29982_18194# 0.225f
C5710 col_n[24] a_27462_9520# 0.0283f
C5711 ctop a_28066_7150# 4.11f
C5712 row_n[11] a_20946_13174# 0.0437f
C5713 VDD a_2161_11190# 0.187f
C5714 m2_28840_18014# m3_27968_18146# 0.0341f
C5715 rowon_n[15] a_20034_17190# 0.248f
C5716 col_n[30] a_2275_13198# 0.113f
C5717 a_33998_4138# a_34490_4500# 0.0658f
C5718 a_33086_4138# a_33390_4178# 0.0931f
C5719 row_n[1] a_30986_3134# 0.0437f
C5720 rowoff_n[1] a_16930_3134# 0.202f
C5721 rowon_n[5] a_30074_7150# 0.248f
C5722 vcm a_8898_6146# 0.1f
C5723 a_10998_8154# a_12002_8154# 0.843f
C5724 a_2475_8178# a_21038_8154# 0.316f
C5725 rowoff_n[11] a_2275_13198# 0.151f
C5726 col[7] a_9994_13174# 0.367f
C5727 col[4] a_6890_3134# 0.0682f
C5728 vcm a_30378_16226# 0.155f
C5729 col[14] a_16930_15182# 0.0682f
C5730 m2_1732_3958# ctop 0.0428f
C5731 VDD a_28466_6508# 0.0779f
C5732 col[27] rowoff_n[12] 0.0901f
C5733 ctop a_8990_10162# 4.11f
C5734 col[20] a_2275_10186# 0.0899f
C5735 col_n[22] a_25054_9158# 0.251f
C5736 a_35002_18194# a_35094_18194# 0.0991f
C5737 VDD a_17934_15182# 0.181f
C5738 rowoff_n[6] a_8386_8516# 0.0133f
C5739 m2_2160_6394# row_n[4] 0.0194f
C5740 m2_7180_2378# row_n[0] 0.0128f
C5741 col_n[29] a_31990_11166# 0.0765f
C5742 m3_9896_18146# a_9994_17190# 0.0303f
C5743 row_n[5] a_7986_7150# 0.282f
C5744 a_2275_5166# a_12002_5142# 0.399f
C5745 col_n[2] a_5278_13214# 0.084f
C5746 m3_1864_12122# m3_1864_11118# 0.202f
C5747 m2_31852_946# m3_32988_1078# 0.0341f
C5748 col_n[0] a_2966_3134# 0.251f
C5749 rowon_n[9] a_7894_11166# 0.118f
C5750 vcm a_23958_10162# 0.1f
C5751 a_2475_10186# a_2475_9182# 0.0666f
C5752 rowoff_n[4] a_17422_6508# 0.0133f
C5753 a_29982_15182# a_30378_15222# 0.0313f
C5754 m2_27836_18014# ctop 0.0422f
C5755 VDD a_9390_9520# 0.0779f
C5756 col_n[13] a_16418_7512# 0.0283f
C5757 ctop a_24050_14178# 4.11f
C5758 col_n[5] a_2475_17214# 0.0531f
C5759 a_2275_2154# a_3878_2130# 0.136f
C5760 a_2475_2154# a_4882_2130# 0.264f
C5761 a_2874_2130# a_3366_2492# 0.0658f
C5762 m2_17220_15430# row_n[13] 0.0128f
C5763 m2_23244_11414# row_n[9] 0.0128f
C5764 col_n[10] a_2475_6170# 0.0531f
C5765 m2_29268_7398# row_n[5] 0.0128f
C5766 m2_34864_2954# row_n[1] 0.267f
C5767 a_14010_7150# a_14314_7190# 0.0931f
C5768 rowoff_n[2] a_26458_4500# 0.0133f
C5769 a_2275_7174# a_27062_7150# 0.399f
C5770 a_14922_7150# a_15414_7512# 0.0658f
C5771 rowoff_n[9] a_8990_11166# 0.294f
C5772 vcm a_4882_13174# 0.1f
C5773 a_26058_12170# a_27062_12170# 0.843f
C5774 col[11] rowoff_n[13] 0.0901f
C5775 a_2275_16210# a_5886_16186# 0.136f
C5776 col[3] a_5886_13174# 0.0682f
C5777 VDD a_24450_13536# 0.0779f
C5778 col[0] a_2475_3158# 0.148f
C5779 ctop a_4974_17190# 4.06f
C5780 row_n[8] a_28978_10162# 0.0437f
C5781 rowoff_n[0] a_35494_2492# 0.0133f
C5782 rowoff_n[7] a_18026_9158# 0.294f
C5783 col_n[11] a_14010_7150# 0.251f
C5784 rowon_n[12] a_28066_14178# 0.248f
C5785 a_2275_4162# a_17326_4178# 0.144f
C5786 a_10906_4138# a_10998_4138# 0.326f
C5787 a_2475_4162# a_19942_4138# 0.264f
C5788 m3_1864_3086# ctop 0.21f
C5789 col_n[18] a_20946_9158# 0.0765f
C5790 rowoff_n[13] a_25054_15182# 0.294f
C5791 col_n[7] a_2275_9182# 0.113f
C5792 vcm a_19942_17190# 0.1f
C5793 a_17022_14178# a_17022_13174# 0.843f
C5794 VDD a_16018_7150# 0.483f
C5795 sample a_1957_13198# 0.345f
C5796 m2_2736_1950# m3_2868_1078# 0.0341f
C5797 rowoff_n[5] a_27062_7150# 0.294f
C5798 a_10906_18194# a_11302_18234# 0.0313f
C5799 a_2275_18218# a_20946_18194# 0.136f
C5800 VDD a_5374_16548# 0.0779f
C5801 a_2275_1150# a_10906_1126# 0.136f
C5802 a_5886_1126# a_6282_1166# 0.0313f
C5803 row_n[12] a_5978_14178# 0.282f
C5804 col_n[2] a_5374_5504# 0.0283f
C5805 vcm a_22042_2130# 0.56f
C5806 col_n[12] a_15414_17552# 0.0283f
C5807 a_2275_6170# a_32386_6186# 0.144f
C5808 a_2475_6170# a_35002_6146# 0.264f
C5809 col_n[27] a_2475_8178# 0.0531f
C5810 col[31] a_34090_6146# 0.367f
C5811 row_n[2] a_16018_4138# 0.282f
C5812 a_29982_11166# a_30474_11528# 0.0658f
C5813 a_29070_11166# a_29374_11206# 0.0931f
C5814 VDD a_6282_1166# 0.0149f
C5815 rowon_n[6] a_15926_8154# 0.118f
C5816 m2_25828_18014# a_26058_17190# 0.843f
C5817 m2_17220_17438# a_17022_17190# 0.165f
C5818 a_2475_15206# a_13006_15182# 0.316f
C5819 a_6982_15182# a_7986_15182# 0.843f
C5820 VDD a_31078_11166# 0.483f
C5821 col[12] a_2475_16210# 0.136f
C5822 row_n[4] a_3270_6186# 0.0117f
C5823 col[17] a_2475_5166# 0.136f
C5824 a_2275_3158# a_25966_3134# 0.136f
C5825 a_2475_18218# a_18938_18194# 0.264f
C5826 col_n[26] a_29374_6186# 0.084f
C5827 vcm a_2874_5142# 0.1f
C5828 rowoff_n[11] a_31478_13536# 0.0133f
C5829 a_25966_8154# a_26058_8154# 0.326f
C5830 col_n[10] a_13006_17190# 0.251f
C5831 col_n[7] a_9902_7150# 0.0765f
C5832 a_2275_12194# a_3970_12170# 0.399f
C5833 col_n[24] a_2275_11190# 0.113f
C5834 m2_3740_18014# VDD 1.07f
C5835 row_n[15] a_26970_17190# 0.0437f
C5836 a_2475_17214# a_28066_17190# 0.316f
C5837 VDD a_12002_14178# 0.483f
C5838 rowon_n[0] a_2874_2130# 0.118f
C5839 a_20946_5142# a_21342_5182# 0.0313f
C5840 m2_1732_1950# sample_n 0.0522f
C5841 row_n[0] col[21] 0.0342f
C5842 rowon_n[3] col[28] 0.0323f
C5843 row_n[1] col[23] 0.0342f
C5844 rowon_n[4] col[30] 0.0323f
C5845 rowon_n[2] col[26] 0.0323f
C5846 rowon_n[0] col[22] 0.0323f
C5847 row_n[2] col[25] 0.0342f
C5848 row_n[5] col[31] 0.0342f
C5849 rowon_n[1] col[24] 0.0323f
C5850 ctop col[18] 0.123f
C5851 rowon_n[5] sample_n 0.0692f
C5852 row_n[3] col[27] 0.0342f
C5853 row_n[4] col[29] 0.0342f
C5854 vcm a_18026_9158# 0.56f
C5855 rowoff_n[14] a_13006_16186# 0.294f
C5856 col[14] a_2275_8178# 0.0899f
C5857 col_n[1] a_4370_15544# 0.0283f
C5858 m2_8184_15430# a_7986_15182# 0.165f
C5859 col[20] a_23046_4138# 0.367f
C5860 a_10906_14178# a_11398_14540# 0.0658f
C5861 a_9994_14178# a_10298_14218# 0.0931f
C5862 a_2275_14202# a_19030_14178# 0.399f
C5863 VDD a_3878_8154# 0.181f
C5864 col[30] a_33086_16186# 0.367f
C5865 col[27] a_29982_6146# 0.0682f
C5866 VDD a_27062_18194# 0.0356f
C5867 a_2475_2154# a_33086_2130# 0.316f
C5868 a_17022_2130# a_18026_2130# 0.843f
C5869 m3_15920_18146# VDD 0.0669f
C5870 vcm a_8290_3174# 0.155f
C5871 row_n[9] a_14010_11166# 0.282f
C5872 m2_27260_11414# a_27062_11166# 0.165f
C5873 rowon_n[13] a_13918_15182# 0.118f
C5874 vcm a_33086_13174# 0.56f
C5875 col_n[15] a_18330_4178# 0.084f
C5876 a_2275_11190# a_9294_11206# 0.144f
C5877 a_6890_11166# a_6982_11166# 0.326f
C5878 a_2475_11190# a_11910_11166# 0.264f
C5879 VDD a_29982_3134# 0.181f
C5880 col_n[25] a_28370_16226# 0.084f
C5881 col_n[0] a_2475_15206# 0.0532f
C5882 a_2275_16210# a_34090_16186# 0.399f
C5883 row_n[11] a_2275_13198# 19.2f
C5884 col_n[4] a_2475_4162# 0.0531f
C5885 rowon_n[3] a_23958_5142# 0.118f
C5886 m2_4744_18014# m3_4876_18146# 3.79f
C5887 rowon_n[15] a_1957_17214# 0.0172f
C5888 col_n[6] a_8898_17190# 0.0765f
C5889 m2_7180_14426# rowon_n[12] 0.0322f
C5890 m2_13204_10410# rowon_n[8] 0.0322f
C5891 m3_1864_14130# a_2966_14178# 0.0302f
C5892 m2_19228_6394# rowon_n[4] 0.0322f
C5893 a_7986_4138# a_7986_3134# 0.843f
C5894 row_n[1] a_11302_3174# 0.0117f
C5895 vcm a_23350_7190# 0.155f
C5896 a_2475_8178# a_2966_8154# 0.317f
C5897 a_2161_8178# a_2275_8178# 0.183f
C5898 rowoff_n[12] a_19430_14540# 0.0133f
C5899 col[31] a_2275_10186# 0.0899f
C5900 ctop a_2475_1150# 0.0736f
C5901 vcm a_14010_16186# 0.56f
C5902 a_2475_13198# a_26970_13174# 0.264f
C5903 a_2275_13198# a_24354_13214# 0.144f
C5904 VDD a_10906_6146# 0.181f
C5905 a_25966_18194# a_26458_18556# 0.0658f
C5906 col[9] a_12002_2130# 0.367f
C5907 a_20946_1126# a_21438_1488# 0.0658f
C5908 a_20034_1126# a_20338_1166# 0.0997f
C5909 col[19] a_22042_14178# 0.367f
C5910 row_n[12] a_35002_14178# 0.0437f
C5911 col[16] a_18938_4138# 0.0682f
C5912 vcm a_16930_1126# 0.0989f
C5913 m2_34288_15430# rowon_n[13] 0.0322f
C5914 a_32082_6146# a_33086_6146# 0.843f
C5915 col[26] a_28978_16186# 0.0682f
C5916 col_n[1] a_2275_7174# 0.113f
C5917 m3_10900_18146# m3_11904_18146# 0.202f
C5918 m2_7756_946# m3_6884_1078# 0.0341f
C5919 m2_18224_9406# a_18026_9158# 0.165f
C5920 vcm a_4274_10202# 0.155f
C5921 a_2275_10186# a_17934_10162# 0.136f
C5922 ctop a_17022_5142# 4.11f
C5923 a_21950_15182# a_22042_15182# 0.326f
C5924 col_n[4] a_7286_2170# 0.084f
C5925 VDD a_25966_10162# 0.181f
C5926 col_n[16] a_2475_17214# 0.0531f
C5927 m2_3164_1374# m2_2736_946# 0.165f
C5928 col_n[21] a_2475_6170# 0.0531f
C5929 col_n[14] a_17326_14218# 0.084f
C5930 vcm a_31990_5142# 0.1f
C5931 rowoff_n[2] a_8898_4138# 0.202f
C5932 a_23046_8154# a_23046_7150# 0.843f
C5933 a_2475_7174# a_9994_7150# 0.316f
C5934 rowoff_n[10] a_25966_12170# 0.202f
C5935 col[22] rowoff_n[13] 0.0901f
C5936 row_n[6] a_22042_8154# 0.282f
C5937 col_n[25] a_28466_8516# 0.0283f
C5938 col[6] a_2475_14202# 0.136f
C5939 vcm a_19334_14218# 0.155f
C5940 a_2275_12194# a_32994_12170# 0.136f
C5941 a_16930_12170# a_17326_12210# 0.0313f
C5942 rowon_n[10] a_21950_12170# 0.118f
C5943 VDD a_17422_4500# 0.0779f
C5944 col_n[3] rowoff_n[7] 0.0471f
C5945 vcm rowoff_n[4] 0.533f
C5946 col[11] a_2475_3158# 0.136f
C5947 col_n[0] rowoff_n[3] 0.0471f
C5948 col_n[2] rowoff_n[6] 0.0471f
C5949 sample rowoff_n[2] 0.0775f
C5950 col_n[4] rowoff_n[8] 0.0471f
C5951 col_n[5] rowoff_n[9] 0.0471f
C5952 VDD rowoff_n[1] 1.51f
C5953 col_n[1] rowoff_n[5] 0.0471f
C5954 ctop a_32082_9158# 4.11f
C5955 VDD a_6890_13174# 0.181f
C5956 row_n[8] a_9294_10202# 0.0117f
C5957 rowoff_n[0] a_17934_2130# 0.202f
C5958 rowon_n[0] a_31990_2130# 0.118f
C5959 col[8] a_10998_12170# 0.367f
C5960 m2_9188_7398# a_8990_7150# 0.165f
C5961 col_n[18] a_2275_9182# 0.113f
C5962 col[5] a_7894_2130# 0.0682f
C5963 vcm a_12914_8154# 0.1f
C5964 m2_29844_18014# m2_30272_18442# 0.165f
C5965 a_2475_9182# a_25054_9158# 0.316f
C5966 rowoff_n[13] a_7382_15544# 0.0133f
C5967 a_13006_9158# a_14010_9158# 0.843f
C5968 col[15] a_17934_14178# 0.0682f
C5969 vcm a_35398_18234# 0.161f
C5970 col_n[23] a_26058_8154# 0.251f
C5971 VDD a_32482_8516# 0.0779f
C5972 rowoff_n[5] a_9390_7512# 0.0133f
C5973 ctop a_13006_12170# 4.11f
C5974 row_n[0] a_9902_2130# 0.0437f
C5975 col_n[30] a_32994_10162# 0.0765f
C5976 col[3] a_2275_17214# 0.0899f
C5977 VDD a_21950_17190# 0.181f
C5978 a_31990_2130# a_32082_2130# 0.326f
C5979 col[8] a_2275_6170# 0.0899f
C5980 rowon_n[4] a_8990_6146# 0.248f
C5981 m2_28264_3382# a_28066_3134# 0.165f
C5982 col_n[3] a_6282_12210# 0.084f
C5983 col[6] rowoff_n[14] 0.0901f
C5984 a_2275_6170# a_16018_6146# 0.399f
C5985 rowoff_n[3] a_18426_5504# 0.0133f
C5986 vcm a_27974_12170# 0.1f
C5987 a_3970_11166# a_3970_10162# 0.843f
C5988 VDD a_24050_2130# 0.483f
C5989 m2_6176_13422# row_n[11] 0.0128f
C5990 m2_1732_17010# a_2966_17190# 0.843f
C5991 col[23] a_2475_16210# 0.136f
C5992 m2_12200_9406# row_n[7] 0.0128f
C5993 m2_18224_5390# row_n[3] 0.0128f
C5994 col_n[14] a_17422_6508# 0.0283f
C5995 a_31990_16186# a_32386_16226# 0.0313f
C5996 col[28] a_2475_5166# 0.136f
C5997 VDD a_13406_11528# 0.0779f
C5998 col_n[24] a_27462_18556# 0.0283f
C5999 ctop a_28066_16186# 4.11f
C6000 a_2475_3158# a_8898_3134# 0.264f
C6001 a_2275_3158# a_6282_3174# 0.144f
C6002 rowoff_n[1] a_27462_3496# 0.0133f
C6003 rowoff_n[8] a_9994_10162# 0.294f
C6004 row_n[13] a_20034_15182# 0.282f
C6005 rowoff_n[11] a_13918_13174# 0.202f
C6006 a_16018_8154# a_16322_8194# 0.0931f
C6007 a_16930_8154# a_17422_8516# 0.0658f
C6008 a_2275_8178# a_31078_8154# 0.399f
C6009 vcm a_8898_15182# 0.1f
C6010 a_28066_13174# a_29070_13174# 0.843f
C6011 VDD a_4974_5142# 0.483f
C6012 col[4] a_6890_12170# 0.0682f
C6013 row_n[3] a_30074_5142# 0.282f
C6014 row_n[15] a_7286_17230# 0.0117f
C6015 m2_33284_14426# row_n[12] 0.0128f
C6016 rowon_n[7] a_29982_9158# 0.118f
C6017 a_2275_17214# a_9902_17190# 0.136f
C6018 VDD a_28466_15544# 0.0779f
C6019 rowoff_n[6] a_19030_8154# 0.294f
C6020 col_n[12] a_15014_6146# 0.251f
C6021 VDD col_n[6] 5.17f
C6022 vcm col_n[3] 1.94f
C6023 row_n[0] sample_n 0.061f
C6024 col[11] col[12] 0.0355f
C6025 sw col[31] 0.04f
C6026 ctop col[29] 0.123f
C6027 col_n[19] a_21950_8154# 0.0765f
C6028 col[25] a_2275_8178# 0.0899f
C6029 a_2475_5166# a_23958_5142# 0.264f
C6030 a_12914_5142# a_13006_5142# 0.326f
C6031 row_n[5] a_17326_7190# 0.0117f
C6032 a_2275_5166# a_21342_5182# 0.144f
C6033 m3_2868_2082# m3_2868_1078# 0.202f
C6034 rowoff_n[15] a_29982_17190# 0.202f
C6035 rowoff_n[4] a_28066_6146# 0.294f
C6036 col_n[0] a_2966_12170# 0.251f
C6037 m2_5748_946# a_5886_1126# 0.225f
C6038 m2_12776_946# a_2475_1150# 0.286f
C6039 a_19030_15182# a_19030_14178# 0.843f
C6040 VDD a_20034_9158# 0.483f
C6041 row_n[7] a_7894_9158# 0.0437f
C6042 rowon_n[11] a_6982_13174# 0.248f
C6043 col_n[3] a_6378_4500# 0.0283f
C6044 VDD a_9390_18556# 0.0858f
C6045 a_7894_2130# a_8290_2170# 0.0313f
C6046 col_n[13] a_16418_16548# 0.0283f
C6047 a_2275_2154# a_14922_2130# 0.136f
C6048 m2_5748_946# VDD 1f
C6049 vcm a_26058_4138# 0.56f
C6050 rowon_n[1] a_17022_3134# 0.248f
C6051 a_2966_7150# a_2966_6146# 0.843f
C6052 col_n[10] a_2475_15206# 0.0531f
C6053 a_31990_12170# a_32482_12532# 0.0658f
C6054 a_31078_12170# a_31382_12210# 0.0931f
C6055 col_n[15] a_2475_4162# 0.0531f
C6056 m2_5748_18014# a_5978_18194# 0.0249f
C6057 a_8990_16186# a_9994_16186# 0.843f
C6058 a_2475_16210# a_17022_16186# 0.316f
C6059 a_24354_1166# m2_23820_946# 0.087f
C6060 a_2275_4162# a_29982_4138# 0.136f
C6061 col_n[27] a_30378_5182# 0.084f
C6062 col_n[1] a_3970_4138# 0.251f
C6063 col[0] a_2475_12194# 0.148f
C6064 col_n[11] a_14010_16186# 0.251f
C6065 col[5] a_2475_1150# 0.136f
C6066 vcm a_6982_7150# 0.56f
C6067 col_n[8] a_10906_6146# 0.0765f
C6068 a_27974_9158# a_28066_9158# 0.326f
C6069 row_n[10] a_28066_12170# 0.282f
C6070 col_n[18] a_20946_18194# 0.0762f
C6071 rowon_n[14] a_27974_16186# 0.118f
C6072 a_2275_13198# a_7986_13174# 0.399f
C6073 col_n[7] a_2275_18218# 0.113f
C6074 VDD a_16018_16186# 0.483f
C6075 col_n[12] a_2275_7174# 0.113f
C6076 a_2475_1150# a_22042_1126# 0.0299f
C6077 row_n[12] a_15318_14218# 0.0117f
C6078 vcm a_31382_2170# 0.155f
C6079 a_22954_6146# a_23350_6186# 0.0313f
C6080 col_n[2] a_5374_14540# 0.0283f
C6081 vcm a_22042_11166# 0.56f
C6082 row_n[2] a_25358_4178# 0.0117f
C6083 col[21] a_24050_3134# 0.367f
C6084 col_n[27] a_2475_17214# 0.0531f
C6085 row_n[14] a_5886_16186# 0.0437f
C6086 VDD a_18938_1126# 0.403f
C6087 col[31] a_34090_15182# 0.367f
C6088 col[2] a_2275_4162# 0.0899f
C6089 col[28] a_30986_5142# 0.0682f
C6090 a_2275_15206# a_23046_15182# 0.399f
C6091 a_12002_15182# a_12306_15222# 0.0931f
C6092 a_12914_15182# a_13406_15544# 0.0658f
C6093 row_n[4] a_15926_6146# 0.0437f
C6094 a_19030_3134# a_20034_3134# 0.843f
C6095 rowon_n[8] a_15014_10162# 0.248f
C6096 col[17] a_2475_14202# 0.136f
C6097 vcm a_12306_5182# 0.155f
C6098 col_n[15] rowoff_n[8] 0.0471f
C6099 col_n[16] a_19334_3174# 0.084f
C6100 col_n[8] rowoff_n[1] 0.0471f
C6101 col_n[16] rowoff_n[9] 0.0471f
C6102 col_n[13] rowoff_n[6] 0.0471f
C6103 col_n[10] rowoff_n[3] 0.0471f
C6104 col_n[12] rowoff_n[5] 0.0471f
C6105 col_n[14] rowoff_n[7] 0.0471f
C6106 col_n[11] rowoff_n[4] 0.0471f
C6107 col[22] a_2475_3158# 0.136f
C6108 col_n[7] rowoff_n[0] 0.0471f
C6109 col_n[9] rowoff_n[2] 0.0471f
C6110 col_n[26] a_29374_15222# 0.084f
C6111 vcm a_2874_14178# 0.1f
C6112 m2_2160_8402# rowon_n[6] 0.0219f
C6113 a_2275_12194# a_13310_12210# 0.144f
C6114 m2_8184_4386# rowon_n[2] 0.0322f
C6115 a_2475_12194# a_15926_12170# 0.264f
C6116 a_8898_12170# a_8990_12170# 0.326f
C6117 VDD a_33998_5142# 0.181f
C6118 rowon_n[10] a_3878_12170# 0.118f
C6119 m2_25252_18442# VDD 0.0456f
C6120 col_n[7] a_9902_16186# 0.0765f
C6121 col_n[29] a_2275_9182# 0.113f
C6122 a_9994_5142# a_9994_4138# 0.843f
C6123 vcm a_27366_9198# 0.155f
C6124 m2_11772_18014# m2_12776_18014# 0.843f
C6125 a_2275_9182# a_6890_9158# 0.136f
C6126 rowon_n[2] a_2161_4162# 0.0177f
C6127 ctop a_5978_3134# 4.11f
C6128 vcm a_18026_18194# 0.165f
C6129 m2_17220_17438# rowon_n[15] 0.0322f
C6130 m3_29976_1078# a_30074_2130# 0.0302f
C6131 a_2275_14202# a_28370_14218# 0.144f
C6132 col[14] a_2275_17214# 0.0899f
C6133 a_2475_14202# a_30986_14178# 0.264f
C6134 m2_23244_13422# rowon_n[11] 0.0322f
C6135 VDD a_14922_8154# 0.181f
C6136 m2_29268_9406# rowon_n[7] 0.0322f
C6137 col[19] a_2275_6170# 0.0899f
C6138 m2_34864_4962# rowon_n[3] 0.231f
C6139 col[20] a_23046_13174# 0.367f
C6140 m2_24824_946# vcm 0.353f
C6141 col[17] rowoff_n[14] 0.0901f
C6142 col[17] a_19942_3134# 0.0682f
C6143 VDD a_3878_17190# 0.181f
C6144 a_22954_2130# a_23446_2492# 0.0658f
C6145 a_22042_2130# a_22346_2170# 0.0931f
C6146 col[27] a_29982_15182# 0.0682f
C6147 vcm rowoff_n[10] 0.533f
C6148 vcm a_20946_3134# 0.1f
C6149 row_n[9] a_23350_11206# 0.0117f
C6150 a_33998_7150# a_34394_7190# 0.0313f
C6151 m2_34864_10986# a_35398_11206# 0.087f
C6152 vcm a_8290_12210# 0.155f
C6153 m2_14784_946# col_n[12] 0.331f
C6154 a_2275_11190# a_21950_11166# 0.136f
C6155 VDD a_6378_2492# 0.0779f
C6156 col_n[5] a_8290_1166# 0.0839f
C6157 m2_24824_18014# a_25054_18194# 0.0249f
C6158 ctop a_21038_7150# 4.11f
C6159 a_23958_16186# a_24050_16186# 0.326f
C6160 col_n[15] a_18330_13214# 0.084f
C6161 row_n[11] a_13918_13174# 0.0437f
C6162 VDD a_29982_12170# 0.181f
C6163 m2_18800_18014# m3_19936_18146# 0.0341f
C6164 rowon_n[15] a_13006_17190# 0.248f
C6165 col_n[4] a_2475_13198# 0.0531f
C6166 row_n[1] a_23958_3134# 0.0437f
C6167 rowoff_n[1] a_9902_3134# 0.202f
C6168 col_n[9] a_2475_2154# 0.0531f
C6169 row_n[13] a_1957_15206# 0.187f
C6170 col_n[26] a_29470_7512# 0.0283f
C6171 vcm a_34394_7190# 0.155f
C6172 rowon_n[5] a_23046_7150# 0.248f
C6173 a_2475_8178# a_14010_8154# 0.316f
C6174 a_25054_9158# a_25054_8154# 0.843f
C6175 rowoff_n[12] a_30074_14178# 0.294f
C6176 m2_34864_946# m2_34864_1950# 0.843f
C6177 vcm a_23350_16226# 0.155f
C6178 a_18938_13174# a_19334_13214# 0.0313f
C6179 VDD a_21438_6508# 0.0779f
C6180 VDD col_n[17] 4.83f
C6181 vcm col_n[14] 1.94f
C6182 col[1] rowoff_n[15] 0.0901f
C6183 ctop a_2475_10186# 0.0488f
C6184 m2_7756_18014# col_n[5] 0.243f
C6185 VDD a_10906_15182# 0.181f
C6186 col[9] a_12002_11166# 0.367f
C6187 col[6] a_8898_1126# 0.0682f
C6188 a_2275_5166# a_4974_5142# 0.399f
C6189 a_2874_5142# a_3270_5182# 0.0313f
C6190 a_3878_5142# a_3970_5142# 0.326f
C6191 m2_22816_946# m3_22948_1078# 3.79f
C6192 col[16] a_18938_13174# 0.0682f
C6193 vcm a_16930_10162# 0.1f
C6194 col_n[1] a_2275_16210# 0.113f
C6195 a_2475_10186# a_29070_10162# 0.316f
C6196 a_15014_10162# a_16018_10162# 0.843f
C6197 row_n[14] a_34090_16186# 0.282f
C6198 m2_14208_16434# a_14010_16186# 0.165f
C6199 col_n[24] a_27062_7150# 0.251f
C6200 rowoff_n[4] a_10394_6508# 0.0133f
C6201 col_n[6] a_2275_5166# 0.113f
C6202 m2_13780_18014# ctop 0.0422f
C6203 VDD a_1957_9182# 0.196f
C6204 col_n[31] a_33998_9158# 0.0765f
C6205 ctop a_17022_14178# 4.11f
C6206 col_n[4] a_7286_11206# 0.084f
C6207 a_33998_3134# a_34090_3134# 0.326f
C6208 col[0] a_2966_9158# 0.367f
C6209 col_n[21] a_2475_15206# 0.0531f
C6210 m2_1732_6970# row_n[5] 0.292f
C6211 m2_7180_3382# row_n[1] 0.0128f
C6212 m2_34864_946# col_n[31] 0.308f
C6213 col_n[26] a_2475_4162# 0.0531f
C6214 a_2275_7174# a_20034_7150# 0.399f
C6215 rowoff_n[2] a_19430_4500# 0.0133f
C6216 rowoff_n[9] a_2475_11190# 3.9f
C6217 m2_33284_12418# a_33086_12170# 0.165f
C6218 row_n[6] a_31382_8194# 0.0117f
C6219 vcm a_31990_14178# 0.1f
C6220 col_n[15] a_18426_5504# 0.0283f
C6221 a_5978_12170# a_5978_11166# 0.843f
C6222 VDD a_28066_4138# 0.483f
C6223 col_n[25] a_28466_17552# 0.0283f
C6224 VDD a_17422_13536# 0.0779f
C6225 col[11] a_2475_12194# 0.136f
C6226 row_n[8] a_21950_10162# 0.0437f
C6227 rowoff_n[7] a_10998_9158# 0.294f
C6228 col[16] a_2475_1150# 0.136f
C6229 rowoff_n[0] a_28466_2492# 0.0133f
C6230 rowon_n[12] a_21038_14178# 0.248f
C6231 a_2475_4162# a_12914_4138# 0.264f
C6232 a_2275_4162# a_10298_4178# 0.144f
C6233 m3_1864_17142# ctop 0.21f
C6234 col_n[0] a_2874_1126# 0.0765f
C6235 m2_16216_16434# row_n[14] 0.0128f
C6236 m2_22240_12418# row_n[10] 0.0128f
C6237 m2_28264_8402# row_n[6] 0.0128f
C6238 a_18938_9158# a_19430_9520# 0.0658f
C6239 a_18026_9158# a_18330_9198# 0.0931f
C6240 a_2275_9182# a_35094_9158# 0.0924f
C6241 rowoff_n[13] a_18026_15182# 0.294f
C6242 m2_34288_4386# row_n[2] 0.0128f
C6243 m2_5172_14426# a_4974_14178# 0.165f
C6244 rowon_n[2] a_31078_4138# 0.248f
C6245 col_n[18] a_2275_18218# 0.113f
C6246 col[5] a_7894_11166# 0.0682f
C6247 vcm a_12914_17190# 0.1f
C6248 a_30074_14178# a_31078_14178# 0.843f
C6249 col_n[23] a_2275_7174# 0.113f
C6250 VDD a_8990_7150# 0.483f
C6251 rowoff_n[5] a_20034_7150# 0.294f
C6252 col_n[13] a_16018_5142# 0.251f
C6253 a_2275_18218# a_13918_18194# 0.136f
C6254 VDD a_32482_17552# 0.0779f
C6255 col_n[23] a_26058_17190# 0.251f
C6256 a_2874_1126# a_2966_1126# 0.0991f
C6257 col_n[20] a_22954_7150# 0.0765f
C6258 m2_1732_1950# a_2161_2154# 0.0454f
C6259 m2_2736_1950# a_2475_2154# 0.287f
C6260 vcm a_15014_2130# 0.56f
C6261 a_2275_6170# a_25358_6186# 0.144f
C6262 a_2475_6170# a_27974_6146# 0.264f
C6263 a_14922_6146# a_15014_6146# 0.326f
C6264 col[8] a_2275_15206# 0.0899f
C6265 m2_24248_10410# a_24050_10162# 0.165f
C6266 col[13] a_2275_4162# 0.0899f
C6267 row_n[2] a_8990_4138# 0.282f
C6268 rowoff_n[3] a_29070_5142# 0.294f
C6269 rowon_n[6] a_8898_8154# 0.118f
C6270 a_21038_16186# a_21038_15182# 0.843f
C6271 a_3878_15182# a_4370_15544# 0.0658f
C6272 a_2966_15182# a_3270_15222# 0.0931f
C6273 a_2475_15206# a_5978_15182# 0.316f
C6274 col_n[4] a_7382_3496# 0.0283f
C6275 VDD a_24050_11166# 0.483f
C6276 col_n[14] a_17422_15544# 0.0283f
C6277 m2_1732_5966# col[0] 0.0137f
C6278 col[28] a_2475_14202# 0.136f
C6279 a_9902_3134# a_10298_3174# 0.0313f
C6280 a_2275_3158# a_18938_3134# 0.136f
C6281 col_n[23] rowoff_n[5] 0.0471f
C6282 col_n[22] rowoff_n[4] 0.0471f
C6283 col_n[27] rowoff_n[9] 0.0471f
C6284 col_n[24] rowoff_n[6] 0.0471f
C6285 col_n[26] rowoff_n[8] 0.0471f
C6286 col_n[21] rowoff_n[3] 0.0471f
C6287 col_n[19] rowoff_n[1] 0.0471f
C6288 a_2475_18218# a_11910_18194# 0.264f
C6289 col_n[25] rowoff_n[7] 0.0471f
C6290 col_n[18] rowoff_n[0] 0.0471f
C6291 col_n[20] rowoff_n[2] 0.0471f
C6292 m2_34864_4962# a_2475_5166# 0.282f
C6293 a_32082_1126# a_2275_1150# 0.0924f
C6294 row_n[13] a_29374_15222# 0.0117f
C6295 vcm a_30074_6146# 0.56f
C6296 rowoff_n[11] a_24450_13536# 0.0133f
C6297 col_n[4] a_2475_18218# 0.0529f
C6298 a_33998_13174# a_34490_13536# 0.0658f
C6299 a_33086_13174# a_33390_13214# 0.0931f
C6300 a_29470_1488# VDD 0.0977f
C6301 row_n[15] a_19942_17190# 0.0437f
C6302 a_2475_17214# a_21038_17190# 0.316f
C6303 a_10998_17190# a_12002_17190# 0.843f
C6304 VDD a_4974_14178# 0.483f
C6305 col_n[2] a_4974_3134# 0.251f
C6306 col_n[28] a_31382_4178# 0.084f
C6307 col_n[12] a_15014_15182# 0.251f
C6308 a_2275_5166# a_33998_5142# 0.136f
C6309 row_n[5] a_29982_7150# 0.0437f
C6310 col_n[9] a_11910_5142# 0.0765f
C6311 m2_15212_8402# a_15014_8154# 0.165f
C6312 rowon_n[9] a_29070_11166# 0.248f
C6313 a_30986_1126# a_31382_1166# 0.0313f
C6314 vcm a_10998_9158# 0.56f
C6315 col_n[19] a_21950_17190# 0.0765f
C6316 col[25] a_2275_17214# 0.0899f
C6317 a_29982_10162# a_30074_10162# 0.326f
C6318 rowoff_n[14] a_5978_16186# 0.294f
C6319 col[30] a_2275_6170# 0.0899f
C6320 m2_1732_15002# a_2275_15206# 0.191f
C6321 m2_34864_946# a_2275_1150# 0.281f
C6322 col[28] rowoff_n[14] 0.0901f
C6323 a_2275_14202# a_12002_14178# 0.399f
C6324 m2_34864_16006# ctop 0.0422f
C6325 col_n[11] rowoff_n[10] 0.0471f
C6326 VDD a_20034_18194# 0.0356f
C6327 a_2475_2154# a_26058_2130# 0.316f
C6328 a_31078_3134# a_31078_2130# 0.843f
C6329 col_n[3] a_6378_13536# 0.0283f
C6330 m2_34288_4386# a_34090_4138# 0.165f
C6331 m2_28840_946# VDD 1f
C6332 vcm a_2275_3158# 6.49f
C6333 row_n[9] a_6982_11166# 0.282f
C6334 a_24962_7150# a_25358_7190# 0.0313f
C6335 rowoff_n[9] a_30986_11166# 0.202f
C6336 col[22] a_25054_2130# 0.367f
C6337 rowon_n[13] a_6890_15182# 0.118f
C6338 vcm a_26058_13174# 0.56f
C6339 a_2874_11166# a_3366_11528# 0.0658f
C6340 a_2275_11190# a_3878_11166# 0.136f
C6341 a_2475_11190# a_4882_11166# 0.264f
C6342 VDD a_22954_3134# 0.181f
C6343 col[29] a_31990_4138# 0.0682f
C6344 m2_11772_18014# a_12306_18234# 0.087f
C6345 m2_33860_18014# a_2275_18218# 0.28f
C6346 ctop a_2966_7150# 4.06f
C6347 col_n[15] a_2475_13198# 0.0531f
C6348 a_14010_16186# a_14314_16226# 0.0931f
C6349 a_2275_16210# a_27062_16186# 0.399f
C6350 a_14922_16186# a_15414_16548# 0.0658f
C6351 rowon_n[3] a_16930_5142# 0.118f
C6352 col_n[20] a_2475_2154# 0.0531f
C6353 a_21038_4138# a_22042_4138# 0.843f
C6354 row_n[1] a_4274_3174# 0.0117f
C6355 col_n[17] a_20338_2170# 0.0839f
C6356 m2_6176_6394# a_5978_6146# 0.165f
C6357 vcm a_16322_7190# 0.155f
C6358 col_n[1] a_3970_13174# 0.251f
C6359 col_n[27] a_30378_14218# 0.084f
C6360 rowoff_n[12] a_12402_14540# 0.0133f
C6361 col_n[12] col_n[13] 0.0101f
C6362 vcm col_n[25] 1.94f
C6363 VDD col_n[28] 5.17f
C6364 col[12] rowoff_n[15] 0.0901f
C6365 col[5] a_2475_10186# 0.136f
C6366 col[22] col[23] 0.0355f
C6367 ctop a_29070_2130# 4.06f
C6368 vcm a_6982_16186# 0.56f
C6369 a_2475_13198# a_19942_13174# 0.264f
C6370 a_10906_13174# a_10998_13174# 0.326f
C6371 col_n[8] a_10906_15182# 0.0765f
C6372 a_2275_13198# a_17326_13214# 0.144f
C6373 VDD a_3366_6508# 0.0779f
C6374 m2_29844_18014# a_2475_18218# 0.286f
C6375 row_n[12] a_27974_14178# 0.0437f
C6376 vcm a_9902_1126# 0.0989f
C6377 m2_6176_15430# rowon_n[13] 0.0322f
C6378 col_n[12] a_2275_16210# 0.113f
C6379 a_12002_6146# a_12002_5142# 0.843f
C6380 m2_12200_11414# rowon_n[9] 0.0322f
C6381 m2_18224_7398# rowon_n[5] 0.0322f
C6382 col_n[17] a_2275_5166# 0.113f
C6383 m2_24248_3382# rowon_n[1] 0.0322f
C6384 vcm a_31382_11206# 0.155f
C6385 a_2275_10186# a_10906_10162# 0.136f
C6386 a_5886_10162# a_6282_10202# 0.0313f
C6387 m2_34864_17010# a_34090_17190# 0.843f
C6388 ctop a_9994_5142# 4.11f
C6389 col[21] a_24050_12170# 0.367f
C6390 a_2475_15206# a_35002_15182# 0.264f
C6391 a_2275_15206# a_32386_15222# 0.144f
C6392 VDD a_18938_10162# 0.181f
C6393 col[18] a_20946_2130# 0.0682f
C6394 col[28] a_30986_14178# 0.0682f
C6395 col[2] a_2275_13198# 0.0899f
C6396 a_24050_3134# a_24354_3174# 0.0931f
C6397 a_24962_3134# a_25454_3496# 0.0658f
C6398 col[7] a_2275_2154# 0.0899f
C6399 vcm a_24962_5142# 0.1f
C6400 m2_1732_10986# m2_2160_11414# 0.165f
C6401 a_2475_7174# a_2874_7150# 0.264f
C6402 a_1957_7174# a_2275_7174# 0.158f
C6403 rowoff_n[10] a_18938_12170# 0.202f
C6404 m2_33284_16434# rowon_n[14] 0.0322f
C6405 row_n[6] a_15014_8154# 0.282f
C6406 vcm a_12306_14218# 0.155f
C6407 a_2275_12194# a_25966_12170# 0.136f
C6408 rowon_n[10] a_14922_12170# 0.118f
C6409 col_n[16] a_19334_12210# 0.084f
C6410 col[22] a_2475_12194# 0.136f
C6411 VDD a_10394_4500# 0.0779f
C6412 col[27] a_2475_1150# 0.136f
C6413 ctop a_25054_9158# 4.11f
C6414 a_25966_17190# a_26058_17190# 0.326f
C6415 VDD a_33998_14178# 0.181f
C6416 row_n[8] a_3878_10162# 0.0437f
C6417 rowon_n[0] a_24962_2130# 0.118f
C6418 rowoff_n[0] a_10906_2130# 0.202f
C6419 rowon_n[12] a_2966_14178# 0.248f
C6420 col_n[27] a_30474_6508# 0.0283f
C6421 m2_15788_946# ctop 0.0428f
C6422 col_n[29] a_2275_18218# 0.113f
C6423 vcm a_5886_8154# 0.1f
C6424 m2_22816_18014# m2_23244_18442# 0.165f
C6425 a_2475_9182# a_18026_9158# 0.316f
C6426 a_27062_10162# a_27062_9158# 0.843f
C6427 rowoff_n[14] a_35002_16186# 0.202f
C6428 vcm a_27366_18234# 0.16f
C6429 a_20946_14178# a_21342_14218# 0.0313f
C6430 VDD a_25454_8516# 0.0779f
C6431 rowoff_n[5] a_1957_7174# 0.0219f
C6432 ctop a_5978_12170# 4.11f
C6433 VDD a_14922_17190# 0.181f
C6434 row_n[0] a_2161_2154# 0.0221f
C6435 col[10] a_13006_10162# 0.367f
C6436 col[19] a_2275_15206# 0.0899f
C6437 rowon_n[4] a_2475_6170# 0.31f
C6438 col[17] a_19942_12170# 0.0682f
C6439 m3_34568_1078# VDD 0.0111f
C6440 col[24] a_2275_4162# 0.0899f
C6441 row_n[9] a_34394_11206# 0.0117f
C6442 a_5886_6146# a_6378_6508# 0.0658f
C6443 a_2275_6170# a_8990_6146# 0.399f
C6444 a_4974_6146# a_5278_6186# 0.0931f
C6445 rowon_n[13] a_35094_15182# 0.0141f
C6446 col_n[25] a_28066_6146# 0.251f
C6447 rowoff_n[3] a_11398_5504# 0.0133f
C6448 vcm a_20946_12170# 0.1f
C6449 a_2475_11190# a_33086_11166# 0.316f
C6450 a_17022_11166# a_18026_11166# 0.843f
C6451 VDD a_17022_2130# 0.483f
C6452 m2_30848_18014# a_31382_18234# 0.087f
C6453 VDD a_6378_11528# 0.0779f
C6454 col_n[31] rowoff_n[2] 0.0471f
C6455 col_n[29] rowoff_n[0] 0.0471f
C6456 col_n[5] a_8290_10202# 0.084f
C6457 col_n[30] rowoff_n[1] 0.0471f
C6458 m2_33860_18014# m3_32988_18146# 0.0341f
C6459 ctop a_21038_16186# 4.11f
C6460 col_n[15] a_2475_18218# 0.0529f
C6461 rowoff_n[1] a_20434_3496# 0.0133f
C6462 rowoff_n[8] a_2874_10162# 0.202f
C6463 row_n[13] a_13006_15182# 0.282f
C6464 m2_34864_15002# m2_34864_13998# 0.843f
C6465 a_2275_8178# a_24050_8154# 0.399f
C6466 rowoff_n[11] a_6890_13174# 0.202f
C6467 col_n[16] a_19430_4500# 0.0283f
C6468 col_n[9] a_2475_11190# 0.0531f
C6469 vcm a_34394_16226# 0.155f
C6470 col_n[26] a_29470_16548# 0.0283f
C6471 a_7986_13174# a_7986_12170# 0.843f
C6472 VDD a_32082_6146# 0.483f
C6473 row_n[3] a_23046_5142# 0.282f
C6474 rowon_n[7] a_22954_9158# 0.118f
C6475 a_2161_17214# a_2275_17214# 0.183f
C6476 m2_5172_14426# row_n[12] 0.0128f
C6477 a_2475_17214# a_2966_17190# 0.317f
C6478 m2_11196_10410# row_n[8] 0.0128f
C6479 rowoff_n[6] a_12002_8154# 0.294f
C6480 VDD a_21438_15544# 0.0779f
C6481 a_2475_2154# m2_34864_1950# 0.282f
C6482 m2_17220_6394# row_n[4] 0.0128f
C6483 m3_12908_18146# a_13006_17190# 0.0303f
C6484 a_2275_5166# a_14314_5182# 0.144f
C6485 a_2475_5166# a_16930_5142# 0.264f
C6486 row_n[5] a_10298_7190# 0.0117f
C6487 m2_24824_946# col_n[22] 0.331f
C6488 col[6] a_8898_10162# 0.0682f
C6489 rowoff_n[15] a_22954_17190# 0.202f
C6490 a_20946_10162# a_21438_10524# 0.0658f
C6491 a_20034_10162# a_20338_10202# 0.0931f
C6492 rowoff_n[4] a_21038_6146# 0.294f
C6493 col_n[14] a_17022_4138# 0.251f
C6494 a_32082_15182# a_33086_15182# 0.843f
C6495 col_n[22] rowoff_n[10] 0.0471f
C6496 m2_22816_18014# col[20] 0.347f
C6497 VDD a_13006_9158# 0.483f
C6498 col_n[24] a_27062_16186# 0.251f
C6499 col_n[6] a_2275_14202# 0.113f
C6500 col_n[21] a_23958_6146# 0.0765f
C6501 VDD a_1957_18218# 0.4f
C6502 col_n[11] a_2275_3158# 0.113f
C6503 col_n[31] a_33998_18194# 0.0762f
C6504 a_2275_2154# a_7894_2130# 0.136f
C6505 m2_32280_15430# row_n[13] 0.0128f
C6506 vcm a_19030_4138# 0.56f
C6507 rowon_n[1] a_9994_3134# 0.248f
C6508 a_16930_7150# a_17022_7150# 0.326f
C6509 a_2275_7174# a_29374_7190# 0.144f
C6510 a_2475_7174# a_31990_7150# 0.264f
C6511 rowoff_n[2] a_30074_4138# 0.294f
C6512 col_n[26] a_2475_13198# 0.0531f
C6513 col_n[31] a_2475_2154# 0.0531f
C6514 col_n[5] a_8386_2492# 0.0283f
C6515 a_23046_17190# a_23046_16186# 0.843f
C6516 a_2475_16210# a_9994_16186# 0.316f
C6517 col_n[15] a_18426_14540# 0.0283f
C6518 VDD a_28066_13174# 0.483f
C6519 a_2275_4162# a_22954_4138# 0.136f
C6520 a_11910_4138# a_12306_4178# 0.0313f
C6521 VDD row_n[12] 3.29f
C6522 col_n[2] rowon_n[14] 0.111f
C6523 col_n[1] row_n[14] 0.298f
C6524 m3_11904_1078# ctop 0.21f
C6525 col_n[4] rowon_n[15] 0.111f
C6526 vcm rowon_n[13] 0.65f
C6527 col_n[3] row_n[15] 0.298f
C6528 col_n[0] row_n[13] 0.298f
C6529 sample rowon_n[12] 0.0935f
C6530 col[23] rowoff_n[15] 0.0901f
C6531 col[16] a_2475_10186# 0.136f
C6532 vcm a_34090_8154# 0.56f
C6533 row_n[10] a_21038_12170# 0.282f
C6534 col_n[0] a_2874_10162# 0.0765f
C6535 col_n[6] rowoff_n[11] 0.0471f
C6536 rowon_n[14] a_20946_16186# 0.118f
C6537 col_n[3] a_5978_2130# 0.251f
C6538 col_n[29] a_32386_3174# 0.084f
C6539 row_n[0] a_31078_2130# 0.282f
C6540 VDD a_8990_16186# 0.483f
C6541 col_n[23] a_2275_16210# 0.113f
C6542 row_n[12] a_8290_14218# 0.0117f
C6543 a_2475_1150# a_15014_1126# 0.0299f
C6544 col_n[13] a_16018_14178# 0.251f
C6545 rowon_n[4] a_30986_6146# 0.118f
C6546 col_n[28] a_2275_5166# 0.113f
C6547 col_n[10] a_12914_4138# 0.0765f
C6548 vcm a_24354_2170# 0.155f
C6549 col_n[20] a_22954_16186# 0.0765f
C6550 m2_13780_946# m2_14784_946# 0.843f
C6551 vcm a_15014_11166# 0.56f
C6552 row_n[2] a_18330_4178# 0.0117f
C6553 a_31990_11166# a_32082_11166# 0.326f
C6554 VDD a_11910_1126# 0.405f
C6555 m2_20232_17438# a_20034_17190# 0.165f
C6556 col[13] a_2275_13198# 0.0899f
C6557 a_2275_15206# a_16018_15182# 0.399f
C6558 col[18] a_2275_2154# 0.0899f
C6559 rowon_n[0] m2_29268_2378# 0.0322f
C6560 row_n[4] a_8898_6146# 0.0437f
C6561 col_n[4] a_7382_12532# 0.0283f
C6562 a_2475_3158# a_30074_3134# 0.316f
C6563 a_33086_4138# a_33086_3134# 0.843f
C6564 col_n[1] a_3878_2130# 0.0765f
C6565 rowon_n[8] a_7986_10162# 0.248f
C6566 rowoff_n[8] a_31990_10162# 0.202f
C6567 vcm a_5278_5182# 0.155f
C6568 rowoff_n[11] a_35094_13174# 0.0135f
C6569 a_26970_8154# a_27366_8194# 0.0313f
C6570 col[30] a_32994_3134# 0.0682f
C6571 vcm a_30074_15182# 0.56f
C6572 a_2275_12194# a_6282_12210# 0.144f
C6573 a_2475_12194# a_8898_12170# 0.264f
C6574 VDD a_26970_5142# 0.181f
C6575 m2_11196_18442# VDD 0.0456f
C6576 a_16930_17190# a_17422_17552# 0.0658f
C6577 a_16018_17190# a_16322_17230# 0.0931f
C6578 a_2275_17214# a_31078_17190# 0.399f
C6579 col_n[3] a_2475_9182# 0.0531f
C6580 col_n[18] a_21342_1166# 0.0839f
C6581 a_23046_5142# a_24050_5142# 0.843f
C6582 col_n[28] a_31382_13214# 0.084f
C6583 col_n[2] a_4974_12170# 0.251f
C6584 m2_4744_18014# m2_5748_18014# 0.843f
C6585 vcm a_20338_9198# 0.155f
C6586 a_35002_10162# a_35398_10202# 0.0313f
C6587 col_n[9] a_11910_14178# 0.0765f
C6588 m2_11196_15430# a_10998_15182# 0.165f
C6589 ctop a_33086_4138# 4.11f
C6590 vcm a_10998_18194# 0.165f
C6591 a_2475_14202# a_23958_14178# 0.264f
C6592 a_2275_14202# a_21342_14218# 0.144f
C6593 a_12914_14178# a_13006_14178# 0.326f
C6594 VDD a_7894_8154# 0.181f
C6595 row_n[7] a_29070_9158# 0.282f
C6596 col[30] a_2275_15206# 0.0899f
C6597 m2_1732_8978# rowon_n[7] 0.236f
C6598 m2_7180_5390# rowon_n[3] 0.0322f
C6599 rowon_n[11] a_28978_13174# 0.118f
C6600 VDD a_29374_18234# 0.019f
C6601 m3_30980_18146# VDD 0.0911f
C6602 row_n[9] a_16322_11206# 0.0117f
C6603 vcm a_13918_3134# 0.1f
C6604 a_14010_7150# a_14010_6146# 0.843f
C6605 m2_30272_11414# a_30074_11166# 0.165f
C6606 vcm a_2275_12194# 6.49f
C6607 a_7894_11166# a_8290_11206# 0.0313f
C6608 a_2275_11190# a_14922_11166# 0.136f
C6609 VDD a_33486_3496# 0.0779f
C6610 row_n[8] rowoff_n[7] 0.085f
C6611 col[22] a_25054_11166# 0.367f
C6612 col_n[5] a_2275_1150# 0.113f
C6613 m2_34864_10986# VDD 0.772f
C6614 col[19] a_21950_1126# 0.0682f
C6615 ctop a_14010_7150# 4.11f
C6616 a_2966_16186# a_2966_15182# 0.843f
C6617 row_n[11] a_6890_13174# 0.0437f
C6618 col[29] a_31990_13174# 0.0682f
C6619 VDD a_22954_12170# 0.181f
C6620 col_n[26] a_2475_18218# 0.0529f
C6621 m2_9764_18014# m3_9896_18146# 3.79f
C6622 rowon_n[15] a_5978_17190# 0.248f
C6623 ctop a_2966_16186# 4.06f
C6624 m2_22240_14426# rowon_n[12] 0.0322f
C6625 m2_28264_10410# rowon_n[8] 0.0322f
C6626 m2_34288_6394# rowon_n[4] 0.0322f
C6627 a_26058_4138# a_26362_4178# 0.0931f
C6628 a_26970_4138# a_27462_4500# 0.0658f
C6629 col_n[20] a_2475_11190# 0.0531f
C6630 rowoff_n[1] a_2161_3158# 0.0226f
C6631 row_n[1] a_16930_3134# 0.0437f
C6632 rowon_n[5] a_16018_7150# 0.248f
C6633 vcm a_28978_7150# 0.1f
C6634 rowoff_n[12] a_23046_14178# 0.294f
C6635 a_2475_8178# a_6982_8154# 0.316f
C6636 a_3970_8154# a_4974_8154# 0.843f
C6637 m2_1732_12994# a_1957_13198# 0.245f
C6638 col_n[17] a_20338_11206# 0.084f
C6639 vcm a_16322_16226# 0.155f
C6640 a_2275_13198# a_29982_13174# 0.136f
C6641 VDD a_14410_6508# 0.0779f
C6642 ctop a_29070_11166# 4.11f
C6643 a_27974_18194# a_28066_18194# 0.0991f
C6644 col[10] a_2475_8178# 0.136f
C6645 VDD a_3366_15544# 0.0779f
C6646 a_22954_1126# a_23046_1126# 0.0991f
C6647 col_n[28] a_31478_5504# 0.0283f
C6648 m2_12776_946# m3_11904_1078# 0.0341f
C6649 m3_1864_18146# m3_1864_17142# 0.202f
C6650 m2_21236_9406# a_21038_9158# 0.165f
C6651 vcm a_9902_10162# 0.1f
C6652 a_2475_10186# a_22042_10162# 0.316f
C6653 a_29070_11166# a_29070_10162# 0.843f
C6654 row_n[14] a_27062_16186# 0.282f
C6655 col_n[17] a_2275_14202# 0.113f
C6656 rowoff_n[4] a_2966_6146# 0.294f
C6657 col_n[22] a_2275_3158# 0.113f
C6658 a_22954_15182# a_23350_15222# 0.0313f
C6659 VDD a_29470_10524# 0.0779f
C6660 col[11] a_14010_9158# 0.367f
C6661 ctop a_9994_14178# 4.11f
C6662 col[18] a_20946_11166# 0.0682f
C6663 col_n[26] a_29070_5142# 0.251f
C6664 a_2275_7174# a_13006_7150# 0.399f
C6665 rowoff_n[2] a_12402_4500# 0.0133f
C6666 a_7894_7150# a_8386_7512# 0.0658f
C6667 a_6982_7150# a_7286_7190# 0.0931f
C6668 col[7] a_2275_11190# 0.0899f
C6669 rowoff_n[10] a_29470_12532# 0.0133f
C6670 m2_28840_18014# vcm 0.353f
C6671 row_n[6] a_24354_8194# 0.0117f
C6672 vcm a_24962_14178# 0.1f
C6673 a_19030_12170# a_20034_12170# 0.843f
C6674 VDD a_21038_4138# 0.483f
C6675 col_n[6] a_9294_9198# 0.084f
C6676 VDD a_10394_13536# 0.0779f
C6677 col_n[12] row_n[14] 0.298f
C6678 col_n[13] rowon_n[14] 0.111f
C6679 col_n[11] rowon_n[13] 0.111f
C6680 col_n[14] row_n[15] 0.298f
C6681 col_n[9] rowon_n[12] 0.111f
C6682 col_n[8] row_n[12] 0.298f
C6683 col_n[5] rowon_n[10] 0.111f
C6684 sample row_n[7] 0.423f
C6685 col_n[4] row_n[10] 0.298f
C6686 col_n[6] row_n[11] 0.298f
C6687 col_n[1] rowon_n[8] 0.111f
C6688 vcm row_n[8] 0.616f
C6689 col_n[7] rowon_n[11] 0.111f
C6690 col_n[23] col_n[24] 0.0101f
C6691 col_n[10] row_n[13] 0.298f
C6692 col_n[2] row_n[9] 0.298f
C6693 col_n[0] rowon_n[7] 0.111f
C6694 VDD rowon_n[6] 3.04f
C6695 col_n[3] rowon_n[9] 0.111f
C6696 col_n[15] rowon_n[15] 0.111f
C6697 col[27] a_2475_10186# 0.136f
C6698 row_n[8] a_14922_10162# 0.0437f
C6699 rowoff_n[0] a_21438_2492# 0.0133f
C6700 rowoff_n[7] a_3970_9158# 0.294f
C6701 rowon_n[12] a_14010_14178# 0.248f
C6702 a_2475_4162# a_5886_4138# 0.264f
C6703 a_2275_4162# a_3270_4178# 0.144f
C6704 m3_7888_18146# ctop 0.209f
C6705 col_n[17] a_20434_3496# 0.0283f
C6706 col_n[17] rowoff_n[11] 0.0471f
C6707 m2_12200_7398# a_12002_7150# 0.165f
C6708 rowoff_n[13] a_10998_15182# 0.294f
C6709 col_n[27] a_30474_15544# 0.0283f
C6710 a_2275_9182# a_28066_9158# 0.399f
C6711 m2_6176_4386# row_n[2] 0.0128f
C6712 row_n[10] a_2966_12170# 0.281f
C6713 rowon_n[2] a_24050_4138# 0.248f
C6714 vcm a_5886_17190# 0.1f
C6715 m3_19936_1078# a_20034_1126# 3.24f
C6716 rowon_n[14] a_2275_16210# 1.79f
C6717 a_9994_14178# a_9994_13174# 0.843f
C6718 VDD a_2475_7174# 26.1f
C6719 rowoff_n[5] a_13006_7150# 0.294f
C6720 a_2275_18218# a_6890_18194# 0.136f
C6721 VDD a_25454_17552# 0.0779f
C6722 a_32994_2130# a_33390_2170# 0.0313f
C6723 col[0] a_2874_7150# 0.0682f
C6724 m2_31276_3382# a_31078_3134# 0.165f
C6725 vcm a_7986_2130# 0.56f
C6726 a_2275_6170# a_18330_6186# 0.144f
C6727 a_2475_6170# a_20946_6146# 0.264f
C6728 col[7] a_9902_9158# 0.0682f
C6729 col[24] a_2275_13198# 0.0899f
C6730 rowoff_n[3] a_22042_5142# 0.294f
C6731 row_n[2] a_2475_4162# 0.405f
C6732 a_22042_11166# a_22346_11206# 0.0931f
C6733 a_22954_11166# a_23446_11528# 0.0658f
C6734 col_n[15] a_18026_3134# 0.251f
C6735 col[29] a_2275_2154# 0.0899f
C6736 m2_15212_17438# row_n[15] 0.0128f
C6737 m2_21236_13422# row_n[11] 0.0128f
C6738 col_n[25] a_28066_15182# 0.251f
C6739 m2_27260_9406# row_n[7] 0.0128f
C6740 m2_33284_5390# row_n[3] 0.0128f
C6741 col_n[22] a_24962_5142# 0.0765f
C6742 row_n[11] a_35094_13174# 0.0123f
C6743 a_33998_16186# a_34394_16226# 0.0313f
C6744 VDD a_17022_11166# 0.483f
C6745 m2_1732_16006# m3_1864_17142# 0.0341f
C6746 rowon_n[15] a_35002_17190# 0.118f
C6747 col_n[1] rowoff_n[12] 0.0471f
C6748 a_2275_3158# a_11910_3134# 0.136f
C6749 a_2475_18218# a_4882_18194# 0.264f
C6750 rowoff_n[1] a_31078_3134# 0.294f
C6751 a_25054_1126# a_2275_1150# 0.0924f
C6752 row_n[13] a_22346_15222# 0.0117f
C6753 vcm a_23046_6146# 0.56f
C6754 a_18938_8154# a_19030_8154# 0.326f
C6755 a_2275_8178# a_33390_8194# 0.144f
C6756 rowoff_n[11] a_17422_13536# 0.0133f
C6757 col_n[6] a_9390_1488# 0.0283f
C6758 col_n[16] a_19430_13536# 0.0283f
C6759 row_n[3] a_32386_5182# 0.0117f
C6760 row_n[15] a_12914_17190# 0.0437f
C6761 col_n[14] a_2475_9182# 0.0531f
C6762 a_2475_17214# a_14010_17190# 0.316f
C6763 VDD a_32082_15182# 0.483f
C6764 a_13918_5142# a_14314_5182# 0.0313f
C6765 a_2275_5166# a_26970_5142# 0.136f
C6766 row_n[5] a_22954_7150# 0.0437f
C6767 rowon_n[9] a_22042_11166# 0.248f
C6768 vcm a_3970_9158# 0.56f
C6769 rowoff_n[15] a_33486_17552# 0.0133f
C6770 col[4] a_2475_6170# 0.136f
C6771 a_2275_14202# a_4974_14178# 0.399f
C6772 m2_6752_946# a_7286_1166# 0.087f
C6773 a_3878_14178# a_3970_14178# 0.326f
C6774 a_2874_14178# a_3270_14218# 0.0313f
C6775 m2_21812_946# a_2475_1150# 0.286f
C6776 col_n[30] a_33390_2170# 0.084f
C6777 col_n[14] a_17022_13174# 0.251f
C6778 col_n[11] a_13918_3134# 0.0765f
C6779 VDD a_13006_18194# 0.0356f
C6780 a_9994_2130# a_10998_2130# 0.843f
C6781 a_2475_2154# a_19030_2130# 0.316f
C6782 col_n[21] a_23958_15182# 0.0765f
C6783 m2_13204_1374# VDD 0.0194f
C6784 col_n[11] a_2275_12194# 0.113f
C6785 vcm a_28370_4178# 0.155f
C6786 rowoff_n[9] a_23958_11166# 0.202f
C6787 row_n[4] rowoff_n[4] 0.209f
C6788 m2_1732_17010# sample_n 0.0522f
C6789 col_n[16] a_2275_1150# 0.0948f
C6790 vcm a_19030_13174# 0.56f
C6791 a_33998_12170# a_34090_12170# 0.326f
C6792 VDD a_15926_3134# 0.181f
C6793 m2_19804_18014# a_2275_18218# 0.28f
C6794 a_2275_16210# a_20034_16186# 0.399f
C6795 rowon_n[3] a_9902_5142# 0.118f
C6796 col_n[31] a_2475_11190# 0.0531f
C6797 col_n[5] a_8386_11528# 0.0283f
C6798 a_27974_1126# m2_27836_946# 0.225f
C6799 col[1] a_2275_9182# 0.0899f
C6800 rowoff_n[7] a_32994_9158# 0.202f
C6801 a_2475_4162# a_34090_4138# 0.316f
C6802 col[31] a_33998_2130# 0.0682f
C6803 vcm a_9294_7190# 0.155f
C6804 a_28978_9158# a_29374_9198# 0.0313f
C6805 rowoff_n[12] a_5374_14540# 0.0133f
C6806 row_n[10] a_30378_12210# 0.0117f
C6807 vcm a_34090_17190# 0.56f
C6808 ctop a_22042_2130# 4.06f
C6809 a_2475_13198# a_12914_13174# 0.264f
C6810 a_2275_13198# a_10298_13214# 0.144f
C6811 col[21] a_2475_8178# 0.136f
C6812 VDD a_30986_7150# 0.181f
C6813 a_2275_18218# a_35094_18194# 0.0924f
C6814 a_18938_18194# a_19430_18556# 0.0658f
C6815 m2_15788_18014# a_2475_18218# 0.286f
C6816 row_n[12] a_20946_14178# 0.0437f
C6817 a_13918_1126# a_14410_1488# 0.0658f
C6818 col_n[3] a_5978_11166# 0.251f
C6819 col_n[29] a_32386_12210# 0.084f
C6820 vcm a_2161_1150# 0.0169f
C6821 a_25054_6146# a_26058_6146# 0.843f
C6822 col_n[28] a_2275_14202# 0.113f
C6823 col_n[10] a_12914_13174# 0.0765f
C6824 vcm a_24354_11206# 0.155f
C6825 row_n[2] a_30986_4138# 0.0437f
C6826 a_2874_10162# a_2966_10162# 0.326f
C6827 VDD a_22442_1488# 0.0977f
C6828 rowon_n[6] a_30074_8154# 0.248f
C6829 a_2275_15206# a_25358_15222# 0.144f
C6830 a_14922_15182# a_15014_15182# 0.326f
C6831 a_2475_15206# a_27974_15182# 0.264f
C6832 VDD a_11910_10162# 0.181f
C6833 m2_1732_12994# m3_1864_14130# 0.0341f
C6834 col[18] a_2275_11190# 0.0899f
C6835 a_2475_18218# a_33086_18194# 0.0299f
C6836 vcm a_17934_5142# 0.1f
C6837 rowoff_n[10] a_11910_12170# 0.202f
C6838 col_n[1] a_3878_11166# 0.0765f
C6839 a_16018_8154# a_16018_7150# 0.843f
C6840 a_31078_1126# vcm 0.165f
C6841 col[23] a_26058_10162# 0.367f
C6842 m2_5172_16434# rowon_n[14] 0.0322f
C6843 m2_11196_12418# rowon_n[10] 0.0322f
C6844 row_n[6] a_7986_8154# 0.282f
C6845 vcm a_5278_14218# 0.155f
C6846 m2_17220_8402# rowon_n[6] 0.0322f
C6847 a_2275_12194# a_18938_12170# 0.136f
C6848 a_9902_12170# a_10298_12210# 0.0313f
C6849 m2_23244_4386# rowon_n[2] 0.0322f
C6850 VDD a_2966_4138# 0.485f
C6851 rowon_n[10] a_7894_12170# 0.118f
C6852 col_n[16] rowon_n[10] 0.111f
C6853 col_n[4] rowon_n[4] 0.111f
C6854 col_n[0] row_n[2] 0.298f
C6855 col_n[12] rowon_n[8] 0.111f
C6856 col_n[11] row_n[8] 0.298f
C6857 col_n[2] rowon_n[3] 0.111f
C6858 col_n[25] row_n[15] 0.298f
C6859 col_n[20] rowon_n[12] 0.111f
C6860 col_n[3] row_n[4] 0.298f
C6861 col_n[7] row_n[6] 0.298f
C6862 col_n[26] rowon_n[15] 0.111f
C6863 sample rowon_n[1] 0.0935f
C6864 col_n[23] row_n[14] 0.298f
C6865 col_n[18] rowon_n[11] 0.111f
C6866 col_n[1] row_n[3] 0.298f
C6867 col_n[14] rowon_n[9] 0.111f
C6868 col_n[17] row_n[11] 0.298f
C6869 col_n[22] rowon_n[13] 0.111f
C6870 col_n[21] row_n[13] 0.298f
C6871 col_n[13] row_n[9] 0.298f
C6872 col_n[5] row_n[5] 0.298f
C6873 col_n[24] rowon_n[14] 0.111f
C6874 col_n[9] row_n[7] 0.298f
C6875 col_n[6] rowon_n[5] 0.111f
C6876 VDD row_n[1] 3.29f
C6877 col_n[15] row_n[10] 0.298f
C6878 col[30] a_32994_12170# 0.0682f
C6879 col_n[10] rowon_n[7] 0.111f
C6880 col_n[19] row_n[12] 0.298f
C6881 vcm rowon_n[2] 0.65f
C6882 col_n[8] rowon_n[6] 0.111f
C6883 m2_32856_18014# VDD 0.993f
C6884 ctop a_18026_9158# 4.11f
C6885 VDD a_26970_14178# 0.181f
C6886 col_n[28] rowoff_n[11] 0.0471f
C6887 rowon_n[0] a_17934_2130# 0.118f
C6888 rowoff_n[0] a_3366_2492# 0.0133f
C6889 a_28978_5142# a_29470_5504# 0.0658f
C6890 a_28066_5142# a_28370_5182# 0.0931f
C6891 col_n[18] a_21342_10202# 0.084f
C6892 vcm a_32994_9158# 0.1f
C6893 m2_15788_18014# m2_16216_18442# 0.165f
C6894 col_n[8] a_2475_7174# 0.0531f
C6895 a_2475_9182# a_10998_9158# 0.316f
C6896 a_5978_9158# a_6982_9158# 0.843f
C6897 rowoff_n[14] a_27974_16186# 0.202f
C6898 vcm a_20338_18234# 0.16f
C6899 m3_32988_1078# a_33086_2130# 0.0302f
C6900 m2_32280_17438# rowon_n[15] 0.0322f
C6901 a_2275_14202# a_33998_14178# 0.136f
C6902 VDD a_18426_8516# 0.0779f
C6903 ctop a_33086_13174# 4.11f
C6904 col_n[29] a_32482_4500# 0.0283f
C6905 VDD a_7894_17190# 0.181f
C6906 a_24962_2130# a_25054_2130# 0.326f
C6907 m3_6884_1078# VDD 0.0157f
C6908 row_n[9] a_28978_11166# 0.0437f
C6909 a_2475_6170# a_2275_6170# 2.76f
C6910 a_1957_6170# a_2161_6170# 0.115f
C6911 m2_34864_11990# vcm 0.395f
C6912 rowon_n[13] a_28066_15182# 0.248f
C6913 rowoff_n[3] a_4370_5504# 0.0133f
C6914 vcm a_13918_12170# 0.1f
C6915 a_2475_11190# a_26058_11166# 0.316f
C6916 a_31078_12170# a_31078_11166# 0.843f
C6917 VDD a_9994_2130# 0.483f
C6918 col[12] a_15014_8154# 0.367f
C6919 a_24962_16186# a_25358_16226# 0.0313f
C6920 VDD a_33486_12532# 0.0779f
C6921 m2_23820_18014# m3_24956_18146# 0.0341f
C6922 col_n[12] rowoff_n[12] 0.0471f
C6923 col_n[5] a_2275_10186# 0.113f
C6924 col[19] a_21950_10162# 0.0682f
C6925 ctop a_14010_16186# 4.11f
C6926 col_n[27] a_30074_4138# 0.251f
C6927 rowoff_n[1] a_13406_3496# 0.0133f
C6928 row_n[13] a_5978_15182# 0.282f
C6929 a_2275_8178# a_17022_8154# 0.399f
C6930 a_9902_8154# a_10394_8516# 0.0658f
C6931 a_8990_8154# a_9294_8194# 0.0931f
C6932 col_n[25] a_2475_9182# 0.0531f
C6933 vcm a_28978_16186# 0.1f
C6934 col_n[7] a_10298_8194# 0.084f
C6935 a_21038_13174# a_22042_13174# 0.843f
C6936 VDD a_25054_6146# 0.483f
C6937 row_n[3] a_16018_5142# 0.282f
C6938 rowon_n[7] a_15926_9158# 0.118f
C6939 VDD a_14410_15544# 0.0779f
C6940 rowoff_n[6] a_4974_8154# 0.294f
C6941 col[10] a_2475_17214# 0.136f
C6942 col_n[18] a_21438_2492# 0.0283f
C6943 a_2275_5166# a_7286_5182# 0.144f
C6944 row_n[5] a_3270_7190# 0.0117f
C6945 a_5886_5142# a_5978_5142# 0.326f
C6946 a_2475_5166# a_9902_5142# 0.264f
C6947 col[15] a_2475_6170# 0.136f
C6948 col_n[28] a_31478_14540# 0.0283f
C6949 m2_27836_946# m3_27968_1078# 3.79f
C6950 a_2275_10186# a_32082_10162# 0.399f
C6951 rowoff_n[15] a_15926_17190# 0.202f
C6952 m2_17220_16434# a_17022_16186# 0.165f
C6953 rowoff_n[4] a_14010_6146# 0.294f
C6954 a_12002_15182# a_12002_14178# 0.843f
C6955 VDD a_5978_9158# 0.483f
C6956 m2_1732_9982# m3_1864_11118# 0.0341f
C6957 col[1] a_3970_6146# 0.367f
C6958 col_n[22] a_2275_12194# 0.113f
C6959 rowon_n[0] rowoff_n[0] 20.2f
C6960 ctop rowoff_n[4] 0.177f
C6961 col_n[27] a_2275_1150# 0.113f
C6962 m2_4168_15430# row_n[13] 0.0128f
C6963 m2_10192_11414# row_n[9] 0.0128f
C6964 col[8] a_10906_8154# 0.0682f
C6965 m2_16216_7398# row_n[5] 0.0128f
C6966 m2_22240_3382# row_n[1] 0.0128f
C6967 vcm a_12002_4138# 0.56f
C6968 a_2275_7174# a_22346_7190# 0.144f
C6969 rowon_n[1] a_2874_3134# 0.118f
C6970 a_2475_7174# a_24962_7150# 0.264f
C6971 rowoff_n[2] a_23046_4138# 0.294f
C6972 col_n[16] a_19030_2130# 0.25f
C6973 m2_1732_2954# sample 0.2f
C6974 col_n[26] a_29070_14178# 0.251f
C6975 a_24962_12170# a_25454_12532# 0.0658f
C6976 a_24050_12170# a_24354_12210# 0.0931f
C6977 col_n[23] a_25966_4138# 0.0765f
C6978 m2_1732_13998# VDD 0.856f
C6979 col[12] a_2275_9182# 0.0899f
C6980 a_1957_16210# a_2275_16210# 0.158f
C6981 a_2475_16210# a_2874_16186# 0.264f
C6982 VDD a_21038_13174# 0.483f
C6983 col_n[6] a_9294_18234# 0.084f
C6984 rowoff_n[0] a_32082_2130# 0.294f
C6985 a_2275_4162# a_15926_4138# 0.136f
C6986 m2_8760_946# col_n[6] 0.331f
C6987 m3_34996_10114# ctop 0.209f
C6988 m2_31276_16434# row_n[14] 0.0128f
C6989 vcm a_27062_8154# 0.56f
C6990 a_20946_9158# a_21038_9158# 0.326f
C6991 m2_8184_14426# a_7986_14178# 0.165f
C6992 col_n[17] a_20434_12532# 0.0283f
C6993 row_n[10] a_14010_12170# 0.282f
C6994 rowon_n[14] a_13918_16186# 0.118f
C6995 row_n[0] a_24050_2130# 0.282f
C6996 VDD a_2475_16210# 26.1f
C6997 a_2475_1150# a_7986_1126# 0.0299f
C6998 row_n[12] a_2275_14202# 19.2f
C6999 col_n[2] a_2475_5166# 0.0531f
C7000 rowon_n[4] a_23958_6146# 0.118f
C7001 m2_5172_2378# a_4974_2130# 0.165f
C7002 vcm a_17326_2170# 0.155f
C7003 a_2275_6170# a_30986_6146# 0.136f
C7004 a_15926_6146# a_16322_6186# 0.0313f
C7005 col[0] a_2874_16186# 0.0682f
C7006 m2_6752_946# m2_7756_946# 0.843f
C7007 m2_27260_10410# a_27062_10162# 0.165f
C7008 row_n[2] a_11302_4178# 0.0117f
C7009 vcm a_7986_11166# 0.56f
C7010 col[7] a_9902_18194# 0.0682f
C7011 VDD a_4882_1126# 0.405f
C7012 a_5886_15182# a_6378_15544# 0.0658f
C7013 a_4974_15182# a_5278_15222# 0.0931f
C7014 a_2275_15206# a_8990_15182# 0.399f
C7015 col_n[15] a_18026_12170# 0.251f
C7016 col[29] a_2275_11190# 0.0899f
C7017 col_n[12] a_14922_2130# 0.0765f
C7018 col_n[22] a_24962_14178# 0.0765f
C7019 a_12002_3134# a_13006_3134# 0.843f
C7020 a_2475_3158# a_23046_3134# 0.316f
C7021 rowoff_n[8] a_24962_10162# 0.202f
C7022 row_n[13] a_35002_15182# 0.0437f
C7023 vcm a_32386_6186# 0.155f
C7024 rowoff_n[11] a_28066_13174# 0.294f
C7025 col_n[28] row_n[11] 0.298f
C7026 col_n[29] rowon_n[11] 0.111f
C7027 col_n[13] rowon_n[3] 0.111f
C7028 col_n[10] row_n[2] 0.298f
C7029 col_n[6] row_n[0] 0.298f
C7030 col_n[30] row_n[12] 0.298f
C7031 col_n[14] row_n[4] 0.298f
C7032 col_n[7] rowon_n[0] 0.111f
C7033 col_n[16] row_n[5] 0.298f
C7034 col_n[12] row_n[3] 0.298f
C7035 col_n[26] row_n[10] 0.298f
C7036 col_n[18] row_n[6] 0.298f
C7037 col_n[3] ctop 0.0594f
C7038 col_n[15] rowon_n[4] 0.111f
C7039 col_n[24] row_n[9] 0.298f
C7040 col_n[25] rowon_n[9] 0.111f
C7041 col_n[19] rowon_n[6] 0.111f
C7042 vcm en_bit_n[2] 0.0193f
C7043 col_n[31] rowon_n[12] 0.111f
C7044 VDD col[0] 10.5f
C7045 col_n[22] row_n[8] 0.298f
C7046 col_n[11] rowon_n[2] 0.111f
C7047 rowon_n[14] row_n[14] 18.9f
C7048 col_n[27] rowon_n[10] 0.111f
C7049 col_n[23] rowon_n[8] 0.111f
C7050 col_n[20] row_n[7] 0.298f
C7051 col_n[21] rowon_n[7] 0.111f
C7052 col_n[9] rowon_n[1] 0.111f
C7053 col_n[17] rowon_n[5] 0.111f
C7054 col_n[8] row_n[1] 0.298f
C7055 col_n[0] a_2275_8178# 0.113f
C7056 vcm a_23046_15182# 0.56f
C7057 VDD a_19942_5142# 0.181f
C7058 row_n[12] rowoff_n[11] 0.085f
C7059 a_33086_1126# VDD 0.0352f
C7060 col_n[6] a_9390_10524# 0.0283f
C7061 a_2275_17214# a_24050_17190# 0.399f
C7062 rowoff_n[6] a_33998_8154# 0.202f
C7063 col_n[19] a_2475_7174# 0.0531f
C7064 m3_29976_1078# m3_30980_1078# 0.202f
C7065 m2_18224_8402# a_18026_8154# 0.165f
C7066 vcm a_13310_9198# 0.155f
C7067 a_32994_1126# a_33390_1166# 0.0313f
C7068 a_30986_10162# a_31382_10202# 0.0313f
C7069 vcm a_3970_18194# 0.165f
C7070 ctop a_26058_4138# 4.11f
C7071 a_2275_14202# a_14314_14218# 0.144f
C7072 a_2475_14202# a_16930_14178# 0.264f
C7073 row_n[7] a_22042_9158# 0.282f
C7074 VDD a_35002_9158# 0.258f
C7075 col[4] a_2475_15206# 0.136f
C7076 m2_1732_6970# m3_1864_8106# 0.0341f
C7077 rowon_n[11] a_21950_13174# 0.118f
C7078 col[9] a_2475_4162# 0.136f
C7079 VDD a_22346_18234# 0.019f
C7080 col_n[30] a_33390_11206# 0.084f
C7081 col_n[4] a_6982_10162# 0.251f
C7082 a_15926_2130# a_16418_2492# 0.0658f
C7083 a_15014_2130# a_15318_2170# 0.0931f
C7084 a_2275_2154# a_29070_2130# 0.399f
C7085 col_n[11] a_13918_12170# 0.0765f
C7086 m3_2868_18146# VDD 0.0853f
C7087 vcm a_6890_3134# 0.1f
C7088 row_n[9] a_9294_11206# 0.0117f
C7089 rowoff_n[9] a_34490_11528# 0.0133f
C7090 rowon_n[1] a_31990_3134# 0.118f
C7091 a_27062_7150# a_28066_7150# 0.843f
C7092 vcm a_28370_13214# 0.155f
C7093 a_2275_11190# a_7894_11166# 0.136f
C7094 col_n[23] rowoff_n[12] 0.0471f
C7095 col_n[16] a_2275_10186# 0.113f
C7096 VDD a_26458_3496# 0.0779f
C7097 m2_15788_18014# a_15926_18194# 0.225f
C7098 ctop a_6982_7150# 4.11f
C7099 a_2475_16210# a_31990_16186# 0.264f
C7100 a_2275_16210# a_29374_16226# 0.144f
C7101 a_16930_16186# a_17022_16186# 0.326f
C7102 VDD a_15926_12170# 0.181f
C7103 m2_6176_6394# rowon_n[4] 0.0322f
C7104 m2_11196_2378# rowon_n[0] 0.0322f
C7105 row_n[1] a_9902_3134# 0.0437f
C7106 col[1] a_2275_18218# 0.0899f
C7107 m2_9188_6394# a_8990_6146# 0.165f
C7108 col[24] a_27062_9158# 0.367f
C7109 vcm a_21950_7150# 0.1f
C7110 col[6] a_2275_7174# 0.0899f
C7111 rowon_n[5] a_8990_7150# 0.248f
C7112 a_18026_9158# a_18026_8154# 0.843f
C7113 rowoff_n[12] a_16018_14178# 0.294f
C7114 col[31] a_33998_11166# 0.0682f
C7115 vcm a_9294_16226# 0.155f
C7116 a_11910_13174# a_12306_13214# 0.0313f
C7117 a_2275_13198# a_22954_13174# 0.136f
C7118 VDD a_7382_6508# 0.0779f
C7119 ctop a_22042_11166# 4.11f
C7120 col[21] a_2475_17214# 0.136f
C7121 VDD a_30986_16186# 0.181f
C7122 col[26] a_2475_6170# 0.136f
C7123 col_n[19] a_22346_9198# 0.084f
C7124 m2_21236_15430# rowon_n[13] 0.0322f
C7125 a_30986_6146# a_31478_6508# 0.0658f
C7126 a_30074_6146# a_30378_6186# 0.0931f
C7127 m2_27260_11414# rowon_n[9] 0.0322f
C7128 m2_33284_7398# rowon_n[5] 0.0322f
C7129 vcm a_2161_10186# 0.0169f
C7130 col_n[7] rowoff_n[13] 0.0471f
C7131 a_7986_10162# a_8990_10162# 0.843f
C7132 a_2475_10186# a_15014_10162# 0.316f
C7133 row_n[14] a_20034_16186# 0.282f
C7134 m2_1732_16006# a_2966_16186# 0.843f
C7135 col[8] rowoff_n[7] 0.0901f
C7136 col_n[30] a_33486_3496# 0.0283f
C7137 col[4] rowoff_n[3] 0.0901f
C7138 col[6] rowoff_n[5] 0.0901f
C7139 col[7] rowoff_n[6] 0.0901f
C7140 col[9] rowoff_n[8] 0.0901f
C7141 col[10] rowoff_n[9] 0.0901f
C7142 col[2] rowoff_n[1] 0.0901f
C7143 col[1] rowoff_n[0] 0.0901f
C7144 col[5] rowoff_n[4] 0.0901f
C7145 col[3] rowoff_n[2] 0.0901f
C7146 VDD a_22442_10524# 0.0779f
C7147 row_n[4] a_30074_6146# 0.282f
C7148 a_26970_3134# a_27062_3134# 0.326f
C7149 rowon_n[8] a_29982_10162# 0.118f
C7150 rowoff_n[10] a_22442_12532# 0.0133f
C7151 rowoff_n[2] a_5374_4500# 0.0133f
C7152 a_2275_7174# a_5978_7150# 0.399f
C7153 m2_14784_18014# vcm 0.353f
C7154 col[23] a_2275_9182# 0.0899f
C7155 row_n[6] a_17326_8194# 0.0117f
C7156 vcm a_17934_14178# 0.1f
C7157 col[13] a_16018_7150# 0.367f
C7158 a_33086_13174# a_33086_12170# 0.843f
C7159 a_2475_12194# a_30074_12170# 0.316f
C7160 VDD a_14010_4138# 0.483f
C7161 col[20] a_22954_9158# 0.0682f
C7162 row_n[0] m2_27260_2378# 0.0128f
C7163 a_26970_17190# a_27366_17230# 0.0313f
C7164 VDD a_2966_13174# 0.485f
C7165 row_n[8] a_7894_10162# 0.0437f
C7166 col_n[28] a_31078_3134# 0.251f
C7167 rowoff_n[0] a_14410_2492# 0.0133f
C7168 rowon_n[12] a_6982_14178# 0.248f
C7169 m2_24824_946# ctop 0.0428f
C7170 a_2275_9182# a_21038_9158# 0.399f
C7171 a_10998_9158# a_11302_9198# 0.0931f
C7172 a_11910_9158# a_12402_9520# 0.0658f
C7173 col_n[8] a_11302_7190# 0.084f
C7174 rowoff_n[13] a_3970_15182# 0.294f
C7175 rowon_n[2] a_17022_4138# 0.248f
C7176 ctop rowoff_n[10] 0.177f
C7177 vcm a_32994_18194# 0.101f
C7178 col_n[8] a_2475_16210# 0.0531f
C7179 a_23046_14178# a_24050_14178# 0.843f
C7180 VDD a_29070_8154# 0.483f
C7181 rowoff_n[5] a_5978_7150# 0.294f
C7182 m2_1732_3958# m3_1864_5094# 0.0341f
C7183 col_n[13] a_2475_5166# 0.0531f
C7184 VDD a_18426_17552# 0.0779f
C7185 col_n[19] a_22442_1488# 0.0283f
C7186 col_n[29] a_32482_13536# 0.0283f
C7187 vcm a_35094_3134# 0.165f
C7188 a_2275_6170# a_11302_6186# 0.144f
C7189 a_7894_6146# a_7986_6146# 0.326f
C7190 a_2475_6170# a_13918_6146# 0.264f
C7191 rowoff_n[3] a_15014_5142# 0.294f
C7192 col[3] a_2475_2154# 0.136f
C7193 m2_34864_18014# a_35002_18194# 0.225f
C7194 m2_11772_18014# a_12002_17190# 0.843f
C7195 m2_5172_5390# row_n[3] 0.0128f
C7196 row_n[11] a_28066_13174# 0.282f
C7197 a_14010_16186# a_14010_15182# 0.843f
C7198 col[2] a_4974_5142# 0.367f
C7199 VDD a_9994_11166# 0.483f
C7200 col[12] a_15014_17190# 0.367f
C7201 rowon_n[15] a_27974_17190# 0.118f
C7202 col[9] a_11910_7150# 0.0682f
C7203 col_n[17] row_n[0] 0.297f
C7204 col_n[14] ctop 0.0597f
C7205 col_n[21] row_n[2] 0.298f
C7206 vcm col[8] 5.46f
C7207 col_n[18] rowon_n[0] 0.111f
C7208 col_n[4] col[4] 0.489f
C7209 col_n[31] row_n[7] 0.298f
C7210 col_n[19] row_n[1] 0.298f
C7211 col_n[28] rowon_n[5] 0.111f
C7212 col_n[30] rowon_n[6] 0.111f
C7213 VDD col[11] 3.83f
C7214 a_2275_3158# a_4882_3134# 0.136f
C7215 col_n[23] row_n[3] 0.298f
C7216 col_n[20] rowon_n[1] 0.111f
C7217 col_n[24] rowon_n[3] 0.111f
C7218 col_n[26] rowon_n[4] 0.111f
C7219 a_2966_3134# a_3970_3134# 0.843f
C7220 col_n[25] row_n[4] 0.298f
C7221 col_n[29] row_n[6] 0.298f
C7222 col_n[27] row_n[5] 0.298f
C7223 col_n[22] rowon_n[2] 0.111f
C7224 rowoff_n[1] a_24050_3134# 0.294f
C7225 col_n[17] a_20034_1126# 0.303f
C7226 col_n[10] a_2275_8178# 0.113f
C7227 row_n[13] a_15318_15222# 0.0117f
C7228 vcm a_16018_6146# 0.56f
C7229 rowoff_n[11] a_10394_13536# 0.0133f
C7230 col_n[27] a_30074_13174# 0.251f
C7231 a_2475_8178# a_28978_8154# 0.264f
C7232 a_2275_8178# a_26362_8194# 0.144f
C7233 col_n[24] a_26970_3134# 0.0765f
C7234 a_26058_13174# a_26362_13214# 0.0931f
C7235 a_26970_13174# a_27462_13536# 0.0658f
C7236 VDD a_35398_6186# 0.0882f
C7237 row_n[3] a_25358_5182# 0.0117f
C7238 col_n[7] a_10298_17230# 0.084f
C7239 row_n[15] a_5886_17190# 0.0437f
C7240 m2_20232_14426# row_n[12] 0.0128f
C7241 a_3970_17190# a_4974_17190# 0.843f
C7242 a_2475_17214# a_6982_17190# 0.316f
C7243 m2_26256_10410# row_n[8] 0.0128f
C7244 VDD a_25054_15182# 0.483f
C7245 col_n[30] a_2475_7174# 0.0531f
C7246 m2_32280_6394# row_n[4] 0.0128f
C7247 col[0] a_2275_5166# 0.099f
C7248 m3_15920_18146# a_16018_17190# 0.0303f
C7249 row_n[5] a_15926_7150# 0.0437f
C7250 a_2275_5166# a_19942_5142# 0.136f
C7251 m3_34996_5094# m3_34996_4090# 0.202f
C7252 col_n[18] a_21438_11528# 0.0283f
C7253 rowon_n[9] a_15014_11166# 0.248f
C7254 vcm a_31078_10162# 0.56f
C7255 a_22954_10162# a_23046_10162# 0.326f
C7256 rowoff_n[15] a_26458_17552# 0.0133f
C7257 col[15] a_2475_15206# 0.136f
C7258 col[20] a_2475_4162# 0.136f
C7259 m2_4744_946# a_2275_1150# 0.28f
C7260 rowon_n[11] a_3878_13174# 0.118f
C7261 m3_34996_12122# a_34090_12170# 0.0303f
C7262 VDD a_5978_18194# 0.0356f
C7263 a_2475_2154# a_12002_2130# 0.316f
C7264 a_24050_3134# a_24050_2130# 0.843f
C7265 col[1] a_3970_15182# 0.367f
C7266 vcm a_21342_4178# 0.155f
C7267 a_2275_7174# a_35002_7150# 0.136f
C7268 a_17934_7150# a_18330_7190# 0.0313f
C7269 col_n[27] a_2275_10186# 0.113f
C7270 rowoff_n[9] a_16930_11166# 0.202f
C7271 col[8] a_10906_17190# 0.0682f
C7272 m2_1732_15002# vcm 0.316f
C7273 vcm a_12002_13174# 0.56f
C7274 col_n[16] a_19030_11166# 0.251f
C7275 VDD a_8898_3134# 0.181f
C7276 m2_3740_18014# a_3878_18194# 0.225f
C7277 m2_5748_18014# a_2275_18218# 0.28f
C7278 col_n[13] a_15926_1126# 0.0765f
C7279 a_7894_16186# a_8386_16548# 0.0658f
C7280 a_6982_16186# a_7286_16226# 0.0931f
C7281 a_2275_16210# a_13006_16186# 0.399f
C7282 rowon_n[3] a_2161_5166# 0.0177f
C7283 col_n[23] a_25966_13174# 0.0765f
C7284 col[12] a_2275_18218# 0.0899f
C7285 rowoff_n[7] a_25966_9158# 0.202f
C7286 col[17] a_2275_7174# 0.0899f
C7287 a_2475_4162# a_27062_4138# 0.316f
C7288 a_14010_4138# a_15014_4138# 0.843f
C7289 m3_26964_1078# ctop 0.21f
C7290 vcm a_3878_7150# 0.1f
C7291 rowoff_n[13] a_32994_15182# 0.202f
C7292 row_n[10] a_23350_12210# 0.0117f
C7293 col_n[7] a_10394_9520# 0.0283f
C7294 ctop a_15014_2130# 4.06f
C7295 vcm a_27062_17190# 0.56f
C7296 a_2275_13198# a_3270_13214# 0.144f
C7297 a_2475_13198# a_5886_13174# 0.264f
C7298 VDD a_23958_7150# 0.181f
C7299 rowoff_n[5] a_35002_7150# 0.202f
C7300 m2_1732_18014# a_2475_18218# 0.139f
C7301 a_2275_18218# a_28066_18194# 0.0924f
C7302 row_n[0] a_33390_2170# 0.0117f
C7303 row_n[12] a_13918_14178# 0.0437f
C7304 a_2275_1150# a_18026_1126# 0.399f
C7305 col_n[18] rowoff_n[13] 0.0471f
C7306 vcm a_29982_2130# 0.1f
C7307 m2_34864_5966# m2_35292_6394# 0.165f
C7308 a_4974_6146# a_4974_5142# 0.843f
C7309 col_n[2] a_2475_14202# 0.0531f
C7310 m2_34864_9982# a_35398_10202# 0.087f
C7311 row_n[2] a_23958_4138# 0.0437f
C7312 vcm a_17326_11206# 0.155f
C7313 col_n[7] a_2475_3158# 0.0531f
C7314 col[15] rowoff_n[3] 0.0901f
C7315 col[19] rowoff_n[7] 0.0901f
C7316 col[21] rowoff_n[9] 0.0901f
C7317 col[18] rowoff_n[6] 0.0901f
C7318 a_32994_11166# a_33390_11206# 0.0313f
C7319 col[12] rowoff_n[0] 0.0901f
C7320 col[13] rowoff_n[1] 0.0901f
C7321 col[16] rowoff_n[4] 0.0901f
C7322 col[17] rowoff_n[5] 0.0901f
C7323 col[14] rowoff_n[2] 0.0901f
C7324 col[20] rowoff_n[8] 0.0901f
C7325 row_n[14] a_1957_16210# 0.187f
C7326 VDD a_15414_1488# 0.0977f
C7327 rowon_n[6] a_23046_8154# 0.248f
C7328 m2_23244_17438# a_23046_17190# 0.165f
C7329 m2_30848_18014# a_31078_17190# 0.843f
C7330 ctop a_30074_6146# 4.11f
C7331 a_2475_15206# a_20946_15182# 0.264f
C7332 a_2275_15206# a_18330_15222# 0.144f
C7333 VDD a_4882_10162# 0.181f
C7334 col_n[5] a_7986_9158# 0.251f
C7335 col_n[12] a_14922_11166# 0.0765f
C7336 a_17022_3134# a_17326_3174# 0.0931f
C7337 a_2275_3158# a_33086_3134# 0.399f
C7338 a_17934_3134# a_18426_3496# 0.0658f
C7339 a_2475_18218# a_26058_18194# 0.0299f
C7340 rowoff_n[8] a_35494_10524# 0.0133f
C7341 a_24354_1166# a_23958_1126# 0.0313f
C7342 vcm a_10906_5142# 0.1f
C7343 a_29070_8154# a_30074_8154# 0.843f
C7344 rowoff_n[10] a_4882_12170# 0.202f
C7345 a_24050_1126# vcm 0.165f
C7346 m2_16792_18014# col[14] 0.347f
C7347 vcm a_32386_15222# 0.155f
C7348 a_2275_12194# a_11910_12170# 0.136f
C7349 VDD a_30474_5504# 0.0779f
C7350 col_n[0] a_2275_17214# 0.113f
C7351 m2_18800_18014# VDD 1.1f
C7352 ctop a_10998_9158# 4.11f
C7353 row_n[15] a_34090_17190# 0.282f
C7354 a_2275_17214# a_33390_17230# 0.144f
C7355 a_18938_17190# a_19030_17190# 0.326f
C7356 col_n[4] a_2275_6170# 0.113f
C7357 VDD a_19942_14178# 0.181f
C7358 col_n[2] rowoff_n[14] 0.0471f
C7359 rowon_n[0] a_10906_2130# 0.118f
C7360 col[25] a_28066_8154# 0.367f
C7361 col[5] rowoff_n[10] 0.0901f
C7362 vcm a_25966_9158# 0.1f
C7363 col_n[19] a_2475_16210# 0.0531f
C7364 m2_8760_18014# m2_9188_18442# 0.165f
C7365 a_2475_9182# a_3970_9158# 0.316f
C7366 a_2275_9182# a_2966_9158# 0.399f
C7367 rowoff_n[14] a_20946_16186# 0.202f
C7368 a_20034_10162# a_20034_9158# 0.843f
C7369 col_n[24] a_2475_5166# 0.0531f
C7370 m2_14208_15430# a_14010_15182# 0.165f
C7371 vcm a_13310_18234# 0.16f
C7372 ctop a_2275_3158# 0.0683f
C7373 m2_22816_946# a_23046_1126# 0.0249f
C7374 a_13918_14178# a_14314_14218# 0.0313f
C7375 m3_34996_2082# a_34090_2130# 0.0303f
C7376 m2_4168_17438# rowon_n[15] 0.0322f
C7377 a_2275_14202# a_26970_14178# 0.136f
C7378 m2_10192_13422# rowon_n[11] 0.0322f
C7379 row_n[7] a_31382_9198# 0.0117f
C7380 VDD a_11398_8516# 0.0779f
C7381 m2_16216_9406# rowon_n[7] 0.0322f
C7382 m2_22240_5390# rowon_n[3] 0.0322f
C7383 m2_16792_946# vcm 0.353f
C7384 ctop a_26058_13174# 4.11f
C7385 VDD a_35002_18194# 0.419f
C7386 col_n[20] a_23350_8194# 0.084f
C7387 col[9] a_2475_13198# 0.136f
C7388 row_n[9] a_21950_11166# 0.0437f
C7389 a_32994_7150# a_33486_7512# 0.0658f
C7390 col[14] a_2475_2154# 0.136f
C7391 a_32082_7150# a_32386_7190# 0.0931f
C7392 m2_33284_11414# a_33086_11166# 0.165f
C7393 rowon_n[13] a_21038_15182# 0.248f
C7394 vcm a_6890_12170# 0.1f
C7395 a_2475_11190# a_19030_11166# 0.316f
C7396 a_9994_11166# a_10998_11166# 0.843f
C7397 VDD a_2874_2130# 0.182f
C7398 col_n[31] a_34490_2492# 0.0283f
C7399 rowon_n[3] a_31078_5142# 0.248f
C7400 VDD a_26458_12532# 0.0779f
C7401 vcm col[19] 5.46f
C7402 VDD col[22] 3.83f
C7403 col_n[9] col[10] 7.13f
C7404 col_n[31] rowon_n[1] 0.111f
C7405 col_n[30] row_n[1] 0.298f
C7406 col_n[28] row_n[0] 0.298f
C7407 col_n[29] rowon_n[0] 0.111f
C7408 col_n[25] ctop 0.0595f
C7409 m2_14784_18014# m3_14916_18146# 3.79f
C7410 m2_32856_18014# col_n[30] 0.243f
C7411 col_n[21] a_2275_8178# 0.113f
C7412 ctop a_6982_16186# 4.11f
C7413 a_28978_4138# a_29070_4138# 0.326f
C7414 rowoff_n[1] a_6378_3496# 0.0133f
C7415 a_2275_8178# a_9994_8154# 0.399f
C7416 col[14] a_17022_6146# 0.367f
C7417 m2_5172_13422# a_4974_13174# 0.165f
C7418 vcm a_21950_16186# 0.1f
C7419 col[6] a_2275_16210# 0.0899f
C7420 col[21] a_23958_8154# 0.0682f
C7421 a_2475_13198# a_34090_13174# 0.316f
C7422 VDD a_18026_6146# 0.483f
C7423 row_n[3] a_8990_5142# 0.282f
C7424 col[11] a_2275_5166# 0.0899f
C7425 rowon_n[7] a_8898_9158# 0.118f
C7426 a_28978_18194# a_29374_18234# 0.0313f
C7427 col_n[29] a_32082_2130# 0.251f
C7428 VDD a_7382_15544# 0.0779f
C7429 col[26] a_2475_15206# 0.136f
C7430 col_n[9] a_12306_6186# 0.084f
C7431 m3_25960_18146# m3_26964_18146# 0.202f
C7432 m2_24248_9406# a_24050_9158# 0.165f
C7433 col[31] a_2475_4162# 0.136f
C7434 col_n[19] a_22346_18234# 0.084f
C7435 rowoff_n[15] a_8898_17190# 0.202f
C7436 a_13006_10162# a_13310_10202# 0.0931f
C7437 a_2275_10186# a_25054_10162# 0.399f
C7438 a_13918_10162# a_14410_10524# 0.0658f
C7439 row_n[14] a_29374_16226# 0.0117f
C7440 rowoff_n[4] a_6982_6146# 0.294f
C7441 a_25054_15182# a_26058_15182# 0.843f
C7442 VDD a_33086_10162# 0.483f
C7443 col_n[30] a_33486_12532# 0.0283f
C7444 col_n[1] a_2475_1150# 0.0486f
C7445 m2_34864_3958# a_2475_4162# 0.282f
C7446 vcm a_4974_4138# 0.56f
C7447 rowoff_n[10] a_33086_12170# 0.294f
C7448 a_2275_7174# a_15318_7190# 0.144f
C7449 rowoff_n[2] a_16018_4138# 0.294f
C7450 a_9902_7150# a_9994_7150# 0.326f
C7451 a_2475_7174# a_17934_7150# 0.264f
C7452 row_n[6] a_29982_8154# 0.0437f
C7453 col[3] a_5978_4138# 0.367f
C7454 rowon_n[10] a_29070_12170# 0.248f
C7455 col[23] a_2275_18218# 0.0899f
C7456 col[13] a_16018_16186# 0.367f
C7457 col[28] a_2275_7174# 0.0899f
C7458 a_16018_17190# a_16018_16186# 0.843f
C7459 VDD a_14010_13174# 0.483f
C7460 col[10] a_12914_6146# 0.0682f
C7461 col[20] a_22954_18194# 0.0682f
C7462 rowoff_n[0] a_25054_2130# 0.294f
C7463 a_4882_4138# a_5278_4178# 0.0313f
C7464 a_2275_4162# a_8898_4138# 0.136f
C7465 m3_22948_18146# ctop 0.209f
C7466 col_n[28] a_31078_12170# 0.251f
C7467 m2_15212_7398# a_15014_7150# 0.165f
C7468 col_n[25] a_27974_2130# 0.0765f
C7469 m2_3164_16434# row_n[14] 0.0128f
C7470 m2_9188_12418# row_n[10] 0.0128f
C7471 vcm a_20034_8154# 0.56f
C7472 a_2275_9182# a_30378_9198# 0.144f
C7473 m2_15212_8402# row_n[6] 0.0128f
C7474 a_2475_9182# a_32994_9158# 0.264f
C7475 m2_1732_4962# rowoff_n[3] 0.415f
C7476 m2_21236_4386# row_n[2] 0.0128f
C7477 row_n[10] a_6982_12170# 0.282f
C7478 m2_1732_13998# a_2275_14202# 0.191f
C7479 col_n[8] a_11302_16226# 0.084f
C7480 a_28066_14178# a_28370_14218# 0.0931f
C7481 a_28978_14178# a_29470_14540# 0.0658f
C7482 rowon_n[14] a_6890_16186# 0.118f
C7483 col[1] a_3878_4138# 0.0682f
C7484 col_n[29] rowoff_n[13] 0.0471f
C7485 row_n[0] a_17022_2130# 0.282f
C7486 VDD a_29070_17190# 0.484f
C7487 col_n[13] a_2475_14202# 0.0531f
C7488 rowon_n[4] a_16930_6146# 0.118f
C7489 m2_34288_3382# a_34090_3134# 0.165f
C7490 col_n[18] a_2475_3158# 0.0531f
C7491 col[29] rowoff_n[6] 0.0901f
C7492 col[27] rowoff_n[4] 0.0901f
C7493 col[23] rowoff_n[0] 0.0901f
C7494 col[25] rowoff_n[2] 0.0901f
C7495 col[31] rowoff_n[8] 0.0901f
C7496 col[28] rowoff_n[5] 0.0901f
C7497 col[24] rowoff_n[1] 0.0901f
C7498 col_n[19] a_22442_10524# 0.0283f
C7499 col[30] rowoff_n[7] 0.0901f
C7500 vcm a_10298_2170# 0.155f
C7501 col[26] rowoff_n[3] 0.0901f
C7502 sample_n rowoff_n[9] 0.14f
C7503 a_2275_6170# a_23958_6146# 0.136f
C7504 row_n[2] a_4274_4178# 0.0117f
C7505 vcm a_35094_12170# 0.165f
C7506 col[9] a_2475_18218# 0.136f
C7507 a_24962_11166# a_25054_11166# 0.326f
C7508 VDD a_31990_2130# 0.181f
C7509 m2_30272_17438# row_n[15] 0.0128f
C7510 m2_35292_13422# row_n[11] 0.0128f
C7511 a_1957_15206# a_2161_15206# 0.115f
C7512 a_2475_15206# a_2275_15206# 2.76f
C7513 col[3] a_2475_11190# 0.136f
C7514 col[2] a_4974_14178# 0.367f
C7515 a_26058_4138# a_26058_3134# 0.843f
C7516 a_2475_3158# a_16018_3134# 0.316f
C7517 rowoff_n[8] a_17934_10162# 0.202f
C7518 col[9] a_11910_16186# 0.0682f
C7519 m2_6176_5390# a_5978_5142# 0.165f
C7520 a_29982_1126# a_2475_1150# 0.264f
C7521 a_27366_1166# a_2275_1150# 0.145f
C7522 row_n[13] a_27974_15182# 0.0437f
C7523 vcm a_25358_6186# 0.155f
C7524 rowoff_n[11] a_21038_13174# 0.294f
C7525 a_19942_8154# a_20338_8194# 0.0313f
C7526 col_n[10] a_2275_17214# 0.113f
C7527 col_n[17] a_20034_10162# 0.251f
C7528 vcm a_16018_15182# 0.56f
C7529 col_n[15] a_2275_6170# 0.113f
C7530 VDD a_12914_5142# 0.181f
C7531 col_n[24] a_26970_12170# 0.0765f
C7532 col_n[13] rowoff_n[14] 0.0471f
C7533 a_26058_1126# VDD 0.035f
C7534 a_9902_17190# a_10394_17552# 0.0658f
C7535 a_8990_17190# a_9294_17230# 0.0931f
C7536 a_2275_17214# a_17022_17190# 0.399f
C7537 rowoff_n[6] a_26970_8154# 0.202f
C7538 VDD a_35398_15222# 0.0882f
C7539 col[16] rowoff_n[10] 0.0901f
C7540 col_n[30] a_2475_16210# 0.0531f
C7541 col[0] a_2275_14202# 0.099f
C7542 a_16018_5142# a_17022_5142# 0.843f
C7543 a_2475_5166# a_31078_5142# 0.316f
C7544 m3_15920_1078# m3_16924_1078# 0.202f
C7545 col[5] a_2275_3158# 0.0899f
C7546 vcm a_6282_9198# 0.155f
C7547 col_n[8] a_11398_8516# 0.0283f
C7548 rowoff_n[14] a_2275_16210# 0.151f
C7549 m2_34864_16006# a_34090_16186# 0.843f
C7550 ctop a_19030_4138# 4.11f
C7551 m2_27836_946# a_2275_1150# 0.28f
C7552 m2_10768_946# a_10906_1126# 0.225f
C7553 a_2475_14202# a_9902_14178# 0.264f
C7554 a_5886_14178# a_5978_14178# 0.326f
C7555 a_2275_14202# a_7286_14218# 0.144f
C7556 row_n[7] a_15014_9158# 0.282f
C7557 VDD a_27974_9158# 0.181f
C7558 col[20] a_2475_13198# 0.136f
C7559 rowon_n[11] a_14922_13174# 0.118f
C7560 VDD a_15318_18234# 0.019f
C7561 col[25] a_2475_2154# 0.136f
C7562 a_2275_2154# a_22042_2130# 0.399f
C7563 m2_22240_1374# VDD 0.0194f
C7564 vcm a_33998_4138# 0.1f
C7565 row_n[9] a_3878_11166# 0.0437f
C7566 rowon_n[1] a_24962_3134# 0.118f
C7567 a_6982_7150# a_6982_6146# 0.843f
C7568 rowoff_n[9] a_27462_11528# 0.0133f
C7569 rowon_n[13] a_2966_15182# 0.248f
C7570 vcm a_21342_13214# 0.155f
C7571 sample sample_n 11.3f
C7572 rowon_n[6] rowon_n[5] 0.0632f
C7573 vcm col[30] 5.46f
C7574 col_n[15] col[15] 0.413f
C7575 VDD a_19430_3496# 0.0779f
C7576 VDD rowoff_n[15] 1.51f
C7577 col_n[31] analog_in 0.134f
C7578 rowon_n[13] ctop 0.203f
C7579 m2_10768_18014# a_10998_18194# 0.0249f
C7580 col_n[6] a_8990_8154# 0.251f
C7581 ctop a_34090_8154# 4.06f
C7582 a_2475_16210# a_24962_16186# 0.264f
C7583 a_2275_16210# a_22346_16226# 0.144f
C7584 VDD a_8898_12170# 0.181f
C7585 a_29374_1166# m2_28840_946# 0.087f
C7586 col_n[13] a_15926_10162# 0.0765f
C7587 col[0] rowoff_n[11] 0.0901f
C7588 a_19942_4138# a_20434_4500# 0.0658f
C7589 a_19030_4138# a_19334_4178# 0.0931f
C7590 row_n[1] a_2161_3158# 0.0221f
C7591 col[17] a_2275_16210# 0.0899f
C7592 rowon_n[5] a_2475_7174# 0.31f
C7593 vcm a_14922_7150# 0.1f
C7594 a_31078_9158# a_32082_9158# 0.843f
C7595 rowoff_n[12] a_8990_14178# 0.294f
C7596 col[22] a_2275_5166# 0.0899f
C7597 row_n[10] a_34394_12210# 0.0117f
C7598 vcm a_3878_16186# 0.1f
C7599 a_2275_13198# a_15926_13174# 0.136f
C7600 rowon_n[14] a_35094_16186# 0.0141f
C7601 VDD a_34490_7512# 0.0779f
C7602 ctop a_15014_11166# 4.11f
C7603 col_n[7] a_10394_18556# 0.0283f
C7604 a_20946_18194# a_21038_18194# 0.0991f
C7605 VDD a_23958_16186# 0.181f
C7606 a_15926_1126# a_16018_1126# 0.0991f
C7607 col[26] a_29070_7150# 0.367f
C7608 m2_5172_7398# rowon_n[5] 0.0322f
C7609 m2_29844_946# m2_30848_946# 0.843f
C7610 m2_11196_3382# rowon_n[1] 0.0322f
C7611 vcm a_29982_11166# 0.1f
C7612 a_2475_10186# a_7986_10162# 0.316f
C7613 a_22042_11166# a_22042_10162# 0.843f
C7614 row_n[14] a_13006_16186# 0.282f
C7615 col_n[7] a_2475_12194# 0.0531f
C7616 a_15926_15182# a_16322_15222# 0.0313f
C7617 a_2275_15206# a_30986_15182# 0.136f
C7618 VDD a_15414_10524# 0.0779f
C7619 col_n[12] a_2475_1150# 0.0531f
C7620 col_n[21] a_24354_7190# 0.084f
C7621 ctop a_30074_15182# 4.11f
C7622 row_n[4] a_23046_6146# 0.282f
C7623 rowon_n[8] a_22954_10162# 0.118f
C7624 col_n[2] a_4882_8154# 0.0765f
C7625 a_35002_8154# a_35494_8516# 0.0658f
C7626 rowoff_n[10] a_15414_12532# 0.0133f
C7627 a_35398_1166# vcm 0.161f
C7628 a_28978_1126# col_n[26] 0.0777f
C7629 m2_20232_16434# rowon_n[14] 0.0322f
C7630 m2_26256_12418# rowon_n[10] 0.0322f
C7631 row_n[6] a_10298_8194# 0.0117f
C7632 m2_32280_8402# rowon_n[6] 0.0322f
C7633 vcm a_10906_14178# 0.1f
C7634 a_2475_12194# a_23046_12170# 0.316f
C7635 a_12002_12170# a_13006_12170# 0.843f
C7636 VDD a_6982_4138# 0.483f
C7637 VDD a_30474_14540# 0.0779f
C7638 m2_33860_946# col[31] 0.274f
C7639 rowoff_n[0] a_7382_2492# 0.0133f
C7640 col_n[4] a_2275_15206# 0.113f
C7641 a_30986_5142# a_31078_5142# 0.326f
C7642 col[15] a_18026_5142# 0.367f
C7643 col_n[9] a_2275_4162# 0.113f
C7644 vcm a_1957_8178# 0.139f
C7645 col[25] a_28066_17190# 0.367f
C7646 rowoff_n[14] a_31478_16548# 0.0133f
C7647 a_2275_9182# a_14010_9158# 0.399f
C7648 col[22] a_24962_7150# 0.0682f
C7649 rowon_n[2] a_9994_4138# 0.248f
C7650 vcm a_25966_18194# 0.101f
C7651 VDD a_22042_8154# 0.483f
C7652 col_n[24] a_2475_14202# 0.0531f
C7653 ctop a_2275_12194# 0.0683f
C7654 col_n[29] a_2475_3158# 0.0531f
C7655 VDD a_11398_17552# 0.0779f
C7656 analog_in a_2275_1150# 0.0504f
C7657 a_25966_2130# a_26362_2170# 0.0313f
C7658 col_n[10] a_13310_5182# 0.084f
C7659 m3_21944_1078# VDD 0.0157f
C7660 vcm a_28066_3134# 0.56f
C7661 col[20] a_2475_18218# 0.136f
C7662 col_n[20] a_23350_17230# 0.084f
C7663 a_2275_6170# a_4274_6186# 0.144f
C7664 a_2475_6170# a_6890_6146# 0.264f
C7665 rowoff_n[3] a_7986_5142# 0.294f
C7666 a_15014_11166# a_15318_11206# 0.0931f
C7667 a_2275_11190# a_29070_11166# 0.399f
C7668 a_15926_11166# a_16418_11528# 0.0658f
C7669 col[14] a_2475_11190# 0.136f
C7670 m2_29844_18014# a_30074_18194# 0.0249f
C7671 a_27062_16186# a_28066_16186# 0.843f
C7672 row_n[11] a_21038_13174# 0.282f
C7673 VDD a_2874_11166# 0.182f
C7674 col_n[31] a_34490_11528# 0.0283f
C7675 m2_28840_18014# m3_29976_18146# 0.0341f
C7676 rowon_n[15] a_20946_17190# 0.118f
C7677 row_n[1] a_31078_3134# 0.282f
C7678 rowoff_n[1] a_17022_3134# 0.294f
C7679 col_n[21] a_2275_17214# 0.113f
C7680 row_n[13] a_8290_15222# 0.0117f
C7681 vcm a_8990_6146# 0.56f
C7682 col_n[26] a_2275_6170# 0.113f
C7683 rowon_n[5] a_30986_7150# 0.118f
C7684 a_2275_8178# a_19334_8194# 0.144f
C7685 a_2475_8178# a_21950_8154# 0.264f
C7686 a_11910_8154# a_12002_8154# 0.326f
C7687 rowoff_n[11] a_2966_13174# 0.294f
C7688 col[4] a_6982_3134# 0.367f
C7689 col_n[24] rowoff_n[14] 0.0471f
C7690 col[14] a_17022_15182# 0.367f
C7691 row_n[3] a_18330_5182# 0.0117f
C7692 col[11] a_13918_5142# 0.0682f
C7693 col[27] rowoff_n[10] 0.0901f
C7694 col[21] a_23958_17190# 0.0682f
C7695 VDD a_18026_15182# 0.483f
C7696 col[11] a_2275_14202# 0.0899f
C7697 m2_4168_6394# row_n[4] 0.0128f
C7698 m2_9188_2378# row_n[0] 0.0128f
C7699 col_n[29] a_32082_11166# 0.251f
C7700 col[16] a_2275_3158# 0.0899f
C7701 a_2275_5166# a_12914_5142# 0.136f
C7702 row_n[5] a_8898_7150# 0.0437f
C7703 a_6890_5142# a_7286_5182# 0.0313f
C7704 m3_34996_12122# m3_34996_11118# 0.202f
C7705 m2_32856_946# m3_32988_1078# 3.79f
C7706 rowon_n[9] a_7986_11166# 0.248f
C7707 vcm a_24050_10162# 0.56f
C7708 a_2275_10186# a_35398_10202# 0.145f
C7709 rowoff_n[15] a_19430_17552# 0.0133f
C7710 col_n[9] a_12306_15222# 0.084f
C7711 m2_20232_16434# a_20034_16186# 0.165f
C7712 col[31] a_2475_13198# 0.136f
C7713 a_30986_15182# a_31478_15544# 0.0658f
C7714 a_30074_15182# a_30378_15222# 0.0931f
C7715 m2_21812_946# a_22042_2130# 0.843f
C7716 m2_28840_18014# ctop 0.0422f
C7717 m2_19228_15430# row_n[13] 0.0128f
C7718 col_n[20] a_23446_9520# 0.0283f
C7719 a_2475_2154# a_4974_2130# 0.316f
C7720 m2_25252_11414# row_n[9] 0.0128f
C7721 m2_31276_7398# row_n[5] 0.0128f
C7722 vcm a_14314_4178# 0.155f
C7723 a_2275_7174# a_27974_7150# 0.136f
C7724 rowon_n[14] col[7] 0.0323f
C7725 row_n[12] col[2] 0.0342f
C7726 row_n[13] col[4] 0.0342f
C7727 rowon_n[12] col[3] 0.0323f
C7728 rowon_n[13] col[5] 0.0323f
C7729 rowon_n[11] col[1] 0.0323f
C7730 rowon_n[15] col[9] 0.0323f
C7731 col_n[20] col[21] 7.13f
C7732 col_n[1] a_2475_10186# 0.0531f
C7733 rowoff_n[9] a_9902_11166# 0.202f
C7734 row_n[8] ctop 0.186f
C7735 col_n[8] rowoff_n[15] 0.0471f
C7736 row_n[15] col[8] 0.0342f
C7737 rowon_n[3] row_n[3] 18.9f
C7738 row_n[14] col[6] 0.0342f
C7739 row_n[11] col[0] 0.0322f
C7740 vcm a_4974_13174# 0.56f
C7741 a_26970_12170# a_27062_12170# 0.326f
C7742 col[11] rowoff_n[11] 0.0901f
C7743 a_2275_16210# a_5978_16186# 0.399f
C7744 col[3] a_5978_13174# 0.367f
C7745 row_n[8] a_29070_10162# 0.282f
C7746 rowoff_n[7] a_18938_9158# 0.202f
C7747 col[28] a_2275_16210# 0.0899f
C7748 col[10] a_12914_15182# 0.0682f
C7749 rowon_n[12] a_28978_14178# 0.118f
C7750 a_28066_5142# a_28066_4138# 0.843f
C7751 a_2475_4162# a_20034_4138# 0.316f
C7752 col_n[18] a_21038_9158# 0.251f
C7753 vcm a_29374_8194# 0.155f
C7754 a_21950_9158# a_22346_9198# 0.0313f
C7755 rowoff_n[13] a_25966_15182# 0.202f
C7756 row_n[10] a_16322_12210# 0.0117f
C7757 m2_11196_14426# a_10998_14178# 0.165f
C7758 col_n[25] a_27974_11166# 0.0765f
C7759 ctop a_7986_2130# 4.06f
C7760 vcm a_20034_17190# 0.56f
C7761 VDD a_16930_7150# 0.181f
C7762 rowoff_n[5] a_27974_7150# 0.202f
C7763 col_n[3] a_2275_2154# 0.113f
C7764 a_2275_18218# a_21038_18194# 0.0924f
C7765 a_11910_18194# a_12402_18556# 0.0658f
C7766 row_n[0] a_26362_2170# 0.0117f
C7767 a_6890_1126# a_7382_1488# 0.0658f
C7768 row_n[12] a_6890_14178# 0.0437f
C7769 a_2275_1150# a_10998_1126# 0.0924f
C7770 col[1] a_3878_13174# 0.0682f
C7771 m2_8184_2378# a_7986_2130# 0.165f
C7772 vcm a_22954_2130# 0.1f
C7773 a_2475_6170# a_35094_6146# 0.0299f
C7774 a_18026_6146# a_19030_6146# 0.843f
C7775 col_n[9] a_12402_7512# 0.0283f
C7776 m2_10768_946# m2_11196_1374# 0.165f
C7777 m2_30272_10410# a_30074_10162# 0.165f
C7778 col_n[18] a_2475_12194# 0.0531f
C7779 vcm a_10298_11206# 0.155f
C7780 row_n[2] a_16930_4138# 0.0437f
C7781 VDD a_8386_1488# 0.0977f
C7782 col_n[23] a_2475_1150# 0.0531f
C7783 rowon_n[6] a_16018_8154# 0.248f
C7784 ctop a_23046_6146# 4.11f
C7785 a_2275_15206# a_11302_15222# 0.144f
C7786 a_7894_15182# a_7986_15182# 0.326f
C7787 a_2475_15206# a_13918_15182# 0.264f
C7788 VDD a_31990_11166# 0.181f
C7789 a_2475_18218# a_19030_18194# 0.0299f
C7790 a_2275_3158# a_26058_3134# 0.399f
C7791 rowoff_n[8] a_28466_10524# 0.0133f
C7792 col[8] a_2475_9182# 0.136f
C7793 a_8990_8154# a_8990_7150# 0.843f
C7794 m2_1732_11990# a_1957_12194# 0.245f
C7795 col_n[7] a_9994_7150# 0.251f
C7796 vcm a_25358_15222# 0.155f
C7797 a_2966_12170# a_3970_12170# 0.843f
C7798 a_2275_12194# a_4882_12170# 0.136f
C7799 VDD a_23446_5504# 0.0779f
C7800 m2_4744_18014# VDD 0.993f
C7801 col_n[14] a_16930_9158# 0.0765f
C7802 row_n[15] a_27062_17190# 0.282f
C7803 ctop a_3970_9158# 4.11f
C7804 a_2275_17214# a_26362_17230# 0.144f
C7805 a_2475_17214# a_28978_17190# 0.264f
C7806 col_n[15] a_2275_15206# 0.113f
C7807 VDD a_12914_14178# 0.181f
C7808 col_n[20] a_2275_4162# 0.113f
C7809 a_21038_5142# a_21342_5182# 0.0931f
C7810 a_21950_5142# a_22442_5504# 0.0658f
C7811 m2_21236_8402# a_21038_8154# 0.165f
C7812 vcm a_18938_9158# 0.1f
C7813 m2_1732_18014# m2_2160_18442# 0.165f
C7814 a_33086_10162# a_34090_10162# 0.843f
C7815 rowoff_n[14] a_13918_16186# 0.202f
C7816 col[5] a_2275_12194# 0.0899f
C7817 vcm a_6282_18234# 0.16f
C7818 col_n[8] a_11398_17552# 0.0283f
C7819 a_2275_14202# a_19942_14178# 0.136f
C7820 row_n[7] a_24354_9198# 0.0117f
C7821 VDD a_4370_8516# 0.0779f
C7822 col[10] a_2275_1150# 0.0899f
C7823 col_n[31] a_34394_8194# 0.084f
C7824 col[27] a_30074_6146# 0.367f
C7825 ctop a_19030_13174# 4.11f
C7826 col[31] a_2475_18218# 0.136f
C7827 VDD a_27974_18194# 0.343f
C7828 a_17934_2130# a_18026_2130# 0.326f
C7829 a_2275_2154# a_31382_2170# 0.144f
C7830 a_2475_2154# a_33998_2130# 0.264f
C7831 m3_17928_18146# VDD 0.0313f
C7832 row_n[9] a_14922_11166# 0.0437f
C7833 col[25] a_2475_11190# 0.136f
C7834 rowon_n[13] a_14010_15182# 0.248f
C7835 vcm a_33998_13174# 0.1f
C7836 a_2475_11190# a_12002_11166# 0.316f
C7837 a_24050_12170# a_24050_11166# 0.843f
C7838 VDD a_30074_3134# 0.483f
C7839 m2_16792_18014# a_17326_18234# 0.087f
C7840 row_n[11] a_2966_13174# 0.281f
C7841 col_n[22] a_25358_6186# 0.084f
C7842 a_17934_16186# a_18330_16226# 0.0313f
C7843 a_2275_16210# a_35002_16186# 0.136f
C7844 rowon_n[3] a_24050_5142# 0.248f
C7845 VDD a_19430_12532# 0.0779f
C7846 m2_5748_18014# m3_4876_18146# 0.0341f
C7847 rowon_n[15] a_2275_17214# 1.79f
C7848 col_n[6] a_8990_17190# 0.251f
C7849 ctop a_34090_17190# 4.02f
C7850 m2_9188_14426# rowon_n[12] 0.0322f
C7851 col_n[3] a_5886_7150# 0.0765f
C7852 m2_15212_10410# rowon_n[8] 0.0322f
C7853 m2_21236_6394# rowon_n[4] 0.0322f
C7854 row_n[14] rowoff_n[14] 0.209f
C7855 m2_12200_6394# a_12002_6146# 0.165f
C7856 a_2275_8178# a_2874_8154# 0.136f
C7857 a_2475_8178# a_3878_8154# 0.264f
C7858 vcm a_14922_16186# 0.1f
C7859 a_14010_13174# a_15014_13174# 0.843f
C7860 a_2475_13198# a_27062_13174# 0.316f
C7861 VDD a_10998_6146# 0.483f
C7862 col[22] a_2275_14202# 0.0899f
C7863 row_n[3] a_2475_5166# 0.405f
C7864 col[27] a_2275_3158# 0.0899f
C7865 VDD a_34490_16548# 0.0779f
C7866 row_n[12] a_35094_14178# 0.0123f
C7867 col[16] a_19030_4138# 0.367f
C7868 vcm a_17022_1126# 0.165f
C7869 m2_35292_15430# rowon_n[13] 0.0322f
C7870 a_32994_6146# a_33086_6146# 0.326f
C7871 col[26] a_29070_16186# 0.367f
C7872 m3_11904_18146# m3_12908_18146# 0.202f
C7873 m2_7756_946# m3_8892_1078# 0.0341f
C7874 col[23] a_25966_6146# 0.0682f
C7875 a_2275_10186# a_18026_10162# 0.399f
C7876 row_n[14] a_22346_16226# 0.0117f
C7877 a_4974_15182# a_4974_14178# 0.843f
C7878 VDD a_26058_10162# 0.483f
C7879 m2_1732_1950# col[0] 0.0137f
C7880 row_n[4] a_32386_6186# 0.0117f
C7881 col_n[11] a_14314_4178# 0.084f
C7882 rowon_n[9] col[8] 0.0323f
C7883 row_n[11] col[11] 0.0342f
C7884 rowon_n[8] col[6] 0.0323f
C7885 row_n[13] col[15] 0.0342f
C7886 row_n[10] col[9] 0.0342f
C7887 rowon_n[13] col[16] 0.0323f
C7888 col_n[19] rowoff_n[15] 0.0471f
C7889 row_n[8] col[5] 0.0342f
C7890 rowon_n[5] col[0] 0.0318f
C7891 row_n[14] col[17] 0.0342f
C7892 rowon_n[10] col[10] 0.0323f
C7893 rowon_n[12] col[14] 0.0323f
C7894 row_n[6] col[1] 0.0342f
C7895 rowon_n[11] col[12] 0.0323f
C7896 rowon_n[2] ctop 0.203f
C7897 col_n[12] a_2475_10186# 0.0531f
C7898 rowon_n[7] col[4] 0.0323f
C7899 col_n[26] col[26] 0.542f
C7900 rowon_n[14] col[18] 0.0323f
C7901 rowon_n[6] col[2] 0.0323f
C7902 row_n[15] col[19] 0.0342f
C7903 row_n[9] col[7] 0.0342f
C7904 row_n[7] col[3] 0.0342f
C7905 rowon_n[15] col[20] 0.0323f
C7906 row_n[12] col[13] 0.0342f
C7907 a_27974_3134# a_28370_3174# 0.0313f
C7908 col_n[21] a_24354_16226# 0.084f
C7909 vcm a_32082_5142# 0.56f
C7910 a_2275_7174# a_8290_7190# 0.144f
C7911 a_2475_7174# a_10906_7150# 0.264f
C7912 rowoff_n[2] a_8990_4138# 0.294f
C7913 rowoff_n[10] a_26058_12170# 0.294f
C7914 col_n[2] a_4882_17190# 0.0765f
C7915 col[22] rowoff_n[11] 0.0901f
C7916 row_n[6] a_22954_8154# 0.0437f
C7917 a_17022_12170# a_17326_12210# 0.0931f
C7918 a_2275_12194# a_33086_12170# 0.399f
C7919 a_17934_12170# a_18426_12532# 0.0658f
C7920 rowon_n[10] a_22042_12170# 0.248f
C7921 col[2] a_2475_7174# 0.136f
C7922 a_29070_17190# a_30074_17190# 0.843f
C7923 VDD a_6982_13174# 0.483f
C7924 rowon_n[0] a_32082_2130# 0.248f
C7925 rowoff_n[0] a_18026_2130# 0.294f
C7926 a_2475_4162# a_1957_4162# 0.0734f
C7927 col[5] a_7986_2130# 0.367f
C7928 vcm a_13006_8154# 0.56f
C7929 a_2275_9182# a_23350_9198# 0.144f
C7930 a_13918_9158# a_14010_9158# 0.326f
C7931 a_2475_9182# a_25966_9158# 0.264f
C7932 col[15] a_18026_14178# 0.367f
C7933 col_n[9] a_2275_13198# 0.113f
C7934 col[12] a_14922_4138# 0.0682f
C7935 vcm a_1957_17214# 0.139f
C7936 col_n[14] a_2275_2154# 0.113f
C7937 m2_34864_11990# ctop 0.0422f
C7938 col[22] a_24962_16186# 0.0682f
C7939 a_2275_18218# a_2966_18194# 0.0924f
C7940 row_n[0] a_9994_2130# 0.282f
C7941 VDD a_22042_17190# 0.484f
C7942 col_n[30] a_33086_10162# 0.251f
C7943 rowon_n[4] a_9902_6146# 0.118f
C7944 col_n[29] a_2475_12194# 0.0531f
C7945 col[6] rowoff_n[12] 0.0901f
C7946 vcm a_3270_2170# 0.16f
C7947 a_8898_6146# a_9294_6186# 0.0313f
C7948 a_2275_6170# a_16930_6146# 0.136f
C7949 col_n[10] a_13310_14218# 0.084f
C7950 vcm a_28066_12170# 0.56f
C7951 VDD a_24962_2130# 0.181f
C7952 m2_2160_17438# row_n[15] 0.0194f
C7953 m2_8184_13422# row_n[11] 0.0128f
C7954 m2_3164_17438# a_2966_17190# 0.165f
C7955 m2_14208_9406# row_n[7] 0.0128f
C7956 m2_20232_5390# row_n[3] 0.0128f
C7957 row_n[11] a_30378_13214# 0.0117f
C7958 a_32994_16186# a_33486_16548# 0.0658f
C7959 a_32082_16186# a_32386_16226# 0.0931f
C7960 m2_1732_946# m2_2160_1374# 0.165f
C7961 col[19] a_2475_9182# 0.136f
C7962 col_n[21] a_24450_8516# 0.0283f
C7963 a_4974_3134# a_5978_3134# 0.843f
C7964 a_2475_3158# a_8990_3134# 0.316f
C7965 rowoff_n[8] a_10906_10162# 0.202f
C7966 row_n[13] a_20946_15182# 0.0437f
C7967 vcm a_18330_6186# 0.155f
C7968 a_2275_8178# a_31990_8154# 0.136f
C7969 rowoff_n[11] a_14010_13174# 0.294f
C7970 sample a_2161_2154# 0.0858f
C7971 vcm a_8990_15182# 0.56f
C7972 col_n[26] a_2275_15206# 0.113f
C7973 m3_2868_1078# m2_1732_946# 0.0341f
C7974 a_28978_13174# a_29070_13174# 0.326f
C7975 VDD a_5886_5142# 0.181f
C7976 row_n[3] a_30986_5142# 0.0437f
C7977 col_n[31] a_2275_4162# 0.113f
C7978 col[4] a_6982_12170# 0.367f
C7979 a_2275_17214# a_9994_17190# 0.399f
C7980 m2_34864_13998# row_n[12] 0.267f
C7981 rowon_n[7] a_30074_9158# 0.248f
C7982 rowoff_n[6] a_19942_8154# 0.202f
C7983 col[11] a_13918_14178# 0.0682f
C7984 m3_18932_18146# a_19030_17190# 0.0303f
C7985 col_n[19] a_22042_8154# 0.251f
C7986 a_30074_6146# a_30074_5142# 0.843f
C7987 a_2475_5166# a_24050_5142# 0.316f
C7988 m3_1864_1078# m3_2868_1078# 0.202f
C7989 col[16] a_2275_12194# 0.0899f
C7990 vcm a_33390_10202# 0.155f
C7991 col_n[26] a_28978_10162# 0.0765f
C7992 a_23958_10162# a_24354_10202# 0.0313f
C7993 col[21] a_2275_1150# 0.0899f
C7994 rowoff_n[15] a_30074_17190# 0.294f
C7995 rowoff_n[4] a_28978_6146# 0.202f
C7996 ctop a_12002_4138# 4.11f
C7997 m2_5748_946# a_5978_1126# 0.0249f
C7998 m2_13780_946# a_2475_1150# 0.286f
C7999 VDD a_20946_9158# 0.181f
C8000 row_n[7] a_7986_9158# 0.282f
C8001 rowon_n[11] a_7894_13174# 0.118f
C8002 VDD a_8290_18234# 0.019f
C8003 a_2275_2154# a_15014_2130# 0.399f
C8004 a_7986_2130# a_8290_2170# 0.0931f
C8005 a_8898_2130# a_9390_2492# 0.0658f
C8006 col_n[10] a_13406_6508# 0.0283f
C8007 m2_6752_946# VDD 1f
C8008 vcm a_26970_4138# 0.1f
C8009 m2_1732_8978# m2_2160_9406# 0.165f
C8010 rowoff_n[9] a_20434_11528# 0.0133f
C8011 rowon_n[1] a_17934_3134# 0.118f
C8012 a_20034_7150# a_21038_7150# 0.843f
C8013 col_n[20] a_23446_18556# 0.0283f
C8014 vcm a_14314_13214# 0.155f
C8015 VDD a_12402_3496# 0.0779f
C8016 col_n[6] a_2475_8178# 0.0531f
C8017 ctop a_27062_8154# 4.11f
C8018 a_2275_16210# a_15318_16226# 0.144f
C8019 a_2475_16210# a_17934_16186# 0.264f
C8020 a_9902_16186# a_9994_16186# 0.326f
C8021 rowoff_n[7] a_29470_9520# 0.0133f
C8022 a_2275_4162# a_30074_4138# 0.399f
C8023 vcm a_7894_7150# 0.1f
C8024 col_n[8] a_10998_6146# 0.251f
C8025 a_10998_9158# a_10998_8154# 0.843f
C8026 rowoff_n[12] a_2475_14202# 3.9f
C8027 row_n[10] a_28978_12170# 0.0437f
C8028 vcm a_29374_17230# 0.155f
C8029 rowon_n[14] a_28066_16186# 0.248f
C8030 a_2275_13198# a_8898_13174# 0.136f
C8031 a_4882_13174# a_5278_13214# 0.0313f
C8032 col_n[15] a_17934_8154# 0.0765f
C8033 VDD a_27462_7512# 0.0779f
C8034 ctop a_7986_11166# 4.11f
C8035 a_2275_18218# a_30378_18234# 0.145f
C8036 VDD a_16930_16186# 0.181f
C8037 a_2275_1150# a_20338_1166# 0.126f
C8038 a_2475_1150# a_22954_1126# 0.264f
C8039 col_n[3] a_2275_11190# 0.113f
C8040 a_23958_6146# a_24450_6508# 0.0658f
C8041 a_23046_6146# a_23350_6186# 0.0931f
C8042 m2_22816_946# m2_23820_946# 0.843f
C8043 vcm a_22954_11166# 0.1f
C8044 col_n[9] a_12402_16548# 0.0283f
C8045 row_n[14] a_5978_16186# 0.282f
C8046 VDD a_19030_1126# 0.992f
C8047 m2_26256_17438# a_26058_17190# 0.165f
C8048 col[28] a_31078_5142# 0.367f
C8049 a_2275_15206# a_23958_15182# 0.136f
C8050 row_n[15] col[30] 0.0342f
C8051 row_n[3] col[6] 0.0342f
C8052 rowon_n[3] col[7] 0.0323f
C8053 row_n[6] col[12] 0.0342f
C8054 rowon_n[11] col[23] 0.0323f
C8055 row_n[8] col[16] 0.0342f
C8056 rowon_n[0] col[1] 0.0323f
C8057 rowon_n[15] col[31] 0.0323f
C8058 row_n[9] col[18] 0.0342f
C8059 col_n[30] rowoff_n[15] 0.0471f
C8060 rowon_n[5] col[11] 0.0323f
C8061 rowon_n[8] col[17] 0.0323f
C8062 rowon_n[7] col[15] 0.0323f
C8063 row_n[5] col[10] 0.0342f
C8064 row_n[0] col[0] 0.0322f
C8065 rowon_n[12] col[25] 0.0323f
C8066 rowon_n[6] col[13] 0.0323f
C8067 row_n[4] col[8] 0.0342f
C8068 row_n[1] col[2] 0.0342f
C8069 sw analog_in 0.905f
C8070 row_n[14] col[28] 0.0342f
C8071 rowon_n[13] col[27] 0.0323f
C8072 row_n[2] col[4] 0.0342f
C8073 row_n[11] col[22] 0.0342f
C8074 rowon_n[14] col[29] 0.0323f
C8075 rowon_n[10] col[21] 0.0323f
C8076 rowon_n[2] col[5] 0.0323f
C8077 row_n[10] col[20] 0.0342f
C8078 rowon_n[1] col[3] 0.0323f
C8079 row_n[7] col[14] 0.0342f
C8080 row_n[12] col[24] 0.0342f
C8081 row_n[13] col[26] 0.0342f
C8082 rowon_n[9] col[19] 0.0323f
C8083 rowon_n[4] col[9] 0.0323f
C8084 col_n[23] a_2475_10186# 0.0531f
C8085 VDD a_8386_10524# 0.0779f
C8086 ctop a_23046_15182# 4.11f
C8087 row_n[4] a_16018_6146# 0.282f
C8088 a_19942_3134# a_20034_3134# 0.326f
C8089 rowon_n[8] a_15926_10162# 0.118f
C8090 a_2275_3158# a_2275_2154# 0.0715f
C8091 m2_34864_12994# m2_34864_11990# 0.843f
C8092 rowoff_n[10] a_8386_12532# 0.0133f
C8093 a_26362_1166# vcm 0.16f
C8094 row_n[6] a_3270_8194# 0.0117f
C8095 m2_4168_8402# rowon_n[6] 0.0322f
C8096 col[13] a_2475_7174# 0.136f
C8097 a_26058_13174# a_26058_12170# 0.843f
C8098 m2_10192_4386# rowon_n[2] 0.0322f
C8099 a_2475_12194# a_16018_12170# 0.316f
C8100 VDD a_34090_5142# 0.483f
C8101 col_n[23] a_26362_5182# 0.084f
C8102 m2_26256_18442# VDD 0.0456f
C8103 col_n[7] a_9994_16186# 0.251f
C8104 a_19942_17190# a_20338_17230# 0.0313f
C8105 col_n[4] a_6890_6146# 0.0765f
C8106 VDD a_23446_14540# 0.0779f
C8107 a_2874_1126# m2_2736_946# 0.225f
C8108 col_n[14] a_16930_18194# 0.0762f
C8109 col_n[20] a_2275_13198# 0.113f
C8110 col_n[25] a_2275_2154# 0.113f
C8111 a_2275_9182# a_6982_9158# 0.399f
C8112 a_3970_9158# a_4274_9198# 0.0931f
C8113 a_4882_9158# a_5374_9520# 0.0658f
C8114 rowoff_n[14] a_24450_16548# 0.0133f
C8115 m2_17220_15430# a_17022_15182# 0.165f
C8116 rowon_n[2] a_2874_4138# 0.118f
C8117 vcm a_18938_18194# 0.101f
C8118 m2_19228_17438# rowon_n[15] 0.0322f
C8119 a_16018_14178# a_17022_14178# 0.843f
C8120 a_2475_14202# a_31078_14178# 0.316f
C8121 m2_25252_13422# rowon_n[11] 0.0322f
C8122 VDD a_15014_8154# 0.483f
C8123 m2_31276_9406# rowon_n[7] 0.0322f
C8124 m2_25828_946# vcm 0.353f
C8125 col[17] a_20034_3134# 0.367f
C8126 col[10] a_2275_10186# 0.0899f
C8127 col[17] rowoff_n[12] 0.0901f
C8128 VDD a_4370_17552# 0.0779f
C8129 col_n[31] a_34394_17230# 0.084f
C8130 col[27] a_30074_15182# 0.367f
C8131 col[24] a_26970_5142# 0.0682f
C8132 vcm a_21038_3134# 0.56f
C8133 a_35002_7150# a_35094_7150# 0.0991f
C8134 a_34090_7150# a_34394_7190# 0.0931f
C8135 a_2275_11190# a_22042_11166# 0.399f
C8136 col[30] a_2475_9182# 0.136f
C8137 row_n[11] a_14010_13174# 0.282f
C8138 a_6982_16186# a_6982_15182# 0.843f
C8139 VDD a_30074_12170# 0.483f
C8140 m2_19804_18014# m3_19936_18146# 3.79f
C8141 col_n[12] a_15318_3174# 0.084f
C8142 rowon_n[15] a_13918_17190# 0.118f
C8143 col_n[22] a_25358_15222# 0.084f
C8144 a_29982_4138# a_30378_4178# 0.0313f
C8145 rowoff_n[1] a_9994_3134# 0.294f
C8146 row_n[1] a_24050_3134# 0.282f
C8147 col_n[3] a_5886_16186# 0.0765f
C8148 row_n[13] a_2275_15206# 19.2f
C8149 rowon_n[5] a_23958_7150# 0.118f
C8150 vcm a_2475_6170# 1.08f
C8151 rowoff_n[12] a_30986_14178# 0.202f
C8152 a_2275_8178# a_12306_8194# 0.144f
C8153 a_2475_8178# a_14922_8154# 0.264f
C8154 m2_8184_13422# a_7986_13174# 0.165f
C8155 a_19030_13174# a_19334_13214# 0.0931f
C8156 a_19942_13174# a_20434_13536# 0.0658f
C8157 row_n[3] a_11302_5182# 0.0117f
C8158 col[1] rowoff_n[13] 0.0901f
C8159 m3_1864_8106# a_2966_8154# 0.0302f
C8160 VDD a_10998_15182# 0.483f
C8161 col[27] a_2275_12194# 0.0899f
C8162 m2_10768_18014# col[8] 0.347f
C8163 a_2275_5166# a_5886_5142# 0.136f
C8164 col[16] a_19030_13174# 0.367f
C8165 m2_23820_946# m3_22948_1078# 0.0341f
C8166 m2_27260_9406# a_27062_9158# 0.165f
C8167 col[13] a_15926_3134# 0.0682f
C8168 vcm a_17022_10162# 0.56f
C8169 a_2275_10186# a_27366_10202# 0.144f
C8170 a_15926_10162# a_16018_10162# 0.326f
C8171 a_2475_10186# a_29982_10162# 0.264f
C8172 rowoff_n[15] a_12402_17552# 0.0133f
C8173 row_n[14] a_35002_16186# 0.0437f
C8174 col[23] a_25966_15182# 0.0682f
C8175 VDD a_2275_9182# 1.96f
C8176 m2_14784_18014# ctop 0.0422f
C8177 col_n[31] a_34090_9158# 0.251f
C8178 col_n[1] a_4274_1166# 0.0572f
C8179 a_17022_3134# a_17022_2130# 0.843f
C8180 m2_3164_7398# row_n[5] 0.0128f
C8181 col_n[11] a_14314_13214# 0.084f
C8182 m2_9188_3382# row_n[1] 0.0128f
C8183 vcm a_7286_4178# 0.155f
C8184 a_2275_7174# a_20946_7150# 0.136f
C8185 a_10906_7150# a_11302_7190# 0.0313f
C8186 rowoff_n[9] a_2161_11190# 0.0226f
C8187 col_n[17] a_2475_8178# 0.0531f
C8188 vcm a_32082_14178# 0.56f
C8189 VDD a_28978_4138# 0.181f
C8190 col_n[22] a_25454_7512# 0.0283f
C8191 a_35002_17190# a_35494_17552# 0.0658f
C8192 row_n[8] a_22042_10162# 0.282f
C8193 col[2] a_2475_16210# 0.136f
C8194 rowoff_n[7] a_11910_9158# 0.202f
C8195 rowon_n[12] a_21950_14178# 0.118f
C8196 a_2475_4162# a_13006_4138# 0.316f
C8197 col[7] a_2475_5166# 0.136f
C8198 a_6982_4138# a_7986_4138# 0.843f
C8199 m3_1864_16138# ctop 0.21f
C8200 m2_18224_7398# a_18026_7150# 0.165f
C8201 col_n[0] a_3366_1488# 0.0283f
C8202 m2_18224_16434# row_n[14] 0.0128f
C8203 m2_24248_12418# row_n[10] 0.0128f
C8204 vcm a_22346_8194# 0.155f
C8205 rowoff_n[13] a_18938_15182# 0.202f
C8206 a_2275_9182# a_34394_9198# 0.144f
C8207 m2_30272_8402# row_n[6] 0.0128f
C8208 m2_35292_4386# row_n[2] 0.0128f
C8209 row_n[10] a_9294_12210# 0.0117f
C8210 rowon_n[2] a_31990_4138# 0.118f
C8211 col[5] a_7986_11166# 0.367f
C8212 m2_26832_18014# col_n[24] 0.243f
C8213 vcm a_13006_17190# 0.56f
C8214 col[2] a_4882_1126# 0.0682f
C8215 a_30986_14178# a_31078_14178# 0.326f
C8216 VDD a_9902_7150# 0.181f
C8217 rowoff_n[5] a_20946_7150# 0.202f
C8218 col[12] a_14922_13174# 0.0682f
C8219 col_n[14] a_2275_11190# 0.113f
C8220 a_2275_18218# a_14010_18194# 0.0924f
C8221 row_n[0] a_19334_2170# 0.0117f
C8222 a_2275_1150# a_3970_1126# 0.399f
C8223 col_n[20] a_23046_7150# 0.251f
C8224 vcm a_15926_2130# 0.1f
C8225 col_n[27] a_29982_9158# 0.0765f
C8226 a_32082_7150# a_32082_6146# 0.843f
C8227 a_2475_6170# a_28066_6146# 0.316f
C8228 rowoff_n[3] a_29982_5142# 0.202f
C8229 vcm a_3270_11206# 0.155f
C8230 row_n[2] a_9902_4138# 0.0437f
C8231 row_n[7] col[25] 0.0342f
C8232 row_n[10] col[31] 0.0342f
C8233 rowon_n[4] col[20] 0.0323f
C8234 row_n[9] col[29] 0.0342f
C8235 row_n[4] col[19] 0.0342f
C8236 rowon_n[9] col[30] 0.0323f
C8237 rowon_n[6] col[24] 0.0323f
C8238 row_n[3] col[17] 0.0342f
C8239 row_n[1] col[13] 0.0342f
C8240 ctop col[8] 0.123f
C8241 row_n[8] col[27] 0.0342f
C8242 rowon_n[3] col[18] 0.0323f
C8243 row_n[0] col[11] 0.0342f
C8244 row_n[2] col[15] 0.0342f
C8245 rowon_n[10] sample_n 0.0692f
C8246 rowon_n[2] col[16] 0.0323f
C8247 a_25966_11166# a_26362_11206# 0.0313f
C8248 rowon_n[8] col[28] 0.0323f
C8249 row_n[6] col[23] 0.0342f
C8250 rowon_n[1] col[14] 0.0323f
C8251 row_n[5] col[21] 0.0342f
C8252 rowon_n[7] col[26] 0.0323f
C8253 rowon_n[0] col[12] 0.0323f
C8254 rowon_n[5] col[22] 0.0323f
C8255 VDD a_35494_2492# 0.106f
C8256 col[4] a_2275_8178# 0.0899f
C8257 rowon_n[6] a_8990_8154# 0.248f
C8258 m2_34864_6970# VDD 0.772f
C8259 ctop a_16018_6146# 4.11f
C8260 a_2275_15206# a_4274_15222# 0.144f
C8261 a_2475_15206# a_6890_15182# 0.264f
C8262 VDD a_24962_11166# 0.181f
C8263 col_n[11] a_14410_5504# 0.0283f
C8264 a_10906_3134# a_11398_3496# 0.0658f
C8265 a_2275_3158# a_19030_3134# 0.399f
C8266 a_9994_3134# a_10298_3174# 0.0931f
C8267 a_2475_18218# a_12002_18194# 0.0299f
C8268 rowoff_n[8] a_21438_10524# 0.0133f
C8269 col_n[21] a_24450_17552# 0.0283f
C8270 a_32994_1126# a_2275_1150# 0.136f
C8271 m2_9188_5390# a_8990_5142# 0.165f
C8272 col[24] a_2475_7174# 0.136f
C8273 vcm a_30986_6146# 0.1f
C8274 a_22042_8154# a_23046_8154# 0.843f
C8275 vcm a_18330_15222# 0.155f
C8276 VDD a_16418_5504# 0.0779f
C8277 sample a_2161_11190# 0.0858f
C8278 a_28370_1166# VDD 0.0149f
C8279 row_n[15] a_20034_17190# 0.282f
C8280 ctop a_31078_10162# 4.11f
C8281 a_11910_17190# a_12002_17190# 0.326f
C8282 a_2475_17214# a_21950_17190# 0.264f
C8283 a_2275_17214# a_19334_17230# 0.144f
C8284 rowoff_n[6] a_30474_8516# 0.0133f
C8285 VDD a_5886_14178# 0.181f
C8286 col_n[31] a_2275_13198# 0.113f
C8287 row_n[5] a_30074_7150# 0.282f
C8288 a_2275_5166# a_34090_5142# 0.399f
C8289 col_n[9] a_12002_5142# 0.251f
C8290 rowon_n[9] a_29982_11166# 0.118f
C8291 vcm a_11910_9158# 0.1f
C8292 col_n[19] a_22042_17190# 0.251f
C8293 a_31990_1126# a_32482_1488# 0.0658f
C8294 rowoff_n[14] a_6890_16186# 0.202f
C8295 a_13006_10162# a_13006_9158# 0.843f
C8296 col_n[16] a_18938_7150# 0.0765f
C8297 m2_1732_15002# a_2966_15182# 0.843f
C8298 col[21] a_2275_10186# 0.0899f
C8299 m2_11772_946# a_12306_1166# 0.087f
C8300 a_6890_14178# a_7286_14218# 0.0313f
C8301 col[28] rowoff_n[12] 0.0901f
C8302 a_2275_14202# a_12914_14178# 0.136f
C8303 m2_1732_15002# ctop 0.0428f
C8304 row_n[7] a_17326_9198# 0.0117f
C8305 VDD a_31478_9520# 0.0779f
C8306 ctop a_12002_13174# 4.11f
C8307 VDD a_20946_18194# 0.343f
C8308 a_2475_2154# a_26970_2130# 0.264f
C8309 a_2275_2154# a_24354_2170# 0.144f
C8310 m2_29844_946# VDD 1f
C8311 vcm a_2966_3134# 0.56f
C8312 row_n[9] a_7894_11166# 0.0437f
C8313 rowoff_n[9] a_31078_11166# 0.294f
C8314 a_25966_7150# a_26458_7512# 0.0658f
C8315 a_25054_7150# a_25358_7190# 0.0931f
C8316 col_n[10] a_13406_15544# 0.0283f
C8317 rowon_n[13] a_6982_15182# 0.248f
C8318 vcm a_26970_13174# 0.1f
C8319 a_2475_11190# a_4974_11166# 0.316f
C8320 VDD a_23046_3134# 0.483f
C8321 col[29] a_32082_4138# 0.367f
C8322 m2_34864_18014# a_2275_18218# 0.278f
C8323 a_2275_16210# a_27974_16186# 0.136f
C8324 VDD a_12402_12532# 0.0779f
C8325 rowon_n[3] a_17022_5142# 0.248f
C8326 a_32994_1126# m2_32856_946# 0.225f
C8327 col_n[6] a_2475_17214# 0.0531f
C8328 ctop a_27062_17190# 4.06f
C8329 col_n[11] a_2475_6170# 0.0531f
C8330 a_21950_4138# a_22042_4138# 0.326f
C8331 col_n[24] a_27366_4178# 0.084f
C8332 col[12] rowoff_n[13] 0.0901f
C8333 vcm a_7894_16186# 0.1f
C8334 a_28066_14178# a_28066_13174# 0.843f
C8335 a_2475_13198# a_20034_13174# 0.316f
C8336 col_n[8] a_10998_15182# 0.251f
C8337 VDD a_3970_6146# 0.483f
C8338 col_n[5] a_7894_5142# 0.0765f
C8339 col[1] a_2475_3158# 0.136f
C8340 m2_30848_18014# a_2475_18218# 0.286f
C8341 col_n[15] a_17934_17190# 0.0765f
C8342 a_21950_18194# a_22346_18234# 0.0313f
C8343 VDD a_27462_16548# 0.0779f
C8344 a_16930_1126# a_17326_1166# 0.0313f
C8345 row_n[12] a_28066_14178# 0.282f
C8346 vcm a_9994_1126# 0.165f
C8347 m2_8184_15430# rowon_n[13] 0.0322f
C8348 m2_14208_11414# rowon_n[9] 0.0322f
C8349 m2_20232_7398# rowon_n[5] 0.0322f
C8350 m2_26256_3382# rowon_n[1] 0.0322f
C8351 m2_33860_946# m2_34864_946# 0.512f
C8352 col_n[8] a_2275_9182# 0.113f
C8353 a_2275_10186# a_10998_10162# 0.399f
C8354 a_5978_10162# a_6282_10202# 0.0931f
C8355 a_6890_10162# a_7382_10524# 0.0658f
C8356 row_n[14] a_15318_16226# 0.0117f
C8357 m2_34864_17010# a_35002_17190# 0.225f
C8358 a_2475_15206# a_35094_15182# 0.0299f
C8359 m2_4744_946# a_4974_2130# 0.843f
C8360 a_18026_15182# a_19030_15182# 0.843f
C8361 VDD a_19030_10162# 0.483f
C8362 col[18] a_21038_2130# 0.367f
C8363 col[28] a_31078_14178# 0.367f
C8364 row_n[4] a_25358_6186# 0.0117f
C8365 col[25] a_27974_4138# 0.0682f
C8366 col_n[28] a_2475_8178# 0.0531f
C8367 vcm a_25054_5142# 0.56f
C8368 rowoff_n[10] a_19030_12170# 0.294f
C8369 rowoff_n[2] a_2475_4162# 3.9f
C8370 m2_34864_16006# rowon_n[14] 0.231f
C8371 row_n[6] a_15926_8154# 0.0437f
C8372 a_2275_12194# a_26058_12170# 0.399f
C8373 rowon_n[10] a_15014_12170# 0.248f
C8374 col_n[13] a_16322_2170# 0.084f
C8375 col[13] a_2475_16210# 0.136f
C8376 a_8990_17190# a_8990_16186# 0.843f
C8377 VDD a_34090_14178# 0.483f
C8378 col_n[23] a_26362_14218# 0.084f
C8379 col[18] a_2475_5166# 0.136f
C8380 rowoff_n[0] a_10998_2130# 0.294f
C8381 rowon_n[0] a_25054_2130# 0.248f
C8382 col_n[4] a_6890_15182# 0.0765f
C8383 rowon_n[12] a_3878_14178# 0.118f
C8384 a_31990_5142# a_32386_5182# 0.0313f
C8385 m2_16792_946# ctop 0.0435f
C8386 vcm a_5978_8154# 0.56f
C8387 a_2275_9182# a_16322_9198# 0.144f
C8388 a_2475_9182# a_18938_9158# 0.264f
C8389 rowoff_n[14] a_35094_16186# 0.0135f
C8390 col_n[25] a_2275_11190# 0.113f
C8391 a_21950_14178# a_22442_14540# 0.0658f
C8392 a_21038_14178# a_21342_14218# 0.0931f
C8393 rowoff_n[5] a_2275_7174# 0.151f
C8394 row_n[0] a_2874_2130# 0.0436f
C8395 VDD a_15014_17190# 0.484f
C8396 a_28066_2130# a_29070_2130# 0.843f
C8397 rowon_n[4] a_2161_6170# 0.0177f
C8398 col[17] a_20034_12170# 0.367f
C8399 row_n[2] col[26] 0.0342f
C8400 rowon_n[1] col[25] 0.0323f
C8401 row_n[1] col[24] 0.0342f
C8402 ctop col[19] 0.123f
C8403 col[6] col[7] 0.0355f
C8404 en_bit_n[2] col[16] 0.142f
C8405 row_n[0] col[22] 0.0342f
C8406 rowon_n[4] col[31] 0.0323f
C8407 vcm a_30378_3174# 0.155f
C8408 rowon_n[3] col[29] 0.0323f
C8409 rowon_n[0] col[23] 0.0323f
C8410 row_n[4] col[30] 0.0342f
C8411 row_n[3] col[28] 0.0342f
C8412 row_n[5] sample_n 0.0596f
C8413 rowon_n[2] col[27] 0.0323f
C8414 col[14] a_16930_2130# 0.0682f
C8415 a_2275_6170# a_9902_6146# 0.136f
C8416 m2_1732_12994# sample_n 0.0522f
C8417 col[15] a_2275_8178# 0.0899f
C8418 col[24] a_26970_14178# 0.0682f
C8419 vcm a_21038_12170# 0.56f
C8420 a_2475_11190# a_33998_11166# 0.264f
C8421 a_2275_11190# a_31382_11206# 0.144f
C8422 a_17934_11166# a_18026_11166# 0.326f
C8423 VDD a_17934_2130# 0.181f
C8424 row_n[11] a_23350_13214# 0.0117f
C8425 m2_33860_18014# m3_34996_18146# 0.0341f
C8426 col_n[12] a_15318_12210# 0.084f
C8427 a_19030_4138# a_19030_3134# 0.843f
C8428 row_n[1] a_33390_3174# 0.0117f
C8429 rowoff_n[8] a_3366_10524# 0.0133f
C8430 row_n[13] a_13918_15182# 0.0437f
C8431 vcm a_11302_6186# 0.155f
C8432 a_12914_8154# a_13310_8194# 0.0313f
C8433 rowoff_n[11] a_6982_13174# 0.294f
C8434 a_2275_8178# a_24962_8154# 0.136f
C8435 vcm a_2475_15206# 1.08f
C8436 VDD a_32994_6146# 0.181f
C8437 col_n[23] a_26458_6508# 0.0283f
C8438 col_n[5] a_2475_4162# 0.0531f
C8439 row_n[3] a_23958_5142# 0.0437f
C8440 row_n[15] a_1957_17214# 0.187f
C8441 rowon_n[7] a_23046_9158# 0.248f
C8442 a_2275_17214# a_2874_17190# 0.136f
C8443 m2_7180_14426# row_n[12] 0.0128f
C8444 a_2475_17214# a_3878_17190# 0.264f
C8445 rowoff_n[6] a_12914_8154# 0.202f
C8446 m2_13204_10410# row_n[8] 0.0128f
C8447 m2_19228_6394# row_n[4] 0.0128f
C8448 a_8990_5142# a_9994_5142# 0.843f
C8449 a_2475_5166# a_17022_5142# 0.316f
C8450 m2_34864_8978# a_35398_9198# 0.087f
C8451 col[6] a_8990_10162# 0.367f
C8452 vcm a_26362_10202# 0.155f
C8453 en_C0_n a_2475_1150# 0.0162f
C8454 rowoff_n[15] a_23046_17190# 0.294f
C8455 m2_23244_16434# a_23046_16186# 0.165f
C8456 rowoff_n[4] a_21950_6146# 0.202f
C8457 col[13] a_15926_12170# 0.0682f
C8458 ctop a_4974_4138# 4.11f
C8459 m2_27836_946# col[25] 0.425f
C8460 a_32994_15182# a_33086_15182# 0.326f
C8461 VDD a_13918_9158# 0.181f
C8462 col_n[21] a_24050_6146# 0.251f
C8463 VDD a_2275_18218# 22.9f
C8464 a_2275_2154# a_7986_2130# 0.399f
C8465 m2_34288_15430# row_n[13] 0.0128f
C8466 col_n[28] a_30986_8154# 0.0765f
C8467 col_n[2] a_2275_7174# 0.113f
C8468 vcm a_19942_4138# 0.1f
C8469 rowon_n[1] a_10906_3134# 0.118f
C8470 rowoff_n[2] a_30986_4138# 0.202f
C8471 a_34090_8154# a_34090_7150# 0.843f
C8472 rowoff_n[9] a_13406_11528# 0.0133f
C8473 col_n[1] a_4274_10202# 0.084f
C8474 a_2475_7174# a_32082_7150# 0.316f
C8475 vcm a_7286_13214# 0.155f
C8476 a_27974_12170# a_28370_12210# 0.0313f
C8477 VDD a_5374_3496# 0.0779f
C8478 col_n[17] a_2475_17214# 0.0531f
C8479 ctop a_20034_8154# 4.11f
C8480 a_2475_16210# a_10906_16186# 0.264f
C8481 a_2275_16210# a_8290_16226# 0.144f
C8482 col_n[22] a_2475_6170# 0.0531f
C8483 VDD a_28978_13174# 0.181f
C8484 col_n[12] a_15414_4500# 0.0283f
C8485 row_n[8] a_31382_10202# 0.0117f
C8486 rowoff_n[7] a_22442_9520# 0.0133f
C8487 col_n[22] a_25454_16548# 0.0283f
C8488 a_12002_4138# a_12306_4178# 0.0931f
C8489 a_2275_4162# a_23046_4138# 0.399f
C8490 a_12914_4138# a_13406_4500# 0.0658f
C8491 m3_13912_1078# ctop 0.21f
C8492 col[23] rowoff_n[13] 0.0901f
C8493 vcm a_35002_8154# 0.101f
C8494 col[7] a_2475_14202# 0.136f
C8495 rowoff_n[13] a_29470_15544# 0.0133f
C8496 a_24050_9158# a_25054_9158# 0.843f
C8497 m2_14208_14426# a_14010_14178# 0.165f
C8498 row_n[10] a_21950_12170# 0.0437f
C8499 sample rowoff_n[1] 0.0775f
C8500 col_n[2] rowoff_n[5] 0.0471f
C8501 col[12] a_2475_3158# 0.136f
C8502 col_n[4] rowoff_n[7] 0.0471f
C8503 vcm rowoff_n[3] 0.533f
C8504 col_n[5] rowoff_n[8] 0.0471f
C8505 col_n[3] rowoff_n[6] 0.0471f
C8506 col_n[0] rowoff_n[2] 0.0471f
C8507 col_n[1] rowoff_n[4] 0.0471f
C8508 VDD rowoff_n[0] 1.51f
C8509 col_n[0] a_3366_10524# 0.0283f
C8510 col_n[6] rowoff_n[9] 0.0471f
C8511 vcm a_22346_17230# 0.155f
C8512 a_2475_13198# a_1957_13198# 0.0734f
C8513 rowon_n[14] a_21038_16186# 0.248f
C8514 VDD a_20434_7512# 0.0779f
C8515 rowoff_n[5] a_31478_7512# 0.0133f
C8516 col[2] a_4882_10162# 0.0682f
C8517 a_13918_18194# a_14010_18194# 0.0991f
C8518 a_2275_18218# a_23350_18234# 0.145f
C8519 row_n[0] a_31990_2130# 0.0437f
C8520 VDD a_9902_16186# 0.181f
C8521 a_2475_1150# a_15926_1126# 0.264f
C8522 a_2275_1150# a_13310_1166# 0.145f
C8523 a_8898_1126# a_8990_1126# 0.0991f
C8524 rowon_n[4] a_31078_6146# 0.248f
C8525 m2_11196_2378# a_10998_2130# 0.165f
C8526 col_n[10] a_13006_4138# 0.251f
C8527 col_n[19] a_2275_9182# 0.113f
C8528 col_n[20] a_23046_16186# 0.251f
C8529 m2_34864_7974# vcm 0.395f
C8530 col_n[17] a_19942_6146# 0.0765f
C8531 m2_33284_10410# a_33086_10162# 0.165f
C8532 vcm a_15926_11166# 0.1f
C8533 a_15014_11166# a_15014_10162# 0.843f
C8534 col_n[27] a_29982_18194# 0.0762f
C8535 VDD a_12002_1126# 0.035f
C8536 a_8898_15182# a_9294_15222# 0.0313f
C8537 a_2275_15206# a_16930_15182# 0.136f
C8538 VDD a_35494_11528# 0.106f
C8539 col[4] a_2275_17214# 0.0899f
C8540 m2_34864_15002# m3_34996_16138# 0.0341f
C8541 rowon_n[0] m2_31276_2378# 0.0322f
C8542 ctop a_16018_15182# 4.11f
C8543 row_n[4] a_8990_6146# 0.282f
C8544 col[9] a_2275_6170# 0.0899f
C8545 col[7] rowoff_n[14] 0.0901f
C8546 a_2475_3158# a_30986_3134# 0.264f
C8547 a_2275_3158# a_28370_3174# 0.144f
C8548 col_n[1] a_4370_2492# 0.0283f
C8549 rowon_n[8] a_8898_10162# 0.118f
C8550 rowoff_n[8] a_32082_10162# 0.294f
C8551 col_n[11] a_14410_14540# 0.0283f
C8552 a_27974_8154# a_28466_8516# 0.0658f
C8553 a_27062_8154# a_27366_8194# 0.0931f
C8554 col[30] a_33086_3134# 0.367f
C8555 m2_5172_12418# a_4974_12170# 0.165f
C8556 col[24] a_2475_16210# 0.136f
C8557 vcm a_30986_15182# 0.1f
C8558 a_4974_12170# a_5978_12170# 0.843f
C8559 a_2475_12194# a_8990_12170# 0.316f
C8560 VDD a_27062_5142# 0.483f
C8561 col[29] a_2475_5166# 0.136f
C8562 m2_12200_18442# VDD 0.0456f
C8563 row_n[15] a_29374_17230# 0.0117f
C8564 a_2275_17214# a_31990_17190# 0.136f
C8565 VDD a_16418_14540# 0.0779f
C8566 rowon_n[0] m2_20232_2378# 0.0322f
C8567 a_23958_5142# a_24050_5142# 0.326f
C8568 m2_24248_8402# a_24050_8154# 0.165f
C8569 col_n[25] a_28370_3174# 0.084f
C8570 col_n[0] a_2475_2154# 0.0532f
C8571 rowoff_n[14] a_17422_16548# 0.0133f
C8572 col_n[9] a_12002_14178# 0.251f
C8573 col_n[6] a_8898_4138# 0.0765f
C8574 vcm a_11910_18194# 0.101f
C8575 a_2475_14202# a_24050_14178# 0.316f
C8576 a_30074_15182# a_30074_14178# 0.843f
C8577 row_n[7] a_29982_9158# 0.0437f
C8578 col_n[16] a_18938_16186# 0.0765f
C8579 VDD a_7986_8154# 0.483f
C8580 m2_3164_9406# rowon_n[7] 0.0322f
C8581 m2_9188_5390# rowon_n[3] 0.0322f
C8582 rowon_n[11] a_29070_13174# 0.248f
C8583 VDD col_n[7] 5.17f
C8584 vcm col_n[4] 1.94f
C8585 VDD a_31478_18556# 0.0858f
C8586 ctop col[30] 0.125f
C8587 col[26] a_2275_8178# 0.0899f
C8588 a_18938_2130# a_19334_2170# 0.0313f
C8589 m2_34864_2954# a_2475_3158# 0.282f
C8590 m3_32988_18146# VDD 0.0277f
C8591 vcm a_14010_3134# 0.56f
C8592 vcm a_2966_12170# 0.56f
C8593 a_2275_11190# a_15014_11166# 0.399f
C8594 a_7986_11166# a_8290_11206# 0.0931f
C8595 a_8898_11166# a_9390_11528# 0.0658f
C8596 m2_20808_18014# a_20946_18194# 0.225f
C8597 m2_1732_9982# VDD 0.856f
C8598 a_20034_16186# a_21038_16186# 0.843f
C8599 row_n[11] a_6982_13174# 0.282f
C8600 col[29] a_32082_13174# 0.367f
C8601 VDD a_23046_12170# 0.483f
C8602 m2_10768_18014# m3_9896_18146# 0.0341f
C8603 col[26] a_28978_3134# 0.0682f
C8604 rowon_n[15] a_6890_17190# 0.118f
C8605 m2_24248_14426# rowon_n[12] 0.0322f
C8606 m2_30272_10410# rowon_n[8] 0.0322f
C8607 m2_35292_6394# rowon_n[4] 0.0322f
C8608 rowoff_n[1] a_2874_3134# 0.202f
C8609 row_n[1] a_17022_3134# 0.282f
C8610 m2_15212_6394# a_15014_6146# 0.165f
C8611 col_n[11] a_2475_15206# 0.0531f
C8612 rowon_n[5] a_16930_7150# 0.118f
C8613 vcm a_29070_7150# 0.56f
C8614 a_3878_8154# a_4274_8194# 0.0313f
C8615 a_4882_8154# a_4974_8154# 0.326f
C8616 a_2275_8178# a_5278_8194# 0.144f
C8617 a_2475_8178# a_7894_8154# 0.264f
C8618 rowoff_n[12] a_23958_14178# 0.202f
C8619 col_n[16] a_2475_4162# 0.0531f
C8620 m2_1732_12994# a_2275_13198# 0.191f
C8621 col_n[14] a_17326_1166# 0.0839f
C8622 a_2275_13198# a_30074_13174# 0.399f
C8623 col_n[24] a_27366_13214# 0.084f
C8624 row_n[3] a_4274_5182# 0.0117f
C8625 VDD a_3970_15182# 0.483f
C8626 col_n[5] a_7894_14178# 0.0765f
C8627 col[1] a_2475_12194# 0.136f
C8628 vcm a_19334_1166# 0.155f
C8629 col[6] a_2475_1150# 0.136f
C8630 m2_12776_946# m3_13912_1078# 0.0341f
C8631 vcm a_9994_10162# 0.56f
C8632 a_2275_10186# a_20338_10202# 0.144f
C8633 a_2475_10186# a_22954_10162# 0.264f
C8634 rowoff_n[15] a_5374_17552# 0.0133f
C8635 row_n[14] a_27974_16186# 0.0437f
C8636 rowoff_n[4] a_3878_6146# 0.202f
C8637 a_23046_15182# a_23350_15222# 0.0931f
C8638 col_n[8] a_2275_18218# 0.113f
C8639 a_23958_15182# a_24450_15544# 0.0658f
C8640 m2_34864_11990# m3_34996_13126# 0.0341f
C8641 col_n[13] a_2275_7174# 0.113f
C8642 col[18] a_21038_11166# 0.367f
C8643 a_30074_3134# a_31078_3134# 0.843f
C8644 col[15] a_17934_1126# 0.0699f
C8645 m2_6176_4386# a_5978_4138# 0.165f
C8646 vcm a_35398_5182# 0.161f
C8647 col[25] a_27974_13174# 0.0682f
C8648 a_2275_7174# a_13918_7150# 0.136f
C8649 col_n[28] a_2475_17214# 0.0531f
C8650 m2_29844_18014# vcm 0.353f
C8651 col_n[0] a_3270_7190# 0.084f
C8652 vcm a_25054_14178# 0.56f
C8653 a_19942_12170# a_20034_12170# 0.326f
C8654 a_2275_12194# a_2275_11190# 0.0715f
C8655 VDD a_21950_4138# 0.181f
C8656 col[3] a_2275_4162# 0.0899f
C8657 col_n[13] a_16322_11206# 0.084f
C8658 row_n[8] a_15014_10162# 0.282f
C8659 rowoff_n[7] a_4882_9158# 0.202f
C8660 col[18] a_2475_14202# 0.136f
C8661 rowon_n[12] a_14922_14178# 0.118f
C8662 a_2966_4138# a_3270_4178# 0.0931f
C8663 a_21038_5142# a_21038_4138# 0.843f
C8664 a_2475_4162# a_5978_4138# 0.316f
C8665 a_3878_4138# a_4370_4500# 0.0658f
C8666 m3_9896_18146# ctop 0.209f
C8667 col_n[14] rowoff_n[6] 0.0471f
C8668 col[23] a_2475_3158# 0.136f
C8669 col_n[17] rowoff_n[9] 0.0471f
C8670 col_n[9] rowoff_n[1] 0.0471f
C8671 col_n[12] rowoff_n[4] 0.0471f
C8672 col_n[15] rowoff_n[7] 0.0471f
C8673 col_n[10] rowoff_n[2] 0.0471f
C8674 col_n[16] rowoff_n[8] 0.0471f
C8675 col_n[11] rowoff_n[3] 0.0471f
C8676 col_n[8] rowoff_n[0] 0.0471f
C8677 col_n[13] rowoff_n[5] 0.0471f
C8678 m2_33860_18014# m2_34864_18014# 0.843f
C8679 vcm a_15318_8194# 0.155f
C8680 m2_2160_8402# row_n[6] 0.0194f
C8681 a_2275_9182# a_28978_9158# 0.136f
C8682 a_14922_9158# a_15318_9198# 0.0313f
C8683 rowoff_n[13] a_11910_15182# 0.202f
C8684 m2_8184_4386# row_n[2] 0.0128f
C8685 col_n[24] a_27462_5504# 0.0283f
C8686 row_n[10] a_3878_12170# 0.0437f
C8687 m2_34864_15002# a_34090_15182# 0.843f
C8688 rowon_n[2] a_24962_4138# 0.118f
C8689 ctop a_28066_3134# 4.11f
C8690 vcm a_5978_17190# 0.56f
C8691 rowon_n[14] a_2966_16186# 0.248f
C8692 VDD a_2161_7174# 0.187f
C8693 rowoff_n[5] a_13918_7150# 0.202f
C8694 a_2275_18218# a_6982_18194# 0.0924f
C8695 a_4882_18194# a_5374_18556# 0.0658f
C8696 col_n[30] a_2275_9182# 0.113f
C8697 row_n[0] a_12306_2170# 0.0117f
C8698 a_33998_2130# a_34490_2492# 0.0658f
C8699 a_33086_2130# a_33390_2170# 0.0931f
C8700 vcm a_8898_2130# 0.1f
C8701 a_2475_6170# a_21038_6146# 0.316f
C8702 col[7] a_9994_9158# 0.367f
C8703 a_10998_6146# a_12002_6146# 0.843f
C8704 row_n[2] a_2161_4162# 0.0221f
C8705 rowoff_n[3] a_22954_5142# 0.202f
C8706 vcm a_30378_12210# 0.155f
C8707 col[14] a_16930_11166# 0.0682f
C8708 m2_17220_17438# row_n[15] 0.0128f
C8709 VDD a_28466_2492# 0.0779f
C8710 col[15] a_2275_17214# 0.0899f
C8711 rowon_n[6] a_2475_8178# 0.31f
C8712 m2_23244_13422# row_n[11] 0.0128f
C8713 m2_16792_18014# a_17022_17190# 0.843f
C8714 m2_29268_9406# row_n[7] 0.0128f
C8715 m2_34864_4962# row_n[3] 0.267f
C8716 ctop a_8990_6146# 4.11f
C8717 col[20] a_2275_6170# 0.0899f
C8718 a_35002_16186# a_35094_16186# 0.0991f
C8719 row_n[11] a_34394_13214# 0.0117f
C8720 a_34090_16186# a_34394_16226# 0.0931f
C8721 col_n[22] a_25054_5142# 0.251f
C8722 VDD a_17934_11166# 0.181f
C8723 m2_1732_16006# m3_1864_16138# 3.79f
C8724 col[18] rowoff_n[14] 0.0901f
C8725 rowon_n[15] a_35094_17190# 0.0141f
C8726 col_n[29] a_31990_7150# 0.0765f
C8727 a_2275_3158# a_12002_3134# 0.399f
C8728 a_2475_18218# a_4974_18194# 0.0299f
C8729 col_n[1] rowoff_n[10] 0.0471f
C8730 rowoff_n[1] a_31990_3134# 0.202f
C8731 rowoff_n[8] a_14410_10524# 0.0133f
C8732 col_n[2] a_5278_9198# 0.084f
C8733 a_25966_1126# a_2275_1150# 0.136f
C8734 vcm a_23958_6146# 0.1f
C8735 a_2475_8178# a_2475_7174# 0.0666f
C8736 vcm a_11302_15222# 0.155f
C8737 a_29982_13174# a_30378_13214# 0.0313f
C8738 VDD a_9390_5504# 0.0779f
C8739 col_n[13] a_16418_3496# 0.0283f
C8740 ctop a_24050_10162# 4.11f
C8741 row_n[15] a_13006_17190# 0.282f
C8742 a_2475_17214# a_14922_17190# 0.264f
C8743 a_2275_17214# a_12306_17230# 0.144f
C8744 rowoff_n[6] a_23446_8516# 0.0133f
C8745 VDD a_32994_15182# 0.181f
C8746 col_n[23] a_26458_15544# 0.0283f
C8747 col_n[5] a_2475_13198# 0.0531f
C8748 m3_21944_18146# a_22042_17190# 0.0303f
C8749 col_n[10] a_2475_2154# 0.0531f
C8750 a_14922_5142# a_15414_5504# 0.0658f
C8751 a_2275_5166# a_27062_5142# 0.399f
C8752 row_n[5] a_23046_7150# 0.282f
C8753 a_14010_5142# a_14314_5182# 0.0931f
C8754 rowon_n[9] a_22954_11166# 0.118f
C8755 vcm a_4882_9158# 0.1f
C8756 a_26058_10162# a_27062_10162# 0.843f
C8757 rowoff_n[4] a_32482_6508# 0.0133f
C8758 VDD col_n[18] 5.17f
C8759 col_n[7] col_n[8] 0.0101f
C8760 vcm col_n[15] 1.93f
C8761 m2_22816_946# a_2475_1150# 0.286f
C8762 col[17] col[18] 0.0337f
C8763 a_2275_14202# a_5886_14178# 0.136f
C8764 col[2] rowoff_n[15] 0.0901f
C8765 row_n[7] a_10298_9198# 0.0117f
C8766 VDD a_24450_9520# 0.0779f
C8767 col[3] a_5886_9158# 0.0682f
C8768 m2_34864_8978# m3_34996_10114# 0.0341f
C8769 ctop a_4974_13174# 4.11f
C8770 col_n[11] a_14010_3134# 0.251f
C8771 VDD a_13918_18194# 0.343f
C8772 a_10906_2130# a_10998_2130# 0.326f
C8773 a_2275_2154# a_17326_2170# 0.144f
C8774 a_2475_2154# a_19942_2130# 0.264f
C8775 col_n[21] a_24050_15182# 0.251f
C8776 m2_14208_1374# VDD 0.0194f
C8777 col_n[18] a_20946_5142# 0.0765f
C8778 rowoff_n[9] a_24050_11166# 0.294f
C8779 col_n[2] a_2275_16210# 0.113f
C8780 col_n[28] a_30986_17190# 0.0765f
C8781 col_n[7] a_2275_5166# 0.113f
C8782 vcm a_19942_13174# 0.1f
C8783 a_17022_12170# a_17022_11166# 0.843f
C8784 VDD a_16018_3134# 0.483f
C8785 sample a_1957_9182# 0.345f
C8786 m2_20808_18014# a_2275_18218# 0.28f
C8787 a_10906_16186# a_11302_16226# 0.0313f
C8788 a_2275_16210# a_20946_16186# 0.136f
C8789 rowon_n[3] a_9994_5142# 0.248f
C8790 VDD a_5374_12532# 0.0779f
C8791 a_28066_1126# m2_27836_946# 0.0249f
C8792 col_n[2] a_5374_1488# 0.0283f
C8793 ctop a_20034_17190# 4.06f
C8794 rowoff_n[7] a_33086_9158# 0.294f
C8795 col_n[22] a_2475_15206# 0.0531f
C8796 col_n[12] a_15414_13536# 0.0283f
C8797 col_n[27] a_2475_4162# 0.0531f
C8798 a_2275_4162# a_32386_4178# 0.144f
C8799 a_2475_4162# a_35002_4138# 0.264f
C8800 col[31] a_34090_2130# 0.365f
C8801 m2_1732_16006# m2_1732_15002# 0.843f
C8802 a_29982_9158# a_30474_9520# 0.0658f
C8803 a_29070_9158# a_29374_9198# 0.0931f
C8804 vcm a_35002_17190# 0.101f
C8805 a_2475_13198# a_13006_13174# 0.316f
C8806 a_6982_13174# a_7986_13174# 0.843f
C8807 VDD a_31078_7150# 0.483f
C8808 col[12] a_2475_12194# 0.136f
C8809 m2_16792_18014# a_2475_18218# 0.286f
C8810 a_2275_18218# a_34394_18234# 0.145f
C8811 VDD a_20434_16548# 0.0779f
C8812 col[17] a_2475_1150# 0.136f
C8813 row_n[12] a_21038_14178# 0.282f
C8814 col_n[26] a_29374_2170# 0.084f
C8815 vcm a_2874_1126# 0.0989f
C8816 a_25966_6146# a_26058_6146# 0.326f
C8817 col_n[10] a_13006_13174# 0.251f
C8818 m2_26832_946# m2_27260_1374# 0.165f
C8819 col_n[7] a_9902_3134# 0.0765f
C8820 col_n[19] a_2275_18218# 0.113f
C8821 row_n[2] a_31078_4138# 0.282f
C8822 a_2275_10186# a_3970_10162# 0.399f
C8823 row_n[14] a_8290_16226# 0.0117f
C8824 VDD a_21342_1166# 0.0149f
C8825 col_n[17] a_19942_15182# 0.0765f
C8826 rowon_n[6] a_30986_8154# 0.118f
C8827 col_n[24] a_2275_7174# 0.113f
C8828 m2_29268_17438# a_29070_17190# 0.165f
C8829 a_32082_16186# a_32082_15182# 0.843f
C8830 a_2475_15206# a_28066_15182# 0.316f
C8831 VDD a_12002_10162# 0.483f
C8832 m2_1732_12994# m3_1864_13126# 3.79f
C8833 row_n[4] a_18330_6186# 0.0117f
C8834 a_20946_3134# a_21342_3174# 0.0313f
C8835 a_2475_18218# a_33998_18194# 0.264f
C8836 col[9] a_2275_15206# 0.0899f
C8837 vcm a_18026_5142# 0.56f
C8838 col[14] a_2275_4162# 0.0899f
C8839 col_n[1] a_4370_11528# 0.0283f
C8840 rowoff_n[10] a_12002_12170# 0.294f
C8841 a_31990_1126# vcm 0.0989f
C8842 m2_7180_16434# rowon_n[14] 0.0322f
C8843 row_n[6] a_8898_8154# 0.0437f
C8844 m2_13204_12418# rowon_n[10] 0.0322f
C8845 m2_19228_8402# rowon_n[6] 0.0322f
C8846 a_9994_12170# a_10298_12210# 0.0931f
C8847 a_2275_12194# a_19030_12170# 0.399f
C8848 a_10906_12170# a_11398_12532# 0.0658f
C8849 m2_25252_4386# rowon_n[2] 0.0322f
C8850 rowon_n[10] a_7986_12170# 0.248f
C8851 VDD a_3878_4138# 0.181f
C8852 col[30] a_33086_12170# 0.367f
C8853 m2_33860_18014# VDD 1f
C8854 col[27] a_29982_2130# 0.0682f
C8855 a_22042_17190# a_23046_17190# 0.843f
C8856 col[29] a_2475_14202# 0.136f
C8857 VDD a_27062_14178# 0.483f
C8858 col_n[26] rowoff_n[7] 0.0471f
C8859 col_n[25] rowoff_n[6] 0.0471f
C8860 col_n[20] rowoff_n[1] 0.0471f
C8861 col_n[22] rowoff_n[3] 0.0471f
C8862 col_n[19] rowoff_n[0] 0.0471f
C8863 col_n[27] rowoff_n[8] 0.0471f
C8864 col_n[28] rowoff_n[9] 0.0471f
C8865 col_n[21] rowoff_n[2] 0.0471f
C8866 col_n[24] rowoff_n[5] 0.0471f
C8867 col_n[23] rowoff_n[4] 0.0471f
C8868 rowon_n[0] a_18026_2130# 0.248f
C8869 rowoff_n[0] a_3970_2130# 0.294f
C8870 m2_1732_17010# col[0] 0.0137f
C8871 col_n[5] a_2475_18218# 0.0529f
C8872 vcm a_33086_9158# 0.56f
C8873 a_6890_9158# a_6982_9158# 0.326f
C8874 rowoff_n[14] a_28066_16186# 0.294f
C8875 a_2475_9182# a_11910_9158# 0.264f
C8876 a_2275_9182# a_9294_9198# 0.144f
C8877 m2_20232_15430# a_20034_15182# 0.165f
C8878 col_n[25] a_28370_12210# 0.084f
C8879 col_n[0] a_2475_11190# 0.0532f
C8880 a_2275_14202# a_34090_14178# 0.399f
C8881 m2_34288_17438# rowon_n[15] 0.0322f
C8882 m2_34864_5966# m3_34996_7102# 0.0341f
C8883 col_n[6] a_8898_13174# 0.0765f
C8884 VDD a_7986_17190# 0.484f
C8885 m3_8892_1078# VDD 0.0157f
C8886 vcm a_23350_3174# 0.155f
C8887 row_n[9] a_29070_11166# 0.282f
C8888 col[26] a_2275_17214# 0.0899f
C8889 a_2161_6170# a_2275_6170# 0.183f
C8890 a_2475_6170# a_2966_6146# 0.317f
C8891 m2_1732_10986# vcm 0.316f
C8892 rowon_n[13] a_28978_15182# 0.118f
C8893 col[31] a_2275_6170# 0.0899f
C8894 vcm a_14010_12170# 0.56f
C8895 a_2275_11190# a_24354_11206# 0.144f
C8896 a_2475_11190# a_26970_11166# 0.264f
C8897 VDD a_10906_2130# 0.181f
C8898 col[29] rowoff_n[14] 0.0901f
C8899 row_n[11] a_16322_13214# 0.0117f
C8900 a_25054_16186# a_25358_16226# 0.0931f
C8901 a_25966_16186# a_26458_16548# 0.0658f
C8902 col_n[12] rowoff_n[10] 0.0471f
C8903 m2_24824_18014# m3_24956_18146# 3.79f
C8904 col[19] a_22042_10162# 0.367f
C8905 a_32082_4138# a_33086_4138# 0.843f
C8906 col[26] a_28978_12170# 0.0682f
C8907 col_n[1] a_2275_3158# 0.113f
C8908 row_n[1] a_26362_3174# 0.0117f
C8909 row_n[13] a_6890_15182# 0.0437f
C8910 vcm a_4274_6186# 0.155f
C8911 rowoff_n[12] a_34490_14540# 0.0133f
C8912 a_2275_8178# a_17934_8154# 0.136f
C8913 m2_11196_13422# a_10998_13174# 0.165f
C8914 vcm a_29070_16186# 0.56f
C8915 a_21950_13174# a_22042_13174# 0.326f
C8916 VDD a_25966_6146# 0.181f
C8917 col_n[16] a_2475_13198# 0.0531f
C8918 row_n[3] a_16930_5142# 0.0437f
C8919 col_n[21] a_2475_2154# 0.0531f
C8920 col_n[14] a_17326_10202# 0.084f
C8921 rowon_n[7] a_16018_9158# 0.248f
C8922 rowoff_n[6] a_5886_8154# 0.202f
C8923 m2_34864_3958# m2_35292_4386# 0.165f
C8924 a_23046_6146# a_23046_5142# 0.843f
C8925 a_2475_5166# a_9994_5142# 0.316f
C8926 m2_28840_946# m3_27968_1078# 0.0341f
C8927 m2_30272_9406# a_30074_9158# 0.165f
C8928 vcm col_n[26] 1.94f
C8929 col_n[25] a_28466_4500# 0.0283f
C8930 VDD col_n[29] 5.17f
C8931 vcm a_19334_10202# 0.155f
C8932 col[13] rowoff_n[15] 0.0901f
C8933 col[6] a_2475_10186# 0.136f
C8934 a_16930_10162# a_17326_10202# 0.0313f
C8935 rowoff_n[15] a_16018_17190# 0.294f
C8936 a_2275_10186# a_32994_10162# 0.136f
C8937 rowoff_n[4] a_14922_6146# 0.202f
C8938 ctop a_32082_5142# 4.11f
C8939 VDD a_6890_9158# 0.181f
C8940 m2_1732_9982# m3_1864_10114# 3.79f
C8941 col_n[13] a_2275_16210# 0.113f
C8942 m2_6176_15430# row_n[13] 0.0128f
C8943 col[8] a_10998_8154# 0.367f
C8944 m2_12200_11414# row_n[9] 0.0128f
C8945 m2_18224_7398# row_n[5] 0.0128f
C8946 col_n[18] a_2275_5166# 0.113f
C8947 m2_24248_3382# row_n[1] 0.0128f
C8948 vcm a_12914_4138# 0.1f
C8949 a_13006_7150# a_14010_7150# 0.843f
C8950 a_2475_7174# a_25054_7150# 0.316f
C8951 rowoff_n[2] a_23958_4138# 0.202f
C8952 rowoff_n[9] a_6378_11528# 0.0133f
C8953 col[15] a_17934_10162# 0.0682f
C8954 m2_1732_10986# a_1957_11190# 0.245f
C8955 vcm a_35398_14218# 0.161f
C8956 col_n[23] a_26058_4138# 0.251f
C8957 VDD a_32482_4500# 0.0779f
C8958 col_n[0] a_3270_16226# 0.084f
C8959 ctop a_13006_8154# 4.11f
C8960 col_n[30] a_32994_6146# 0.0765f
C8961 col[3] a_2275_13198# 0.0899f
C8962 VDD a_21950_13174# 0.181f
C8963 col[8] a_2275_2154# 0.0899f
C8964 row_n[8] a_24354_10202# 0.0117f
C8965 col_n[3] a_6282_8194# 0.084f
C8966 rowoff_n[0] a_32994_2130# 0.202f
C8967 rowoff_n[7] a_15414_9520# 0.0133f
C8968 a_2275_4162# a_16018_4138# 0.399f
C8969 m3_34996_9110# ctop 0.209f
C8970 m2_21236_7398# a_21038_7150# 0.165f
C8971 a_30378_1166# col_n[27] 0.084f
C8972 m2_33284_16434# row_n[14] 0.0128f
C8973 vcm a_27974_8154# 0.1f
C8974 a_3970_9158# a_3970_8154# 0.843f
C8975 rowoff_n[13] a_22442_15544# 0.0133f
C8976 m2_11772_946# col[9] 0.425f
C8977 col[23] a_2475_12194# 0.136f
C8978 row_n[10] a_14922_12170# 0.0437f
C8979 col_n[14] a_17422_2492# 0.0283f
C8980 vcm a_15318_17230# 0.155f
C8981 rowon_n[14] a_14010_16186# 0.248f
C8982 col[28] a_2475_1150# 0.136f
C8983 a_31990_14178# a_32386_14218# 0.0313f
C8984 VDD a_13406_7512# 0.0779f
C8985 m2_34864_2954# m3_34996_4090# 0.0341f
C8986 rowoff_n[5] a_24450_7512# 0.0133f
C8987 col_n[24] a_27462_14540# 0.0283f
C8988 ctop a_28066_12170# 4.11f
C8989 a_2275_18218# a_16322_18234# 0.145f
C8990 row_n[0] a_24962_2130# 0.0437f
C8991 VDD a_2161_16210# 0.187f
C8992 a_2475_1150# a_8898_1126# 0.264f
C8993 row_n[12] a_2966_14178# 0.281f
C8994 a_2275_1150# a_6282_1166# 0.145f
C8995 rowon_n[4] a_24050_6146# 0.248f
C8996 col_n[30] a_2275_18218# 0.113f
C8997 a_16018_6146# a_16322_6186# 0.0931f
C8998 a_16930_6146# a_17422_6508# 0.0658f
C8999 a_2275_6170# a_31078_6146# 0.399f
C9000 vcm a_8898_11166# 0.1f
C9001 rowoff_n[3] a_33486_5504# 0.0133f
C9002 m2_2736_18014# col_n[0] 0.243f
C9003 a_28066_11166# a_29070_11166# 0.843f
C9004 VDD a_4974_1126# 0.0349f
C9005 col[4] a_6890_8154# 0.0682f
C9006 a_2275_15206# a_9902_15182# 0.136f
C9007 VDD a_28466_11528# 0.0779f
C9008 m2_4744_18014# col[2] 0.347f
C9009 a_30986_1126# col[28] 0.0682f
C9010 col_n[12] a_15014_2130# 0.251f
C9011 col[20] a_2275_15206# 0.0899f
C9012 ctop a_8990_15182# 4.11f
C9013 row_n[4] a_2475_6170# 0.405f
C9014 col_n[22] a_25054_14178# 0.251f
C9015 col[25] a_2275_4162# 0.0899f
C9016 col_n[19] a_21950_4138# 0.0765f
C9017 a_12914_3134# a_13006_3134# 0.326f
C9018 a_2275_3158# a_21342_3174# 0.144f
C9019 a_2475_3158# a_23958_3134# 0.264f
C9020 rowoff_n[8] a_25054_10162# 0.294f
C9021 m2_12200_5390# a_12002_5142# 0.165f
C9022 col_n[29] a_31990_16186# 0.0765f
C9023 row_n[13] a_35094_15182# 0.0123f
C9024 rowoff_n[11] a_28978_13174# 0.202f
C9025 col_n[2] a_5278_18234# 0.084f
C9026 col_n[0] a_2966_8154# 0.251f
C9027 vcm a_23958_15182# 0.1f
C9028 a_19030_13174# a_19030_12170# 0.843f
C9029 VDD a_20034_5142# 0.483f
C9030 a_35002_1126# VDD 0.482f
C9031 col_n[30] rowoff_n[0] 0.0471f
C9032 col_n[31] rowoff_n[1] 0.0471f
C9033 row_n[15] a_22346_17230# 0.0117f
C9034 a_2275_17214# a_24962_17190# 0.136f
C9035 a_12914_17190# a_13310_17230# 0.0313f
C9036 rowoff_n[6] a_34090_8154# 0.294f
C9037 VDD a_9390_14540# 0.0779f
C9038 col_n[13] a_16418_12532# 0.0283f
C9039 col_n[16] a_2475_18218# 0.0529f
C9040 a_2966_5142# a_2966_4138# 0.843f
C9041 row_n[5] a_32386_7190# 0.0117f
C9042 col_n[10] a_2475_11190# 0.0531f
C9043 m3_30980_1078# m3_31984_1078# 0.202f
C9044 a_35002_1126# a_35094_1126# 0.0991f
C9045 a_31078_10162# a_31382_10202# 0.0931f
C9046 rowoff_n[14] a_10394_16548# 0.0133f
C9047 a_31990_10162# a_32482_10524# 0.0658f
C9048 vcm a_4882_18194# 0.101f
C9049 a_2475_14202# a_17022_14178# 0.316f
C9050 m2_15788_946# a_15926_1126# 0.225f
C9051 a_8990_14178# a_9994_14178# 0.843f
C9052 row_n[7] a_22954_9158# 0.0437f
C9053 m2_1732_6970# m3_1864_7102# 3.79f
C9054 rowon_n[11] a_22042_13174# 0.248f
C9055 col[3] a_5886_18194# 0.0682f
C9056 VDD a_24450_18556# 0.0858f
C9057 a_2275_2154# a_29982_2130# 0.136f
C9058 col[0] a_2475_8178# 0.148f
C9059 col_n[11] a_14010_12170# 0.251f
C9060 m3_4876_18146# VDD 0.0277f
C9061 vcm a_6982_3134# 0.56f
C9062 col_n[8] a_10906_2130# 0.0765f
C9063 rowon_n[1] a_32082_3134# 0.248f
C9064 a_27974_7150# a_28066_7150# 0.326f
C9065 m2_20808_18014# col_n[18] 0.243f
C9066 col_n[18] a_20946_14178# 0.0765f
C9067 a_2275_11190# a_7986_11166# 0.399f
C9068 col_n[23] rowoff_n[10] 0.0471f
C9069 m2_15788_18014# a_16018_18194# 0.0249f
C9070 col_n[7] a_2275_14202# 0.113f
C9071 a_2475_16210# a_32082_16186# 0.316f
C9072 a_34090_17190# a_34090_16186# 0.843f
C9073 VDD a_16018_12170# 0.483f
C9074 col_n[12] a_2275_3158# 0.113f
C9075 sample a_1957_18218# 0.345f
C9076 m2_1046_19620# m3_1046_19620# 0.25f
C9077 m2_2160_10410# rowon_n[8] 0.0219f
C9078 m2_8184_6394# rowon_n[4] 0.0322f
C9079 m2_13204_2378# rowon_n[0] 0.0322f
C9080 a_22954_4138# a_23350_4178# 0.0313f
C9081 col_n[2] a_5374_10524# 0.0283f
C9082 row_n[1] a_9994_3134# 0.282f
C9083 rowon_n[5] a_9902_7150# 0.118f
C9084 vcm a_22042_7150# 0.56f
C9085 rowoff_n[12] a_16930_14178# 0.202f
C9086 col_n[27] a_2475_13198# 0.0531f
C9087 col[31] a_34090_11166# 0.367f
C9088 a_12002_13174# a_12306_13214# 0.0931f
C9089 a_2275_13198# a_23046_13174# 0.399f
C9090 a_12914_13174# a_13406_13536# 0.0658f
C9091 VDD a_31078_16186# 0.483f
C9092 row_n[12] a_30378_14218# 0.0117f
C9093 a_19030_1126# a_20034_1126# 0.843f
C9094 col_n[3] rowon_n[14] 0.111f
C9095 col_n[5] rowon_n[15] 0.111f
C9096 col_n[1] rowon_n[13] 0.111f
C9097 vcm row_n[13] 0.616f
C9098 VDD rowon_n[11] 3.04f
C9099 sample row_n[12] 0.423f
C9100 col_n[2] row_n[14] 0.298f
C9101 col_n[18] col_n[19] 0.0101f
C9102 col_n[4] row_n[15] 0.298f
C9103 col_n[0] rowon_n[12] 0.111f
C9104 col[24] rowoff_n[15] 0.0901f
C9105 col[17] a_2475_10186# 0.136f
C9106 col[28] col[29] 0.0355f
C9107 vcm a_12306_1166# 0.16f
C9108 m2_23244_15430# rowon_n[13] 0.0322f
C9109 m2_29268_11414# rowon_n[9] 0.0322f
C9110 m2_34864_6970# rowon_n[5] 0.231f
C9111 vcm a_2874_10162# 0.1f
C9112 col_n[26] a_29374_11206# 0.084f
C9113 col_n[7] rowoff_n[11] 0.0471f
C9114 a_8898_10162# a_8990_10162# 0.326f
C9115 a_2275_10186# a_13310_10202# 0.144f
C9116 a_2475_10186# a_15926_10162# 0.264f
C9117 row_n[14] a_20946_16186# 0.0437f
C9118 m2_3164_16434# a_2966_16186# 0.165f
C9119 col_n[7] a_9902_12170# 0.0765f
C9120 col_n[24] a_2275_16210# 0.113f
C9121 row_n[4] a_30986_6146# 0.0437f
C9122 col_n[29] a_2275_5166# 0.113f
C9123 a_9994_3134# a_9994_2130# 0.843f
C9124 rowon_n[8] a_30074_10162# 0.248f
C9125 m2_34864_10986# rowoff_n[9] 0.278f
C9126 vcm a_27366_5182# 0.155f
C9127 a_2275_7174# a_6890_7150# 0.136f
C9128 m2_15788_18014# vcm 0.353f
C9129 vcm a_18026_14178# 0.56f
C9130 a_2275_12194# a_28370_12210# 0.144f
C9131 a_2475_12194# a_30986_12170# 0.264f
C9132 col[14] a_2275_13198# 0.0899f
C9133 VDD a_14922_4138# 0.181f
C9134 col[19] a_2275_2154# 0.0899f
C9135 col[20] a_23046_9158# 0.367f
C9136 a_27062_17190# a_27366_17230# 0.0931f
C9137 row_n[0] m2_29268_2378# 0.0128f
C9138 a_27974_17190# a_28466_17552# 0.0658f
C9139 VDD a_3878_13174# 0.181f
C9140 row_n[8] a_7986_10162# 0.282f
C9141 col[27] a_29982_11166# 0.0682f
C9142 rowon_n[12] a_7894_14178# 0.118f
C9143 a_33998_5142# a_34394_5182# 0.0313f
C9144 m2_25828_946# ctop 0.0428f
C9145 vcm a_8290_8194# 0.155f
C9146 m2_26832_18014# m2_27836_18014# 0.843f
C9147 rowoff_n[13] a_4882_15182# 0.202f
C9148 a_2275_9182# a_21950_9158# 0.136f
C9149 rowon_n[2] a_17934_4138# 0.118f
C9150 vcm a_33086_18194# 0.165f
C9151 ctop a_21038_3134# 4.11f
C9152 col_n[15] a_18330_9198# 0.084f
C9153 a_23958_14178# a_24050_14178# 0.326f
C9154 VDD a_29982_8154# 0.181f
C9155 m2_1732_3958# m3_1864_4090# 3.79f
C9156 rowoff_n[5] a_6890_7150# 0.202f
C9157 row_n[0] a_5278_2170# 0.0117f
C9158 col_n[4] a_2475_9182# 0.0531f
C9159 vcm a_34394_3174# 0.155f
C9160 col_n[26] a_29470_3496# 0.0283f
C9161 a_2475_6170# a_14010_6146# 0.316f
C9162 a_25054_7150# a_25054_6146# 0.843f
C9163 vcm a_23350_12210# 0.155f
C9164 rowoff_n[3] a_15926_5142# 0.202f
C9165 a_18938_11166# a_19334_11206# 0.0313f
C9166 VDD a_21438_2492# 0.0779f
C9167 m2_33860_18014# a_34394_18234# 0.087f
C9168 m2_34864_18014# a_35094_18194# 0.0249f
C9169 m2_1732_8978# row_n[7] 0.292f
C9170 col[31] a_2275_15206# 0.0899f
C9171 ctop a_2475_6170# 0.0488f
C9172 m2_7180_5390# row_n[3] 0.0128f
C9173 row_n[11] a_28978_13174# 0.0437f
C9174 VDD a_10906_11166# 0.181f
C9175 rowon_n[15] a_28066_17190# 0.248f
C9176 col[9] a_12002_7150# 0.367f
C9177 a_3878_3134# a_3970_3134# 0.326f
C9178 a_2874_3134# a_3270_3174# 0.0313f
C9179 a_2275_3158# a_4974_3134# 0.399f
C9180 rowoff_n[8] a_7382_10524# 0.0133f
C9181 rowoff_n[1] a_24962_3134# 0.202f
C9182 col[16] a_18938_9158# 0.0682f
C9183 m2_34864_16006# rowoff_n[14] 0.278f
C9184 vcm a_16930_6146# 0.1f
C9185 a_15014_8154# a_16018_8154# 0.843f
C9186 a_2475_8178# a_29070_8154# 0.316f
C9187 col_n[1] a_2275_12194# 0.113f
C9188 col_n[24] a_27062_3134# 0.251f
C9189 rowon_n[7] rowoff_n[7] 20.2f
C9190 col_n[6] a_2275_1150# 0.113f
C9191 vcm a_4274_15222# 0.155f
C9192 VDD a_1957_5166# 0.196f
C9193 col_n[31] a_33998_5142# 0.0765f
C9194 col_n[27] a_2475_18218# 0.0529f
C9195 ctop a_17022_10162# 4.11f
C9196 row_n[15] a_5978_17190# 0.282f
C9197 a_2475_17214# a_7894_17190# 0.264f
C9198 a_2275_17214# a_5278_17230# 0.144f
C9199 m2_22240_14426# row_n[12] 0.0128f
C9200 a_4882_17190# a_4974_17190# 0.326f
C9201 a_3878_17190# a_4274_17230# 0.0313f
C9202 col_n[4] a_7286_7190# 0.084f
C9203 m2_28264_10410# row_n[8] 0.0128f
C9204 rowoff_n[6] a_16418_8516# 0.0133f
C9205 VDD a_25966_15182# 0.181f
C9206 m2_34288_6394# row_n[4] 0.0128f
C9207 col[0] a_2966_5142# 0.367f
C9208 col_n[21] a_2475_11190# 0.0531f
C9209 row_n[5] a_16018_7150# 0.282f
C9210 a_2275_5166# a_20034_5142# 0.399f
C9211 m3_1864_4090# m3_1864_3086# 0.202f
C9212 rowon_n[9] a_15926_11166# 0.118f
C9213 vcm a_31990_10162# 0.1f
C9214 a_24962_1126# a_25454_1488# 0.0658f
C9215 a_5978_10162# a_5978_9158# 0.843f
C9216 en_C0_n a_4274_1166# 0.0266f
C9217 m2_26256_16434# a_26058_16186# 0.165f
C9218 rowoff_n[4] a_25454_6508# 0.0133f
C9219 col_n[25] a_28466_13536# 0.0283f
C9220 m3_4876_1078# a_4974_2130# 0.0302f
C9221 m2_5748_946# a_2275_1150# 0.28f
C9222 m2_26832_946# a_27062_2130# 0.843f
C9223 VDD a_17422_9520# 0.0779f
C9224 row_n[7] a_3270_9198# 0.0117f
C9225 col[11] a_2475_8178# 0.136f
C9226 ctop a_32082_14178# 4.11f
C9227 VDD a_6890_18194# 0.343f
C9228 a_2275_2154# a_10298_2170# 0.144f
C9229 a_2475_2154# a_12914_2130# 0.264f
C9230 a_18026_7150# a_18330_7190# 0.0931f
C9231 rowoff_n[2] a_34490_4500# 0.0133f
C9232 a_2275_7174# a_35094_7150# 0.0924f
C9233 rowoff_n[9] a_17022_11166# 0.294f
C9234 a_18938_7150# a_19430_7512# 0.0658f
C9235 col[8] a_10998_17190# 0.367f
C9236 col[5] a_7894_7150# 0.0682f
C9237 col_n[18] a_2275_14202# 0.113f
C9238 vcm a_12914_13174# 0.1f
C9239 a_30074_12170# a_31078_12170# 0.843f
C9240 VDD a_8990_3134# 0.483f
C9241 col_n[23] a_2275_3158# 0.113f
C9242 m2_6752_18014# a_2275_18218# 0.28f
C9243 m2_2736_18014# a_3270_18234# 0.087f
C9244 a_2275_16210# a_13918_16186# 0.136f
C9245 VDD a_32482_13536# 0.0779f
C9246 col_n[23] a_26058_13174# 0.251f
C9247 rowon_n[3] a_2874_5142# 0.118f
C9248 col_n[20] a_22954_3134# 0.0765f
C9249 ctop a_13006_17190# 4.06f
C9250 rowoff_n[7] a_26058_9158# 0.294f
C9251 col_n[30] a_32994_15182# 0.0765f
C9252 a_2275_4162# a_25358_4178# 0.144f
C9253 a_14922_4138# a_15014_4138# 0.326f
C9254 a_2475_4162# a_27974_4138# 0.264f
C9255 m3_28972_1078# ctop 0.21f
C9256 col[8] a_2275_11190# 0.0899f
C9257 col_n[3] a_6282_17230# 0.084f
C9258 rowoff_n[13] a_33086_15182# 0.294f
C9259 m2_17220_14426# a_17022_14178# 0.165f
C9260 vcm a_27974_17190# 0.1f
C9261 a_21038_14178# a_21038_13174# 0.843f
C9262 a_2966_13174# a_3270_13214# 0.0931f
C9263 a_2475_13198# a_5978_13174# 0.316f
C9264 a_3878_13174# a_4370_13536# 0.0658f
C9265 VDD a_24050_7150# 0.483f
C9266 rowoff_n[5] a_35094_7150# 0.0135f
C9267 col_n[4] rowon_n[9] 0.111f
C9268 col_n[11] row_n[13] 0.298f
C9269 col_n[12] rowon_n[13] 0.111f
C9270 sample rowon_n[6] 0.0935f
C9271 col_n[5] row_n[10] 0.298f
C9272 VDD row_n[6] 3.29f
C9273 col_n[1] row_n[8] 0.298f
C9274 col_n[15] row_n[15] 0.298f
C9275 col_n[13] row_n[14] 0.298f
C9276 col_n[7] row_n[11] 0.298f
C9277 vcm rowon_n[7] 0.65f
C9278 col_n[0] row_n[7] 0.298f
C9279 col_n[8] rowon_n[11] 0.111f
C9280 col_n[6] rowon_n[10] 0.111f
C9281 col_n[2] rowon_n[8] 0.111f
C9282 col_n[16] rowon_n[15] 0.111f
C9283 col_n[3] row_n[9] 0.298f
C9284 col_n[14] rowon_n[14] 0.111f
C9285 col_n[9] row_n[12] 0.298f
C9286 col_n[10] rowon_n[12] 0.111f
C9287 col_n[14] a_17422_11528# 0.0283f
C9288 m2_2736_18014# a_2475_18218# 0.287f
C9289 a_14922_18194# a_15318_18234# 0.0313f
C9290 a_2275_18218# a_28978_18194# 0.136f
C9291 col[28] a_2475_10186# 0.136f
C9292 VDD a_13406_16548# 0.0779f
C9293 a_9902_1126# a_10298_1166# 0.0313f
C9294 row_n[12] a_14010_14178# 0.282f
C9295 a_2275_1150# a_18938_1126# 0.138f
C9296 m2_14208_2378# a_14010_2130# 0.165f
C9297 col_n[18] rowoff_n[11] 0.0471f
C9298 vcm a_30074_2130# 0.56f
C9299 row_n[2] a_24050_4138# 0.282f
C9300 a_33086_11166# a_33390_11206# 0.0931f
C9301 a_33998_11166# a_34490_11528# 0.0658f
C9302 row_n[14] a_2275_16210# 19.2f
C9303 VDD a_14314_1166# 0.0149f
C9304 rowon_n[6] a_23958_8154# 0.118f
C9305 a_2475_15206# a_21038_15182# 0.316f
C9306 a_10998_15182# a_12002_15182# 0.843f
C9307 VDD a_4974_10162# 0.483f
C9308 col[4] a_6890_17190# 0.0682f
C9309 row_n[4] a_11302_6186# 0.0117f
C9310 col_n[12] a_15014_11166# 0.251f
C9311 a_2475_18218# a_26970_18194# 0.264f
C9312 a_2275_3158# a_33998_3134# 0.136f
C9313 col_n[9] a_11910_1126# 0.0765f
C9314 m2_1732_11990# rowoff_n[10] 0.415f
C9315 vcm a_10998_5142# 0.56f
C9316 col_n[19] a_21950_13174# 0.0765f
C9317 col[25] a_2275_13198# 0.0899f
C9318 rowoff_n[10] a_4974_12170# 0.294f
C9319 a_29982_8154# a_30074_8154# 0.326f
C9320 m2_34864_946# sw_n 0.01f
C9321 m2_21812_946# col[19] 0.425f
C9322 a_24962_1126# vcm 0.0989f
C9323 m2_8184_12418# a_7986_12170# 0.165f
C9324 col[30] a_2275_2154# 0.0899f
C9325 a_2275_12194# a_12002_12170# 0.399f
C9326 m2_19804_18014# VDD 1.06f
C9327 col_n[0] a_2966_17190# 0.251f
C9328 row_n[15] a_35002_17190# 0.0437f
C9329 a_2475_17214# a_2475_16210# 0.0666f
C9330 VDD a_20034_14178# 0.483f
C9331 col_n[2] rowoff_n[12] 0.0471f
C9332 col_n[3] a_6378_9520# 0.0283f
C9333 rowon_n[0] a_10998_2130# 0.248f
C9334 a_24962_5142# a_25358_5182# 0.0313f
C9335 m2_27260_8402# a_27062_8154# 0.165f
C9336 vcm a_26058_9158# 0.56f
C9337 rowoff_n[14] a_21038_16186# 0.294f
C9338 a_2874_9158# a_3366_9520# 0.0658f
C9339 a_2275_9182# a_3878_9158# 0.136f
C9340 a_2475_9182# a_4882_9158# 0.264f
C9341 ctop a_2966_3134# 4.02f
C9342 col_n[15] a_2475_9182# 0.0531f
C9343 a_2275_14202# a_27062_14178# 0.399f
C9344 m2_6176_17438# rowon_n[15] 0.0322f
C9345 a_14010_14178# a_14314_14218# 0.0931f
C9346 a_14922_14178# a_15414_14540# 0.0658f
C9347 m2_12200_13422# rowon_n[11] 0.0322f
C9348 m2_18224_9406# rowon_n[7] 0.0322f
C9349 m2_24248_5390# rowon_n[3] 0.0322f
C9350 VDD a_35094_18194# 0.0356f
C9351 a_21038_2130# a_22042_2130# 0.843f
C9352 row_n[9] a_22042_11166# 0.282f
C9353 vcm a_16322_3174# 0.155f
C9354 col_n[1] a_3970_9158# 0.251f
C9355 col_n[27] a_30378_10202# 0.084f
C9356 col[0] a_2475_17214# 0.148f
C9357 rowon_n[13] a_21950_15182# 0.118f
C9358 col[5] a_2475_6170# 0.136f
C9359 vcm a_6982_12170# 0.56f
C9360 col_n[8] a_10906_11166# 0.0765f
C9361 a_2275_11190# a_17326_11206# 0.144f
C9362 a_2475_11190# a_19942_11166# 0.264f
C9363 a_10906_11166# a_10998_11166# 0.326f
C9364 VDD a_3366_2492# 0.0779f
C9365 m2_21812_18014# a_22346_18234# 0.087f
C9366 row_n[11] a_9294_13214# 0.0117f
C9367 rowon_n[3] a_31990_5142# 0.118f
C9368 m2_15788_18014# m3_14916_18146# 0.0341f
C9369 col_n[12] a_2275_12194# 0.113f
C9370 m2_1732_1950# rowoff_n[0] 0.415f
C9371 a_12002_4138# a_12002_3134# 0.843f
C9372 row_n[1] a_19334_3174# 0.0117f
C9373 row_n[4] rowoff_n[3] 0.085f
C9374 col_n[17] a_2275_1150# 0.0947f
C9375 m2_18224_6394# a_18026_6146# 0.165f
C9376 m2_1732_17010# rowoff_n[15] 0.415f
C9377 vcm a_31382_7190# 0.155f
C9378 a_5886_8154# a_6282_8194# 0.0313f
C9379 rowoff_n[12] a_27462_14540# 0.0133f
C9380 a_2275_8178# a_10906_8154# 0.136f
C9381 vcm a_22042_16186# 0.56f
C9382 col[21] a_24050_8154# 0.367f
C9383 a_2475_13198# a_35002_13174# 0.264f
C9384 a_2275_13198# a_32386_13214# 0.144f
C9385 VDD a_18938_6146# 0.181f
C9386 row_n[3] a_9902_5142# 0.0437f
C9387 rowon_n[7] a_8990_9158# 0.248f
C9388 col[28] a_30986_10162# 0.0682f
C9389 col[2] a_2275_9182# 0.0899f
C9390 a_29982_18194# a_30474_18556# 0.0658f
C9391 a_2475_5166# a_2874_5142# 0.264f
C9392 a_1957_5166# a_2275_5166# 0.158f
C9393 m3_26964_18146# m3_27968_18146# 0.202f
C9394 vcm a_12306_10202# 0.155f
C9395 a_2275_10186# a_25966_10162# 0.136f
C9396 rowoff_n[15] a_8990_17190# 0.294f
C9397 col_n[16] a_19334_8194# 0.084f
C9398 col[22] a_2475_8178# 0.136f
C9399 rowoff_n[4] a_7894_6146# 0.202f
C9400 ctop a_25054_5142# 4.11f
C9401 a_25966_15182# a_26058_15182# 0.326f
C9402 VDD a_33998_10162# 0.181f
C9403 col_n[27] a_30474_2492# 0.0283f
C9404 m2_9188_4386# a_8990_4138# 0.165f
C9405 col_n[29] a_2275_14202# 0.113f
C9406 vcm a_5886_4138# 0.1f
C9407 rowoff_n[2] a_16930_4138# 0.202f
C9408 rowoff_n[10] a_33998_12170# 0.202f
C9409 a_2475_7174# a_18026_7150# 0.316f
C9410 a_27062_8154# a_27062_7150# 0.843f
C9411 row_n[6] a_30074_8154# 0.282f
C9412 vcm a_27366_14218# 0.155f
C9413 a_20946_12170# a_21342_12210# 0.0313f
C9414 VDD a_25454_4500# 0.0779f
C9415 rowon_n[10] a_29982_12170# 0.118f
C9416 ctop a_5978_8154# 4.11f
C9417 col[10] a_13006_6146# 0.367f
C9418 VDD a_14922_13174# 0.181f
C9419 col[19] a_2275_11190# 0.0899f
C9420 row_n[8] a_17326_10202# 0.0117f
C9421 rowoff_n[7] a_8386_9520# 0.0133f
C9422 rowoff_n[0] a_25966_2130# 0.202f
C9423 col[17] a_19942_8154# 0.0682f
C9424 a_4974_4138# a_5278_4178# 0.0931f
C9425 a_2275_4162# a_8990_4138# 0.399f
C9426 a_5886_4138# a_6378_4500# 0.0658f
C9427 m3_24956_18146# ctop 0.209f
C9428 m2_5172_16434# row_n[14] 0.0128f
C9429 col_n[25] a_28066_2130# 0.251f
C9430 m2_11196_12418# row_n[10] 0.0128f
C9431 vcm a_20946_8154# 0.1f
C9432 a_17022_9158# a_18026_9158# 0.843f
C9433 a_2475_9182# a_33086_9158# 0.316f
C9434 m2_17220_8402# row_n[6] 0.0128f
C9435 rowoff_n[13] a_15414_15544# 0.0133f
C9436 m2_23244_4386# row_n[2] 0.0128f
C9437 m2_1732_13998# a_2966_14178# 0.843f
C9438 row_n[10] a_7894_12170# 0.0437f
C9439 col_n[3] rowon_n[3] 0.111f
C9440 col_n[19] rowon_n[11] 0.111f
C9441 col_n[24] row_n[14] 0.298f
C9442 sample row_n[1] 0.423f
C9443 col_n[12] row_n[8] 0.298f
C9444 col_n[14] row_n[9] 0.298f
C9445 col_n[27] rowon_n[15] 0.111f
C9446 col_n[29] col_n[30] 0.0161f
C9447 VDD rowon_n[0] 3.04f
C9448 col_n[11] rowon_n[7] 0.111f
C9449 col_n[9] rowon_n[6] 0.111f
C9450 col_n[22] row_n[13] 0.298f
C9451 col_n[8] row_n[6] 0.298f
C9452 col_n[18] row_n[11] 0.298f
C9453 col_n[15] rowon_n[9] 0.111f
C9454 col_n[23] rowon_n[13] 0.111f
C9455 col_n[0] rowon_n[1] 0.111f
C9456 col_n[10] row_n[7] 0.298f
C9457 col_n[4] row_n[4] 0.298f
C9458 col_n[5] rowon_n[4] 0.111f
C9459 col_n[13] rowon_n[8] 0.111f
C9460 col_n[16] row_n[10] 0.298f
C9461 col_n[26] row_n[15] 0.298f
C9462 col_n[1] rowon_n[2] 0.111f
C9463 col_n[25] rowon_n[14] 0.111f
C9464 vcm row_n[2] 0.616f
C9465 col_n[17] rowon_n[10] 0.111f
C9466 col_n[2] row_n[3] 0.298f
C9467 col_n[20] row_n[12] 0.298f
C9468 col_n[7] rowon_n[5] 0.111f
C9469 col_n[6] row_n[5] 0.298f
C9470 col_n[21] rowon_n[12] 0.111f
C9471 vcm a_8290_17230# 0.155f
C9472 rowon_n[14] a_6982_16186# 0.248f
C9473 VDD a_6378_7512# 0.0779f
C9474 rowoff_n[5] a_17422_7512# 0.0133f
C9475 col_n[5] a_8290_6186# 0.084f
C9476 ctop a_21038_12170# 4.11f
C9477 col_n[29] rowoff_n[11] 0.0471f
C9478 a_6890_18194# a_6982_18194# 0.0991f
C9479 a_2275_18218# a_9294_18234# 0.145f
C9480 col_n[15] a_18330_18234# 0.084f
C9481 row_n[0] a_17934_2130# 0.0437f
C9482 VDD a_29982_17190# 0.181f
C9483 rowon_n[4] a_17022_6146# 0.248f
C9484 a_2275_6170# a_24050_6146# 0.399f
C9485 col_n[9] a_2475_7174# 0.0531f
C9486 vcm a_34394_12210# 0.155f
C9487 rowoff_n[3] a_26458_5504# 0.0133f
C9488 col_n[26] a_29470_12532# 0.0283f
C9489 a_7986_11166# a_7986_10162# 0.843f
C9490 VDD a_32082_2130# 0.483f
C9491 m2_32280_17438# row_n[15] 0.0128f
C9492 m2_34864_17010# a_2275_17214# 0.278f
C9493 a_2161_15206# a_2275_15206# 0.183f
C9494 a_2475_15206# a_2966_15182# 0.317f
C9495 VDD a_21438_11528# 0.0779f
C9496 ctop a_2475_15206# 0.0488f
C9497 a_2475_3158# a_16930_3134# 0.264f
C9498 a_2275_3158# a_14314_3174# 0.144f
C9499 rowoff_n[8] a_18026_10162# 0.294f
C9500 rowoff_n[1] a_35494_3496# 0.0133f
C9501 col[9] a_12002_16186# 0.367f
C9502 a_30074_1126# a_2475_1150# 0.0299f
C9503 row_n[13] a_28066_15182# 0.282f
C9504 col[6] a_8898_6146# 0.0682f
C9505 a_20946_8154# a_21438_8516# 0.0658f
C9506 rowoff_n[11] a_21950_13174# 0.202f
C9507 a_20034_8154# a_20338_8194# 0.0931f
C9508 col[16] a_18938_18194# 0.0682f
C9509 vcm a_16930_15182# 0.1f
C9510 a_32082_13174# a_33086_13174# 0.843f
C9511 VDD a_13006_5142# 0.483f
C9512 col_n[24] a_27062_12170# 0.251f
C9513 col_n[13] rowoff_n[12] 0.0471f
C9514 a_26970_1126# VDD 0.405f
C9515 col_n[6] a_2275_10186# 0.113f
C9516 col_n[21] a_23958_2130# 0.0765f
C9517 row_n[15] a_15318_17230# 0.0117f
C9518 a_2275_17214# a_17934_17190# 0.136f
C9519 rowoff_n[6] a_27062_8154# 0.294f
C9520 VDD a_1957_14202# 0.196f
C9521 col_n[31] a_33998_14178# 0.0765f
C9522 m3_24956_18146# a_25054_17190# 0.0303f
C9523 col_n[4] a_7286_16226# 0.084f
C9524 a_2275_5166# a_29374_5182# 0.144f
C9525 row_n[5] a_25358_7190# 0.0117f
C9526 a_16930_5142# a_17022_5142# 0.326f
C9527 a_2475_5166# a_31990_5142# 0.264f
C9528 col[0] a_2966_14178# 0.367f
C9529 m3_16924_1078# m3_17928_1078# 0.202f
C9530 col_n[26] a_2475_9182# 0.0531f
C9531 rowoff_n[14] a_2966_16186# 0.294f
C9532 m2_34864_16006# a_35002_16186# 0.225f
C9533 a_23046_15182# a_23046_14178# 0.843f
C9534 m2_10768_946# a_10998_1126# 0.0249f
C9535 m2_28840_946# a_2275_1150# 0.28f
C9536 a_2475_14202# a_9994_14178# 0.316f
C9537 col_n[15] a_18426_10524# 0.0283f
C9538 row_n[7] a_15926_9158# 0.0437f
C9539 VDD a_28066_9158# 0.483f
C9540 rowon_n[11] a_15014_13174# 0.248f
C9541 VDD a_17422_18556# 0.0858f
C9542 col[11] a_2475_17214# 0.136f
C9543 a_2275_2154# a_22954_2130# 0.136f
C9544 a_11910_2130# a_12306_2170# 0.0313f
C9545 col[16] a_2475_6170# 0.136f
C9546 m2_23244_1374# VDD 0.0194f
C9547 vcm a_34090_4138# 0.56f
C9548 m3_34568_1078# col_n[31] 0.0456f
C9549 rowon_n[1] a_25054_3134# 0.248f
C9550 rowon_n[13] a_3878_15182# 0.118f
C9551 col_n[0] a_2874_6146# 0.0765f
C9552 VDD rowoff_n[13] 1.51f
C9553 col[5] a_7894_16186# 0.0682f
C9554 a_2475_16210# a_25054_16186# 0.316f
C9555 m3_34996_6098# a_34090_6146# 0.0303f
C9556 a_13006_16186# a_14010_16186# 0.843f
C9557 VDD a_8990_12170# 0.483f
C9558 col_n[23] a_2275_12194# 0.113f
C9559 col_n[13] a_16018_10162# 0.251f
C9560 col[0] rowoff_n[9] 0.0901f
C9561 ctop rowoff_n[3] 0.177f
C9562 row_n[0] rowoff_n[0] 0.209f
C9563 col_n[28] a_2275_1150# 0.113f
C9564 col_n[20] a_22954_12170# 0.0765f
C9565 row_n[1] a_2874_3134# 0.0436f
C9566 vcm a_15014_7150# 0.56f
C9567 rowon_n[5] a_2161_7174# 0.0177f
C9568 rowoff_n[12] a_9902_14178# 0.202f
C9569 a_31990_9158# a_32082_9158# 0.326f
C9570 col[13] a_2275_9182# 0.0899f
C9571 m2_1732_13998# sample 0.2f
C9572 a_2275_13198# a_16018_13174# 0.399f
C9573 m2_34864_7974# ctop 0.0422f
C9574 col_n[4] a_7382_8516# 0.0283f
C9575 VDD a_24050_16186# 0.483f
C9576 row_n[12] a_23350_14218# 0.0117f
C9577 a_31478_1488# col_n[28] 0.0283f
C9578 vcm a_5278_1166# 0.16f
C9579 a_26970_6146# a_27366_6186# 0.0313f
C9580 m2_1732_10986# rowon_n[9] 0.236f
C9581 m2_7180_7398# rowon_n[5] 0.0322f
C9582 m2_13204_3382# rowon_n[1] 0.0322f
C9583 vcm a_30074_11166# 0.56f
C9584 row_n[2] a_33390_4178# 0.0117f
C9585 a_2275_10186# a_6282_10202# 0.144f
C9586 a_2475_10186# a_8898_10162# 0.264f
C9587 row_n[14] a_13918_16186# 0.0437f
C9588 m2_32280_17438# a_32082_17190# 0.165f
C9589 a_2275_15206# a_31078_15182# 0.399f
C9590 a_16930_15182# a_17422_15544# 0.0658f
C9591 a_16018_15182# a_16322_15222# 0.0931f
C9592 row_n[4] a_23958_6146# 0.0437f
C9593 col_n[3] a_2475_5166# 0.0531f
C9594 a_23046_3134# a_24050_3134# 0.843f
C9595 rowon_n[8] a_23046_10162# 0.248f
C9596 col_n[2] a_4974_8154# 0.251f
C9597 col_n[28] a_31382_9198# 0.084f
C9598 vcm a_20338_5182# 0.155f
C9599 a_35002_8154# a_35398_8194# 0.0313f
C9600 col_n[9] a_11910_10162# 0.0765f
C9601 m2_1732_18014# vcm 0.32f
C9602 m2_22240_16434# rowon_n[14] 0.0322f
C9603 m2_28264_12418# rowon_n[10] 0.0322f
C9604 m2_34288_8402# rowon_n[6] 0.0322f
C9605 vcm a_10998_14178# 0.56f
C9606 a_2475_12194# a_23958_12170# 0.264f
C9607 a_12914_12170# a_13006_12170# 0.326f
C9608 a_2275_12194# a_21342_12210# 0.144f
C9609 VDD a_7894_4138# 0.181f
C9610 col[30] a_2275_11190# 0.0899f
C9611 a_14010_5142# a_14010_4138# 0.843f
C9612 col_n[16] rowon_n[4] 0.111f
C9613 col_n[31] row_n[12] 0.298f
C9614 col_n[3] a_6378_18556# 0.0283f
C9615 col_n[29] row_n[11] 0.298f
C9616 m2_34864_7974# a_35398_8194# 0.087f
C9617 col_n[11] row_n[2] 0.298f
C9618 col_n[8] rowon_n[0] 0.111f
C9619 col_n[20] rowon_n[6] 0.111f
C9620 col_n[9] row_n[1] 0.298f
C9621 col_n[24] rowon_n[8] 0.111f
C9622 col_n[25] row_n[9] 0.298f
C9623 col_n[28] rowon_n[10] 0.111f
C9624 col_n[27] row_n[10] 0.298f
C9625 col_n[30] rowon_n[11] 0.111f
C9626 col_n[12] rowon_n[2] 0.111f
C9627 col_n[23] row_n[8] 0.298f
C9628 col_n[21] row_n[7] 0.298f
C9629 col_n[22] rowon_n[7] 0.111f
C9630 col_n[10] rowon_n[1] 0.111f
C9631 col_n[4] ctop 0.0594f
C9632 col_n[13] row_n[3] 0.298f
C9633 rowon_n[14] rowon_n[13] 0.0632f
C9634 vcm en_bit_n[0] 0.0193f
C9635 col_n[18] rowon_n[5] 0.111f
C9636 col_n[14] rowon_n[3] 0.111f
C9637 col_n[15] row_n[4] 0.298f
C9638 col_n[26] rowon_n[9] 0.111f
C9639 VDD col[1] 3.83f
C9640 col_n[19] row_n[6] 0.298f
C9641 col_n[17] row_n[5] 0.298f
C9642 col_n[7] row_n[0] 0.298f
C9643 vcm a_2275_8178# 6.49f
C9644 m2_19804_18014# m2_20808_18014# 0.843f
C9645 a_2275_9182# a_14922_9158# 0.136f
C9646 a_7894_9158# a_8290_9198# 0.0313f
C9647 col[22] a_25054_7150# 0.367f
C9648 m2_23244_15430# a_23046_15182# 0.165f
C9649 rowon_n[2] a_10906_4138# 0.118f
C9650 rowon_n[11] rowoff_n[11] 20.2f
C9651 vcm a_26058_18194# 0.165f
C9652 ctop a_14010_3134# 4.11f
C9653 a_2966_14178# a_2966_13174# 0.843f
C9654 VDD a_22954_8154# 0.181f
C9655 col[29] a_31990_9158# 0.0682f
C9656 ctop a_2966_12170# 4.06f
C9657 a_26058_2130# a_26362_2170# 0.0931f
C9658 a_26970_2130# a_27462_2492# 0.0658f
C9659 col_n[20] a_2475_7174# 0.0531f
C9660 m3_23952_1078# VDD 0.0157f
C9661 m2_1732_6970# m2_2160_7398# 0.165f
C9662 row_n[9] a_31382_11206# 0.0117f
C9663 vcm a_28978_3134# 0.1f
C9664 a_3970_6146# a_4974_6146# 0.843f
C9665 a_2475_6170# a_6982_6146# 0.316f
C9666 col_n[17] a_20338_7190# 0.084f
C9667 rowoff_n[3] a_8898_5142# 0.202f
C9668 vcm a_16322_12210# 0.155f
C9669 a_2275_11190# a_29982_11166# 0.136f
C9670 VDD a_14410_2492# 0.0779f
C9671 col[5] a_2475_15206# 0.136f
C9672 ctop a_29070_7150# 4.11f
C9673 row_n[11] a_21950_13174# 0.0437f
C9674 a_27974_16186# a_28066_16186# 0.326f
C9675 col[10] a_2475_4162# 0.136f
C9676 VDD a_3366_11528# 0.0779f
C9677 a_24962_1126# col_n[22] 0.0765f
C9678 m2_29844_18014# m3_29976_18146# 3.79f
C9679 rowon_n[15] a_21038_17190# 0.248f
C9680 row_n[1] a_31990_3134# 0.0437f
C9681 rowoff_n[1] a_17934_3134# 0.202f
C9682 vcm a_9902_6146# 0.1f
C9683 rowon_n[5] a_31078_7150# 0.248f
C9684 rowoff_n[11] a_3878_13174# 0.202f
C9685 a_2475_8178# a_22042_8154# 0.316f
C9686 a_29070_9158# a_29070_8154# 0.843f
C9687 col_n[17] a_2275_10186# 0.113f
C9688 m2_14208_13422# a_14010_13174# 0.165f
C9689 col_n[24] rowoff_n[12] 0.0471f
C9690 vcm a_31382_16226# 0.155f
C9691 a_22954_13174# a_23350_13214# 0.0313f
C9692 VDD a_29470_6508# 0.0779f
C9693 col[11] a_14010_5142# 0.367f
C9694 ctop a_9994_10162# 4.11f
C9695 col[21] a_24050_17190# 0.367f
C9696 rowoff_n[6] a_9390_8516# 0.0133f
C9697 VDD a_18938_15182# 0.181f
C9698 m2_6176_6394# row_n[4] 0.0128f
C9699 col[18] a_20946_7150# 0.0682f
C9700 m2_11196_2378# row_n[0] 0.0128f
C9701 col[2] a_2275_18218# 0.0899f
C9702 row_n[5] a_8990_7150# 0.282f
C9703 a_2275_5166# a_13006_5142# 0.399f
C9704 a_7894_5142# a_8386_5504# 0.0658f
C9705 col[7] a_2275_7174# 0.0899f
C9706 a_6982_5142# a_7286_5182# 0.0931f
C9707 m2_33284_9406# a_33086_9158# 0.165f
C9708 m3_1864_11118# m3_1864_10114# 0.202f
C9709 m2_33860_946# m3_32988_1078# 0.0341f
C9710 rowon_n[9] a_8898_11166# 0.118f
C9711 vcm a_24962_10162# 0.1f
C9712 a_19030_10162# a_20034_10162# 0.843f
C9713 rowoff_n[4] a_18426_6508# 0.0133f
C9714 col_n[6] a_9294_5182# 0.084f
C9715 m2_33860_946# analog_in 1.11f
C9716 VDD a_10394_9520# 0.0779f
C9717 m2_29844_18014# ctop 0.0422f
C9718 col_n[16] a_19334_17230# 0.084f
C9719 col[22] a_2475_17214# 0.136f
C9720 col[27] a_2475_6170# 0.136f
C9721 ctop a_25054_14178# 4.11f
C9722 m2_21236_15430# row_n[13] 0.0128f
C9723 a_2475_2154# a_5886_2130# 0.264f
C9724 a_2275_2154# a_3270_2170# 0.145f
C9725 m2_27260_11414# row_n[9] 0.0128f
C9726 m2_33284_7398# row_n[5] 0.0128f
C9727 m2_34864_10986# m2_34864_9982# 0.843f
C9728 col_n[8] rowoff_n[13] 0.0471f
C9729 rowoff_n[2] a_27462_4500# 0.0133f
C9730 a_2275_7174# a_28066_7150# 0.399f
C9731 col_n[27] a_30474_11528# 0.0283f
C9732 rowoff_n[9] a_9994_11166# 0.294f
C9733 m2_5172_11414# a_4974_11166# 0.165f
C9734 vcm a_5886_13174# 0.1f
C9735 a_9994_12170# a_9994_11166# 0.843f
C9736 VDD a_2475_3158# 26.1f
C9737 col[9] rowoff_n[7] 0.0901f
C9738 col[3] rowoff_n[1] 0.0901f
C9739 col[4] rowoff_n[2] 0.0901f
C9740 col[6] rowoff_n[4] 0.0901f
C9741 col[11] rowoff_n[9] 0.0901f
C9742 col[2] rowoff_n[0] 0.0901f
C9743 col[8] rowoff_n[6] 0.0901f
C9744 col[7] rowoff_n[5] 0.0901f
C9745 col[5] rowoff_n[3] 0.0901f
C9746 col[10] rowoff_n[8] 0.0901f
C9747 a_2275_16210# a_6890_16186# 0.136f
C9748 VDD a_25454_13536# 0.0779f
C9749 col[0] a_2874_3134# 0.0682f
C9750 row_n[8] a_29982_10162# 0.0437f
C9751 ctop a_5978_17190# 4.06f
C9752 rowoff_n[7] a_19030_9158# 0.294f
C9753 col[10] a_13006_15182# 0.367f
C9754 rowon_n[12] a_29070_14178# 0.248f
C9755 col[7] a_9902_5142# 0.0682f
C9756 a_2475_4162# a_20946_4138# 0.264f
C9757 a_2275_4162# a_18330_4178# 0.144f
C9758 m3_34996_2082# ctop 0.209f
C9759 m2_24248_7398# a_24050_7150# 0.165f
C9760 col[17] a_19942_17190# 0.0682f
C9761 col[24] a_2275_9182# 0.0899f
C9762 rowoff_n[13] a_26058_15182# 0.294f
C9763 a_22042_9158# a_22346_9198# 0.0931f
C9764 a_22954_9158# a_23446_9520# 0.0658f
C9765 col_n[25] a_28066_11166# 0.251f
C9766 vcm a_20946_17190# 0.1f
C9767 a_33998_14178# a_34394_14218# 0.0313f
C9768 VDD a_17022_7150# 0.483f
C9769 rowoff_n[5] a_28066_7150# 0.294f
C9770 a_2275_18218# a_21950_18194# 0.136f
C9771 VDD a_6378_16548# 0.0779f
C9772 col_n[5] a_8290_15222# 0.084f
C9773 a_2275_1150# a_11910_1126# 0.136f
C9774 row_n[12] a_6982_14178# 0.282f
C9775 vcm a_23046_2130# 0.56f
C9776 a_18938_6146# a_19030_6146# 0.326f
C9777 a_2275_6170# a_33390_6186# 0.144f
C9778 row_n[2] a_17022_4138# 0.282f
C9779 VDD a_7286_1166# 0.0149f
C9780 col_n[16] a_19430_9520# 0.0283f
C9781 col_n[9] a_2475_16210# 0.0531f
C9782 rowon_n[6] a_16930_8154# 0.118f
C9783 col_n[14] a_2475_5166# 0.0531f
C9784 a_25054_16186# a_25054_15182# 0.843f
C9785 a_2475_15206# a_14010_15182# 0.316f
C9786 VDD a_32082_11166# 0.483f
C9787 row_n[4] a_4274_6186# 0.0117f
C9788 a_2275_3158# a_26970_3134# 0.136f
C9789 a_13918_3134# a_14314_3174# 0.0313f
C9790 a_2475_18218# a_19942_18194# 0.264f
C9791 m2_15212_5390# a_15014_5142# 0.165f
C9792 vcm a_3970_5142# 0.56f
C9793 rowoff_n[11] a_32482_13536# 0.0133f
C9794 col[4] a_2475_2154# 0.136f
C9795 m2_1732_11990# a_2275_12194# 0.191f
C9796 col[6] a_8898_15182# 0.0682f
C9797 a_3878_12170# a_3970_12170# 0.326f
C9798 a_2874_12170# a_3270_12210# 0.0313f
C9799 a_2275_12194# a_4974_12170# 0.399f
C9800 m2_5748_18014# VDD 1f
C9801 col_n[14] a_17022_9158# 0.251f
C9802 row_n[15] a_27974_17190# 0.0437f
C9803 a_15014_17190# a_16018_17190# 0.843f
C9804 a_2475_17214# a_29070_17190# 0.316f
C9805 VDD a_13006_14178# 0.483f
C9806 vcm col[9] 5.46f
C9807 col_n[4] col[5] 7.13f
C9808 col_n[29] rowon_n[5] 0.111f
C9809 col_n[26] row_n[4] 0.298f
C9810 col_n[20] row_n[1] 0.298f
C9811 col_n[24] row_n[3] 0.298f
C9812 col_n[21] rowon_n[1] 0.111f
C9813 col_n[28] row_n[5] 0.298f
C9814 col_n[25] rowon_n[3] 0.111f
C9815 col_n[22] row_n[2] 0.298f
C9816 col_n[21] a_23958_11166# 0.0765f
C9817 VDD col[12] 3.83f
C9818 col_n[31] rowon_n[6] 0.111f
C9819 col_n[27] rowon_n[4] 0.111f
C9820 col_n[23] rowon_n[2] 0.111f
C9821 col_n[19] rowon_n[0] 0.111f
C9822 rowon_n[11] row_n[11] 18.9f
C9823 col_n[15] ctop 0.0624f
C9824 col_n[18] row_n[0] 0.298f
C9825 col_n[30] row_n[6] 0.298f
C9826 rowon_n[0] a_3970_2130# 0.248f
C9827 col_n[11] a_2275_8178# 0.113f
C9828 vcm a_19030_9158# 0.56f
C9829 rowoff_n[14] a_14010_16186# 0.294f
C9830 a_33998_10162# a_34090_10162# 0.326f
C9831 a_2275_14202# a_20034_14178# 0.399f
C9832 m2_16792_946# a_17326_1166# 0.087f
C9833 col_n[31] a_2475_7174# 0.0531f
C9834 col_n[5] a_8386_7512# 0.0283f
C9835 col[1] a_2275_5166# 0.0899f
C9836 VDD a_28066_18194# 0.0356f
C9837 a_2475_2154# a_34090_2130# 0.316f
C9838 m2_6176_3382# a_5978_3134# 0.165f
C9839 m3_19936_18146# VDD 0.0666f
C9840 m2_5748_946# col[3] 0.425f
C9841 vcm a_9294_3174# 0.155f
C9842 row_n[9] a_15014_11166# 0.282f
C9843 a_28978_7150# a_29374_7190# 0.0313f
C9844 rowon_n[13] a_14922_15182# 0.118f
C9845 col[16] a_2475_15206# 0.136f
C9846 vcm a_34090_13174# 0.56f
C9847 col[21] a_2475_4162# 0.136f
C9848 a_2275_11190# a_10298_11206# 0.144f
C9849 a_2475_11190# a_12914_11166# 0.264f
C9850 VDD a_30986_3134# 0.181f
C9851 col_n[0] a_2874_15182# 0.0765f
C9852 a_2275_16210# a_35094_16186# 0.0924f
C9853 a_18026_16186# a_18330_16226# 0.0931f
C9854 a_18938_16186# a_19430_16548# 0.0658f
C9855 row_n[11] a_3878_13174# 0.0437f
C9856 rowon_n[3] a_24962_5142# 0.118f
C9857 m2_5748_18014# m3_6884_18146# 0.0341f
C9858 rowon_n[15] a_2966_17190# 0.248f
C9859 m2_11196_14426# rowon_n[12] 0.0322f
C9860 col_n[29] a_32386_8194# 0.084f
C9861 m2_17220_10410# rowon_n[8] 0.0322f
C9862 col_n[3] a_5978_7150# 0.251f
C9863 m2_23244_6394# rowon_n[4] 0.0322f
C9864 a_25054_4138# a_26058_4138# 0.843f
C9865 col_n[28] a_2275_10186# 0.113f
C9866 row_n[1] a_12306_3174# 0.0117f
C9867 col_n[10] a_12914_9158# 0.0765f
C9868 vcm a_24354_7190# 0.155f
C9869 rowoff_n[12] a_20434_14540# 0.0133f
C9870 a_2874_8154# a_2966_8154# 0.326f
C9871 m2_34864_13998# a_34090_14178# 0.843f
C9872 vcm a_15014_16186# 0.56f
C9873 a_2275_13198# a_25358_13214# 0.144f
C9874 a_2475_13198# a_27974_13174# 0.264f
C9875 a_14922_13174# a_15014_13174# 0.326f
C9876 VDD a_11910_6146# 0.181f
C9877 row_n[3] a_2161_5166# 0.0221f
C9878 col[13] a_2275_18218# 0.0899f
C9879 rowon_n[7] a_2475_9182# 0.31f
C9880 col[18] a_2275_7174# 0.0899f
C9881 row_n[12] a_34394_14218# 0.0117f
C9882 col_n[4] a_7382_17552# 0.0283f
C9883 vcm a_17934_1126# 0.0983f
C9884 a_16018_6146# a_16018_5142# 0.843f
C9885 col_n[1] a_3878_7150# 0.0765f
C9886 m3_12908_18146# m3_13912_18146# 0.202f
C9887 col[23] a_26058_6146# 0.367f
C9888 m2_8760_946# m3_8892_1078# 3.79f
C9889 vcm a_5278_10202# 0.155f
C9890 rowoff_n[15] a_2475_17214# 3.9f
C9891 a_2275_10186# a_18938_10162# 0.136f
C9892 a_9902_10162# a_10298_10202# 0.0313f
C9893 col[30] a_32994_8154# 0.0682f
C9894 m2_34864_2954# VDD 0.766f
C9895 ctop a_18026_5142# 4.11f
C9896 m2_9764_946# a_9994_2130# 0.843f
C9897 VDD a_26970_10162# 0.181f
C9898 m2_2736_1950# col[0] 0.359f
C9899 col_n[19] rowoff_n[13] 0.0471f
C9900 a_28066_3134# a_28370_3174# 0.0931f
C9901 a_28978_3134# a_29470_3496# 0.0658f
C9902 col_n[3] a_2475_14202# 0.0531f
C9903 col_n[18] a_21342_6186# 0.084f
C9904 vcm a_32994_5142# 0.1f
C9905 rowoff_n[10] a_26970_12170# 0.202f
C9906 rowoff_n[2] a_9902_4138# 0.202f
C9907 col_n[8] a_2475_3158# 0.0531f
C9908 a_5978_7150# a_6982_7150# 0.843f
C9909 a_2475_7174# a_10998_7150# 0.316f
C9910 col[22] rowoff_n[9] 0.0901f
C9911 col[15] rowoff_n[2] 0.0901f
C9912 col[14] rowoff_n[1] 0.0901f
C9913 col[21] rowoff_n[8] 0.0901f
C9914 col[18] rowoff_n[5] 0.0901f
C9915 col[13] rowoff_n[0] 0.0901f
C9916 col[19] rowoff_n[6] 0.0901f
C9917 col[20] rowoff_n[7] 0.0901f
C9918 col[17] rowoff_n[4] 0.0901f
C9919 col[16] rowoff_n[3] 0.0901f
C9920 col_n[2] a_4974_17190# 0.251f
C9921 col_n[28] a_31382_18234# 0.084f
C9922 row_n[6] a_23046_8154# 0.282f
C9923 vcm a_20338_14218# 0.155f
C9924 a_2275_12194# a_33998_12170# 0.136f
C9925 VDD a_18426_4500# 0.0779f
C9926 rowon_n[10] a_22954_12170# 0.118f
C9927 ctop a_33086_9158# 4.11f
C9928 a_29982_17190# a_30074_17190# 0.326f
C9929 VDD a_7894_13174# 0.181f
C9930 m2_14784_18014# col_n[12] 0.243f
C9931 row_n[8] a_10298_10202# 0.0117f
C9932 rowon_n[0] a_32994_2130# 0.118f
C9933 rowoff_n[0] a_18938_2130# 0.202f
C9934 a_1957_4162# a_2161_4162# 0.115f
C9935 a_2475_4162# a_2275_4162# 2.76f
C9936 vcm a_13918_8154# 0.1f
C9937 m2_30848_18014# m2_31276_18442# 0.165f
C9938 a_31078_10162# a_31078_9158# 0.843f
C9939 rowoff_n[13] a_8386_15544# 0.0133f
C9940 a_2475_9182# a_26058_9158# 0.316f
C9941 col[12] a_15014_4138# 0.367f
C9942 vcm a_2275_17214# 6.49f
C9943 a_24962_14178# a_25358_14218# 0.0313f
C9944 m3_16924_1078# a_18026_1126# 0.0341f
C9945 VDD a_33486_8516# 0.0779f
C9946 m2_1732_10986# ctop 0.0428f
C9947 col[22] a_25054_16186# 0.367f
C9948 rowoff_n[5] a_10394_7512# 0.0133f
C9949 col_n[5] a_2275_6170# 0.113f
C9950 col[19] a_21950_6146# 0.0682f
C9951 ctop a_14010_12170# 4.11f
C9952 col_n[3] rowoff_n[14] 0.0471f
C9953 a_2275_18218# a_3878_18194# 0.136f
C9954 a_2874_18194# a_3366_18556# 0.0658f
C9955 row_n[0] a_10906_2130# 0.0437f
C9956 VDD a_22954_17190# 0.181f
C9957 col[29] a_31990_18194# 0.0682f
C9958 rowon_n[4] a_9994_6146# 0.248f
C9959 col[6] rowoff_n[10] 0.0901f
C9960 a_2275_6170# a_17022_6146# 0.399f
C9961 a_8990_6146# a_9294_6186# 0.0931f
C9962 a_9902_6146# a_10394_6508# 0.0658f
C9963 col_n[20] a_2475_16210# 0.0531f
C9964 col_n[25] a_2475_5166# 0.0531f
C9965 vcm a_28978_12170# 0.1f
C9966 rowoff_n[3] a_19430_5504# 0.0133f
C9967 col_n[7] a_10298_4178# 0.084f
C9968 a_21038_11166# a_22042_11166# 0.843f
C9969 VDD a_25054_2130# 0.483f
C9970 m2_4168_17438# row_n[15] 0.0128f
C9971 col_n[17] a_20338_16226# 0.084f
C9972 m2_10192_13422# row_n[11] 0.0128f
C9973 m2_16216_9406# row_n[7] 0.0128f
C9974 m2_22240_5390# row_n[3] 0.0128f
C9975 VDD a_14410_11528# 0.0779f
C9976 ctop a_29070_16186# 4.11f
C9977 col[10] a_2475_13198# 0.136f
C9978 a_2275_3158# a_7286_3174# 0.144f
C9979 a_2475_3158# a_9902_3134# 0.264f
C9980 a_5886_3134# a_5978_3134# 0.326f
C9981 rowoff_n[1] a_28466_3496# 0.0133f
C9982 col[15] a_2475_2154# 0.136f
C9983 rowoff_n[8] a_10998_10162# 0.294f
C9984 col_n[28] a_31478_10524# 0.0283f
C9985 row_n[13] a_21038_15182# 0.282f
C9986 rowoff_n[11] a_14922_13174# 0.202f
C9987 a_2275_8178# a_32082_8154# 0.399f
C9988 vcm a_9902_15182# 0.1f
C9989 m3_2868_1078# m2_2736_946# 3.79f
C9990 a_12002_13174# a_12002_12170# 0.843f
C9991 VDD a_5978_5142# 0.483f
C9992 row_n[3] a_31078_5142# 0.282f
C9993 col_n[26] ctop 0.0594f
C9994 VDD col[23] 3.83f
C9995 col_n[29] row_n[0] 0.298f
C9996 vcm col[20] 5.46f
C9997 col_n[31] row_n[1] 0.298f
C9998 col_n[30] rowon_n[0] 0.111f
C9999 col_n[10] col[10] 0.489f
C10000 col[1] a_3970_2130# 0.367f
C10001 row_n[15] a_8290_17230# 0.0117f
C10002 rowon_n[7] a_30986_9158# 0.118f
C10003 col_n[22] a_2275_8178# 0.113f
C10004 a_5886_17190# a_6282_17230# 0.0313f
C10005 a_2275_17214# a_10906_17190# 0.136f
C10006 rowoff_n[6] a_20034_8154# 0.294f
C10007 VDD a_29470_15544# 0.0779f
C10008 col[11] a_14010_14178# 0.367f
C10009 col[8] a_10906_4138# 0.0682f
C10010 col[18] a_20946_16186# 0.0682f
C10011 row_n[5] a_18330_7190# 0.0117f
C10012 a_2475_5166# a_24962_5142# 0.264f
C10013 a_2275_5166# a_22346_5182# 0.144f
C10014 m3_2868_1078# m3_3872_1078# 0.125f
C10015 a_26970_1126# a_27062_1126# 0.0991f
C10016 col_n[26] a_29070_10162# 0.251f
C10017 a_24962_10162# a_25454_10524# 0.0658f
C10018 a_24050_10162# a_24354_10202# 0.0931f
C10019 col[7] a_2275_16210# 0.0899f
C10020 rowoff_n[15] a_30986_17190# 0.202f
C10021 m2_29268_16434# a_29070_16186# 0.165f
C10022 rowoff_n[4] a_29070_6146# 0.294f
C10023 col[12] a_2275_5166# 0.0899f
C10024 m2_14784_946# a_2475_1150# 0.286f
C10025 a_2475_14202# a_2874_14178# 0.264f
C10026 m3_7888_1078# a_7986_2130# 0.0302f
C10027 a_1957_14202# a_2275_14202# 0.158f
C10028 row_n[7] a_8898_9158# 0.0437f
C10029 VDD a_21038_9158# 0.483f
C10030 col_n[6] a_9294_14218# 0.084f
C10031 rowon_n[11] a_7986_13174# 0.248f
C10032 VDD a_10394_18556# 0.0858f
C10033 a_2275_2154# a_15926_2130# 0.136f
C10034 col[27] a_2475_15206# 0.136f
C10035 m2_7756_946# VDD 1f
C10036 vcm a_27062_4138# 0.56f
C10037 rowon_n[1] a_18026_3134# 0.248f
C10038 a_20946_7150# a_21038_7150# 0.326f
C10039 col_n[17] a_20434_8516# 0.0283f
C10040 m2_6752_18014# a_6890_18194# 0.225f
C10041 a_2475_16210# a_18026_16186# 0.316f
C10042 a_27062_17190# a_27062_16186# 0.843f
C10043 VDD a_2475_12194# 26.1f
C10044 col_n[2] a_2475_1150# 0.0531f
C10045 sample_n m2_1732_946# 0.0523f
C10046 a_2275_4162# a_30986_4138# 0.136f
C10047 a_15926_4138# a_16322_4178# 0.0313f
C10048 col[0] a_2874_12170# 0.0682f
C10049 vcm a_7986_7150# 0.56f
C10050 col[7] a_9902_14178# 0.0682f
C10051 rowoff_n[12] a_2161_14202# 0.0226f
C10052 row_n[10] a_29070_12170# 0.282f
C10053 m2_20232_14426# a_20034_14178# 0.165f
C10054 col[24] a_2275_18218# 0.0899f
C10055 rowon_n[14] a_28978_16186# 0.118f
C10056 col_n[15] a_18026_8154# 0.251f
C10057 a_5886_13174# a_6378_13536# 0.0658f
C10058 a_2275_13198# a_8990_13174# 0.399f
C10059 a_4974_13174# a_5278_13214# 0.0931f
C10060 col[29] a_2275_7174# 0.0899f
C10061 col_n[22] a_24962_10162# 0.0765f
C10062 VDD a_17022_16186# 0.483f
C10063 a_2475_1150# a_23046_1126# 0.0299f
C10064 row_n[12] a_16322_14218# 0.0117f
C10065 m2_17220_2378# a_17022_2130# 0.165f
C10066 vcm a_32386_2170# 0.155f
C10067 m2_1732_8978# sample_n 0.0522f
C10068 col_n[0] a_2275_4162# 0.113f
C10069 row_n[2] a_26362_4178# 0.0117f
C10070 vcm a_23046_11166# 0.56f
C10071 row_n[14] a_6890_16186# 0.0437f
C10072 VDD a_19942_1126# 0.404f
C10073 col_n[6] a_9390_6508# 0.0283f
C10074 a_2275_15206# a_24050_15182# 0.399f
C10075 col_n[16] a_19430_18556# 0.0283f
C10076 col_n[30] rowoff_n[13] 0.0471f
C10077 col_n[14] a_2475_14202# 0.0531f
C10078 row_n[4] a_16930_6146# 0.0437f
C10079 col_n[19] a_2475_3158# 0.0531f
C10080 col[27] rowoff_n[3] 0.0901f
C10081 rowon_n[8] a_16018_10162# 0.248f
C10082 sample_n rowoff_n[8] 0.14f
C10083 col[24] rowoff_n[0] 0.0901f
C10084 col[29] rowoff_n[5] 0.0901f
C10085 col[25] rowoff_n[1] 0.0901f
C10086 col[26] rowoff_n[2] 0.0901f
C10087 col[31] rowoff_n[7] 0.0901f
C10088 col[30] rowoff_n[6] 0.0901f
C10089 col[28] rowoff_n[4] 0.0901f
C10090 vcm a_13310_5182# 0.155f
C10091 a_30986_8154# a_31382_8194# 0.0313f
C10092 col[10] a_2475_18218# 0.136f
C10093 m2_11196_12418# a_10998_12170# 0.165f
C10094 m2_6176_8402# rowon_n[6] 0.0322f
C10095 vcm a_3970_14178# 0.56f
C10096 m2_12200_4386# rowon_n[2] 0.0322f
C10097 a_2475_12194# a_16930_12170# 0.264f
C10098 a_2275_12194# a_14314_12210# 0.144f
C10099 VDD a_35002_5142# 0.258f
C10100 col[4] a_2475_11190# 0.136f
C10101 m2_27260_18442# VDD 0.0456f
C10102 a_20034_17190# a_20338_17230# 0.0931f
C10103 a_20946_17190# a_21438_17552# 0.0658f
C10104 col_n[4] a_6982_6146# 0.251f
C10105 col_n[30] a_33390_7190# 0.084f
C10106 col_n[11] a_13918_8154# 0.0765f
C10107 a_27062_5142# a_28066_5142# 0.843f
C10108 m2_30272_8402# a_30074_8154# 0.165f
C10109 col_n[11] a_2275_17214# 0.113f
C10110 vcm a_28370_9198# 0.155f
C10111 m2_12776_18014# m2_13780_18014# 0.843f
C10112 a_2275_9182# a_7894_9158# 0.136f
C10113 col_n[16] a_2275_6170# 0.113f
C10114 vcm a_19030_18194# 0.165f
C10115 col_n[14] rowoff_n[14] 0.0471f
C10116 ctop a_6982_3134# 4.11f
C10117 m2_21236_17438# rowon_n[15] 0.0322f
C10118 a_16930_14178# a_17022_14178# 0.326f
C10119 a_2275_14202# a_29374_14218# 0.144f
C10120 a_2475_14202# a_31990_14178# 0.264f
C10121 m2_27260_13422# rowon_n[11] 0.0322f
C10122 VDD a_15926_8154# 0.181f
C10123 m2_33284_9406# rowon_n[7] 0.0322f
C10124 m2_26832_946# vcm 0.353f
C10125 col[17] rowoff_n[10] 0.0901f
C10126 col_n[5] a_8386_16548# 0.0283f
C10127 col_n[31] a_2475_16210# 0.0531f
C10128 col[1] a_2275_14202# 0.0899f
C10129 col[24] a_27062_5142# 0.367f
C10130 col[6] a_2275_3158# 0.0899f
C10131 vcm a_21950_3134# 0.1f
C10132 row_n[9] a_24354_11206# 0.0117f
C10133 a_18026_7150# a_18026_6146# 0.843f
C10134 m2_1732_9982# a_1957_10186# 0.245f
C10135 col[31] a_33998_7150# 0.0682f
C10136 vcm a_9294_12210# 0.155f
C10137 a_11910_11166# a_12306_11206# 0.0313f
C10138 a_2275_11190# a_22954_11166# 0.136f
C10139 VDD a_7382_2492# 0.0779f
C10140 m2_25828_18014# a_25966_18194# 0.225f
C10141 ctop a_22042_7150# 4.11f
C10142 row_n[11] a_14922_13174# 0.0437f
C10143 col[21] a_2475_13198# 0.136f
C10144 VDD a_30986_12170# 0.181f
C10145 m2_20808_18014# m3_19936_18146# 0.0341f
C10146 col[26] a_2475_2154# 0.136f
C10147 rowon_n[15] a_14010_17190# 0.248f
C10148 col_n[19] a_22346_5182# 0.084f
C10149 a_30074_4138# a_30378_4178# 0.0931f
C10150 a_30986_4138# a_31478_4500# 0.0658f
C10151 rowoff_n[1] a_10906_3134# 0.202f
C10152 row_n[1] a_24962_3134# 0.0437f
C10153 col_n[3] a_5978_16186# 0.251f
C10154 m2_21236_6394# a_21038_6146# 0.165f
C10155 col_n[29] a_32386_17230# 0.084f
C10156 row_n[13] a_2966_15182# 0.281f
C10157 vcm a_2161_6170# 0.0169f
C10158 rowon_n[5] a_24050_7150# 0.248f
C10159 rowoff_n[12] a_31078_14178# 0.294f
C10160 a_2475_8178# a_15014_8154# 0.316f
C10161 a_7986_8154# a_8990_8154# 0.843f
C10162 col_n[15] col[16] 7.13f
C10163 row_n[13] ctop 0.186f
C10164 vcm col[31] 5.19f
C10165 sample rowoff_n[15] 0.0786f
C10166 col_n[10] a_12914_18194# 0.0762f
C10167 vcm a_24354_16226# 0.155f
C10168 VDD a_22442_6508# 0.0779f
C10169 col[1] rowoff_n[11] 0.0901f
C10170 a_31990_18194# a_32082_18194# 0.0991f
C10171 rowoff_n[6] a_1957_8178# 0.0219f
C10172 VDD a_11910_15182# 0.181f
C10173 col[18] a_2275_16210# 0.0899f
C10174 row_n[5] a_2475_7174# 0.405f
C10175 a_2275_5166# a_5978_5142# 0.399f
C10176 m2_34864_3958# vcm 0.408f
C10177 col[23] a_2275_5166# 0.0899f
C10178 m2_23820_946# m3_24956_1078# 0.0341f
C10179 col[13] a_16018_3134# 0.367f
C10180 vcm a_17934_10162# 0.1f
C10181 col_n[1] a_3878_16186# 0.0765f
C10182 a_33086_11166# a_33086_10162# 0.843f
C10183 a_2475_10186# a_30074_10162# 0.316f
C10184 row_n[14] a_35094_16186# 0.0123f
C10185 col[23] a_26058_15182# 0.367f
C10186 rowoff_n[4] a_11398_6508# 0.0133f
C10187 col[20] a_22954_5142# 0.0682f
C10188 a_26970_15182# a_27366_15222# 0.0313f
C10189 VDD a_2966_9158# 0.485f
C10190 m2_15788_18014# ctop 0.0422f
C10191 col[30] a_32994_17190# 0.0682f
C10192 ctop a_18026_14178# 4.11f
C10193 m2_12200_4386# a_12002_4138# 0.165f
C10194 m2_5172_7398# row_n[5] 0.0128f
C10195 m2_11196_3382# row_n[1] 0.0128f
C10196 rowoff_n[2] a_20434_4500# 0.0133f
C10197 col_n[8] a_11302_3174# 0.084f
C10198 a_10998_7150# a_11302_7190# 0.0931f
C10199 a_2275_7174# a_21038_7150# 0.399f
C10200 a_11910_7150# a_12402_7512# 0.0658f
C10201 rowoff_n[9] a_2874_11166# 0.202f
C10202 row_n[6] a_32386_8194# 0.0117f
C10203 col_n[18] a_21342_15222# 0.084f
C10204 vcm a_32994_14178# 0.1f
C10205 col_n[8] a_2475_12194# 0.0531f
C10206 a_23046_12170# a_24050_12170# 0.843f
C10207 VDD a_29070_4138# 0.483f
C10208 col_n[13] a_2475_1150# 0.0531f
C10209 a_35002_17190# a_35398_17230# 0.0313f
C10210 VDD a_18426_13536# 0.0779f
C10211 row_n[8] a_22954_10162# 0.0437f
C10212 m3_1864_15134# a_2966_15182# 0.0302f
C10213 rowoff_n[7] a_12002_9158# 0.294f
C10214 rowoff_n[0] a_29470_2492# 0.0133f
C10215 col_n[29] a_32482_9520# 0.0283f
C10216 rowon_n[12] a_22042_14178# 0.248f
C10217 a_7894_4138# a_7986_4138# 0.326f
C10218 a_2475_4162# a_13918_4138# 0.264f
C10219 a_2275_4162# a_11302_4178# 0.144f
C10220 m3_1864_15134# ctop 0.21f
C10221 m2_20232_16434# row_n[14] 0.0128f
C10222 m2_26256_12418# row_n[10] 0.0128f
C10223 m2_32280_8402# row_n[6] 0.0128f
C10224 rowoff_n[13] a_19030_15182# 0.294f
C10225 m2_31852_946# col_n[29] 0.357f
C10226 rowon_n[2] a_32082_4138# 0.248f
C10227 vcm a_13918_17190# 0.1f
C10228 a_14010_14178# a_14010_13174# 0.843f
C10229 VDD a_9994_7150# 0.483f
C10230 rowoff_n[5] a_21038_7150# 0.294f
C10231 col[12] a_15014_13174# 0.367f
C10232 a_7894_18194# a_8290_18234# 0.0313f
C10233 a_2275_18218# a_14922_18194# 0.136f
C10234 col[9] a_11910_3134# 0.0682f
C10235 m2_29844_18014# col[27] 0.347f
C10236 VDD a_33486_17552# 0.0779f
C10237 col_n[5] a_2275_15206# 0.113f
C10238 a_2275_1150# a_4882_1126# 0.136f
C10239 col[19] a_21950_15182# 0.0682f
C10240 m2_2736_1950# a_2874_2130# 0.225f
C10241 col_n[10] a_2275_4162# 0.113f
C10242 vcm a_16018_2130# 0.56f
C10243 a_2475_6170# a_28978_6146# 0.264f
C10244 col_n[27] a_30074_9158# 0.251f
C10245 a_2275_6170# a_26362_6186# 0.144f
C10246 rowoff_n[3] a_30074_5142# 0.294f
C10247 row_n[2] a_9994_4138# 0.282f
C10248 a_26970_11166# a_27462_11528# 0.0658f
C10249 a_26058_11166# a_26362_11206# 0.0931f
C10250 VDD a_35398_2170# 0.0882f
C10251 rowon_n[6] a_9902_8154# 0.118f
C10252 m2_21812_18014# a_22042_17190# 0.843f
C10253 col_n[25] a_2475_14202# 0.0531f
C10254 m2_1732_5966# VDD 0.856f
C10255 col_n[7] a_10298_13214# 0.084f
C10256 a_2475_15206# a_6982_15182# 0.316f
C10257 a_3970_15182# a_4974_15182# 0.843f
C10258 col_n[30] a_2475_3158# 0.0531f
C10259 VDD a_25054_11166# 0.483f
C10260 col[0] a_2275_1150# 0.099f
C10261 col[21] a_2475_18218# 0.136f
C10262 a_2475_18218# a_12914_18194# 0.264f
C10263 a_2275_3158# a_19942_3134# 0.136f
C10264 a_33086_1126# a_2275_1150# 0.0924f
C10265 col_n[18] a_21438_7512# 0.0283f
C10266 row_n[13] a_30378_15222# 0.0117f
C10267 vcm a_31078_6146# 0.56f
C10268 a_22954_8154# a_23046_8154# 0.326f
C10269 rowoff_n[11] a_25454_13536# 0.0133f
C10270 col[15] a_2475_11190# 0.136f
C10271 a_30474_1488# VDD 0.0977f
C10272 row_n[15] a_20946_17190# 0.0437f
C10273 a_2475_17214# a_22042_17190# 0.316f
C10274 VDD a_5978_14178# 0.483f
C10275 col[1] a_3970_11166# 0.367f
C10276 m3_27968_18146# a_28066_17190# 0.0303f
C10277 col_n[22] a_2275_17214# 0.113f
C10278 col_n[27] a_2275_6170# 0.113f
C10279 a_2275_5166# a_35002_5142# 0.136f
C10280 row_n[5] a_30986_7150# 0.0437f
C10281 a_17934_5142# a_18330_5182# 0.0313f
C10282 col[8] a_10906_13174# 0.0682f
C10283 col_n[25] rowoff_n[14] 0.0471f
C10284 rowon_n[9] a_30074_11166# 0.248f
C10285 vcm a_12002_9158# 0.56f
C10286 rowoff_n[14] a_6982_16186# 0.294f
C10287 col_n[16] a_19030_7150# 0.251f
C10288 m2_3164_15430# a_2966_15182# 0.165f
C10289 col[28] rowoff_n[10] 0.0901f
C10290 a_2275_14202# a_13006_14178# 0.399f
C10291 a_7894_14178# a_8386_14540# 0.0658f
C10292 a_6982_14178# a_7286_14218# 0.0931f
C10293 col_n[23] a_25966_9158# 0.0765f
C10294 col[12] a_2275_14202# 0.0899f
C10295 col[17] a_2275_3158# 0.0899f
C10296 VDD a_21038_18194# 0.0356f
C10297 a_2475_2154# a_27062_2130# 0.316f
C10298 a_14010_2130# a_15014_2130# 0.843f
C10299 m2_30848_946# VDD 1f
C10300 vcm a_3878_3134# 0.1f
C10301 row_n[9] a_7986_11166# 0.282f
C10302 rowoff_n[9] a_31990_11166# 0.202f
C10303 rowon_n[13] a_7894_15182# 0.118f
C10304 vcm a_27062_13174# 0.56f
C10305 col_n[7] a_10394_5504# 0.0283f
C10306 a_2475_11190# a_5886_11166# 0.264f
C10307 a_2275_11190# a_3270_11206# 0.144f
C10308 VDD a_23958_3134# 0.181f
C10309 col_n[17] a_20434_17552# 0.0283f
C10310 a_2275_16210# a_28066_16186# 0.399f
C10311 rowon_n[3] a_17934_5142# 0.118f
C10312 a_33086_1126# m2_32856_946# 0.0249f
C10313 m2_1732_1950# rowon_n[0] 0.236f
C10314 a_4974_4138# a_4974_3134# 0.843f
C10315 row_n[13] col[5] 0.0342f
C10316 rowon_n[10] col[0] 0.0318f
C10317 col_n[21] col[21] 0.489f
C10318 row_n[14] col[7] 0.0342f
C10319 rowon_n[14] col[8] 0.0323f
C10320 row_n[11] col[1] 0.0342f
C10321 rowon_n[11] col[2] 0.0323f
C10322 col_n[9] rowoff_n[15] 0.0471f
C10323 rowon_n[12] col[4] 0.0323f
C10324 row_n[1] a_5278_3174# 0.0117f
C10325 row_n[15] col[9] 0.0342f
C10326 rowon_n[7] ctop 0.203f
C10327 col_n[2] a_2475_10186# 0.0531f
C10328 row_n[12] col[3] 0.0342f
C10329 rowon_n[13] col[6] 0.0323f
C10330 rowon_n[15] col[10] 0.0323f
C10331 rowon_n[3] rowon_n[2] 0.0632f
C10332 vcm a_17326_7190# 0.155f
C10333 rowoff_n[12] a_13406_14540# 0.0133f
C10334 a_32994_9158# a_33390_9198# 0.0313f
C10335 col[12] rowoff_n[11] 0.0901f
C10336 ctop a_30074_2130# 4.06f
C10337 vcm a_7986_16186# 0.56f
C10338 a_2475_13198# a_20946_13174# 0.264f
C10339 a_2275_13198# a_18330_13214# 0.144f
C10340 VDD a_4882_6146# 0.181f
C10341 col_n[5] a_7986_5142# 0.251f
C10342 col_n[15] a_18026_17190# 0.251f
C10343 m2_31852_18014# a_2475_18218# 0.286f
C10344 a_22954_18194# a_23446_18556# 0.0658f
C10345 col[29] a_2275_16210# 0.0899f
C10346 col_n[12] a_14922_7150# 0.0765f
C10347 row_n[12] a_28978_14178# 0.0437f
C10348 a_17934_1126# a_18426_1488# 0.0664f
C10349 vcm a_10906_1126# 0.0989f
C10350 m2_10192_15430# rowon_n[13] 0.0322f
C10351 a_29070_6146# a_30074_6146# 0.843f
C10352 m2_16216_11414# rowon_n[9] 0.0322f
C10353 m2_22240_7398# rowon_n[5] 0.0322f
C10354 m2_28264_3382# rowon_n[1] 0.0322f
C10355 m2_34864_946# m2_35292_1374# 0.165f
C10356 vcm a_32386_11206# 0.155f
C10357 a_2275_10186# a_11910_10162# 0.136f
C10358 m2_34864_17010# a_35094_17190# 0.0249f
C10359 col_n[0] a_2275_13198# 0.113f
C10360 ctop a_10998_5142# 4.11f
C10361 a_2275_15206# a_33390_15222# 0.144f
C10362 a_18938_15182# a_19030_15182# 0.326f
C10363 col_n[4] a_2275_2154# 0.113f
C10364 VDD a_19942_10162# 0.181f
C10365 col_n[6] a_9390_15544# 0.0283f
C10366 col[25] a_28066_4138# 0.367f
C10367 vcm a_25966_5142# 0.1f
C10368 col_n[19] a_2475_12194# 0.0531f
C10369 rowoff_n[2] a_2161_4162# 0.0226f
C10370 rowoff_n[10] a_19942_12170# 0.202f
C10371 a_2475_7174# a_3970_7150# 0.316f
C10372 a_2275_7174# a_2966_7150# 0.399f
C10373 a_20034_8154# a_20034_7150# 0.843f
C10374 col_n[24] a_2475_1150# 0.0531f
C10375 row_n[6] a_16018_8154# 0.282f
C10376 vcm a_13310_14218# 0.155f
C10377 a_2275_12194# a_26970_12170# 0.136f
C10378 a_13918_12170# a_14314_12210# 0.0313f
C10379 rowon_n[10] a_15926_12170# 0.118f
C10380 VDD a_11398_4500# 0.0779f
C10381 ctop a_26058_9158# 4.11f
C10382 VDD a_35002_14178# 0.258f
C10383 col_n[20] a_23350_4178# 0.084f
C10384 row_n[8] a_3270_10202# 0.0117f
C10385 rowoff_n[0] a_11910_2130# 0.202f
C10386 col[9] a_2475_9182# 0.136f
C10387 rowon_n[0] a_25966_2130# 0.118f
C10388 col_n[30] a_33390_16226# 0.084f
C10389 col_n[4] a_6982_15182# 0.251f
C10390 a_32994_5142# a_33486_5504# 0.0658f
C10391 a_32082_5142# a_32386_5182# 0.0931f
C10392 col_n[11] a_13918_17190# 0.0765f
C10393 vcm a_6890_8154# 0.1f
C10394 m2_23820_18014# m2_24248_18442# 0.165f
C10395 a_9994_9158# a_10998_9158# 0.843f
C10396 a_2475_9182# a_19030_9158# 0.316f
C10397 m2_26256_15430# a_26058_15182# 0.165f
C10398 vcm a_28370_18234# 0.16f
C10399 VDD a_26458_8516# 0.0779f
C10400 col_n[16] a_2275_15206# 0.113f
C10401 rowoff_n[5] a_2966_7150# 0.294f
C10402 col_n[21] a_2275_4162# 0.113f
C10403 ctop a_6982_12170# 4.11f
C10404 VDD a_15926_17190# 0.181f
C10405 a_28978_2130# a_29070_2130# 0.326f
C10406 rowon_n[4] a_2874_6146# 0.118f
C10407 col[14] a_17022_2130# 0.367f
C10408 a_2275_6170# a_9994_6146# 0.399f
C10409 col[24] a_27062_14178# 0.367f
C10410 col[6] a_2275_12194# 0.0899f
C10411 rowoff_n[3] a_12402_5504# 0.0133f
C10412 vcm a_21950_12170# 0.1f
C10413 col[21] a_23958_4138# 0.0682f
C10414 a_2475_11190# a_34090_11166# 0.316f
C10415 VDD a_18026_2130# 0.483f
C10416 col[11] a_2275_1150# 0.0899f
C10417 col[31] a_33998_16186# 0.0682f
C10418 a_28978_16186# a_29374_16226# 0.0313f
C10419 VDD a_7382_11528# 0.0779f
C10420 m2_34864_18014# m3_34996_18146# 3.79f
C10421 ctop a_22042_16186# 4.11f
C10422 col[26] a_2475_11190# 0.136f
C10423 rowoff_n[8] a_3970_10162# 0.294f
C10424 rowoff_n[1] a_21438_3496# 0.0133f
C10425 col_n[9] a_12306_2170# 0.084f
C10426 row_n[13] a_14010_15182# 0.282f
C10427 col_n[19] a_22346_14218# 0.084f
C10428 m2_1732_13998# m2_1732_12994# 0.843f
C10429 rowoff_n[11] a_7894_13174# 0.202f
C10430 a_2275_8178# a_25054_8154# 0.399f
C10431 a_13006_8154# a_13310_8194# 0.0931f
C10432 a_13918_8154# a_14410_8516# 0.0658f
C10433 m2_17220_13422# a_17022_13174# 0.165f
C10434 vcm a_2161_15206# 0.0169f
C10435 a_25054_13174# a_26058_13174# 0.843f
C10436 VDD a_33086_6146# 0.483f
C10437 row_n[3] a_24050_5142# 0.282f
C10438 row_n[15] a_2275_17214# 19.2f
C10439 rowon_n[7] a_23958_9158# 0.118f
C10440 m2_9188_14426# row_n[12] 0.0128f
C10441 a_2874_17190# a_2966_17190# 0.326f
C10442 m2_15212_10410# row_n[8] 0.0128f
C10443 rowoff_n[6] a_13006_8154# 0.294f
C10444 col_n[30] a_33486_8516# 0.0283f
C10445 VDD a_22442_15544# 0.0779f
C10446 m2_21236_6394# row_n[4] 0.0128f
C10447 a_2475_5166# a_17934_5142# 0.264f
C10448 a_2275_5166# a_15318_5182# 0.144f
C10449 a_9902_5142# a_9994_5142# 0.326f
C10450 row_n[5] a_11302_7190# 0.0117f
C10451 rowoff_n[15] a_23958_17190# 0.202f
C10452 col[23] a_2275_14202# 0.0899f
C10453 rowoff_n[4] a_22042_6146# 0.294f
C10454 col[13] a_16018_12170# 0.367f
C10455 col[28] a_2275_3158# 0.0899f
C10456 a_16018_15182# a_16018_14178# 0.843f
C10457 col[10] a_12914_2130# 0.0682f
C10458 VDD a_14010_9158# 0.483f
C10459 col[20] a_22954_14178# 0.0682f
C10460 VDD a_2966_18194# 0.0356f
C10461 a_2275_2154# a_8898_2130# 0.136f
C10462 m2_35292_15430# row_n[13] 0.0128f
C10463 a_4882_2130# a_5278_2170# 0.0313f
C10464 col_n[28] a_31078_8154# 0.251f
C10465 vcm a_20034_4138# 0.56f
C10466 rowon_n[1] a_10998_3134# 0.248f
C10467 rowoff_n[2] a_31078_4138# 0.294f
C10468 a_2475_7174# a_32994_7150# 0.264f
C10469 a_2275_7174# a_30378_7190# 0.144f
C10470 m2_8184_11414# a_7986_11166# 0.165f
C10471 col_n[8] a_11302_12210# 0.084f
C10472 a_28066_12170# a_28370_12210# 0.0931f
C10473 a_28978_12170# a_29470_12532# 0.0658f
C10474 a_5978_16186# a_6982_16186# 0.843f
C10475 a_2475_16210# a_10998_16186# 0.316f
C10476 VDD a_29070_13174# 0.483f
C10477 row_n[15] col[20] 0.0342f
C10478 rowon_n[0] row_n[0] 18.9f
C10479 rowon_n[11] col[13] 0.0323f
C10480 row_n[7] col[4] 0.0342f
C10481 row_n[11] col[12] 0.0342f
C10482 col_n[26] col[27] 7.07f
C10483 row_n[13] col[16] 0.0342f
C10484 rowon_n[14] col[19] 0.0323f
C10485 row_n[6] col[2] 0.0342f
C10486 rowon_n[6] col[3] 0.0323f
C10487 rowon_n[15] col[21] 0.0323f
C10488 row_n[5] col[0] 0.0322f
C10489 col_n[20] rowoff_n[15] 0.0471f
C10490 rowon_n[10] col[11] 0.0323f
C10491 rowon_n[7] col[5] 0.0323f
C10492 rowon_n[13] col[17] 0.0323f
C10493 rowon_n[8] col[7] 0.0323f
C10494 rowon_n[12] col[15] 0.0323f
C10495 rowon_n[5] col[1] 0.0323f
C10496 col_n[13] a_2475_10186# 0.0531f
C10497 row_n[10] col[10] 0.0342f
C10498 row_n[8] col[6] 0.0342f
C10499 row_n[12] col[14] 0.0342f
C10500 row_n[14] col[18] 0.0342f
C10501 row_n[2] ctop 0.186f
C10502 row_n[9] col[8] 0.0342f
C10503 rowon_n[9] col[9] 0.0323f
C10504 m2_1732_12994# col[0] 0.0137f
C10505 col_n[19] a_22442_6508# 0.0283f
C10506 a_2275_4162# a_23958_4138# 0.136f
C10507 m3_15920_1078# ctop 0.21f
C10508 col[23] rowoff_n[11] 0.0901f
C10509 m2_27260_7398# a_27062_7150# 0.165f
C10510 col_n[29] a_32482_18556# 0.0283f
C10511 vcm a_35094_8154# 0.165f
C10512 a_24962_9158# a_25054_9158# 0.326f
C10513 row_n[10] a_22042_12170# 0.282f
C10514 rowon_n[14] a_21950_16186# 0.118f
C10515 a_1957_13198# a_2161_13198# 0.115f
C10516 a_2475_13198# a_2275_13198# 2.76f
C10517 col[3] a_2475_7174# 0.136f
C10518 col[2] a_4974_10162# 0.367f
C10519 row_n[0] a_32082_2130# 0.282f
C10520 VDD a_9994_16186# 0.483f
C10521 a_2475_1150# a_16018_1126# 0.0299f
C10522 row_n[12] a_9294_14218# 0.0117f
C10523 rowon_n[4] a_31990_6146# 0.118f
C10524 col[9] a_11910_12170# 0.0682f
C10525 vcm a_25358_2170# 0.155f
C10526 a_19942_6146# a_20338_6186# 0.0313f
C10527 m2_1732_6970# vcm 0.316f
C10528 m2_14784_946# m2_15788_946# 0.843f
C10529 col_n[17] a_20034_6146# 0.251f
C10530 col_n[10] a_2275_13198# 0.113f
C10531 vcm a_16018_11166# 0.56f
C10532 row_n[2] a_19334_4178# 0.0117f
C10533 col_n[15] a_2275_2154# 0.113f
C10534 VDD a_12914_1126# 0.405f
C10535 col_n[24] a_26970_8154# 0.0765f
C10536 a_8990_15182# a_9294_15222# 0.0931f
C10537 a_2275_15206# a_17022_15182# 0.399f
C10538 a_9902_15182# a_10394_15544# 0.0658f
C10539 VDD a_35398_11206# 0.0882f
C10540 m2_34864_15002# m3_34996_15134# 3.79f
C10541 rowon_n[0] m2_33284_2378# 0.0322f
C10542 row_n[4] a_9902_6146# 0.0437f
C10543 col_n[30] a_2475_12194# 0.0531f
C10544 col[0] a_2275_10186# 0.099f
C10545 a_16018_3134# a_17022_3134# 0.843f
C10546 a_2475_3158# a_31078_3134# 0.316f
C10547 rowon_n[8] a_8990_10162# 0.248f
C10548 col[7] rowoff_n[12] 0.0901f
C10549 rowoff_n[8] a_32994_10162# 0.202f
C10550 m2_18224_5390# a_18026_5142# 0.165f
C10551 vcm a_6282_5182# 0.155f
C10552 col_n[8] a_11398_4500# 0.0283f
C10553 col_n[18] a_21438_16548# 0.0283f
C10554 vcm a_31078_15182# 0.56f
C10555 a_5886_12170# a_5978_12170# 0.326f
C10556 a_2275_12194# a_7286_12210# 0.144f
C10557 a_2475_12194# a_9902_12170# 0.264f
C10558 VDD a_27974_5142# 0.181f
C10559 m2_13204_18442# VDD 0.0456f
C10560 col[20] a_2475_9182# 0.136f
C10561 a_2275_17214# a_32082_17190# 0.399f
C10562 a_6982_5142# a_6982_4138# 0.843f
C10563 m2_5748_18014# m2_6752_18014# 0.843f
C10564 vcm a_21342_9198# 0.155f
C10565 col_n[27] a_2275_15206# 0.113f
C10566 col_n[6] a_8990_4138# 0.251f
C10567 ctop a_34090_4138# 4.06f
C10568 vcm a_12002_18194# 0.165f
C10569 a_2275_14202# a_22346_14218# 0.144f
C10570 a_2475_14202# a_24962_14178# 0.264f
C10571 col_n[16] a_19030_16186# 0.251f
C10572 row_n[7] a_30074_9158# 0.282f
C10573 VDD a_8898_8154# 0.181f
C10574 m2_5172_9406# rowon_n[7] 0.0322f
C10575 m2_11196_5390# rowon_n[3] 0.0322f
C10576 col_n[13] a_15926_6146# 0.0765f
C10577 rowon_n[11] a_29982_13174# 0.118f
C10578 VDD a_30378_18234# 0.019f
C10579 col_n[23] a_25966_18194# 0.0762f
C10580 a_19030_2130# a_19334_2170# 0.0931f
C10581 a_19942_2130# a_20434_2492# 0.0658f
C10582 m2_9188_3382# a_8990_3134# 0.165f
C10583 col[17] a_2275_12194# 0.0899f
C10584 m3_34996_18146# VDD 0.0942f
C10585 row_n[9] a_17326_11206# 0.0117f
C10586 vcm a_14922_3134# 0.1f
C10587 a_31078_7150# a_32082_7150# 0.843f
C10588 col[22] a_2275_1150# 0.0899f
C10589 vcm a_3878_12170# 0.1f
C10590 a_2275_11190# a_15926_11166# 0.136f
C10591 VDD a_34490_3496# 0.0779f
C10592 m2_20808_18014# a_21038_18194# 0.0249f
C10593 ctop a_15014_7150# 4.11f
C10594 col_n[7] a_10394_14540# 0.0283f
C10595 row_n[11] a_7894_13174# 0.0437f
C10596 a_20946_16186# a_21038_16186# 0.326f
C10597 VDD a_23958_12170# 0.181f
C10598 m2_10768_18014# m3_11904_18146# 0.0341f
C10599 col[26] a_29070_3134# 0.367f
C10600 rowon_n[15] a_6982_17190# 0.248f
C10601 m2_26256_14426# rowon_n[12] 0.0322f
C10602 m2_32280_10410# rowon_n[8] 0.0322f
C10603 row_n[1] a_17934_3134# 0.0437f
C10604 rowoff_n[1] a_3366_3496# 0.0133f
C10605 rowon_n[5] a_17022_7150# 0.248f
C10606 vcm a_29982_7150# 0.1f
C10607 rowoff_n[12] a_24050_14178# 0.294f
C10608 a_2475_8178# a_7986_8154# 0.316f
C10609 a_22042_9158# a_22042_8154# 0.843f
C10610 m2_1732_12994# a_2966_13174# 0.843f
C10611 col_n[7] a_2475_8178# 0.0531f
C10612 vcm a_17326_16226# 0.155f
C10613 a_15926_13174# a_16322_13214# 0.0313f
C10614 a_2275_13198# a_30986_13174# 0.136f
C10615 VDD a_15414_6508# 0.0779f
C10616 col_n[21] a_24354_3174# 0.084f
C10617 ctop a_30074_11166# 4.11f
C10618 VDD a_4882_15182# 0.181f
C10619 col_n[5] a_7986_14178# 0.251f
C10620 col_n[2] a_4882_4138# 0.0765f
C10621 col_n[12] a_14922_16186# 0.0765f
C10622 a_35002_6146# a_35494_6508# 0.0658f
C10623 m2_13780_946# m3_13912_1078# 3.79f
C10624 vcm a_10906_10162# 0.1f
C10625 a_2475_10186# a_23046_10162# 0.316f
C10626 a_12002_10162# a_13006_10162# 0.843f
C10627 row_n[14] a_28066_16186# 0.282f
C10628 m2_34864_16006# a_2275_16210# 0.278f
C10629 rowoff_n[4] a_4370_6508# 0.0133f
C10630 VDD a_30474_10524# 0.0779f
C10631 m2_34864_11990# m3_34996_12122# 3.79f
C10632 ctop a_10998_14178# 4.11f
C10633 col_n[4] a_2275_11190# 0.113f
C10634 a_30986_3134# a_31078_3134# 0.326f
C10635 col[15] a_18026_1126# 0.428f
C10636 col[25] a_28066_13174# 0.367f
C10637 vcm a_1957_4162# 0.139f
C10638 rowoff_n[2] a_13406_4500# 0.0133f
C10639 rowoff_n[10] a_30474_12532# 0.0133f
C10640 a_2275_7174# a_14010_7150# 0.399f
C10641 m2_30848_18014# vcm 0.353f
C10642 col[22] a_24962_3134# 0.0682f
C10643 row_n[6] a_25358_8194# 0.0117f
C10644 vcm a_25966_14178# 0.1f
C10645 VDD a_22042_4138# 0.483f
C10646 row_n[8] col[17] 0.0342f
C10647 rowon_n[1] col[4] 0.0323f
C10648 row_n[12] col[25] 0.0342f
C10649 row_n[7] col[15] 0.0342f
C10650 rowon_n[8] col[18] 0.0323f
C10651 rowon_n[12] col[26] 0.0323f
C10652 rowon_n[11] col[24] 0.0323f
C10653 sw_n analog_in 0.0649f
C10654 row_n[13] col[27] 0.0342f
C10655 row_n[4] col[9] 0.0342f
C10656 rowon_n[4] col[10] 0.0323f
C10657 row_n[1] col[3] 0.0342f
C10658 rowon_n[3] col[8] 0.0323f
C10659 rowon_n[15] sample_n 0.0693f
C10660 row_n[10] col[21] 0.0342f
C10661 rowon_n[2] col[6] 0.0323f
C10662 rowon_n[7] col[16] 0.0323f
C10663 col_n[24] a_2475_10186# 0.0531f
C10664 row_n[2] col[5] 0.0342f
C10665 rowon_n[6] col[14] 0.0323f
C10666 rowon_n[5] col[12] 0.0323f
C10667 row_n[15] col[31] 0.0342f
C10668 rowon_n[9] col[20] 0.0323f
C10669 row_n[5] col[11] 0.0342f
C10670 row_n[3] col[7] 0.0342f
C10671 rowon_n[14] col[30] 0.0323f
C10672 col_n[31] rowoff_n[15] 0.0471f
C10673 rowon_n[13] col[28] 0.0323f
C10674 row_n[9] col[19] 0.0342f
C10675 rowon_n[10] col[22] 0.0323f
C10676 row_n[0] col[1] 0.0342f
C10677 row_n[11] col[23] 0.0342f
C10678 row_n[6] col[13] 0.0342f
C10679 rowon_n[0] col[2] 0.0323f
C10680 row_n[14] col[29] 0.0342f
C10681 ctop a_2275_8178# 0.0683f
C10682 a_30986_17190# a_31382_17230# 0.0313f
C10683 VDD a_11398_13536# 0.0779f
C10684 row_n[8] a_15926_10162# 0.0437f
C10685 rowoff_n[0] a_22442_2492# 0.0133f
C10686 rowoff_n[7] a_4974_9158# 0.294f
C10687 col_n[10] a_13310_1166# 0.0839f
C10688 rowon_n[12] a_15014_14178# 0.248f
C10689 a_2475_4162# a_6890_4138# 0.264f
C10690 col_n[20] a_23350_13214# 0.084f
C10691 a_2275_4162# a_4274_4178# 0.144f
C10692 m3_11904_18146# ctop 0.209f
C10693 a_2275_9182# a_29070_9158# 0.399f
C10694 m2_4168_8402# row_n[6] 0.0128f
C10695 a_15014_9158# a_15318_9198# 0.0931f
C10696 a_15926_9158# a_16418_9520# 0.0658f
C10697 col[14] a_2475_7174# 0.136f
C10698 rowoff_n[13] a_12002_15182# 0.294f
C10699 m2_10192_4386# row_n[2] 0.0128f
C10700 m2_34864_15002# a_35002_15182# 0.225f
C10701 rowon_n[2] a_25054_4138# 0.248f
C10702 vcm a_6890_17190# 0.1f
C10703 rowon_n[14] a_3878_16186# 0.118f
C10704 a_27062_14178# a_28066_14178# 0.843f
C10705 VDD a_2874_7150# 0.182f
C10706 col_n[31] a_34490_7512# 0.0283f
C10707 rowoff_n[5] a_14010_7150# 0.294f
C10708 a_2275_18218# a_7894_18194# 0.136f
C10709 VDD a_26458_17552# 0.0779f
C10710 col_n[21] a_2275_13198# 0.113f
C10711 vcm a_8990_2130# 0.56f
C10712 col_n[26] a_2275_2154# 0.113f
C10713 a_2275_6170# a_19334_6186# 0.144f
C10714 a_11910_6146# a_12002_6146# 0.326f
C10715 a_2475_6170# a_21950_6146# 0.264f
C10716 rowoff_n[3] a_23046_5142# 0.294f
C10717 row_n[2] a_2874_4138# 0.0436f
C10718 col[14] a_17022_11166# 0.367f
C10719 m2_19228_17438# row_n[15] 0.0128f
C10720 m2_25252_13422# row_n[11] 0.0128f
C10721 rowon_n[6] a_2161_8178# 0.0177f
C10722 col[11] a_13918_1126# 0.0682f
C10723 m2_31276_9406# row_n[7] 0.0128f
C10724 col[21] a_23958_13174# 0.0682f
C10725 a_18026_16186# a_18026_15182# 0.843f
C10726 VDD a_18026_11166# 0.483f
C10727 col[18] rowoff_n[12] 0.0901f
C10728 col[11] a_2275_10186# 0.0899f
C10729 m2_1732_16006# m3_1864_15134# 0.0341f
C10730 col_n[29] a_32082_7150# 0.251f
C10731 a_6890_3134# a_7286_3174# 0.0313f
C10732 a_2275_3158# a_12914_3134# 0.136f
C10733 a_2475_18218# a_5886_18194# 0.264f
C10734 rowoff_n[1] a_32082_3134# 0.294f
C10735 a_26058_1126# a_2275_1150# 0.0924f
C10736 row_n[13] a_23350_15222# 0.0117f
C10737 vcm a_24050_6146# 0.56f
C10738 m2_15788_946# col_n[13] 0.331f
C10739 rowoff_n[11] a_18426_13536# 0.0133f
C10740 a_2275_8178# a_35398_8194# 0.145f
C10741 col_n[9] a_12306_11206# 0.084f
C10742 col[31] a_2475_9182# 0.136f
C10743 a_30074_13174# a_30378_13214# 0.0931f
C10744 a_30986_13174# a_31478_13536# 0.0658f
C10745 row_n[3] a_33390_5182# 0.0117f
C10746 row_n[15] a_13918_17190# 0.0437f
C10747 a_2475_17214# a_15014_17190# 0.316f
C10748 a_7986_17190# a_8990_17190# 0.843f
C10749 VDD a_33086_15182# 0.483f
C10750 col_n[20] a_23446_5504# 0.0283f
C10751 col_n[30] a_33486_17552# 0.0283f
C10752 row_n[5] a_23958_7150# 0.0437f
C10753 col_n[1] a_2475_6170# 0.0531f
C10754 a_2275_5166# a_27974_5142# 0.136f
C10755 rowon_n[9] a_23046_11166# 0.248f
C10756 vcm a_4974_9158# 0.56f
C10757 a_27974_1126# a_28370_1166# 0.0313f
C10758 rowoff_n[15] a_34490_17552# 0.0133f
C10759 a_26970_10162# a_27062_10162# 0.326f
C10760 m2_32280_16434# a_32082_16186# 0.165f
C10761 m2_31852_946# a_32082_2130# 0.843f
C10762 m2_23820_946# a_2475_1150# 0.286f
C10763 col[2] rowoff_n[13] 0.0901f
C10764 m3_10900_1078# a_10998_2130# 0.0302f
C10765 m2_8760_18014# col_n[6] 0.243f
C10766 a_2275_14202# a_5978_14178# 0.399f
C10767 col[3] a_5978_9158# 0.367f
C10768 m2_34864_8978# m3_34996_9110# 3.79f
C10769 col[28] a_2275_12194# 0.0899f
C10770 col[10] a_12914_11166# 0.0682f
C10771 VDD a_14010_18194# 0.0356f
C10772 a_2475_2154# a_20034_2130# 0.316f
C10773 a_28066_3134# a_28066_2130# 0.843f
C10774 m2_15212_1374# VDD 0.0194f
C10775 col_n[18] a_21038_5142# 0.251f
C10776 vcm a_29374_4178# 0.155f
C10777 rowoff_n[9] a_24962_11166# 0.202f
C10778 a_21950_7150# a_22346_7190# 0.0313f
C10779 col_n[28] a_31078_17190# 0.251f
C10780 col_n[25] a_27974_7150# 0.0765f
C10781 vcm a_20034_13174# 0.56f
C10782 VDD a_16930_3134# 0.181f
C10783 m2_21812_18014# a_2275_18218# 0.28f
C10784 m2_7756_18014# a_8290_18234# 0.087f
C10785 a_2275_16210# a_21038_16186# 0.399f
C10786 a_11910_16186# a_12402_16548# 0.0658f
C10787 a_10998_16186# a_11302_16226# 0.0931f
C10788 rowon_n[3] a_10906_5142# 0.118f
C10789 col[1] a_3878_9158# 0.0682f
C10790 rowoff_n[7] a_33998_9158# 0.202f
C10791 a_18026_4138# a_19030_4138# 0.843f
C10792 a_2475_4162# a_35094_4138# 0.0299f
C10793 col_n[9] a_12402_3496# 0.0283f
C10794 m2_34864_6970# a_35398_7190# 0.087f
C10795 col_n[18] a_2475_8178# 0.0531f
C10796 vcm a_10298_7190# 0.155f
C10797 col_n[19] a_22442_15544# 0.0283f
C10798 rowoff_n[12] a_6378_14540# 0.0133f
C10799 row_n[10] a_31382_12210# 0.0117f
C10800 m2_23244_14426# a_23046_14178# 0.165f
C10801 ctop a_23046_2130# 4.06f
C10802 vcm a_35094_17190# 0.165f
C10803 a_2475_13198# a_13918_13174# 0.264f
C10804 a_2275_13198# a_11302_13214# 0.144f
C10805 a_7894_13174# a_7986_13174# 0.326f
C10806 VDD a_31990_7150# 0.181f
C10807 m2_17796_18014# a_2475_18218# 0.286f
C10808 col[3] a_2475_16210# 0.136f
C10809 row_n[12] a_21950_14178# 0.0437f
C10810 col[8] a_2475_5166# 0.136f
C10811 a_8990_6146# a_8990_5142# 0.843f
C10812 col_n[7] a_9994_3134# 0.251f
C10813 vcm a_25358_11206# 0.155f
C10814 row_n[2] a_31990_4138# 0.0437f
C10815 a_2275_10186# a_4882_10162# 0.136f
C10816 a_2966_10162# a_3970_10162# 0.843f
C10817 VDD a_23446_1488# 0.0977f
C10818 col_n[17] a_20034_15182# 0.251f
C10819 rowon_n[6] a_31078_8154# 0.248f
C10820 ctop a_3970_5142# 4.11f
C10821 col_n[14] a_16930_5142# 0.0765f
C10822 col_n[15] a_2275_11190# 0.113f
C10823 a_2475_15206# a_28978_15182# 0.264f
C10824 a_2275_15206# a_26362_15222# 0.144f
C10825 VDD a_12914_10162# 0.181f
C10826 col_n[24] a_26970_17190# 0.0765f
C10827 m2_1732_12994# m3_1864_12122# 0.0341f
C10828 a_21038_3134# a_21342_3174# 0.0931f
C10829 a_2475_18218# a_34090_18194# 0.0299f
C10830 a_21950_3134# a_22442_3496# 0.0658f
C10831 vcm a_18938_5142# 0.1f
C10832 a_33086_8154# a_34090_8154# 0.843f
C10833 rowoff_n[10] a_12914_12170# 0.202f
C10834 row_n[10] sample_n 0.0596f
C10835 row_n[9] col[30] 0.0342f
C10836 rowon_n[8] col[29] 0.0323f
C10837 rowon_n[1] col[15] 0.0323f
C10838 row_n[3] col[18] 0.0342f
C10839 rowon_n[3] col[19] 0.0323f
C10840 row_n[5] col[22] 0.0342f
C10841 ctop col[9] 0.123f
C10842 row_n[2] col[16] 0.0342f
C10843 row_n[1] col[14] 0.0342f
C10844 rowon_n[5] col[23] 0.0323f
C10845 rowon_n[7] col[27] 0.0323f
C10846 row_n[8] col[28] 0.0342f
C10847 rowon_n[2] col[17] 0.0323f
C10848 row_n[0] col[12] 0.0342f
C10849 row_n[7] col[26] 0.0342f
C10850 col[1] col[2] 0.0337f
C10851 rowon_n[9] col[31] 0.0323f
C10852 rowon_n[6] col[25] 0.0323f
C10853 rowon_n[4] col[21] 0.0323f
C10854 row_n[6] col[24] 0.0342f
C10855 row_n[4] col[20] 0.0342f
C10856 rowon_n[0] col[13] 0.0323f
C10857 a_32082_1126# vcm 0.165f
C10858 m2_14208_12418# a_14010_12170# 0.165f
C10859 m2_9188_16434# rowon_n[14] 0.0322f
C10860 col[5] a_2275_8178# 0.0899f
C10861 row_n[6] a_8990_8154# 0.282f
C10862 m2_15212_12418# rowon_n[10] 0.0322f
C10863 vcm a_6282_14218# 0.155f
C10864 m2_21236_8402# rowon_n[6] 0.0322f
C10865 col_n[8] a_11398_13536# 0.0283f
C10866 m2_27260_4386# rowon_n[2] 0.0322f
C10867 a_2275_12194# a_19942_12170# 0.136f
C10868 VDD a_4370_4500# 0.0779f
C10869 rowon_n[10] a_8898_12170# 0.118f
C10870 col_n[31] a_34394_4178# 0.084f
C10871 m2_34864_18014# VDD 1.4f
C10872 ctop a_19030_9158# 4.11f
C10873 col[27] a_30074_2130# 0.367f
C10874 a_22954_17190# a_23046_17190# 0.326f
C10875 VDD a_27974_14178# 0.181f
C10876 rowoff_n[0] a_4882_2130# 0.202f
C10877 rowon_n[0] a_18938_2130# 0.118f
C10878 col[25] a_2475_7174# 0.136f
C10879 m2_33284_8402# a_33086_8154# 0.165f
C10880 vcm a_33998_9158# 0.1f
C10881 m2_16792_18014# m2_17220_18442# 0.165f
C10882 rowoff_n[14] a_28978_16186# 0.202f
C10883 a_24050_10162# a_24050_9158# 0.843f
C10884 a_2475_9182# a_12002_9158# 0.316f
C10885 vcm a_21342_18234# 0.16f
C10886 a_2275_14202# a_35002_14178# 0.136f
C10887 a_17934_14178# a_18330_14218# 0.0313f
C10888 col_n[22] a_25358_2170# 0.084f
C10889 m2_35292_17438# rowon_n[15] 0.0322f
C10890 VDD a_19430_8516# 0.0779f
C10891 m2_34864_5966# m3_34996_6098# 3.79f
C10892 col_n[6] a_8990_13174# 0.251f
C10893 m2_34864_946# vcm 0.408f
C10894 ctop a_34090_13174# 4.06f
C10895 col_n[3] a_5886_3134# 0.0765f
C10896 VDD a_8898_17190# 0.181f
C10897 analog_in a_34090_2130# 0.0385f
C10898 col_n[13] a_15926_15182# 0.0765f
C10899 m3_10900_1078# VDD 0.0157f
C10900 row_n[9] a_29982_11166# 0.0437f
C10901 a_2475_6170# a_3878_6146# 0.264f
C10902 a_2275_6170# a_2874_6146# 0.136f
C10903 en_bit_n[1] a_18330_1166# 0.0266f
C10904 m2_5172_10410# a_4974_10162# 0.165f
C10905 rowon_n[13] a_29070_15182# 0.248f
C10906 vcm a_14922_12170# 0.1f
C10907 rowoff_n[3] a_5374_5504# 0.0133f
C10908 a_14010_11166# a_15014_11166# 0.843f
C10909 a_2475_11190# a_27062_11166# 0.316f
C10910 col[22] a_2275_10186# 0.0899f
C10911 VDD a_10998_2130# 0.483f
C10912 col[29] rowoff_n[12] 0.0901f
C10913 m2_26832_18014# a_27366_18234# 0.087f
C10914 VDD a_34490_12532# 0.0779f
C10915 m2_25828_18014# m3_24956_18146# 0.0341f
C10916 ctop a_15014_16186# 4.11f
C10917 a_32994_4138# a_33086_4138# 0.326f
C10918 col[26] a_29070_12170# 0.367f
C10919 rowoff_n[1] a_14410_3496# 0.0133f
C10920 col[23] a_25966_2130# 0.0682f
C10921 m2_24248_6394# a_24050_6146# 0.165f
C10922 row_n[13] a_6982_15182# 0.282f
C10923 a_2275_8178# a_18026_8154# 0.399f
C10924 vcm a_29982_16186# 0.1f
C10925 a_4974_13174# a_4974_12170# 0.843f
C10926 VDD a_26058_6146# 0.483f
C10927 row_n[3] a_17022_5142# 0.282f
C10928 col_n[7] a_2475_17214# 0.0531f
C10929 a_32994_18194# a_33390_18234# 0.0313f
C10930 rowon_n[7] a_16930_9158# 0.118f
C10931 VDD a_15414_15544# 0.0779f
C10932 rowoff_n[6] a_5978_8154# 0.294f
C10933 col_n[12] a_2475_6170# 0.0531f
C10934 col_n[21] a_24354_12210# 0.084f
C10935 row_n[5] a_4274_7190# 0.0117f
C10936 a_2275_5166# a_8290_5182# 0.144f
C10937 a_2475_5166# a_10906_5142# 0.264f
C10938 col_n[2] a_4882_13174# 0.0765f
C10939 m2_28840_946# m3_29976_1078# 0.0341f
C10940 col[13] rowoff_n[13] 0.0901f
C10941 a_2275_10186# a_33086_10162# 0.399f
C10942 a_17934_10162# a_18426_10524# 0.0658f
C10943 a_17022_10162# a_17326_10202# 0.0931f
C10944 rowoff_n[15] a_16930_17190# 0.202f
C10945 rowoff_n[4] a_15014_6146# 0.294f
C10946 col[2] a_2475_3158# 0.136f
C10947 a_29070_15182# a_30074_15182# 0.843f
C10948 VDD a_6982_9158# 0.483f
C10949 m2_1732_9982# m3_1864_9110# 0.0341f
C10950 m2_8184_15430# row_n[13] 0.0128f
C10951 a_2475_2154# a_1957_2154# 0.0734f
C10952 m2_14208_11414# row_n[9] 0.0128f
C10953 m2_20232_7398# row_n[5] 0.0128f
C10954 m2_15212_4386# a_15014_4138# 0.165f
C10955 m2_26256_3382# row_n[1] 0.0128f
C10956 vcm a_13006_4138# 0.56f
C10957 rowoff_n[2] a_24050_4138# 0.294f
C10958 rowon_n[1] a_3970_3134# 0.248f
C10959 a_2275_7174# a_23350_7190# 0.144f
C10960 a_2475_7174# a_25966_7150# 0.264f
C10961 a_13918_7150# a_14010_7150# 0.326f
C10962 col_n[9] a_2275_9182# 0.113f
C10963 col[15] a_18026_10162# 0.367f
C10964 m2_1732_10986# a_2275_11190# 0.191f
C10965 vcm a_1957_13198# 0.139f
C10966 col[22] a_24962_12170# 0.0682f
C10967 a_2275_16210# a_2966_16186# 0.399f
C10968 a_2475_16210# a_3970_16186# 0.316f
C10969 a_20034_17190# a_20034_16186# 0.843f
C10970 col_n[30] a_33086_6146# 0.251f
C10971 VDD a_22042_13174# 0.483f
C10972 ctop a_2275_17214# 0.0683f
C10973 rowoff_n[0] a_33086_2130# 0.294f
C10974 col_n[29] a_2475_8178# 0.0531f
C10975 a_2275_4162# a_16930_4138# 0.136f
C10976 a_8898_4138# a_9294_4178# 0.0313f
C10977 m3_34996_8106# ctop 0.209f
C10978 col_n[10] a_13310_10202# 0.084f
C10979 m2_34864_16006# row_n[14] 0.267f
C10980 vcm a_28066_8154# 0.56f
C10981 row_n[10] a_15014_12170# 0.282f
C10982 rowon_n[14] a_14922_16186# 0.118f
C10983 col[14] a_2475_16210# 0.136f
C10984 a_32994_14178# a_33486_14540# 0.0658f
C10985 a_32082_14178# a_32386_14218# 0.0931f
C10986 m2_34864_2954# m3_34996_3086# 3.79f
C10987 col[19] a_2475_5166# 0.136f
C10988 col_n[21] a_24450_4500# 0.0283f
C10989 VDD a_2874_16186# 0.182f
C10990 row_n[0] a_25054_2130# 0.282f
C10991 col_n[31] a_34490_16548# 0.0283f
C10992 a_2475_1150# a_8990_1126# 0.0299f
C10993 row_n[12] a_3878_14178# 0.0437f
C10994 rowon_n[4] a_24962_6146# 0.118f
C10995 vcm a_18330_2170# 0.155f
C10996 a_2275_6170# a_31990_6146# 0.136f
C10997 m2_7756_946# m2_8760_946# 0.843f
C10998 col_n[26] a_2275_11190# 0.113f
C10999 vcm a_8990_11166# 0.56f
C11000 row_n[2] a_12306_4178# 0.0117f
C11001 a_28978_11166# a_29070_11166# 0.326f
C11002 VDD a_5886_1126# 0.405f
C11003 col[4] a_6982_8154# 0.367f
C11004 a_2275_15206# a_9994_15182# 0.399f
C11005 col[11] a_13918_10162# 0.0682f
C11006 row_n[4] a_2161_6170# 0.0221f
C11007 col_n[19] a_22042_4138# 0.251f
C11008 row_n[3] col[29] 0.0342f
C11009 row_n[4] col[31] 0.0342f
C11010 row_n[0] col[23] 0.0342f
C11011 rowon_n[8] a_2475_10186# 0.31f
C11012 rowon_n[3] col[30] 0.0323f
C11013 rowon_n[1] col[26] 0.0323f
C11014 a_2475_3158# a_24050_3134# 0.316f
C11015 row_n[1] col[25] 0.0342f
C11016 row_n[2] col[27] 0.0342f
C11017 rowon_n[4] sample_n 0.0692f
C11018 rowon_n[0] col[24] 0.0323f
C11019 ctop col[20] 0.123f
C11020 rowon_n[2] col[28] 0.0323f
C11021 a_30074_4138# a_30074_3134# 0.843f
C11022 rowoff_n[8] a_25966_10162# 0.202f
C11023 col[16] a_2275_8178# 0.0899f
C11024 col_n[29] a_32082_16186# 0.251f
C11025 row_n[13] a_34394_15222# 0.0117f
C11026 col_n[26] a_28978_6146# 0.0765f
C11027 vcm a_33390_6186# 0.155f
C11028 a_23958_8154# a_24354_8194# 0.0313f
C11029 rowoff_n[11] a_29070_13174# 0.294f
C11030 m2_34864_12994# a_34090_13174# 0.843f
C11031 vcm a_24050_15182# 0.56f
C11032 VDD a_20946_5142# 0.181f
C11033 a_26362_1166# col_n[23] 0.0839f
C11034 a_35094_1126# VDD 0.0351f
C11035 a_13006_17190# a_13310_17230# 0.0931f
C11036 a_2275_17214# a_25054_17190# 0.399f
C11037 a_13918_17190# a_14410_17552# 0.0658f
C11038 rowoff_n[6] a_35002_8154# 0.202f
C11039 col_n[10] a_13406_2492# 0.0283f
C11040 m3_30980_18146# a_31078_17190# 0.0303f
C11041 a_20034_5142# a_21038_5142# 0.843f
C11042 col_n[20] a_23446_14540# 0.0283f
C11043 m3_31984_1078# m3_32988_1078# 0.202f
C11044 vcm a_14314_9198# 0.155f
C11045 col_n[1] a_2475_15206# 0.0531f
C11046 col_n[6] a_2475_4162# 0.0531f
C11047 vcm a_4974_18194# 0.165f
C11048 ctop a_27062_4138# 4.11f
C11049 m2_15788_946# a_16018_1126# 0.0249f
C11050 a_2275_14202# a_15318_14218# 0.144f
C11051 a_9902_14178# a_9994_14178# 0.326f
C11052 a_2475_14202# a_17934_14178# 0.264f
C11053 row_n[7] a_23046_9158# 0.282f
C11054 m2_1732_6970# m3_1864_6098# 0.0341f
C11055 m2_34864_7974# rowoff_n[6] 0.278f
C11056 rowon_n[11] a_22954_13174# 0.118f
C11057 VDD a_23350_18234# 0.019f
C11058 a_2275_2154# a_30074_2130# 0.399f
C11059 m2_25828_946# col_n[23] 0.331f
C11060 m3_6884_18146# VDD 0.0864f
C11061 vcm a_7894_3134# 0.1f
C11062 row_n[9] a_10298_11206# 0.0117f
C11063 rowon_n[1] a_32994_3134# 0.118f
C11064 a_10998_7150# a_10998_6146# 0.843f
C11065 rowoff_n[9] a_35494_11528# 0.0133f
C11066 col_n[8] a_10998_2130# 0.251f
C11067 a_26970_1126# col[24] 0.0682f
C11068 en_bit_n[1] a_2475_1150# 0.0162f
C11069 col_n[18] a_21038_14178# 0.251f
C11070 vcm a_29374_13214# 0.155f
C11071 col_n[15] a_17934_4138# 0.0765f
C11072 a_4882_11166# a_5278_11206# 0.0313f
C11073 a_2275_11190# a_8898_11166# 0.136f
C11074 VDD a_27462_3496# 0.0779f
C11075 m2_23820_18014# col[21] 0.347f
C11076 col_n[25] a_27974_16186# 0.0765f
C11077 ctop a_7986_7150# 4.11f
C11078 a_2275_16210# a_30378_16226# 0.144f
C11079 a_2475_16210# a_32994_16186# 0.264f
C11080 VDD a_16930_12170# 0.181f
C11081 m2_1732_18014# m3_1864_18146# 3.79f
C11082 m2_4168_10410# rowon_n[8] 0.0322f
C11083 col_n[3] a_2275_7174# 0.113f
C11084 m2_10192_6394# rowon_n[4] 0.0322f
C11085 m2_15212_2378# rowon_n[0] 0.0322f
C11086 a_23958_4138# a_24450_4500# 0.0658f
C11087 a_23046_4138# a_23350_4178# 0.0931f
C11088 col[1] a_3878_18194# 0.0682f
C11089 row_n[1] a_10906_3134# 0.0437f
C11090 vcm a_22954_7150# 0.1f
C11091 rowon_n[5] a_9994_7150# 0.248f
C11092 rowoff_n[12] a_17022_14178# 0.294f
C11093 col_n[9] a_12402_12532# 0.0283f
C11094 col_n[18] a_2475_17214# 0.0531f
C11095 vcm a_10298_16226# 0.155f
C11096 a_2275_13198# a_23958_13174# 0.136f
C11097 VDD a_8386_6508# 0.0779f
C11098 col_n[23] a_2475_6170# 0.0531f
C11099 ctop a_23046_11166# 4.11f
C11100 a_24962_18194# a_25054_18194# 0.0991f
C11101 VDD a_31990_16186# 0.181f
C11102 a_19942_1126# a_20034_1126# 0.354f
C11103 col[24] rowoff_n[13] 0.0901f
C11104 m2_25252_15430# rowon_n[13] 0.0322f
C11105 m2_31276_11414# rowon_n[9] 0.0322f
C11106 col[8] a_2475_14202# 0.136f
C11107 m2_4744_946# m3_3872_1078# 0.0341f
C11108 col_n[0] rowoff_n[1] 0.0471f
C11109 col_n[6] rowoff_n[8] 0.0471f
C11110 vcm rowoff_n[2] 0.533f
C11111 col[13] a_2475_3158# 0.136f
C11112 col_n[4] rowoff_n[6] 0.0471f
C11113 col_n[5] rowoff_n[7] 0.0471f
C11114 col_n[1] rowoff_n[3] 0.0471f
C11115 col_n[2] rowoff_n[4] 0.0471f
C11116 col_n[7] rowoff_n[9] 0.0471f
C11117 col_n[3] rowoff_n[5] 0.0471f
C11118 sample rowoff_n[0] 0.0775f
C11119 a_2475_10186# a_16018_10162# 0.316f
C11120 a_26058_11166# a_26058_10162# 0.843f
C11121 row_n[14] a_21038_16186# 0.282f
C11122 col_n[7] a_9994_12170# 0.251f
C11123 a_19942_15182# a_20338_15222# 0.0313f
C11124 col_n[4] a_6890_2130# 0.0765f
C11125 VDD a_23446_10524# 0.0779f
C11126 ctop a_3970_14178# 4.11f
C11127 col_n[14] a_16930_14178# 0.0765f
C11128 row_n[4] a_31078_6146# 0.282f
C11129 rowon_n[8] a_30986_10162# 0.118f
C11130 col_n[20] a_2275_9182# 0.113f
C11131 rowoff_n[10] a_23446_12532# 0.0133f
C11132 rowoff_n[2] a_6378_4500# 0.0133f
C11133 a_3970_7150# a_4274_7190# 0.0931f
C11134 a_4882_7150# a_5374_7512# 0.0658f
C11135 a_2275_7174# a_6982_7150# 0.399f
C11136 m2_16792_18014# vcm 0.353f
C11137 row_n[6] a_18330_8194# 0.0117f
C11138 vcm a_18938_14178# 0.1f
C11139 a_2475_12194# a_31078_12170# 0.316f
C11140 a_16018_12170# a_17022_12170# 0.843f
C11141 VDD a_15014_4138# 0.483f
C11142 col[5] a_2275_17214# 0.0899f
C11143 row_n[0] m2_31276_2378# 0.0128f
C11144 VDD a_4370_13536# 0.0779f
C11145 col[10] a_2275_6170# 0.0899f
C11146 col_n[31] a_34394_13214# 0.084f
C11147 col[8] rowoff_n[14] 0.0901f
C11148 col[27] a_30074_11166# 0.367f
C11149 row_n[8] a_8898_10162# 0.0437f
C11150 rowoff_n[0] a_15414_2492# 0.0133f
C11151 rowon_n[12] a_7986_14178# 0.248f
C11152 a_34090_5142# a_34394_5182# 0.0931f
C11153 a_35002_5142# a_35094_5142# 0.0991f
C11154 m2_26832_946# ctop 0.0428f
C11155 col[25] a_2475_16210# 0.136f
C11156 rowoff_n[13] a_4974_15182# 0.294f
C11157 a_2275_9182# a_22042_9158# 0.399f
C11158 col[30] a_2475_5166# 0.136f
C11159 m2_29268_15430# a_29070_15182# 0.165f
C11160 rowon_n[2] a_18026_4138# 0.248f
C11161 vcm a_33998_18194# 0.101f
C11162 a_6982_14178# a_6982_13174# 0.843f
C11163 VDD a_30074_8154# 0.483f
C11164 m2_1732_3958# m3_1864_3086# 0.0341f
C11165 rowoff_n[5] a_6982_7150# 0.294f
C11166 col_n[22] a_25358_11206# 0.084f
C11167 VDD a_19430_17552# 0.0779f
C11168 row_n[0] m2_20232_2378# 0.0128f
C11169 a_29982_2130# a_30378_2170# 0.0313f
C11170 col_n[3] a_5886_12170# 0.0765f
C11171 vcm a_2475_2154# 1.08f
C11172 a_2475_6170# a_14922_6146# 0.264f
C11173 a_2275_6170# a_12306_6186# 0.144f
C11174 rowoff_n[3] a_16018_5142# 0.294f
C11175 a_19942_11166# a_20434_11528# 0.0658f
C11176 a_19030_11166# a_19334_11206# 0.0931f
C11177 m2_3164_9406# row_n[7] 0.0128f
C11178 m2_9188_5390# row_n[3] 0.0128f
C11179 row_n[11] a_29070_13174# 0.282f
C11180 a_31078_16186# a_32082_16186# 0.843f
C11181 VDD col_n[8] 5.17f
C11182 VDD a_10998_11166# 0.483f
C11183 vcm col_n[5] 1.94f
C11184 col_n[2] col_n[3] 0.0101f
C11185 ctop col[31] 0.456f
C11186 col[12] col[13] 0.0355f
C11187 rowon_n[15] a_28978_17190# 0.118f
C11188 col[27] a_2275_8178# 0.0899f
C11189 a_2275_3158# a_5886_3134# 0.136f
C11190 rowoff_n[1] a_25054_3134# 0.294f
C11191 col[16] a_19030_9158# 0.367f
C11192 row_n[13] a_16322_15222# 0.0117f
C11193 vcm a_17022_6146# 0.56f
C11194 rowoff_n[11] a_11398_13536# 0.0133f
C11195 a_2475_8178# a_29982_8154# 0.264f
C11196 a_2275_8178# a_27366_8194# 0.144f
C11197 a_15926_8154# a_16018_8154# 0.326f
C11198 m2_20232_13422# a_20034_13174# 0.165f
C11199 col[23] a_25966_11166# 0.0682f
C11200 m2_1732_9982# sample 0.2f
C11201 VDD a_2275_5166# 1.96f
C11202 m2_34864_3958# ctop 0.0422f
C11203 col_n[31] a_34090_5142# 0.251f
C11204 row_n[3] a_26362_5182# 0.0117f
C11205 row_n[15] a_6890_17190# 0.0437f
C11206 m2_24248_14426# row_n[12] 0.0128f
C11207 a_2475_17214# a_7986_17190# 0.316f
C11208 VDD a_26058_15182# 0.483f
C11209 m2_30272_10410# row_n[8] 0.0128f
C11210 m2_35292_6394# row_n[4] 0.0128f
C11211 col_n[11] a_14314_9198# 0.084f
C11212 col_n[12] a_2475_15206# 0.0531f
C11213 a_10906_5142# a_11302_5182# 0.0313f
C11214 row_n[5] a_16930_7150# 0.0437f
C11215 a_2275_5166# a_20946_5142# 0.136f
C11216 m3_34996_4090# m3_34996_3086# 0.202f
C11217 col_n[17] a_2475_4162# 0.0531f
C11218 rowon_n[9] a_16018_11166# 0.248f
C11219 vcm a_32082_10162# 0.56f
C11220 rowoff_n[15] a_27462_17552# 0.0133f
C11221 m2_6752_946# a_2275_1150# 0.28f
C11222 col_n[22] a_25454_3496# 0.0283f
C11223 a_35002_15182# a_35494_15544# 0.0658f
C11224 m2_4168_1374# a_3970_1126# 0.165f
C11225 col[2] a_2475_12194# 0.136f
C11226 VDD a_6982_18194# 0.0356f
C11227 a_6982_2130# a_7986_2130# 0.843f
C11228 col[7] a_2475_1150# 0.136f
C11229 a_2475_2154# a_13006_2130# 0.316f
C11230 vcm a_22346_4178# 0.155f
C11231 a_2275_7174# a_34394_7190# 0.144f
C11232 rowoff_n[9] a_17934_11166# 0.202f
C11233 m2_11196_11414# a_10998_11166# 0.165f
C11234 col[5] a_7986_7150# 0.367f
C11235 vcm a_13006_13174# 0.56f
C11236 a_30986_12170# a_31078_12170# 0.326f
C11237 VDD a_9902_3134# 0.181f
C11238 col_n[9] a_2275_18218# 0.113f
C11239 m2_7756_18014# a_2275_18218# 0.28f
C11240 col[12] a_14922_9158# 0.0682f
C11241 col_n[14] a_2275_7174# 0.113f
C11242 a_2275_16210# a_14010_16186# 0.399f
C11243 col_n[20] a_23046_3134# 0.251f
C11244 col[16] a_17934_1126# 0.011f
C11245 rowoff_n[7] a_26970_9158# 0.202f
C11246 col_n[30] a_33086_15182# 0.251f
C11247 col_n[27] a_29982_5142# 0.0765f
C11248 a_32082_5142# a_32082_4138# 0.843f
C11249 a_2475_4162# a_28066_4138# 0.316f
C11250 m3_30980_1078# ctop 0.21f
C11251 m2_30272_7398# a_30074_7150# 0.165f
C11252 col_n[29] a_2475_17214# 0.0531f
C11253 vcm a_3270_7190# 0.155f
C11254 a_25966_9158# a_26362_9198# 0.0313f
C11255 rowoff_n[13] a_33998_15182# 0.202f
C11256 col[4] a_2275_4162# 0.0899f
C11257 row_n[10] a_24354_12210# 0.0117f
C11258 vcm a_28066_17190# 0.56f
C11259 ctop a_16018_2130# 4.06f
C11260 a_2275_13198# a_4274_13214# 0.144f
C11261 a_2475_13198# a_6890_13174# 0.264f
C11262 VDD a_24962_7150# 0.181f
C11263 a_2275_18218# a_29070_18194# 0.0924f
C11264 m2_3740_18014# a_2475_18218# 0.286f
C11265 a_15926_18194# a_16418_18556# 0.0658f
C11266 col_n[11] a_14410_1488# 0.0283f
C11267 row_n[0] a_35398_2170# 0.0117f
C11268 a_10906_1126# a_11398_1488# 0.0658f
C11269 col[19] a_2475_14202# 0.136f
C11270 row_n[12] a_14922_14178# 0.0437f
C11271 a_2275_1150# a_19030_1126# 0.399f
C11272 col_n[21] a_24450_13536# 0.0283f
C11273 col_n[10] rowoff_n[1] 0.0471f
C11274 col[24] a_2475_3158# 0.136f
C11275 col_n[15] rowoff_n[6] 0.0471f
C11276 col_n[16] rowoff_n[7] 0.0471f
C11277 col_n[9] rowoff_n[0] 0.0471f
C11278 col_n[17] rowoff_n[8] 0.0471f
C11279 col_n[14] rowoff_n[5] 0.0471f
C11280 col_n[12] rowoff_n[3] 0.0471f
C11281 col_n[13] rowoff_n[4] 0.0471f
C11282 col_n[18] rowoff_n[9] 0.0471f
C11283 col_n[11] rowoff_n[2] 0.0471f
C11284 vcm a_30986_2130# 0.1f
C11285 m2_1732_4962# m2_2160_5390# 0.165f
C11286 a_22042_6146# a_23046_6146# 0.843f
C11287 m2_1732_8978# a_1957_9182# 0.245f
C11288 vcm a_18330_11206# 0.155f
C11289 row_n[2] a_24962_4138# 0.0437f
C11290 row_n[14] a_2966_16186# 0.281f
C11291 VDD a_16418_1488# 0.0977f
C11292 rowon_n[6] a_24050_8154# 0.248f
C11293 sample a_2161_7174# 0.0858f
C11294 ctop a_31078_6146# 4.11f
C11295 a_11910_15182# a_12002_15182# 0.326f
C11296 a_2275_15206# a_19334_15222# 0.144f
C11297 a_2475_15206# a_21950_15182# 0.264f
C11298 VDD a_5886_10162# 0.181f
C11299 col[4] a_6982_17190# 0.367f
C11300 col_n[31] a_2275_9182# 0.113f
C11301 a_2275_3158# a_34090_3134# 0.399f
C11302 a_2475_18218# a_27062_18194# 0.0299f
C11303 m2_21236_5390# a_21038_5142# 0.165f
C11304 col_n[19] a_22042_13174# 0.251f
C11305 vcm a_11910_5142# 0.1f
C11306 rowoff_n[10] a_5886_12170# 0.202f
C11307 a_13006_8154# a_13006_7150# 0.843f
C11308 a_25054_1126# vcm 0.165f
C11309 col_n[16] a_18938_3134# 0.0765f
C11310 col[16] a_2275_17214# 0.0899f
C11311 row_n[6] a_2475_8178# 0.405f
C11312 vcm a_33390_15222# 0.155f
C11313 col_n[26] a_28978_15182# 0.0765f
C11314 col[21] a_2275_6170# 0.0899f
C11315 a_6890_12170# a_7286_12210# 0.0313f
C11316 a_2275_12194# a_12914_12170# 0.136f
C11317 VDD a_31478_5504# 0.0779f
C11318 col[19] rowoff_n[14] 0.0901f
C11319 m2_20808_18014# VDD 0.993f
C11320 row_n[15] a_35094_17190# 0.0123f
C11321 ctop a_12002_9158# 4.11f
C11322 a_2275_17214# a_35398_17230# 0.145f
C11323 VDD a_20946_14178# 0.181f
C11324 col_n[2] rowoff_n[10] 0.0471f
C11325 rowon_n[0] a_11910_2130# 0.118f
C11326 a_25054_5142# a_25358_5182# 0.0931f
C11327 a_25966_5142# a_26458_5504# 0.0658f
C11328 col_n[10] a_13406_11528# 0.0283f
C11329 vcm a_26970_9158# 0.1f
C11330 m2_9764_18014# m2_10192_18442# 0.165f
C11331 rowoff_n[14] a_21950_16186# 0.202f
C11332 a_2475_9182# a_4974_9158# 0.316f
C11333 vcm a_14314_18234# 0.16f
C11334 m2_8184_17438# rowon_n[15] 0.0322f
C11335 m2_23820_946# a_23958_1126# 0.225f
C11336 a_2275_14202# a_27974_14178# 0.136f
C11337 m2_14208_13422# rowon_n[11] 0.0322f
C11338 VDD a_12402_8516# 0.0779f
C11339 row_n[7] a_32386_9198# 0.0117f
C11340 m2_20232_9406# rowon_n[7] 0.0322f
C11341 m2_26256_5390# rowon_n[3] 0.0322f
C11342 col_n[6] a_2475_13198# 0.0531f
C11343 ctop a_27062_13174# 4.11f
C11344 VDD a_34394_18234# 0.019f
C11345 col_n[11] a_2475_2154# 0.0531f
C11346 a_21950_2130# a_22042_2130# 0.326f
C11347 m2_12200_3382# a_12002_3134# 0.165f
C11348 m2_34864_8978# m2_34864_7974# 0.843f
C11349 row_n[9] a_22954_11166# 0.0437f
C11350 rowon_n[13] a_22042_15182# 0.248f
C11351 vcm a_7894_12170# 0.1f
C11352 vcm col_n[16] 1.93f
C11353 VDD col_n[19] 5.17f
C11354 col_n[8] a_10998_11166# 0.251f
C11355 a_28066_12170# a_28066_11166# 0.843f
C11356 a_2475_11190# a_20034_11166# 0.316f
C11357 VDD a_3970_2130# 0.483f
C11358 col[3] rowoff_n[15] 0.0901f
C11359 col_n[5] a_7894_1126# 0.0765f
C11360 col_n[15] a_17934_13174# 0.0765f
C11361 a_21950_16186# a_22346_16226# 0.0313f
C11362 VDD a_27462_12532# 0.0779f
C11363 rowon_n[3] a_32082_5142# 0.248f
C11364 m2_15788_18014# m3_16924_18146# 0.0341f
C11365 ctop a_7986_16186# 4.11f
C11366 m2_2736_1950# rowoff_n[0] 0.281f
C11367 rowoff_n[1] a_7382_3496# 0.0133f
C11368 col_n[3] a_2275_16210# 0.113f
C11369 col_n[8] a_2275_5166# 0.113f
C11370 a_5978_8154# a_6282_8194# 0.0931f
C11371 a_6890_8154# a_7382_8516# 0.0658f
C11372 a_2275_8178# a_10998_8154# 0.399f
C11373 vcm a_22954_16186# 0.1f
C11374 a_18026_13174# a_19030_13174# 0.843f
C11375 a_2475_13198# a_35094_13174# 0.0299f
C11376 VDD a_19030_6146# 0.483f
C11377 row_n[3] a_9994_5142# 0.282f
C11378 rowon_n[7] a_9902_9158# 0.118f
C11379 col[28] a_31078_10162# 0.367f
C11380 col_n[23] a_2475_15206# 0.0531f
C11381 VDD a_8386_15544# 0.0779f
C11382 col_n[28] a_2475_4162# 0.0531f
C11383 m3_27968_18146# m3_28972_18146# 0.202f
C11384 rowoff_n[15] a_9902_17190# 0.202f
C11385 a_2275_10186# a_26058_10162# 0.399f
C11386 row_n[14] a_30378_16226# 0.0117f
C11387 rowoff_n[4] a_7986_6146# 0.294f
C11388 col[13] a_2475_12194# 0.136f
C11389 m2_14784_946# a_15014_2130# 0.843f
C11390 a_8990_15182# a_8990_14178# 0.843f
C11391 col_n[23] a_26362_10202# 0.084f
C11392 VDD a_34090_10162# 0.483f
C11393 col[18] a_2475_1150# 0.136f
C11394 col_n[4] a_6890_11166# 0.0765f
C11395 a_31990_3134# a_32386_3174# 0.0313f
C11396 vcm a_5978_4138# 0.56f
C11397 rowoff_n[10] a_34090_12170# 0.294f
C11398 rowoff_n[2] a_17022_4138# 0.294f
C11399 a_2275_7174# a_16322_7190# 0.144f
C11400 a_2475_7174# a_18938_7150# 0.264f
C11401 col_n[20] a_2275_18218# 0.113f
C11402 col_n[25] a_2275_7174# 0.113f
C11403 row_n[6] a_30986_8154# 0.0437f
C11404 a_21950_12170# a_22442_12532# 0.0658f
C11405 a_21038_12170# a_21342_12210# 0.0931f
C11406 rowon_n[10] a_30074_12170# 0.248f
C11407 a_33086_17190# a_34090_17190# 0.843f
C11408 VDD a_15014_13174# 0.483f
C11409 rowoff_n[0] a_26058_2130# 0.294f
C11410 col[10] a_2275_15206# 0.0899f
C11411 col[17] a_20034_8154# 0.367f
C11412 a_2275_4162# a_9902_4138# 0.136f
C11413 col[15] a_2275_4162# 0.0899f
C11414 m3_26964_18146# ctop 0.209f
C11415 m2_7180_16434# row_n[14] 0.0128f
C11416 col[24] a_26970_10162# 0.0682f
C11417 m2_13204_12418# row_n[10] 0.0128f
C11418 vcm a_21038_8154# 0.56f
C11419 m2_19228_8402# row_n[6] 0.0128f
C11420 a_2275_9182# a_31382_9198# 0.144f
C11421 a_17934_9158# a_18026_9158# 0.326f
C11422 a_2475_9182# a_33998_9158# 0.264f
C11423 m2_25252_4386# row_n[2] 0.0128f
C11424 row_n[10] a_7986_12170# 0.282f
C11425 m2_3164_14426# a_2966_14178# 0.165f
C11426 rowon_n[14] a_7894_16186# 0.118f
C11427 col[30] a_2475_14202# 0.136f
C11428 col_n[21] rowoff_n[1] 0.0471f
C11429 col_n[23] rowoff_n[3] 0.0471f
C11430 col_n[27] rowoff_n[7] 0.0471f
C11431 col_n[22] rowoff_n[2] 0.0471f
C11432 col_n[20] rowoff_n[0] 0.0471f
C11433 col_n[29] rowoff_n[9] 0.0471f
C11434 col_n[24] rowoff_n[4] 0.0471f
C11435 col_n[26] rowoff_n[6] 0.0471f
C11436 col_n[25] rowoff_n[5] 0.0471f
C11437 col_n[28] rowoff_n[8] 0.0471f
C11438 row_n[0] a_18026_2130# 0.282f
C11439 VDD a_30074_17190# 0.484f
C11440 col_n[12] a_15318_8194# 0.084f
C11441 a_19030_2130# a_19030_1126# 0.843f
C11442 rowon_n[4] a_17934_6146# 0.118f
C11443 col_n[6] a_2475_18218# 0.0529f
C11444 vcm a_11302_2170# 0.155f
C11445 a_2275_6170# a_24962_6146# 0.136f
C11446 a_12914_6146# a_13310_6186# 0.0313f
C11447 row_n[2] a_5278_4178# 0.0117f
C11448 vcm a_2475_11190# 1.08f
C11449 m2_34288_17438# row_n[15] 0.0128f
C11450 col_n[23] a_26458_2492# 0.0283f
C11451 VDD a_32994_2130# 0.181f
C11452 a_2475_15206# a_3878_15182# 0.264f
C11453 a_2275_15206# a_2874_15182# 0.136f
C11454 a_8990_3134# a_9994_3134# 0.843f
C11455 a_2475_3158# a_17022_3134# 0.316f
C11456 rowoff_n[8] a_18938_10162# 0.202f
C11457 col[27] a_2275_17214# 0.0899f
C11458 en_bit_n[2] a_19430_1488# 0.018f
C11459 a_28370_1166# a_2275_1150# 0.145f
C11460 a_30986_1126# a_2475_1150# 0.264f
C11461 row_n[13] a_28978_15182# 0.0437f
C11462 col[6] a_8990_6146# 0.367f
C11463 vcm a_26362_6186# 0.155f
C11464 rowoff_n[11] a_22042_13174# 0.294f
C11465 col[30] rowoff_n[14] 0.0901f
C11466 col[13] a_15926_8154# 0.0682f
C11467 vcm a_17022_15182# 0.56f
C11468 a_32994_13174# a_33086_13174# 0.326f
C11469 VDD a_13918_5142# 0.181f
C11470 a_27062_1126# VDD 0.035f
C11471 col_n[13] rowoff_n[10] 0.0471f
C11472 col_n[21] a_24050_2130# 0.251f
C11473 a_2275_17214# a_18026_17190# 0.399f
C11474 VDD a_2275_14202# 1.96f
C11475 rowoff_n[6] a_27974_8154# 0.202f
C11476 a_21038_2130# m2_21236_2378# 0.165f
C11477 col_n[31] a_34090_14178# 0.251f
C11478 col_n[28] a_30986_4138# 0.0765f
C11479 col_n[2] a_2275_3158# 0.113f
C11480 col_n[1] a_4274_6186# 0.084f
C11481 a_34090_6146# a_34090_5142# 0.843f
C11482 a_2475_5166# a_32082_5142# 0.316f
C11483 m3_34996_2082# m3_34996_1078# 0.202f
C11484 m3_17928_1078# m3_18932_1078# 0.0605f
C11485 col_n[11] a_14314_18234# 0.084f
C11486 vcm a_7286_9198# 0.155f
C11487 rowoff_n[14] a_3878_16186# 0.202f
C11488 a_27974_10162# a_28370_10202# 0.0313f
C11489 col_n[17] a_2475_13198# 0.0531f
C11490 m2_34864_16006# a_35094_16186# 0.0249f
C11491 ctop a_20034_4138# 4.11f
C11492 m3_13912_1078# a_14010_2130# 0.0302f
C11493 a_2475_14202# a_10906_14178# 0.264f
C11494 a_2275_14202# a_8290_14218# 0.144f
C11495 col_n[22] a_2475_2154# 0.0531f
C11496 m2_29844_946# a_2275_1150# 0.28f
C11497 row_n[7] a_16018_9158# 0.282f
C11498 VDD a_28978_9158# 0.181f
C11499 rowon_n[11] a_15926_13174# 0.118f
C11500 col_n[22] a_25454_12532# 0.0283f
C11501 VDD a_16322_18234# 0.019f
C11502 a_2275_2154# a_23046_2130# 0.399f
C11503 a_12002_2130# a_12306_2170# 0.0931f
C11504 a_12914_2130# a_13406_2492# 0.0658f
C11505 m2_24248_1374# VDD 0.0194f
C11506 row_n[9] a_3270_11206# 0.0117f
C11507 vcm col_n[27] 1.94f
C11508 col_n[13] col_n[14] 0.0101f
C11509 VDD col_n[30] 5.18f
C11510 vcm a_35002_4138# 0.101f
C11511 col[14] rowoff_n[15] 0.0901f
C11512 rowon_n[1] a_25966_3134# 0.118f
C11513 col[23] col[24] 0.0355f
C11514 a_24050_7150# a_25054_7150# 0.843f
C11515 col[7] a_2475_10186# 0.136f
C11516 rowoff_n[9] a_28466_11528# 0.0133f
C11517 col_n[0] a_3366_6508# 0.0283f
C11518 vcm a_22346_13214# 0.155f
C11519 a_2475_11190# a_1957_11190# 0.0734f
C11520 VDD a_20434_3496# 0.0779f
C11521 VDD rowoff_n[11] 1.51f
C11522 m2_11772_18014# a_11910_18194# 0.225f
C11523 col[5] a_7986_16186# 0.367f
C11524 col[2] a_4882_6146# 0.0682f
C11525 a_2475_16210# a_25966_16186# 0.264f
C11526 a_13918_16186# a_14010_16186# 0.326f
C11527 a_2275_16210# a_23350_16226# 0.144f
C11528 VDD a_9902_12170# 0.181f
C11529 col[12] a_14922_18194# 0.0682f
C11530 col_n[14] a_2275_16210# 0.113f
C11531 col_n[19] a_2275_5166# 0.113f
C11532 col_n[20] a_23046_12170# 0.251f
C11533 col_n[17] a_19942_2130# 0.0765f
C11534 vcm a_15926_7150# 0.1f
C11535 rowon_n[5] a_2874_7150# 0.118f
C11536 rowoff_n[12] a_9994_14178# 0.294f
C11537 a_15014_9158# a_15014_8154# 0.843f
C11538 col_n[27] a_29982_14178# 0.0765f
C11539 m2_26256_14426# a_26058_14178# 0.165f
C11540 vcm a_3270_16226# 0.155f
C11541 a_2275_13198# a_16930_13174# 0.136f
C11542 a_8898_13174# a_9294_13214# 0.0313f
C11543 VDD a_35494_7512# 0.106f
C11544 m2_1732_6970# ctop 0.0428f
C11545 col[4] a_2275_13198# 0.0899f
C11546 ctop a_16018_11166# 4.11f
C11547 col[9] a_2275_2154# 0.0899f
C11548 VDD a_24962_16186# 0.181f
C11549 m2_9764_946# col_n[7] 0.331f
C11550 col_n[11] a_14410_10524# 0.0283f
C11551 a_27974_6146# a_28466_6508# 0.0658f
C11552 a_27062_6146# a_27366_6186# 0.0931f
C11553 m2_3164_11414# rowon_n[9] 0.0322f
C11554 m2_9188_7398# rowon_n[5] 0.0322f
C11555 m2_30848_946# m2_31852_946# 0.843f
C11556 m2_15212_3382# rowon_n[1] 0.0322f
C11557 col[24] a_2475_12194# 0.136f
C11558 vcm a_30986_11166# 0.1f
C11559 a_4974_10162# a_5978_10162# 0.843f
C11560 a_2475_10186# a_8990_10162# 0.316f
C11561 col[29] a_2475_1150# 0.136f
C11562 row_n[14] a_14010_16186# 0.282f
C11563 a_2275_15206# a_31990_15182# 0.136f
C11564 VDD a_16418_10524# 0.0779f
C11565 sample a_2161_16210# 0.0858f
C11566 rowoff_n[0] m2_34864_1950# 0.278f
C11567 ctop a_31078_15182# 4.11f
C11568 m3_34996_13126# a_34090_13174# 0.0303f
C11569 row_n[4] a_24050_6146# 0.282f
C11570 col_n[31] a_2275_18218# 0.113f
C11571 rowon_n[8] a_23958_10162# 0.118f
C11572 a_23958_3134# a_24050_3134# 0.326f
C11573 rowoff_n[10] a_16418_12532# 0.0133f
C11574 col_n[9] a_12002_10162# 0.251f
C11575 m2_2736_18014# vcm 0.353f
C11576 m2_24248_16434# rowon_n[14] 0.0322f
C11577 m2_17220_12418# a_17022_12170# 0.165f
C11578 m2_30272_12418# rowon_n[10] 0.0322f
C11579 row_n[6] a_11302_8194# 0.0117f
C11580 m2_35292_8402# rowon_n[6] 0.0322f
C11581 vcm a_11910_14178# 0.1f
C11582 a_30074_13174# a_30074_12170# 0.843f
C11583 a_2475_12194# a_24050_12170# 0.316f
C11584 VDD a_7986_4138# 0.483f
C11585 col_n[16] a_18938_12170# 0.0765f
C11586 col[21] a_2275_15206# 0.0899f
C11587 a_23958_17190# a_24354_17230# 0.0313f
C11588 VDD a_31478_14540# 0.0779f
C11589 col[26] a_2275_4162# 0.0899f
C11590 rowoff_n[0] a_8386_2492# 0.0133f
C11591 vcm a_2966_8154# 0.56f
C11592 a_2275_9182# a_15014_9158# 0.399f
C11593 rowoff_n[14] a_32482_16548# 0.0133f
C11594 a_8898_9158# a_9390_9520# 0.0658f
C11595 a_7986_9158# a_8290_9198# 0.0931f
C11596 rowon_n[2] a_10998_4138# 0.248f
C11597 col_n[31] rowoff_n[0] 0.0471f
C11598 a_27462_1488# col_n[24] 0.0283f
C11599 vcm a_26970_18194# 0.101f
C11600 a_20034_14178# a_21038_14178# 0.843f
C11601 col[29] a_32082_9158# 0.367f
C11602 VDD a_23046_8154# 0.483f
C11603 col_n[17] a_2475_18218# 0.0529f
C11604 VDD a_12402_17552# 0.0779f
C11605 m3_25960_1078# VDD 0.0157f
C11606 col_n[11] a_2475_11190# 0.0531f
C11607 vcm a_29070_3134# 0.56f
C11608 a_2275_6170# a_5278_6186# 0.144f
C11609 a_2475_6170# a_7894_6146# 0.264f
C11610 a_3878_6146# a_4274_6186# 0.0313f
C11611 a_4882_6146# a_4974_6146# 0.326f
C11612 m2_8184_10410# a_7986_10162# 0.165f
C11613 rowoff_n[3] a_8990_5142# 0.294f
C11614 a_2275_11190# a_30074_11166# 0.399f
C11615 col_n[24] a_27366_9198# 0.084f
C11616 m2_30848_18014# a_30986_18194# 0.225f
C11617 m2_7756_18014# a_7986_17190# 0.843f
C11618 row_n[11] a_22042_13174# 0.282f
C11619 a_10998_16186# a_10998_15182# 0.843f
C11620 VDD a_3970_11166# 0.483f
C11621 m2_30848_18014# m3_29976_18146# 0.0341f
C11622 col_n[5] a_7894_10162# 0.0765f
C11623 rowon_n[15] a_21950_17190# 0.118f
C11624 col[1] a_2475_8178# 0.136f
C11625 rowoff_n[1] a_18026_3134# 0.294f
C11626 row_n[1] a_32082_3134# 0.282f
C11627 m2_27260_6394# a_27062_6146# 0.165f
C11628 row_n[13] a_9294_15222# 0.0117f
C11629 vcm a_9994_6146# 0.56f
C11630 rowon_n[5] a_31990_7150# 0.118f
C11631 a_2475_8178# a_22954_8154# 0.264f
C11632 a_2275_8178# a_20338_8194# 0.144f
C11633 rowoff_n[11] a_4370_13536# 0.0133f
C11634 col_n[24] rowoff_n[10] 0.0471f
C11635 col_n[8] a_2275_14202# 0.113f
C11636 a_23958_13174# a_24450_13536# 0.0658f
C11637 a_23046_13174# a_23350_13214# 0.0931f
C11638 row_n[3] a_19334_5182# 0.0117f
C11639 col_n[13] a_2275_3158# 0.113f
C11640 VDD a_19030_15182# 0.483f
C11641 m2_2160_10410# row_n[8] 0.0194f
C11642 col[18] a_21038_7150# 0.367f
C11643 m2_8184_6394# row_n[4] 0.0128f
C11644 m2_13204_2378# row_n[0] 0.0128f
C11645 col[25] a_27974_9158# 0.0682f
C11646 row_n[5] a_9902_7150# 0.0437f
C11647 a_2275_5166# a_13918_5142# 0.136f
C11648 col_n[28] a_2475_13198# 0.0531f
C11649 m2_1732_4962# sample_n 0.0522f
C11650 m2_33860_946# m3_34568_1078# 1.07f
C11651 m3_34996_11118# m3_34996_10114# 0.202f
C11652 col_n[0] a_3270_3174# 0.084f
C11653 rowon_n[9] a_8990_11166# 0.248f
C11654 vcm a_25054_10162# 0.56f
C11655 rowoff_n[15] a_20434_17552# 0.0133f
C11656 a_19942_10162# a_20034_10162# 0.326f
C11657 a_2275_10186# a_2275_9182# 0.0715f
C11658 m2_30848_18014# ctop 0.0422f
C11659 col_n[13] a_16322_7190# 0.084f
C11660 col_n[1] row_n[13] 0.298f
C11661 col_n[5] row_n[15] 0.298f
C11662 VDD row_n[11] 3.29f
C11663 col_n[4] rowon_n[14] 0.111f
C11664 col_n[6] rowon_n[15] 0.111f
C11665 col_n[3] row_n[14] 0.298f
C11666 col_n[2] rowon_n[13] 0.111f
C11667 col_n[0] row_n[12] 0.298f
C11668 vcm rowon_n[12] 0.65f
C11669 sample rowon_n[11] 0.0935f
C11670 col[18] a_2475_10186# 0.136f
C11671 col[25] rowoff_n[15] 0.0901f
C11672 a_2475_2154# a_5978_2130# 0.316f
C11673 a_3878_2130# a_4370_2492# 0.0658f
C11674 m2_23244_15430# row_n[13] 0.0128f
C11675 a_21038_3134# a_21038_2130# 0.843f
C11676 m2_29268_11414# row_n[9] 0.0128f
C11677 m2_18224_4386# a_18026_4138# 0.165f
C11678 m2_34864_6970# row_n[5] 0.267f
C11679 vcm a_15318_4178# 0.155f
C11680 rowoff_n[9] a_10906_11166# 0.202f
C11681 a_2275_7174# a_28978_7150# 0.136f
C11682 col_n[8] rowoff_n[11] 0.0471f
C11683 a_14922_7150# a_15318_7190# 0.0313f
C11684 vcm a_5978_13174# 0.56f
C11685 VDD a_2161_3158# 0.187f
C11686 col_n[25] a_2275_16210# 0.113f
C11687 a_2275_16210# a_6982_16186# 0.399f
C11688 a_3970_16186# a_4274_16226# 0.0931f
C11689 a_4882_16186# a_5374_16548# 0.0658f
C11690 col_n[30] a_2275_5166# 0.113f
C11691 row_n[8] a_30074_10162# 0.282f
C11692 rowoff_n[7] a_19942_9158# 0.202f
C11693 rowon_n[12] a_29982_14178# 0.118f
C11694 a_2475_4162# a_21038_4138# 0.316f
C11695 a_10998_4138# a_12002_4138# 0.843f
C11696 col[7] a_9994_5142# 0.367f
C11697 m3_2868_1078# ctop 0.0674f
C11698 col[17] a_20034_17190# 0.367f
C11699 vcm a_30378_8194# 0.155f
C11700 col[14] a_16930_7150# 0.0682f
C11701 rowoff_n[13] a_26970_15182# 0.202f
C11702 col[15] a_2275_13198# 0.0899f
C11703 row_n[10] a_17326_12210# 0.0117f
C11704 ctop a_8990_2130# 4.06f
C11705 col[20] a_2275_2154# 0.0899f
C11706 vcm a_21038_17190# 0.56f
C11707 a_35002_14178# a_35094_14178# 0.0991f
C11708 a_34090_14178# a_34394_14218# 0.0931f
C11709 VDD a_17934_7150# 0.181f
C11710 rowoff_n[5] a_28978_7150# 0.202f
C11711 col_n[29] a_31990_3134# 0.0765f
C11712 a_2275_18218# a_22042_18194# 0.0924f
C11713 row_n[0] a_27366_2170# 0.0117f
C11714 row_n[12] a_7894_14178# 0.0437f
C11715 a_2275_1150# a_12002_1126# 0.0924f
C11716 col_n[2] a_5278_5182# 0.084f
C11717 vcm a_23958_2130# 0.1f
C11718 col_n[12] a_15318_17230# 0.084f
C11719 a_2475_6170# a_2475_5166# 0.0666f
C11720 m2_11772_946# m2_12200_1374# 0.165f
C11721 vcm a_11302_11206# 0.155f
C11722 row_n[2] a_17934_4138# 0.0437f
C11723 a_29982_11166# a_30378_11206# 0.0313f
C11724 VDD a_9390_1488# 0.0977f
C11725 rowon_n[6] a_17022_8154# 0.248f
C11726 m2_26832_18014# a_27062_17190# 0.843f
C11727 ctop a_24050_6146# 4.11f
C11728 a_2475_15206# a_14922_15182# 0.264f
C11729 a_2275_15206# a_12306_15222# 0.144f
C11730 VDD a_32994_11166# 0.181f
C11731 col_n[23] a_26458_11528# 0.0283f
C11732 col_n[5] a_2475_9182# 0.0531f
C11733 a_14010_3134# a_14314_3174# 0.0931f
C11734 a_14922_3134# a_15414_3496# 0.0658f
C11735 a_2275_3158# a_27062_3134# 0.399f
C11736 a_2475_18218# a_20034_18194# 0.0299f
C11737 rowoff_n[8] a_29470_10524# 0.0133f
C11738 vcm a_4882_5142# 0.1f
C11739 a_26058_8154# a_27062_8154# 0.843f
C11740 m2_1732_11990# a_2966_12170# 0.843f
C11741 col[6] a_8990_15182# 0.367f
C11742 vcm a_26362_15222# 0.155f
C11743 a_2275_12194# a_5886_12170# 0.136f
C11744 col[3] a_5886_5142# 0.0682f
C11745 VDD a_24450_5504# 0.0779f
C11746 m2_6752_18014# VDD 1.1f
C11747 ctop a_4974_9158# 4.11f
C11748 col[13] a_15926_17190# 0.0682f
C11749 row_n[15] a_28066_17190# 0.282f
C11750 a_2275_17214# a_27366_17230# 0.144f
C11751 a_15926_17190# a_16018_17190# 0.326f
C11752 a_2475_17214# a_29982_17190# 0.264f
C11753 VDD a_13918_14178# 0.181f
C11754 col_n[21] a_24050_11166# 0.251f
C11755 m3_33992_18146# a_34090_17190# 0.0303f
C11756 rowon_n[0] a_4882_2130# 0.118f
C11757 col_n[18] a_20946_1126# 0.0765f
C11758 col_n[28] a_30986_13174# 0.0765f
C11759 col_n[2] a_2275_12194# 0.113f
C11760 row_n[7] rowoff_n[7] 0.209f
C11761 vcm a_19942_9158# 0.1f
C11762 col_n[7] a_2275_1150# 0.113f
C11763 m2_2736_18014# m2_3164_18442# 0.165f
C11764 col_n[1] a_4274_15222# 0.084f
C11765 rowoff_n[14] a_14922_16186# 0.202f
C11766 a_17022_10162# a_17022_9158# 0.843f
C11767 sample a_1957_5166# 0.345f
C11768 m2_34864_15002# a_2275_15206# 0.278f
C11769 col_n[28] a_2475_18218# 0.0529f
C11770 vcm a_7286_18234# 0.16f
C11771 a_2275_14202# a_20946_14178# 0.136f
C11772 a_10906_14178# a_11302_14218# 0.0313f
C11773 row_n[7] a_25358_9198# 0.0117f
C11774 VDD a_5374_8516# 0.0779f
C11775 m2_4744_946# vcm 0.353f
C11776 ctop a_20034_13174# 4.11f
C11777 col_n[22] a_2475_11190# 0.0531f
C11778 VDD a_28978_18194# 0.343f
C11779 col_n[12] a_15414_9520# 0.0283f
C11780 a_2275_2154# a_32386_2170# 0.144f
C11781 a_2475_2154# a_35002_2130# 0.264f
C11782 m3_21944_18146# VDD 0.0313f
C11783 row_n[9] a_15926_11166# 0.0437f
C11784 a_29070_7150# a_29374_7190# 0.0931f
C11785 a_29982_7150# a_30474_7512# 0.0658f
C11786 rowon_n[13] a_15014_15182# 0.248f
C11787 vcm a_35002_13174# 0.101f
C11788 a_6982_11166# a_7986_11166# 0.843f
C11789 a_2475_11190# a_13006_11166# 0.316f
C11790 VDD a_31078_3134# 0.483f
C11791 col[12] a_2475_8178# 0.136f
C11792 col_n[0] a_3366_15544# 0.0283f
C11793 a_2275_16210# a_34394_16226# 0.144f
C11794 rowon_n[3] a_25054_5142# 0.248f
C11795 VDD a_20434_12532# 0.0779f
C11796 m2_6752_18014# m3_6884_18146# 3.79f
C11797 rowon_n[15] a_3878_17190# 0.118f
C11798 m2_13204_14426# rowon_n[12] 0.0322f
C11799 m2_19228_10410# rowon_n[8] 0.0322f
C11800 col[2] a_4882_15182# 0.0682f
C11801 m2_25252_6394# rowon_n[4] 0.0322f
C11802 a_25966_4138# a_26058_4138# 0.326f
C11803 col_n[10] a_13006_9158# 0.251f
C11804 col_n[19] a_2275_14202# 0.113f
C11805 a_2275_8178# a_3970_8154# 0.399f
C11806 col_n[24] a_2275_3158# 0.113f
C11807 m2_34864_13998# a_35002_14178# 0.225f
C11808 col_n[17] a_19942_11166# 0.0765f
C11809 vcm a_15926_16186# 0.1f
C11810 a_32082_14178# a_32082_13174# 0.843f
C11811 a_2475_13198# a_28066_13174# 0.316f
C11812 VDD a_12002_6146# 0.483f
C11813 row_n[3] a_2874_5142# 0.0436f
C11814 rowon_n[7] a_2161_9182# 0.0177f
C11815 a_25966_18194# a_26362_18234# 0.0313f
C11816 VDD a_35494_16548# 0.106f
C11817 a_20946_1126# a_21342_1166# 0.0313f
C11818 col[9] a_2275_11190# 0.0899f
C11819 vcm a_18026_1126# 0.557f
C11820 col_n[1] a_4370_7512# 0.0283f
C11821 m3_13912_18146# m3_14916_18146# 0.202f
C11822 m2_9764_946# m3_8892_1078# 0.0341f
C11823 a_2275_10186# a_19030_10162# 0.399f
C11824 rowoff_n[15] a_2161_17214# 0.0226f
C11825 a_9994_10162# a_10298_10202# 0.0931f
C11826 a_10906_10162# a_11398_10524# 0.0658f
C11827 row_n[14] a_23350_16226# 0.0117f
C11828 col[30] a_33086_8154# 0.367f
C11829 m2_1732_1950# VDD 0.856f
C11830 col_n[1] rowon_n[7] 0.111f
C11831 vcm row_n[7] 0.616f
C11832 col_n[6] row_n[10] 0.298f
C11833 col_n[0] rowon_n[6] 0.111f
C11834 col_n[24] col_n[25] 0.0103f
C11835 col_n[14] row_n[14] 0.298f
C11836 col_n[13] rowon_n[13] 0.111f
C11837 col_n[17] rowon_n[15] 0.111f
C11838 col_n[11] rowon_n[12] 0.111f
C11839 col_n[2] row_n[8] 0.298f
C11840 col_n[8] row_n[11] 0.298f
C11841 sample row_n[6] 0.423f
C11842 col_n[10] row_n[12] 0.298f
C11843 col_n[7] rowon_n[10] 0.111f
C11844 col_n[3] rowon_n[8] 0.111f
C11845 col_n[5] rowon_n[9] 0.111f
C11846 col_n[15] rowon_n[14] 0.111f
C11847 VDD rowon_n[5] 3.04f
C11848 col_n[12] row_n[13] 0.298f
C11849 col_n[4] row_n[9] 0.298f
C11850 a_22042_15182# a_23046_15182# 0.843f
C11851 col_n[16] row_n[15] 0.298f
C11852 col_n[9] rowon_n[11] 0.111f
C11853 col[29] a_2475_10186# 0.136f
C11854 VDD a_27062_10162# 0.483f
C11855 row_n[4] a_33390_6186# 0.0117f
C11856 col_n[19] rowoff_n[11] 0.0471f
C11857 vcm a_33086_5142# 0.56f
C11858 rowoff_n[2] a_9994_4138# 0.294f
C11859 rowoff_n[10] a_27062_12170# 0.294f
C11860 a_2275_7174# a_9294_7190# 0.144f
C11861 a_6890_7150# a_6982_7150# 0.326f
C11862 a_2475_7174# a_11910_7150# 0.264f
C11863 row_n[6] a_23958_8154# 0.0437f
C11864 col_n[0] a_2475_7174# 0.0532f
C11865 col_n[25] a_28370_8194# 0.084f
C11866 a_2275_12194# a_34090_12170# 0.399f
C11867 rowon_n[10] a_23046_12170# 0.248f
C11868 col_n[6] a_8898_9158# 0.0765f
C11869 a_13006_17190# a_13006_16186# 0.843f
C11870 VDD a_7986_13174# 0.483f
C11871 rowoff_n[0] a_19030_2130# 0.294f
C11872 rowon_n[0] a_33086_2130# 0.248f
C11873 col[26] a_2275_13198# 0.0899f
C11874 a_2475_4162# a_2966_4138# 0.317f
C11875 a_2161_4162# a_2275_4162# 0.183f
C11876 col[31] a_2275_2154# 0.0899f
C11877 m2_17796_18014# col[15] 0.347f
C11878 vcm a_14010_8154# 0.56f
C11879 a_2275_9182# a_24354_9198# 0.144f
C11880 a_2475_9182# a_26970_9158# 0.264f
C11881 m2_32280_15430# a_32082_15182# 0.165f
C11882 vcm a_2966_17190# 0.56f
C11883 a_25054_14178# a_25358_14218# 0.0931f
C11884 a_25966_14178# a_26458_14540# 0.0658f
C11885 col[19] a_22042_6146# 0.367f
C11886 col_n[3] rowoff_n[12] 0.0471f
C11887 VDD a_23046_17190# 0.484f
C11888 row_n[0] a_10998_2130# 0.282f
C11889 a_32082_2130# a_33086_2130# 0.843f
C11890 col[26] a_28978_8154# 0.0682f
C11891 rowon_n[4] a_10906_6146# 0.118f
C11892 vcm a_4274_2170# 0.155f
C11893 a_2275_6170# a_17934_6146# 0.136f
C11894 vcm a_29070_12170# 0.56f
C11895 a_21950_11166# a_22042_11166# 0.326f
C11896 m2_6176_17438# row_n[15] 0.0128f
C11897 VDD a_25966_2130# 0.181f
C11898 col_n[16] a_2475_9182# 0.0531f
C11899 m2_12200_13422# row_n[11] 0.0128f
C11900 m2_4168_17438# a_3970_17190# 0.165f
C11901 m2_18224_9406# row_n[7] 0.0128f
C11902 col_n[14] a_17326_6186# 0.084f
C11903 m2_24248_5390# row_n[3] 0.0128f
C11904 row_n[11] a_31382_13214# 0.0117f
C11905 col_n[24] a_27366_18234# 0.084f
C11906 a_23046_4138# a_23046_3134# 0.843f
C11907 a_2475_3158# a_9994_3134# 0.316f
C11908 a_2475_18218# a_1957_18218# 0.0734f
C11909 col[1] a_2475_17214# 0.136f
C11910 rowoff_n[8] a_11910_10162# 0.202f
C11911 m2_34864_5966# a_35398_6186# 0.087f
C11912 row_n[13] a_21950_15182# 0.0437f
C11913 col[6] a_2475_6170# 0.136f
C11914 vcm a_19334_6186# 0.155f
C11915 a_2275_8178# a_32994_8154# 0.136f
C11916 rowoff_n[11] a_15014_13174# 0.294f
C11917 a_16930_8154# a_17326_8194# 0.0313f
C11918 m2_23244_13422# a_23046_13174# 0.165f
C11919 vcm a_9994_15182# 0.56f
C11920 VDD a_6890_5142# 0.181f
C11921 row_n[3] a_31990_5142# 0.0437f
C11922 m2_33860_18014# col_n[31] 0.243f
C11923 rowon_n[7] a_31078_9158# 0.248f
C11924 a_5978_17190# a_6282_17230# 0.0931f
C11925 a_6890_17190# a_7382_17552# 0.0658f
C11926 a_2275_17214# a_10998_17190# 0.399f
C11927 rowoff_n[6] a_20946_8154# 0.202f
C11928 col_n[13] a_2275_12194# 0.113f
C11929 col[8] a_10998_4138# 0.367f
C11930 rowon_n[3] rowoff_n[3] 20.2f
C11931 col_n[18] a_2275_1150# 0.113f
C11932 col[18] a_21038_16186# 0.367f
C11933 a_2475_5166# a_25054_5142# 0.316f
C11934 a_13006_5142# a_14010_5142# 0.843f
C11935 col[15] a_17934_6146# 0.0682f
C11936 m3_3872_1078# m3_4876_1078# 0.202f
C11937 vcm a_35398_10202# 0.161f
C11938 col[25] a_27974_18194# 0.0682f
C11939 rowoff_n[15] a_31078_17190# 0.294f
C11940 rowoff_n[4] a_29982_6146# 0.202f
C11941 col_n[0] a_3270_12210# 0.084f
C11942 ctop a_13006_4138# 4.11f
C11943 m2_6752_946# a_6890_1126# 0.225f
C11944 m2_15788_946# a_2475_1150# 0.286f
C11945 col_n[30] a_32994_2130# 0.0765f
C11946 VDD a_21950_9158# 0.181f
C11947 col[3] a_2275_9182# 0.0899f
C11948 row_n[7] a_8990_9158# 0.282f
C11949 rowon_n[11] a_8898_13174# 0.118f
C11950 col_n[3] a_6282_4178# 0.084f
C11951 VDD a_9294_18234# 0.019f
C11952 col_n[13] a_16322_16226# 0.084f
C11953 a_2275_2154# a_16018_2130# 0.399f
C11954 m2_8760_946# VDD 1f
C11955 vcm a_27974_4138# 0.1f
C11956 a_3970_7150# a_3970_6146# 0.843f
C11957 rowoff_n[9] a_21438_11528# 0.0133f
C11958 rowon_n[1] a_18938_3134# 0.118f
C11959 col[23] a_2475_8178# 0.136f
C11960 m2_14208_11414# a_14010_11166# 0.165f
C11961 vcm a_15318_13214# 0.155f
C11962 a_31990_12170# a_32386_12210# 0.0313f
C11963 VDD a_13406_3496# 0.0779f
C11964 col_n[24] a_27462_10524# 0.0283f
C11965 m2_6752_18014# a_6982_18194# 0.0249f
C11966 ctop a_28066_8154# 4.11f
C11967 a_2275_16210# a_16322_16226# 0.144f
C11968 a_2475_16210# a_18938_16186# 0.264f
C11969 VDD a_2161_12194# 0.187f
C11970 a_25358_1166# m2_24824_946# 0.087f
C11971 rowoff_n[7] a_30474_9520# 0.0133f
C11972 col_n[30] a_2275_14202# 0.113f
C11973 a_2275_4162# a_31078_4138# 0.399f
C11974 a_16018_4138# a_16322_4178# 0.0931f
C11975 a_16930_4138# a_17422_4500# 0.0658f
C11976 m2_33284_7398# a_33086_7150# 0.165f
C11977 vcm a_8898_7150# 0.1f
C11978 rowoff_n[12] a_2874_14178# 0.202f
C11979 col[7] a_9994_14178# 0.367f
C11980 a_28066_9158# a_29070_9158# 0.843f
C11981 col[4] a_6890_4138# 0.0682f
C11982 row_n[10] a_29982_12170# 0.0437f
C11983 vcm a_30378_17230# 0.155f
C11984 a_2275_13198# a_9902_13174# 0.136f
C11985 rowon_n[14] a_29070_16186# 0.248f
C11986 col[14] a_16930_16186# 0.0682f
C11987 VDD a_28466_7512# 0.0779f
C11988 ctop a_8990_11166# 4.11f
C11989 col[20] a_2275_11190# 0.0899f
C11990 col_n[22] a_25054_10162# 0.251f
C11991 a_2275_18218# a_31382_18234# 0.145f
C11992 a_17934_18194# a_18026_18194# 0.0991f
C11993 VDD a_17934_16186# 0.181f
C11994 a_12914_1126# a_13006_1126# 0.0991f
C11995 a_2275_1150# a_21342_1166# 0.145f
C11996 a_2475_1150# a_23958_1126# 0.264f
C11997 col_n[29] a_31990_12170# 0.0765f
C11998 col_n[2] a_5278_14218# 0.084f
C11999 m2_23820_946# m2_24824_946# 0.843f
C12000 m2_5172_9406# a_4974_9158# 0.165f
C12001 col_n[0] a_2966_4138# 0.251f
C12002 vcm rowon_n[1] 0.65f
C12003 col_n[10] rowon_n[6] 0.111f
C12004 col_n[26] rowon_n[14] 0.111f
C12005 col_n[5] row_n[4] 0.298f
C12006 col_n[24] rowon_n[13] 0.111f
C12007 col_n[0] row_n[1] 0.298f
C12008 vcm a_23958_11166# 0.1f
C12009 col_n[1] row_n[2] 0.298f
C12010 col_n[13] row_n[8] 0.298f
C12011 col_n[4] rowon_n[3] 0.111f
C12012 col_n[15] row_n[9] 0.298f
C12013 col_n[16] rowon_n[9] 0.111f
C12014 col_n[14] rowon_n[8] 0.111f
C12015 col_n[17] row_n[10] 0.298f
C12016 col_n[23] row_n[13] 0.298f
C12017 sample rowon_n[0] 0.0935f
C12018 col_n[21] row_n[12] 0.298f
C12019 col_n[18] rowon_n[10] 0.111f
C12020 col_n[22] rowon_n[12] 0.111f
C12021 col_n[27] row_n[15] 0.298f
C12022 col_n[3] row_n[3] 0.298f
C12023 col_n[6] rowon_n[4] 0.111f
C12024 col_n[8] rowon_n[5] 0.111f
C12025 col_n[2] rowon_n[2] 0.111f
C12026 col_n[9] row_n[6] 0.298f
C12027 col_n[7] row_n[5] 0.298f
C12028 col_n[11] row_n[7] 0.298f
C12029 VDD row_n[0] 3.3f
C12030 col_n[28] rowon_n[15] 0.111f
C12031 col_n[12] rowon_n[7] 0.111f
C12032 col_n[25] row_n[14] 0.298f
C12033 col_n[20] rowon_n[11] 0.111f
C12034 col_n[19] row_n[11] 0.298f
C12035 a_19030_11166# a_19030_10162# 0.843f
C12036 VDD a_20034_1126# 0.994f
C12037 row_n[14] a_6982_16186# 0.282f
C12038 a_2275_15206# a_24962_15182# 0.136f
C12039 a_12914_15182# a_13310_15222# 0.0313f
C12040 col_n[30] rowoff_n[11] 0.0471f
C12041 VDD a_9390_10524# 0.0779f
C12042 col_n[13] a_16418_8516# 0.0283f
C12043 ctop a_24050_15182# 4.11f
C12044 row_n[4] a_17022_6146# 0.282f
C12045 rowon_n[8] a_16930_10162# 0.118f
C12046 m2_24248_5390# a_24050_5142# 0.165f
C12047 col_n[10] a_2475_7174# 0.0531f
C12048 m2_1732_11990# m2_1732_10986# 0.843f
C12049 a_31990_8154# a_32482_8516# 0.0658f
C12050 rowoff_n[10] a_9390_12532# 0.0133f
C12051 a_31078_8154# a_31382_8194# 0.0931f
C12052 a_27366_1166# vcm 0.16f
C12053 m2_2160_12418# rowon_n[10] 0.0219f
C12054 row_n[6] a_4274_8194# 0.0117f
C12055 m2_8184_8402# rowon_n[6] 0.0322f
C12056 vcm a_4882_14178# 0.1f
C12057 m2_14208_4386# rowon_n[2] 0.0322f
C12058 a_8990_12170# a_9994_12170# 0.843f
C12059 a_2475_12194# a_17022_12170# 0.316f
C12060 m2_28264_18442# VDD 0.0456f
C12061 VDD a_24450_14540# 0.0779f
C12062 col[3] a_5886_14178# 0.0682f
C12063 a_3970_1126# m2_2736_946# 0.843f
C12064 col[0] a_2475_4162# 0.148f
C12065 col_n[11] a_14010_8154# 0.251f
C12066 a_27974_5142# a_28066_5142# 0.326f
C12067 col_n[18] a_20946_10162# 0.0765f
C12068 a_2275_9182# a_7986_9158# 0.399f
C12069 rowoff_n[14] a_25454_16548# 0.0133f
C12070 rowon_n[2] a_3970_4138# 0.248f
C12071 col_n[14] rowoff_n[12] 0.0471f
C12072 vcm a_19942_18194# 0.101f
C12073 col_n[7] a_2275_10186# 0.113f
C12074 m2_23244_17438# rowon_n[15] 0.0322f
C12075 a_34090_15182# a_34090_14178# 0.843f
C12076 m3_3872_1078# a_3970_1126# 3.24f
C12077 a_2475_14202# a_32082_14178# 0.316f
C12078 VDD a_16018_8154# 0.483f
C12079 m2_29268_13422# rowon_n[11] 0.0322f
C12080 m2_34864_8978# rowon_n[7] 0.231f
C12081 sample a_1957_14202# 0.345f
C12082 col[0] m2_1732_946# 0.0137f
C12083 m2_27836_946# vcm 0.353f
C12084 VDD a_5374_17552# 0.0779f
C12085 a_22954_2130# a_23350_2170# 0.0313f
C12086 col_n[2] a_5374_6508# 0.0283f
C12087 m2_15212_3382# a_15014_3134# 0.165f
C12088 vcm a_22042_3134# 0.56f
C12089 col_n[12] a_15414_18556# 0.0283f
C12090 col_n[27] a_2475_9182# 0.0531f
C12091 m2_1732_9982# a_2275_10186# 0.191f
C12092 col[31] a_34090_7150# 0.367f
C12093 rowoff_n[3] a_2475_5166# 3.9f
C12094 a_2275_11190# a_23046_11166# 0.399f
C12095 a_12002_11166# a_12306_11206# 0.0931f
C12096 a_12914_11166# a_13406_11528# 0.0658f
C12097 m2_25828_18014# a_26058_18194# 0.0249f
C12098 row_n[11] a_15014_13174# 0.282f
C12099 a_24050_16186# a_25054_16186# 0.843f
C12100 VDD a_31078_12170# 0.483f
C12101 m2_20808_18014# m3_21944_18146# 0.0341f
C12102 col[12] a_2475_17214# 0.136f
C12103 rowon_n[15] a_14922_17190# 0.118f
C12104 m2_1732_8978# col[0] 0.0137f
C12105 col[17] a_2475_6170# 0.136f
C12106 rowoff_n[1] a_10998_3134# 0.294f
C12107 row_n[1] a_25054_3134# 0.282f
C12108 row_n[13] a_3878_15182# 0.0437f
C12109 col_n[26] a_29374_7190# 0.084f
C12110 rowon_n[5] a_24962_7150# 0.118f
C12111 vcm a_2874_6146# 0.1f
C12112 rowoff_n[12] a_31990_14178# 0.202f
C12113 a_2475_8178# a_15926_8154# 0.264f
C12114 a_8898_8154# a_8990_8154# 0.326f
C12115 a_2275_8178# a_13310_8194# 0.144f
C12116 sample rowoff_n[13] 0.0775f
C12117 col_n[7] a_9902_8154# 0.0765f
C12118 row_n[3] a_12306_5182# 0.0117f
C12119 col_n[24] a_2275_12194# 0.113f
C12120 ctop rowoff_n[2] 0.177f
C12121 col[1] rowoff_n[9] 0.0901f
C12122 col[0] rowoff_n[8] 0.0901f
C12123 col_n[29] a_2275_1150# 0.113f
C12124 VDD a_12002_15182# 0.483f
C12125 rowoff_n[6] a_2275_8178# 0.151f
C12126 a_2275_5166# a_6890_5142# 0.136f
C12127 row_n[5] a_2161_7174# 0.0221f
C12128 m2_1732_2954# vcm 0.316f
C12129 m3_34996_18146# m3_34996_17142# 0.202f
C12130 m2_24824_946# m3_24956_1078# 3.79f
C12131 rowon_n[9] a_2475_11190# 0.31f
C12132 vcm a_18026_10162# 0.56f
C12133 col[14] a_2275_9182# 0.0899f
C12134 a_2475_10186# a_30986_10162# 0.264f
C12135 a_2275_10186# a_28370_10202# 0.144f
C12136 col_n[1] a_4370_16548# 0.0283f
C12137 rowoff_n[15] a_13406_17552# 0.0133f
C12138 row_n[14] a_34394_16226# 0.0117f
C12139 col[20] a_23046_5142# 0.367f
C12140 a_27974_15182# a_28466_15544# 0.0658f
C12141 a_27062_15182# a_27366_15222# 0.0931f
C12142 m2_16792_18014# ctop 0.0422f
C12143 VDD a_3878_9158# 0.181f
C12144 col[30] a_33086_17190# 0.367f
C12145 col[27] a_29982_7150# 0.0682f
C12146 a_33998_3134# a_34394_3174# 0.0313f
C12147 m2_1732_10986# row_n[9] 0.292f
C12148 m2_7180_7398# row_n[5] 0.0128f
C12149 m2_13204_3382# row_n[1] 0.0128f
C12150 vcm a_8290_4178# 0.155f
C12151 rowoff_n[9] a_3366_11528# 0.0133f
C12152 a_2275_7174# a_21950_7150# 0.136f
C12153 m2_34864_11990# a_34090_12170# 0.843f
C12154 vcm a_33086_14178# 0.56f
C12155 a_23958_12170# a_24050_12170# 0.326f
C12156 col_n[15] a_18330_5182# 0.084f
C12157 VDD a_29982_4138# 0.181f
C12158 col_n[0] a_2475_16210# 0.0532f
C12159 col_n[25] a_28370_17230# 0.084f
C12160 col_n[4] a_2475_5166# 0.0531f
C12161 col_n[6] a_8898_18194# 0.0762f
C12162 row_n[8] a_23046_10162# 0.282f
C12163 rowoff_n[7] a_12914_9158# 0.202f
C12164 rowon_n[12] a_22954_14178# 0.118f
C12165 a_2475_4162# a_14010_4138# 0.316f
C12166 a_25054_5142# a_25054_4138# 0.843f
C12167 m3_1864_14130# ctop 0.21f
C12168 m2_22240_16434# row_n[14] 0.0128f
C12169 vcm a_23350_8194# 0.155f
C12170 m2_28264_12418# row_n[10] 0.0128f
C12171 a_18938_9158# a_19334_9198# 0.0313f
C12172 rowoff_n[13] a_19942_15182# 0.202f
C12173 m2_34288_8402# row_n[6] 0.0128f
C12174 row_n[10] a_10298_12210# 0.0117f
C12175 rowon_n[2] a_32994_4138# 0.118f
C12176 col[31] a_2275_11190# 0.0899f
C12177 vcm a_14010_17190# 0.56f
C12178 ctop a_2475_2154# 0.0466f
C12179 VDD a_10906_7150# 0.181f
C12180 rowoff_n[5] a_21950_7150# 0.202f
C12181 col[9] a_12002_3134# 0.367f
C12182 a_2275_18218# a_15014_18194# 0.0924f
C12183 a_8898_18194# a_9390_18556# 0.0658f
C12184 row_n[0] a_20338_2170# 0.0117f
C12185 a_2275_1150# a_4974_1126# 0.0924f
C12186 a_3878_1126# a_3970_1126# 0.354f
C12187 col[19] a_22042_15182# 0.367f
C12188 a_2874_1126# a_3270_1166# 0.0313f
C12189 col[16] a_18938_5142# 0.0682f
C12190 col_n[22] row_n[7] 0.298f
C12191 col_n[29] rowon_n[10] 0.111f
C12192 col_n[25] rowon_n[8] 0.111f
C12193 col_n[12] row_n[2] 0.298f
C12194 col_n[5] ctop 0.0594f
C12195 col_n[30] row_n[11] 0.298f
C12196 col_n[10] row_n[1] 0.298f
C12197 col_n[21] rowon_n[6] 0.111f
C12198 col_n[23] rowon_n[7] 0.111f
C12199 col_n[31] rowon_n[11] 0.111f
C12200 col_n[19] rowon_n[5] 0.111f
C12201 col_n[14] row_n[3] 0.298f
C12202 col_n[16] row_n[4] 0.298f
C12203 col_n[15] rowon_n[3] 0.111f
C12204 col_n[13] rowon_n[2] 0.111f
C12205 col_n[26] row_n[9] 0.298f
C12206 VDD col[2] 3.83f
C12207 col_n[9] rowon_n[0] 0.111f
C12208 col_n[20] row_n[6] 0.298f
C12209 col_n[17] rowon_n[4] 0.111f
C12210 col_n[28] row_n[10] 0.298f
C12211 col_n[18] row_n[5] 0.298f
C12212 vcm analog_in 0.0445f
C12213 col_n[0] col[0] 0.489f
C12214 col_n[11] rowon_n[1] 0.111f
C12215 col_n[27] rowon_n[9] 0.111f
C12216 col_n[8] row_n[0] 0.298f
C12217 col_n[24] row_n[8] 0.298f
C12218 vcm a_16930_2130# 0.1f
C12219 a_15014_6146# a_16018_6146# 0.843f
C12220 col_n[1] a_2275_8178# 0.113f
C12221 col[26] a_28978_17190# 0.0682f
C12222 a_2475_6170# a_29070_6146# 0.316f
C12223 m2_4744_946# m2_5172_1374# 0.165f
C12224 rowoff_n[3] a_30986_5142# 0.202f
C12225 vcm a_4274_11206# 0.155f
C12226 row_n[2] a_10906_4138# 0.0437f
C12227 row_n[11] rowoff_n[11] 0.209f
C12228 VDD a_1957_1150# 0.404f
C12229 rowon_n[6] a_9994_8154# 0.248f
C12230 ctop a_17022_6146# 4.11f
C12231 a_2475_15206# a_7894_15182# 0.264f
C12232 a_4882_15182# a_4974_15182# 0.326f
C12233 a_3878_15182# a_4274_15222# 0.0313f
C12234 a_2275_15206# a_5278_15222# 0.144f
C12235 VDD a_25966_11166# 0.181f
C12236 col_n[4] a_7286_3174# 0.084f
C12237 col_n[21] a_2475_7174# 0.0531f
C12238 col_n[14] a_17326_15222# 0.084f
C12239 a_2275_3158# a_20034_3134# 0.399f
C12240 a_2475_18218# a_13006_18194# 0.0299f
C12241 rowoff_n[8] a_22442_10524# 0.0133f
C12242 a_35002_1126# a_2275_1150# 0.136f
C12243 vcm a_31990_6146# 0.1f
C12244 a_5978_8154# a_5978_7150# 0.843f
C12245 col_n[25] a_28466_9520# 0.0283f
C12246 vcm a_19334_15222# 0.155f
C12247 col[6] a_2475_15206# 0.136f
C12248 VDD a_17422_5504# 0.0779f
C12249 col[11] a_2475_4162# 0.136f
C12250 a_29374_1166# VDD 0.0149f
C12251 row_n[15] a_21038_17190# 0.282f
C12252 ctop a_32082_10162# 4.11f
C12253 a_2275_17214# a_20338_17230# 0.144f
C12254 a_2475_17214# a_22954_17190# 0.264f
C12255 rowoff_n[6] a_31478_8516# 0.0133f
C12256 VDD a_6890_14178# 0.181f
C12257 a_24050_2130# m2_24248_2378# 0.165f
C12258 a_18026_5142# a_18330_5182# 0.0931f
C12259 a_18938_5142# a_19430_5504# 0.0658f
C12260 row_n[5] a_31078_7150# 0.282f
C12261 a_2275_5166# a_35094_5142# 0.0924f
C12262 col[8] a_10998_13174# 0.367f
C12263 col[5] a_7894_3134# 0.0682f
C12264 rowon_n[9] a_30986_11166# 0.118f
C12265 col_n[25] rowoff_n[12] 0.0471f
C12266 col_n[18] a_2275_10186# 0.113f
C12267 vcm a_12914_9158# 0.1f
C12268 a_30074_10162# a_31078_10162# 0.843f
C12269 rowoff_n[14] a_7894_16186# 0.202f
C12270 col[15] a_17934_15182# 0.0682f
C12271 m3_16924_1078# a_17022_2130# 0.0302f
C12272 a_2275_14202# a_13918_14178# 0.136f
C12273 col_n[23] a_26058_9158# 0.251f
C12274 row_n[7] a_18330_9198# 0.0117f
C12275 VDD a_32482_9520# 0.0779f
C12276 ctop a_13006_13174# 4.11f
C12277 VDD a_21950_18194# 0.343f
C12278 col[3] a_2275_18218# 0.0899f
C12279 col_n[30] a_32994_11166# 0.0765f
C12280 a_2475_2154# a_27974_2130# 0.264f
C12281 a_2275_2154# a_25358_2170# 0.144f
C12282 a_14922_2130# a_15014_2130# 0.326f
C12283 col[8] a_2275_7174# 0.0899f
C12284 col_n[3] a_6282_13214# 0.084f
C12285 m2_31852_946# VDD 1f
C12286 row_n[9] a_8898_11166# 0.0437f
C12287 rowoff_n[9] a_32082_11166# 0.294f
C12288 rowon_n[13] a_7986_15182# 0.248f
C12289 vcm a_27974_13174# 0.1f
C12290 a_2966_11166# a_3270_11206# 0.0931f
C12291 a_2475_11190# a_5978_11166# 0.316f
C12292 a_21038_12170# a_21038_11166# 0.843f
C12293 a_3878_11166# a_4370_11528# 0.0658f
C12294 VDD a_24050_3134# 0.483f
C12295 col[23] a_2475_17214# 0.136f
C12296 m2_12776_18014# a_13310_18234# 0.087f
C12297 col_n[14] a_17422_7512# 0.0283f
C12298 a_2275_16210# a_28978_16186# 0.136f
C12299 a_14922_16186# a_15318_16226# 0.0313f
C12300 col[28] a_2475_6170# 0.136f
C12301 rowon_n[3] a_18026_5142# 0.248f
C12302 VDD a_13406_12532# 0.0779f
C12303 ctop a_28066_17190# 4.06f
C12304 m2_2736_1950# rowon_n[0] 0.233f
C12305 col_n[9] rowoff_n[13] 0.0471f
C12306 a_33086_9158# a_33390_9198# 0.0931f
C12307 a_33998_9158# a_34490_9520# 0.0658f
C12308 m2_29268_14426# a_29070_14178# 0.165f
C12309 col[8] rowoff_n[5] 0.0901f
C12310 col[6] rowoff_n[3] 0.0901f
C12311 col[3] rowoff_n[0] 0.0901f
C12312 col[12] rowoff_n[9] 0.0901f
C12313 col[9] rowoff_n[6] 0.0901f
C12314 col[10] rowoff_n[7] 0.0901f
C12315 col[7] rowoff_n[4] 0.0901f
C12316 col[4] rowoff_n[1] 0.0901f
C12317 col[11] rowoff_n[8] 0.0901f
C12318 col[5] rowoff_n[2] 0.0901f
C12319 vcm a_8898_16186# 0.1f
C12320 a_2475_13198# a_21038_13174# 0.316f
C12321 a_10998_13174# a_12002_13174# 0.843f
C12322 VDD a_4974_6146# 0.483f
C12323 col[4] a_6890_13174# 0.0682f
C12324 m2_32856_18014# a_2475_18218# 0.286f
C12325 VDD a_28466_16548# 0.0779f
C12326 col_n[12] a_15014_7150# 0.251f
C12327 row_n[12] a_29070_14178# 0.282f
C12328 col_n[19] a_21950_9158# 0.0765f
C12329 m2_12200_15430# rowon_n[13] 0.0322f
C12330 vcm a_10998_1126# 0.165f
C12331 col[25] a_2275_9182# 0.0899f
C12332 m2_18224_11414# rowon_n[9] 0.0322f
C12333 a_29982_6146# a_30074_6146# 0.326f
C12334 m2_24248_7398# rowon_n[5] 0.0322f
C12335 m2_30272_3382# rowon_n[1] 0.0322f
C12336 a_2275_10186# a_12002_10162# 0.399f
C12337 row_n[14] a_16322_16226# 0.0117f
C12338 col_n[0] a_2966_13174# 0.251f
C12339 a_2475_15206# a_2475_14202# 0.0666f
C12340 VDD a_20034_10162# 0.483f
C12341 row_n[4] a_26362_6186# 0.0117f
C12342 col_n[3] a_6378_5504# 0.0283f
C12343 col_n[13] a_16418_17552# 0.0283f
C12344 a_24962_3134# a_25358_3174# 0.0313f
C12345 vcm a_26058_5142# 0.56f
C12346 a_2275_7174# a_3878_7150# 0.136f
C12347 rowoff_n[2] a_2874_4138# 0.202f
C12348 rowoff_n[10] a_20034_12170# 0.294f
C12349 a_2475_7174# a_4882_7150# 0.264f
C12350 a_2874_7150# a_3366_7512# 0.0658f
C12351 m2_20232_12418# a_20034_12170# 0.165f
C12352 col_n[10] a_2475_16210# 0.0531f
C12353 row_n[6] a_16930_8154# 0.0437f
C12354 col_n[15] a_2475_5166# 0.0531f
C12355 a_14922_12170# a_15414_12532# 0.0658f
C12356 a_14010_12170# a_14314_12210# 0.0931f
C12357 a_2275_12194# a_27062_12170# 0.399f
C12358 rowon_n[10] a_16018_12170# 0.248f
C12359 a_26058_17190# a_27062_17190# 0.843f
C12360 rowoff_n[0] a_12002_2130# 0.294f
C12361 rowon_n[0] a_26058_2130# 0.248f
C12362 col_n[27] a_30378_6186# 0.084f
C12363 col[0] a_2475_13198# 0.148f
C12364 col_n[1] a_3970_5142# 0.251f
C12365 col[5] a_2475_2154# 0.136f
C12366 col_n[11] a_14010_17190# 0.251f
C12367 vcm a_6982_8154# 0.56f
C12368 col_n[8] a_10906_7150# 0.0765f
C12369 a_2275_9182# a_17326_9198# 0.144f
C12370 a_2475_9182# a_19942_9158# 0.264f
C12371 a_10906_9158# a_10998_9158# 0.326f
C12372 rowoff_n[5] a_3878_7150# 0.202f
C12373 col_n[22] rowon_n[1] 0.111f
C12374 col_n[31] row_n[6] 0.298f
C12375 col_n[25] row_n[3] 0.298f
C12376 col_n[26] rowon_n[3] 0.111f
C12377 col_n[29] row_n[5] 0.298f
C12378 col_n[30] rowon_n[5] 0.111f
C12379 col_n[24] rowon_n[2] 0.111f
C12380 col_n[28] rowon_n[4] 0.111f
C12381 col_n[27] row_n[4] 0.298f
C12382 col_n[19] row_n[0] 0.298f
C12383 col_n[23] row_n[2] 0.298f
C12384 col_n[5] col[5] 0.489f
C12385 vcm col[10] 5.46f
C12386 VDD col[13] 3.83f
C12387 col_n[16] ctop 0.0619f
C12388 col_n[20] rowon_n[0] 0.111f
C12389 rowon_n[11] rowon_n[10] 0.0632f
C12390 col_n[21] row_n[1] 0.298f
C12391 row_n[0] a_3970_2130# 0.282f
C12392 VDD a_16018_17190# 0.484f
C12393 col_n[12] a_2275_8178# 0.113f
C12394 vcm a_31382_3174# 0.155f
C12395 a_2275_6170# a_10906_6146# 0.136f
C12396 a_5886_6146# a_6282_6186# 0.0313f
C12397 col_n[2] a_5374_15544# 0.0283f
C12398 m2_11196_10410# a_10998_10162# 0.165f
C12399 vcm a_22042_12170# 0.56f
C12400 a_2275_11190# a_32386_11206# 0.144f
C12401 a_2475_11190# a_35002_11166# 0.264f
C12402 col[21] a_24050_4138# 0.367f
C12403 VDD a_18938_2130# 0.181f
C12404 m2_31852_18014# a_32386_18234# 0.087f
C12405 col[31] a_34090_16186# 0.367f
C12406 col[28] a_30986_6146# 0.0682f
C12407 row_n[11] a_24354_13214# 0.0117f
C12408 col[2] a_2275_5166# 0.0899f
C12409 a_29982_16186# a_30474_16548# 0.0658f
C12410 a_29070_16186# a_29374_16226# 0.0931f
C12411 m2_34864_18014# m3_34996_17142# 0.0341f
C12412 a_1957_3158# a_2275_3158# 0.158f
C12413 a_2475_3158# a_2874_3134# 0.264f
C12414 row_n[1] a_35398_3174# 0.0117f
C12415 rowoff_n[8] a_4882_10162# 0.202f
C12416 m2_30272_6394# a_30074_6146# 0.165f
C12417 row_n[13] a_14922_15182# 0.0437f
C12418 col[17] a_2475_15206# 0.136f
C12419 vcm a_12306_6186# 0.155f
C12420 rowoff_n[11] a_7986_13174# 0.294f
C12421 a_2275_8178# a_25966_8154# 0.136f
C12422 col[22] a_2475_4162# 0.136f
C12423 col_n[16] a_19334_4178# 0.084f
C12424 col_n[26] a_29374_16226# 0.084f
C12425 vcm a_2874_15182# 0.1f
C12426 a_25966_13174# a_26058_13174# 0.326f
C12427 VDD a_33998_6146# 0.181f
C12428 row_n[3] a_24962_5142# 0.0437f
C12429 row_n[15] a_2966_17190# 0.281f
C12430 col_n[7] a_9902_17190# 0.0765f
C12431 m2_11196_14426# row_n[12] 0.0128f
C12432 a_2275_17214# a_3970_17190# 0.399f
C12433 rowon_n[7] a_24050_9158# 0.248f
C12434 m2_17220_10410# row_n[8] 0.0128f
C12435 rowoff_n[6] a_13918_8154# 0.202f
C12436 m2_23244_6394# row_n[4] 0.0128f
C12437 col_n[29] a_2275_10186# 0.113f
C12438 a_27062_6146# a_27062_5142# 0.843f
C12439 a_2475_5166# a_18026_5142# 0.316f
C12440 m2_1732_7974# a_1957_8178# 0.245f
C12441 vcm a_27366_10202# 0.155f
C12442 rowoff_n[15] a_24050_17190# 0.294f
C12443 a_20946_10162# a_21342_10202# 0.0313f
C12444 rowoff_n[4] a_22954_6146# 0.202f
C12445 ctop a_5978_4138# 4.11f
C12446 col[14] a_2275_18218# 0.0899f
C12447 VDD a_14922_9158# 0.181f
C12448 row_n[7] a_2475_9182# 0.405f
C12449 col[10] a_13006_2130# 0.367f
C12450 col[19] a_2275_7174# 0.0899f
C12451 col[20] a_23046_14178# 0.367f
C12452 col[17] a_19942_4138# 0.0682f
C12453 VDD a_3878_18194# 0.343f
C12454 a_2275_2154# a_8990_2130# 0.399f
C12455 a_4974_2130# a_5278_2170# 0.0931f
C12456 a_5886_2130# a_6378_2492# 0.0658f
C12457 col[27] a_29982_16186# 0.0682f
C12458 m2_21236_4386# a_21038_4138# 0.165f
C12459 vcm a_20946_4138# 0.1f
C12460 rowoff_n[2] a_31990_4138# 0.202f
C12461 rowon_n[1] a_11910_3134# 0.118f
C12462 a_2475_7174# a_33086_7150# 0.316f
C12463 a_17022_7150# a_18026_7150# 0.843f
C12464 rowoff_n[9] a_14410_11528# 0.0133f
C12465 vcm a_8290_13214# 0.155f
C12466 VDD a_6378_3496# 0.0779f
C12467 col_n[5] a_8290_2170# 0.084f
C12468 m2_1732_18014# a_2161_18218# 0.0454f
C12469 m2_34864_13998# VDD 0.783f
C12470 ctop a_21038_8154# 4.11f
C12471 col_n[15] a_18330_14218# 0.084f
C12472 a_2475_16210# a_11910_16186# 0.264f
C12473 a_6890_16186# a_6982_16186# 0.326f
C12474 a_2275_16210# a_9294_16226# 0.144f
C12475 VDD a_29982_13174# 0.181f
C12476 col_n[20] rowoff_n[13] 0.0471f
C12477 row_n[8] a_32386_10202# 0.0117f
C12478 rowoff_n[7] a_23446_9520# 0.0133f
C12479 col_n[4] a_2475_14202# 0.0531f
C12480 a_2275_4162# a_24050_4138# 0.399f
C12481 m3_17928_1078# ctop 0.354f
C12482 col_n[9] a_2475_3158# 0.0531f
C12483 col[14] rowoff_n[0] 0.0901f
C12484 col[23] rowoff_n[9] 0.0901f
C12485 col[18] rowoff_n[4] 0.0901f
C12486 col[22] rowoff_n[8] 0.0901f
C12487 col[15] rowoff_n[1] 0.0901f
C12488 col[17] rowoff_n[3] 0.0901f
C12489 col[19] rowoff_n[5] 0.0901f
C12490 col[16] rowoff_n[2] 0.0901f
C12491 col[20] rowoff_n[6] 0.0901f
C12492 col[21] rowoff_n[7] 0.0901f
C12493 vcm a_34394_8194# 0.155f
C12494 m2_34864_17010# m2_35292_17438# 0.165f
C12495 col_n[26] a_29470_8516# 0.0283f
C12496 a_7986_9158# a_7986_8154# 0.843f
C12497 rowoff_n[13] a_30474_15544# 0.0133f
C12498 row_n[10] a_22954_12170# 0.0437f
C12499 col[0] a_2475_18218# 0.148f
C12500 vcm a_23350_17230# 0.155f
C12501 rowon_n[14] a_22042_16186# 0.248f
C12502 a_2475_13198# a_2966_13174# 0.317f
C12503 a_2161_13198# a_2275_13198# 0.183f
C12504 VDD a_21438_7512# 0.0779f
C12505 rowoff_n[5] a_32482_7512# 0.0133f
C12506 ctop a_2475_11190# 0.0488f
C12507 a_2275_18218# a_24354_18234# 0.145f
C12508 m3_1864_9110# a_2966_9158# 0.0302f
C12509 row_n[0] a_32994_2130# 0.0437f
C12510 VDD a_10906_16186# 0.181f
C12511 a_2475_1150# a_16930_1126# 0.264f
C12512 a_2275_1150# a_14314_1166# 0.145f
C12513 rowon_n[4] a_32082_6146# 0.248f
C12514 col[9] a_12002_12170# 0.367f
C12515 col[6] a_8898_2130# 0.0682f
C12516 a_20946_6146# a_21438_6508# 0.0658f
C12517 a_20034_6146# a_20338_6186# 0.0931f
C12518 col[16] a_18938_14178# 0.0682f
C12519 vcm a_16930_11166# 0.1f
C12520 col_n[1] a_2275_17214# 0.113f
C12521 a_32082_11166# a_33086_11166# 0.843f
C12522 VDD a_13006_1126# 0.035f
C12523 col_n[24] a_27062_8154# 0.251f
C12524 col_n[6] a_2275_6170# 0.113f
C12525 a_2275_15206# a_17934_15182# 0.136f
C12526 col_n[4] rowoff_n[14] 0.0471f
C12527 VDD a_1957_10186# 0.196f
C12528 m2_34864_15002# m3_34996_14130# 0.0341f
C12529 col_n[31] a_33998_10162# 0.0765f
C12530 rowon_n[0] m2_34864_1950# 0.231f
C12531 ctop a_17022_15182# 4.11f
C12532 row_n[4] a_9994_6146# 0.282f
C12533 col_n[4] a_7286_12210# 0.084f
C12534 col[0] a_2966_10162# 0.367f
C12535 a_2275_3158# a_29374_3174# 0.144f
C12536 col[7] rowoff_n[10] 0.0901f
C12537 a_2475_3158# a_31990_3134# 0.264f
C12538 rowon_n[8] a_9902_10162# 0.118f
C12539 a_16930_3134# a_17022_3134# 0.326f
C12540 rowoff_n[8] a_33086_10162# 0.294f
C12541 col_n[21] a_2475_16210# 0.0531f
C12542 col_n[26] a_2475_5166# 0.0531f
C12543 rowoff_n[10] a_1957_12194# 0.0219f
C12544 vcm a_31990_15182# 0.1f
C12545 a_2475_12194# a_9994_12170# 0.316f
C12546 a_23046_13174# a_23046_12170# 0.843f
C12547 col_n[15] a_18426_6508# 0.0283f
C12548 VDD a_28066_5142# 0.483f
C12549 col_n[25] a_28466_18556# 0.0283f
C12550 m2_14208_18442# VDD 0.0456f
C12551 row_n[15] a_30378_17230# 0.0117f
C12552 a_16930_17190# a_17326_17230# 0.0313f
C12553 a_2275_17214# a_32994_17190# 0.136f
C12554 VDD a_17422_14540# 0.0779f
C12555 col[11] a_2475_13198# 0.136f
C12556 col[16] a_2475_2154# 0.136f
C12557 col_n[0] a_2874_2130# 0.0765f
C12558 rowoff_n[14] a_18426_16548# 0.0133f
C12559 col[5] a_7894_12170# 0.0682f
C12560 col_n[31] rowon_n[0] 0.111f
C12561 vcm col[21] 5.46f
C12562 rowon_n[8] row_n[8] 18.9f
C12563 col_n[27] ctop 0.0595f
C12564 VDD col[24] 3.83f
C12565 vcm a_12914_18194# 0.101f
C12566 col_n[30] row_n[0] 0.298f
C12567 col_n[10] col[11] 7.13f
C12568 a_13006_14178# a_14010_14178# 0.843f
C12569 a_2475_14202# a_25054_14178# 0.316f
C12570 VDD a_8990_8154# 0.483f
C12571 col_n[23] a_2275_8178# 0.113f
C12572 row_n[7] a_30986_9158# 0.0437f
C12573 m2_1732_12994# rowon_n[11] 0.236f
C12574 m2_7180_9406# rowon_n[7] 0.0322f
C12575 m2_13204_5390# rowon_n[3] 0.0322f
C12576 col_n[13] a_16018_6146# 0.251f
C12577 rowon_n[11] a_30074_13174# 0.248f
C12578 VDD a_32482_18556# 0.0858f
C12579 col_n[20] a_22954_8154# 0.0765f
C12580 vcm a_15014_3134# 0.56f
C12581 a_31990_7150# a_32082_7150# 0.326f
C12582 col[8] a_2275_16210# 0.0899f
C12583 col[13] a_2275_5166# 0.0899f
C12584 a_2275_11190# a_16018_11166# 0.399f
C12585 a_3970_16186# a_3970_15182# 0.843f
C12586 row_n[11] a_7986_13174# 0.282f
C12587 VDD a_24050_12170# 0.483f
C12588 col_n[4] a_7382_4500# 0.0283f
C12589 m2_11772_18014# m3_11904_18146# 3.79f
C12590 rowon_n[15] a_7894_17190# 0.118f
C12591 m2_28264_14426# rowon_n[12] 0.0322f
C12592 col_n[14] a_17422_16548# 0.0283f
C12593 col[28] a_2475_15206# 0.136f
C12594 m2_34288_10410# rowon_n[8] 0.0322f
C12595 a_26970_4138# a_27366_4178# 0.0313f
C12596 rowoff_n[1] a_3970_3134# 0.294f
C12597 row_n[1] a_18026_3134# 0.282f
C12598 rowon_n[5] a_17934_7150# 0.118f
C12599 vcm a_30074_7150# 0.56f
C12600 rowoff_n[12] a_24962_14178# 0.202f
C12601 a_2475_8178# a_8898_8154# 0.264f
C12602 a_2275_8178# a_6282_8194# 0.144f
C12603 m2_3164_13422# a_2966_13174# 0.165f
C12604 a_2275_13198# a_31078_13174# 0.399f
C12605 a_16930_13174# a_17422_13536# 0.0658f
C12606 a_16018_13174# a_16322_13214# 0.0931f
C12607 row_n[3] a_5278_5182# 0.0117f
C12608 col_n[3] a_2475_1150# 0.0531f
C12609 VDD a_4974_15182# 0.483f
C12610 col_n[2] a_4974_4138# 0.251f
C12611 col_n[28] a_31382_5182# 0.084f
C12612 vcm a_20338_1166# 0.155f
C12613 col_n[12] a_15014_16186# 0.251f
C12614 a_35002_6146# a_35398_6186# 0.0313f
C12615 col_n[9] a_11910_6146# 0.0765f
C12616 m2_14784_946# m3_13912_1078# 0.0341f
C12617 col[25] a_2275_18218# 0.0899f
C12618 vcm a_10998_10162# 0.56f
C12619 col_n[19] a_21950_18194# 0.0762f
C12620 a_12914_10162# a_13006_10162# 0.326f
C12621 a_2475_10186# a_23958_10162# 0.264f
C12622 a_2275_10186# a_21342_10202# 0.144f
C12623 rowoff_n[15] a_6378_17552# 0.0133f
C12624 row_n[14] a_28978_16186# 0.0437f
C12625 col[30] a_2275_7174# 0.0899f
C12626 m2_2736_18014# ctop 0.0422f
C12627 m2_34864_11990# m3_34996_11118# 0.0341f
C12628 a_14010_3134# a_14010_2130# 0.843f
C12629 col_n[3] a_6378_14540# 0.0283f
C12630 vcm a_2275_4162# 6.49f
C12631 a_7894_7150# a_8290_7190# 0.0313f
C12632 a_2275_7174# a_14922_7150# 0.136f
C12633 m3_34568_1078# sw_n 0.0611f
C12634 col[22] a_25054_3134# 0.367f
C12635 m2_31852_18014# vcm 0.353f
C12636 vcm a_26058_14178# 0.56f
C12637 a_2966_12170# a_2966_11166# 0.843f
C12638 VDD a_22954_4138# 0.181f
C12639 col[29] a_31990_5142# 0.0682f
C12640 col_n[31] rowoff_n[13] 0.0471f
C12641 ctop a_2966_8154# 4.06f
C12642 col_n[15] a_2475_14202# 0.0531f
C12643 a_31078_17190# a_31382_17230# 0.0931f
C12644 a_31990_17190# a_32482_17552# 0.0658f
C12645 col_n[20] a_2475_3158# 0.0531f
C12646 col[26] rowoff_n[1] 0.0901f
C12647 col[28] rowoff_n[3] 0.0901f
C12648 col[30] rowoff_n[5] 0.0901f
C12649 col[29] rowoff_n[4] 0.0901f
C12650 col[27] rowoff_n[2] 0.0901f
C12651 col[31] rowoff_n[6] 0.0901f
C12652 col[25] rowoff_n[0] 0.0901f
C12653 row_n[8] a_16018_10162# 0.282f
C12654 sample_n rowoff_n[7] 0.14f
C12655 rowoff_n[7] a_5886_9158# 0.202f
C12656 rowon_n[12] a_15926_14178# 0.118f
C12657 a_2475_4162# a_6982_4138# 0.316f
C12658 a_3970_4138# a_4974_4138# 0.843f
C12659 m3_13912_18146# ctop 0.209f
C12660 col[11] a_2475_18218# 0.136f
C12661 col_n[17] a_20338_3174# 0.084f
C12662 vcm a_16322_8194# 0.155f
C12663 m2_6176_8402# row_n[6] 0.0128f
C12664 col_n[27] a_30378_15222# 0.084f
C12665 a_2275_9182# a_29982_9158# 0.136f
C12666 col_n[1] a_3970_14178# 0.251f
C12667 rowoff_n[13] a_12914_15182# 0.202f
C12668 m2_12200_4386# row_n[2] 0.0128f
C12669 row_n[10] a_3270_12210# 0.0117f
C12670 m2_34864_15002# a_35094_15182# 0.0249f
C12671 rowon_n[2] a_25966_4138# 0.118f
C12672 col[5] a_2475_11190# 0.136f
C12673 ctop a_29070_3134# 4.11f
C12674 vcm a_6982_17190# 0.56f
C12675 a_27974_14178# a_28066_14178# 0.326f
C12676 col_n[8] a_10906_16186# 0.0765f
C12677 VDD a_3366_7512# 0.0779f
C12678 rowoff_n[5] a_14922_7150# 0.202f
C12679 a_2275_18218# a_7986_18194# 0.0924f
C12680 row_n[0] a_13310_2170# 0.0117f
C12681 col_n[12] a_2275_17214# 0.113f
C12682 vcm a_9902_2130# 0.1f
C12683 a_29070_7150# a_29070_6146# 0.843f
C12684 a_2475_6170# a_22042_6146# 0.316f
C12685 col_n[17] a_2275_6170# 0.113f
C12686 rowoff_n[3] a_23958_5142# 0.202f
C12687 vcm a_31382_12210# 0.155f
C12688 col_n[15] rowoff_n[14] 0.0471f
C12689 a_22954_11166# a_23350_11206# 0.0313f
C12690 VDD a_29470_2492# 0.0779f
C12691 m2_21236_17438# row_n[15] 0.0128f
C12692 m2_7180_17438# a_6982_17190# 0.165f
C12693 m2_27260_13422# row_n[11] 0.0128f
C12694 rowon_n[6] a_2874_8154# 0.118f
C12695 m2_33284_9406# row_n[7] 0.0128f
C12696 ctop a_9994_6146# 4.11f
C12697 col[21] a_24050_13174# 0.367f
C12698 VDD a_18938_11166# 0.181f
C12699 col[18] a_20946_3134# 0.0682f
C12700 col[18] rowoff_n[10] 0.0901f
C12701 col[28] a_30986_15182# 0.0682f
C12702 col[2] a_2275_14202# 0.0899f
C12703 a_2475_18218# a_5978_18194# 0.0299f
C12704 a_7894_3134# a_8386_3496# 0.0658f
C12705 col[7] a_2275_3158# 0.0899f
C12706 a_2275_3158# a_13006_3134# 0.399f
C12707 a_6982_3134# a_7286_3174# 0.0931f
C12708 rowoff_n[8] a_15414_10524# 0.0133f
C12709 rowoff_n[1] a_32994_3134# 0.202f
C12710 a_26970_1126# a_2275_1150# 0.136f
C12711 vcm a_24962_6146# 0.1f
C12712 a_19030_8154# a_20034_8154# 0.843f
C12713 m2_26256_13422# a_26058_13174# 0.165f
C12714 col_n[6] a_9294_1166# 0.0839f
C12715 vcm a_12306_15222# 0.155f
C12716 VDD a_10394_5504# 0.0779f
C12717 col_n[16] a_19334_13214# 0.084f
C12718 col[22] a_2475_13198# 0.136f
C12719 a_22346_1166# VDD 0.0149f
C12720 col[27] a_2475_2154# 0.136f
C12721 ctop a_25054_10162# 4.11f
C12722 row_n[15] a_14010_17190# 0.282f
C12723 a_2275_17214# a_13310_17230# 0.144f
C12724 a_2475_17214# a_15926_17190# 0.264f
C12725 a_8898_17190# a_8990_17190# 0.326f
C12726 VDD a_33998_15182# 0.181f
C12727 rowoff_n[6] a_24450_8516# 0.0133f
C12728 a_2275_5166# a_28066_5142# 0.399f
C12729 row_n[5] a_24050_7150# 0.282f
C12730 col_n[27] a_30474_7512# 0.0283f
C12731 col_n[16] col[16] 0.413f
C12732 rowon_n[15] col[0] 0.0318f
C12733 rowon_n[12] ctop 0.203f
C12734 col_n[0] rowoff_n[15] 0.0471f
C12735 vcm sample_n 1.81f
C12736 rowon_n[9] a_23958_11166# 0.118f
C12737 vcm a_5886_9158# 0.1f
C12738 a_28978_1126# a_29470_1488# 0.0658f
C12739 a_9994_10162# a_9994_9158# 0.843f
C12740 rowoff_n[4] a_33486_6508# 0.0133f
C12741 col[2] rowoff_n[11] 0.0901f
C12742 m2_7756_946# a_8290_1166# 0.087f
C12743 m2_24824_946# a_2475_1150# 0.286f
C12744 a_2275_14202# a_6890_14178# 0.136f
C12745 row_n[7] a_11302_9198# 0.0117f
C12746 VDD a_25454_9520# 0.0779f
C12747 m2_34864_8978# m3_34996_8106# 0.0341f
C12748 ctop a_5978_13174# 4.11f
C12749 col[10] a_13006_11166# 0.367f
C12750 VDD a_14922_18194# 0.343f
C12751 m2_11772_18014# col[9] 0.347f
C12752 a_2275_2154# a_18330_2170# 0.144f
C12753 col[19] a_2275_16210# 0.0899f
C12754 a_2475_2154# a_20946_2130# 0.264f
C12755 col[7] a_9902_1126# 0.0682f
C12756 col[24] a_2275_5166# 0.0899f
C12757 m2_16216_1374# VDD 0.0194f
C12758 col[17] a_19942_13174# 0.0682f
C12759 a_22042_7150# a_22346_7190# 0.0931f
C12760 rowoff_n[9] a_25054_11166# 0.294f
C12761 a_22954_7150# a_23446_7512# 0.0658f
C12762 m2_34864_15002# vcm 0.408f
C12763 m2_17220_11414# a_17022_11166# 0.165f
C12764 col_n[25] a_28066_7150# 0.251f
C12765 vcm a_20946_13174# 0.1f
C12766 a_33998_12170# a_34394_12210# 0.0313f
C12767 VDD a_17022_3134# 0.483f
C12768 m2_22816_18014# a_2275_18218# 0.28f
C12769 a_2275_16210# a_21950_16186# 0.136f
C12770 rowon_n[3] a_10998_5142# 0.248f
C12771 VDD a_6378_12532# 0.0779f
C12772 col_n[5] a_8290_11206# 0.084f
C12773 a_28978_1126# m2_28840_946# 0.225f
C12774 ctop a_21038_17190# 4.06f
C12775 rowoff_n[7] a_34090_9158# 0.294f
C12776 a_18938_4138# a_19030_4138# 0.326f
C12777 a_2275_4162# a_33390_4178# 0.144f
C12778 col_n[16] a_19430_5504# 0.0283f
C12779 col_n[9] a_2475_12194# 0.0531f
C12780 col_n[14] a_2475_1150# 0.0531f
C12781 vcm a_34394_17230# 0.155f
C12782 col_n[26] a_29470_17552# 0.0283f
C12783 a_2475_13198# a_14010_13174# 0.316f
C12784 a_25054_14178# a_25054_13174# 0.843f
C12785 VDD a_32082_7150# 0.483f
C12786 a_18938_18194# a_19334_18234# 0.0313f
C12787 m2_18800_18014# a_2475_18218# 0.286f
C12788 VDD a_21438_16548# 0.0779f
C12789 row_n[12] a_22042_14178# 0.282f
C12790 a_13918_1126# a_14314_1166# 0.0313f
C12791 vcm a_3970_1126# 0.557f
C12792 m2_8184_9406# a_7986_9158# 0.165f
C12793 m2_2160_3382# rowon_n[1] 0.0219f
C12794 m2_27836_946# m2_28264_1374# 0.165f
C12795 row_n[2] a_32082_4138# 0.282f
C12796 col[6] a_8898_11166# 0.0682f
C12797 m2_27836_18014# col_n[25] 0.243f
C12798 a_2874_10162# a_3270_10202# 0.0313f
C12799 a_3878_10162# a_3970_10162# 0.326f
C12800 a_2275_10186# a_4974_10162# 0.399f
C12801 row_n[14] a_9294_16226# 0.0117f
C12802 rowon_n[6] a_31990_8154# 0.118f
C12803 col_n[14] a_17022_5142# 0.251f
C12804 a_2475_15206# a_29070_15182# 0.316f
C12805 a_15014_15182# a_16018_15182# 0.843f
C12806 VDD a_13006_10162# 0.483f
C12807 col_n[24] a_27062_17190# 0.251f
C12808 col_n[6] a_2275_15206# 0.113f
C12809 col_n[21] a_23958_7150# 0.0765f
C12810 row_n[4] a_19334_6186# 0.0117f
C12811 col_n[11] a_2275_4162# 0.113f
C12812 a_2475_18218# a_35002_18194# 0.264f
C12813 m2_27260_5390# a_27062_5142# 0.165f
C12814 vcm a_19030_5142# 0.56f
C12815 rowoff_n[10] a_13006_12170# 0.294f
C12816 a_33998_8154# a_34090_8154# 0.326f
C12817 a_32994_1126# vcm 0.0988f
C12818 m2_11196_16434# rowon_n[14] 0.0322f
C12819 row_n[6] a_9902_8154# 0.0437f
C12820 m2_17220_12418# rowon_n[10] 0.0322f
C12821 m2_1732_5966# sample 0.2f
C12822 m2_23244_8402# rowon_n[6] 0.0322f
C12823 col_n[26] a_2475_14202# 0.0531f
C12824 m2_29268_4386# rowon_n[2] 0.0322f
C12825 a_2275_12194# a_20034_12170# 0.399f
C12826 rowon_n[10] a_8990_12170# 0.248f
C12827 col_n[31] a_2475_3158# 0.0531f
C12828 col_n[5] a_8386_3496# 0.0283f
C12829 m2_1732_17010# VDD 0.856f
C12830 col[1] a_2275_1150# 0.0899f
C12831 col_n[15] a_18426_15544# 0.0283f
C12832 a_5978_17190# a_5978_16186# 0.843f
C12833 VDD a_28066_14178# 0.483f
C12834 col[22] a_2475_18218# 0.136f
C12835 rowon_n[0] a_19030_2130# 0.248f
C12836 rowoff_n[0] a_4974_2130# 0.294f
C12837 a_28978_5142# a_29374_5182# 0.0313f
C12838 m2_4744_946# ctop 0.0435f
C12839 col[16] a_2475_11190# 0.136f
C12840 vcm a_34090_9158# 0.56f
C12841 a_2275_9182# a_10298_9198# 0.144f
C12842 rowoff_n[14] a_29070_16186# 0.294f
C12843 a_2475_9182# a_12914_9158# 0.264f
C12844 col_n[0] a_2874_11166# 0.0765f
C12845 a_18938_14178# a_19430_14540# 0.0658f
C12846 a_18026_14178# a_18330_14218# 0.0931f
C12847 a_2275_14202# a_35094_14178# 0.0924f
C12848 m2_34864_5966# m3_34996_5094# 0.0341f
C12849 col_n[29] a_32386_4178# 0.084f
C12850 col_n[3] a_5978_3134# 0.251f
C12851 VDD a_8990_17190# 0.484f
C12852 col_n[23] a_2275_17214# 0.113f
C12853 a_25054_2130# a_26058_2130# 0.843f
C12854 col_n[13] a_16018_15182# 0.251f
C12855 col_n[28] a_2275_6170# 0.113f
C12856 m2_18224_3382# a_18026_3134# 0.165f
C12857 col_n[10] a_12914_5142# 0.0765f
C12858 m3_12908_1078# VDD 0.0157f
C12859 col_n[26] rowoff_n[14] 0.0471f
C12860 row_n[9] a_30074_11166# 0.282f
C12861 vcm a_24354_3174# 0.155f
C12862 a_2874_6146# a_2966_6146# 0.326f
C12863 col_n[20] a_22954_17190# 0.0765f
C12864 rowon_n[13] a_29982_15182# 0.118f
C12865 vcm a_15014_12170# 0.56f
C12866 a_14922_11166# a_15014_11166# 0.326f
C12867 a_2275_11190# a_25358_11206# 0.144f
C12868 a_2475_11190# a_27974_11166# 0.264f
C12869 col[29] rowoff_n[10] 0.0901f
C12870 VDD a_11910_2130# 0.181f
C12871 col[13] a_2275_14202# 0.0899f
C12872 row_n[11] a_17326_13214# 0.0117f
C12873 col[18] a_2275_3158# 0.0899f
C12874 m2_25828_18014# m3_26964_18146# 0.0341f
C12875 col_n[4] a_7382_13536# 0.0283f
C12876 col_n[1] a_3878_3134# 0.0765f
C12877 a_16018_4138# a_16018_3134# 0.843f
C12878 row_n[1] a_27366_3174# 0.0117f
C12879 col[23] a_26058_2130# 0.367f
C12880 row_n[13] a_7894_15182# 0.0437f
C12881 vcm a_5278_6186# 0.155f
C12882 a_2275_8178# a_18938_8154# 0.136f
C12883 rowoff_n[12] a_35494_14540# 0.0133f
C12884 a_9902_8154# a_10298_8194# 0.0313f
C12885 col[30] a_32994_4138# 0.0682f
C12886 vcm a_30074_16186# 0.56f
C12887 ctop a_18026_1126# 1.07f
C12888 VDD a_26970_6146# 0.181f
C12889 row_n[3] a_17934_5142# 0.0437f
C12890 rowon_n[7] a_17022_9158# 0.248f
C12891 a_33998_18194# a_34490_18556# 0.0658f
C12892 rowoff_n[6] a_6890_8154# 0.202f
C12893 m2_1732_1950# row_n[0] 0.292f
C12894 rowon_n[14] col[9] 0.0323f
C12895 row_n[12] col[4] 0.0342f
C12896 row_n[15] col[10] 0.0342f
C12897 row_n[11] col[2] 0.0342f
C12898 rowon_n[10] col[1] 0.0323f
C12899 row_n[7] ctop 0.186f
C12900 rowon_n[13] col[7] 0.0323f
C12901 rowon_n[12] col[5] 0.0323f
C12902 col_n[21] col[22] 7.13f
C12903 row_n[13] col[6] 0.0342f
C12904 row_n[14] col[8] 0.0342f
C12905 row_n[10] col[0] 0.0322f
C12906 col_n[3] a_2475_10186# 0.0531f
C12907 rowon_n[15] col[11] 0.0323f
C12908 col_n[10] rowoff_n[15] 0.0471f
C12909 rowon_n[11] col[3] 0.0323f
C12910 col_n[18] a_21342_2170# 0.084f
C12911 m2_1732_2954# m2_2160_3382# 0.165f
C12912 a_5978_5142# a_6982_5142# 0.843f
C12913 a_2475_5166# a_10998_5142# 0.316f
C12914 col_n[2] a_4974_13174# 0.251f
C12915 col_n[28] a_31382_14218# 0.084f
C12916 m2_29844_946# m3_29976_1078# 3.79f
C12917 col[13] rowoff_n[11] 0.0901f
C12918 vcm a_20338_10202# 0.155f
C12919 a_2275_10186# a_33998_10162# 0.136f
C12920 rowoff_n[15] a_17022_17190# 0.294f
C12921 col_n[9] a_11910_15182# 0.0765f
C12922 rowoff_n[4] a_15926_6146# 0.202f
C12923 ctop a_33086_5142# 4.11f
C12924 a_29982_15182# a_30074_15182# 0.326f
C12925 VDD a_7894_9158# 0.181f
C12926 col[30] a_2275_16210# 0.0899f
C12927 m2_10192_15430# row_n[13] 0.0128f
C12928 a_2475_2154# a_2275_2154# 2.76f
C12929 a_1957_2154# a_2161_2154# 0.115f
C12930 m2_16216_11414# row_n[9] 0.0128f
C12931 m2_22240_7398# row_n[5] 0.0128f
C12932 m2_28264_3382# row_n[1] 0.0128f
C12933 vcm a_13918_4138# 0.1f
C12934 a_2475_7174# a_26058_7150# 0.316f
C12935 a_31078_8154# a_31078_7150# 0.843f
C12936 rowoff_n[2] a_24962_4138# 0.202f
C12937 rowon_n[1] a_4882_3134# 0.118f
C12938 rowoff_n[9] a_7382_11528# 0.0133f
C12939 m2_1732_10986# a_2966_11166# 0.843f
C12940 vcm a_2275_13198# 6.49f
C12941 a_24962_12170# a_25358_12210# 0.0313f
C12942 VDD a_33486_4500# 0.0779f
C12943 col[22] a_25054_12170# 0.367f
C12944 col_n[5] a_2275_2154# 0.113f
C12945 col[19] a_21950_2130# 0.0682f
C12946 ctop a_14010_8154# 4.11f
C12947 a_2475_16210# a_4882_16186# 0.264f
C12948 a_2874_16186# a_3366_16548# 0.0658f
C12949 a_2275_16210# a_3878_16186# 0.136f
C12950 VDD a_22954_13174# 0.181f
C12951 col[29] a_31990_14178# 0.0682f
C12952 row_n[8] a_25358_10202# 0.0117f
C12953 m2_34864_2954# m2_34864_1950# 0.843f
C12954 ctop a_2966_17190# 4.02f
C12955 rowoff_n[7] a_16418_9520# 0.0133f
C12956 rowoff_n[0] a_33998_2130# 0.202f
C12957 a_9902_4138# a_10394_4500# 0.0658f
C12958 a_8990_4138# a_9294_4178# 0.0931f
C12959 col_n[20] a_2475_12194# 0.0531f
C12960 a_2275_4162# a_17022_4138# 0.399f
C12961 m3_34996_7102# ctop 0.209f
C12962 col_n[25] a_2475_1150# 0.0531f
C12963 vcm a_28978_8154# 0.1f
C12964 rowoff_n[13] a_23446_15544# 0.0133f
C12965 a_21038_9158# a_22042_9158# 0.843f
C12966 m2_34864_4962# rowoff_n[3] 0.278f
C12967 col_n[17] a_20338_12210# 0.084f
C12968 row_n[10] a_15926_12170# 0.0437f
C12969 m2_34864_13998# a_2275_14202# 0.278f
C12970 vcm a_16322_17230# 0.155f
C12971 rowon_n[14] a_15014_16186# 0.248f
C12972 VDD a_14410_7512# 0.0779f
C12973 rowoff_n[5] a_25454_7512# 0.0133f
C12974 ctop a_29070_12170# 4.11f
C12975 a_2275_18218# a_17326_18234# 0.145f
C12976 a_10906_18194# a_10998_18194# 0.0991f
C12977 row_n[0] a_25966_2130# 0.0437f
C12978 col[10] a_2475_9182# 0.136f
C12979 VDD a_3366_16548# 0.0779f
C12980 a_2275_1150# a_7286_1166# 0.145f
C12981 a_5886_1126# a_5978_1126# 0.0991f
C12982 a_2475_1150# a_9902_1126# 0.264f
C12983 rowon_n[4] a_25054_6146# 0.248f
C12984 col_n[28] a_31478_6508# 0.0283f
C12985 m2_34864_6970# m2_34864_5966# 0.843f
C12986 a_2275_6170# a_32082_6146# 0.399f
C12987 rowoff_n[3] a_34490_5504# 0.0133f
C12988 vcm a_9902_11166# 0.1f
C12989 a_12002_11166# a_12002_10162# 0.843f
C12990 VDD a_5978_1126# 0.035f
C12991 col_n[17] a_2275_15206# 0.113f
C12992 col_n[22] a_2275_4162# 0.113f
C12993 a_5886_15182# a_6282_15222# 0.0313f
C12994 a_2275_15206# a_10906_15182# 0.136f
C12995 VDD a_29470_11528# 0.0779f
C12996 col[11] a_14010_10162# 0.367f
C12997 ctop a_9994_15182# 4.11f
C12998 row_n[4] a_2874_6146# 0.0436f
C12999 col[18] a_20946_12170# 0.0682f
C13000 a_2475_3158# a_24962_3134# 0.264f
C13001 a_2275_3158# a_22346_3174# 0.144f
C13002 rowon_n[8] a_2161_10186# 0.0177f
C13003 rowoff_n[8] a_26058_10162# 0.294f
C13004 col_n[26] a_29070_6146# 0.251f
C13005 col[7] a_2275_12194# 0.0899f
C13006 a_24962_8154# a_25454_8516# 0.0658f
C13007 a_24050_8154# a_24354_8194# 0.0931f
C13008 rowoff_n[11] a_29982_13174# 0.202f
C13009 m2_34864_12994# a_35002_13174# 0.225f
C13010 col[12] a_2275_1150# 0.0899f
C13011 vcm a_24962_15182# 0.1f
C13012 a_2475_12194# a_2874_12170# 0.264f
C13013 a_1957_12194# a_2275_12194# 0.158f
C13014 VDD a_21038_5142# 0.483f
C13015 a_33390_1166# VDD 0.0149f
C13016 col_n[6] a_9294_10202# 0.084f
C13017 row_n[15] a_23350_17230# 0.0117f
C13018 a_2275_17214# a_25966_17190# 0.136f
C13019 VDD a_10394_14540# 0.0779f
C13020 rowoff_n[6] a_35094_8154# 0.0135f
C13021 a_27062_2130# m2_27260_2378# 0.165f
C13022 col[27] a_2475_11190# 0.136f
C13023 row_n[5] a_33390_7190# 0.0117f
C13024 a_20946_5142# a_21038_5142# 0.326f
C13025 m3_32988_1078# m3_33992_1078# 0.202f
C13026 col_n[17] a_20434_4500# 0.0283f
C13027 col_n[27] a_30474_16548# 0.0283f
C13028 rowoff_n[14] a_11398_16548# 0.0133f
C13029 m3_33992_1078# analog_in 0.057f
C13030 vcm a_5886_18194# 0.101f
C13031 a_27062_15182# a_27062_14178# 0.843f
C13032 m3_19936_1078# a_20034_2130# 0.0176f
C13033 a_2475_14202# a_18026_14178# 0.316f
C13034 VDD a_2475_8178# 26.1f
C13035 row_n[7] a_23958_9158# 0.0437f
C13036 rowon_n[11] a_23046_13174# 0.248f
C13037 VDD a_25454_18556# 0.0858f
C13038 a_2275_2154# a_30986_2130# 0.136f
C13039 a_15926_2130# a_16322_2170# 0.0313f
C13040 col[0] a_2874_8154# 0.0682f
C13041 m3_8892_18146# VDD 0.0277f
C13042 vcm a_7986_3134# 0.56f
C13043 rowon_n[1] a_33086_3134# 0.248f
C13044 col[7] a_9902_10162# 0.0682f
C13045 col[24] a_2275_14202# 0.0899f
C13046 col_n[15] a_18026_4138# 0.251f
C13047 a_5886_11166# a_6378_11528# 0.0658f
C13048 a_2275_11190# a_8990_11166# 0.399f
C13049 m2_28840_946# col[26] 0.425f
C13050 a_4974_11166# a_5278_11206# 0.0931f
C13051 col[29] a_2275_3158# 0.0899f
C13052 m2_16792_18014# a_16930_18194# 0.225f
C13053 col_n[25] a_28066_16186# 0.251f
C13054 col_n[22] a_24962_6146# 0.0765f
C13055 a_17022_16186# a_18026_16186# 0.843f
C13056 a_2475_16210# a_33086_16186# 0.316f
C13057 VDD a_17022_12170# 0.483f
C13058 m2_2736_18014# m3_1864_18146# 0.0341f
C13059 m2_6176_10410# rowon_n[8] 0.0322f
C13060 m2_12200_6394# rowon_n[4] 0.0322f
C13061 m2_17220_2378# rowon_n[0] 0.0322f
C13062 row_n[1] a_10998_3134# 0.282f
C13063 a_22346_1166# col_n[19] 0.0839f
C13064 rowon_n[5] a_10906_7150# 0.118f
C13065 vcm a_23046_7150# 0.56f
C13066 rowoff_n[12] a_17934_14178# 0.202f
C13067 m2_32280_14426# a_32082_14178# 0.165f
C13068 col_n[6] a_9390_2492# 0.0283f
C13069 a_2275_13198# a_24050_13174# 0.399f
C13070 col_n[16] a_19430_14540# 0.0283f
C13071 rowon_n[10] col[12] 0.0323f
C13072 rowon_n[4] col[0] 0.0318f
C13073 row_n[12] col[15] 0.0342f
C13074 col_n[27] col[27] 0.536f
C13075 rowon_n[9] col[10] 0.0323f
C13076 rowon_n[1] ctop 0.203f
C13077 row_n[14] col[19] 0.0342f
C13078 col_n[14] a_2475_10186# 0.0531f
C13079 row_n[8] col[7] 0.0342f
C13080 rowon_n[12] col[16] 0.0323f
C13081 rowon_n[5] col[2] 0.0323f
C13082 rowon_n[15] col[22] 0.0323f
C13083 row_n[15] col[21] 0.0342f
C13084 rowon_n[14] col[20] 0.0323f
C13085 row_n[5] col[1] 0.0342f
C13086 rowon_n[6] col[4] 0.0323f
C13087 rowon_n[7] col[6] 0.0323f
C13088 row_n[10] col[11] 0.0342f
C13089 row_n[9] col[9] 0.0342f
C13090 rowon_n[8] col[8] 0.0323f
C13091 row_n[6] col[3] 0.0342f
C13092 rowon_n[13] col[18] 0.0323f
C13093 row_n[7] col[5] 0.0342f
C13094 col_n[21] rowoff_n[15] 0.0471f
C13095 row_n[13] col[17] 0.0342f
C13096 rowon_n[11] col[14] 0.0323f
C13097 row_n[11] col[13] 0.0342f
C13098 VDD a_32082_16186# 0.483f
C13099 row_n[12] a_31382_14218# 0.0117f
C13100 col[24] rowoff_n[11] 0.0901f
C13101 vcm a_13310_1166# 0.16f
C13102 m2_27260_15430# rowon_n[13] 0.0322f
C13103 a_30986_6146# a_31382_6186# 0.0313f
C13104 m2_33284_11414# rowon_n[9] 0.0322f
C13105 m2_4744_946# m3_5880_1078# 0.0341f
C13106 vcm a_3970_10162# 0.56f
C13107 a_2475_10186# a_16930_10162# 0.264f
C13108 a_2275_10186# a_14314_10202# 0.144f
C13109 row_n[14] a_21950_16186# 0.0437f
C13110 col[4] a_2475_7174# 0.136f
C13111 m2_4168_16434# a_3970_16186# 0.165f
C13112 a_20946_15182# a_21438_15544# 0.0658f
C13113 a_20034_15182# a_20338_15222# 0.0931f
C13114 col_n[4] a_6982_2130# 0.251f
C13115 col_n[30] a_33390_3174# 0.084f
C13116 col_n[14] a_17022_14178# 0.251f
C13117 row_n[4] a_31990_6146# 0.0437f
C13118 col_n[11] a_13918_4138# 0.0765f
C13119 a_27062_3134# a_28066_3134# 0.843f
C13120 rowon_n[8] a_31078_10162# 0.248f
C13121 col_n[21] a_23958_16186# 0.0765f
C13122 m2_34864_4962# a_35398_5182# 0.087f
C13123 col_n[11] a_2275_13198# 0.113f
C13124 vcm a_28370_5182# 0.155f
C13125 a_2275_7174# a_7894_7150# 0.136f
C13126 col_n[16] a_2275_2154# 0.113f
C13127 m2_17796_18014# vcm 0.353f
C13128 m2_23244_12418# a_23046_12170# 0.165f
C13129 vcm a_19030_14178# 0.56f
C13130 a_2475_12194# a_31990_12170# 0.264f
C13131 a_2275_12194# a_29374_12210# 0.144f
C13132 a_16930_12170# a_17022_12170# 0.326f
C13133 VDD a_15926_4138# 0.181f
C13134 row_n[0] m2_33284_2378# 0.0128f
C13135 col_n[31] a_2475_12194# 0.0531f
C13136 col_n[5] a_8386_12532# 0.0283f
C13137 row_n[8] a_8990_10162# 0.282f
C13138 col[8] rowoff_n[12] 0.0901f
C13139 col[1] a_2275_10186# 0.0899f
C13140 rowon_n[12] a_8898_14178# 0.118f
C13141 a_18026_5142# a_18026_4138# 0.843f
C13142 m2_27836_946# ctop 0.0428f
C13143 col[31] a_33998_3134# 0.0682f
C13144 m2_27836_18014# m2_28840_18014# 0.843f
C13145 vcm a_9294_8194# 0.155f
C13146 a_2275_9182# a_22954_9158# 0.136f
C13147 rowoff_n[13] a_5886_15182# 0.202f
C13148 a_11910_9158# a_12306_9198# 0.0313f
C13149 rowon_n[2] a_18938_4138# 0.118f
C13150 ctop a_22042_3134# 4.11f
C13151 vcm a_34090_18194# 0.165f
C13152 col[21] a_2475_9182# 0.136f
C13153 VDD a_30986_8154# 0.181f
C13154 rowoff_n[5] a_7894_7150# 0.202f
C13155 row_n[0] a_6282_2170# 0.0117f
C13156 a_30074_2130# a_30378_2170# 0.0931f
C13157 a_30986_2130# a_31478_2492# 0.0658f
C13158 col_n[29] a_32386_13214# 0.084f
C13159 col_n[3] a_5978_12170# 0.251f
C13160 vcm a_2161_2154# 0.0169f
C13161 a_2475_6170# a_15014_6146# 0.316f
C13162 a_7986_6146# a_8990_6146# 0.843f
C13163 col_n[28] a_2275_15206# 0.113f
C13164 m2_14208_10410# a_14010_10162# 0.165f
C13165 col_n[10] a_12914_14178# 0.0765f
C13166 rowoff_n[3] a_16930_5142# 0.202f
C13167 vcm a_24354_12210# 0.155f
C13168 VDD a_22442_2492# 0.0779f
C13169 m2_12776_18014# a_13006_17190# 0.843f
C13170 m2_5172_9406# row_n[7] 0.0128f
C13171 m2_11196_5390# row_n[3] 0.0128f
C13172 a_31990_16186# a_32082_16186# 0.326f
C13173 row_n[11] a_29982_13174# 0.0437f
C13174 VDD a_11910_11166# 0.181f
C13175 rowon_n[15] a_29070_17190# 0.248f
C13176 col[18] a_2275_12194# 0.0899f
C13177 a_2275_3158# a_5978_3134# 0.399f
C13178 rowoff_n[8] a_8386_10524# 0.0133f
C13179 rowoff_n[1] a_25966_3134# 0.202f
C13180 m2_33284_6394# a_33086_6146# 0.165f
C13181 col[23] a_2275_1150# 0.0899f
C13182 vcm a_17934_6146# 0.1f
C13183 a_33086_9158# a_33086_8154# 0.843f
C13184 a_2475_8178# a_30074_8154# 0.316f
C13185 col_n[1] a_3878_12170# 0.0765f
C13186 col[23] a_26058_11166# 0.367f
C13187 col[20] a_22954_1126# 0.0682f
C13188 vcm a_5278_15222# 0.155f
C13189 a_26970_13174# a_27366_13214# 0.0313f
C13190 VDD a_2966_5142# 0.485f
C13191 m2_1732_2954# ctop 0.0424f
C13192 col[30] a_32994_13174# 0.0682f
C13193 ctop a_18026_10162# 4.11f
C13194 row_n[15] a_6982_17190# 0.282f
C13195 m2_26256_14426# row_n[12] 0.0128f
C13196 a_2275_17214# a_6282_17230# 0.144f
C13197 a_2475_17214# a_8898_17190# 0.264f
C13198 rowoff_n[6] a_17422_8516# 0.0133f
C13199 VDD a_26970_15182# 0.181f
C13200 m2_32280_10410# row_n[8] 0.0128f
C13201 row_n[5] a_17022_7150# 0.282f
C13202 a_11910_5142# a_12402_5504# 0.0658f
C13203 a_2275_5166# a_21038_5142# 0.399f
C13204 a_10998_5142# a_11302_5182# 0.0931f
C13205 m3_1864_3086# m3_1864_2082# 0.202f
C13206 m2_5172_8402# a_4974_8154# 0.165f
C13207 rowon_n[9] a_16930_11166# 0.118f
C13208 col_n[18] a_21342_11206# 0.084f
C13209 vcm a_32994_10162# 0.1f
C13210 col_n[8] a_2475_8178# 0.0531f
C13211 a_23046_10162# a_24050_10162# 0.843f
C13212 rowoff_n[4] a_26458_6508# 0.0133f
C13213 m2_7756_946# a_2275_1150# 0.28f
C13214 a_35002_15182# a_35398_15222# 0.0313f
C13215 VDD a_18426_9520# 0.0779f
C13216 row_n[7] a_4274_9198# 0.0117f
C13217 ctop a_33086_14178# 4.11f
C13218 col_n[29] a_32482_5504# 0.0283f
C13219 VDD a_7894_18194# 0.343f
C13220 a_7894_2130# a_7986_2130# 0.326f
C13221 a_2475_2154# a_13918_2130# 0.264f
C13222 a_2275_2154# a_11302_2170# 0.144f
C13223 m2_24248_4386# a_24050_4138# 0.165f
C13224 rowoff_n[9] a_18026_11166# 0.294f
C13225 rowoff_n[2] a_35494_4500# 0.0133f
C13226 vcm a_13918_13174# 0.1f
C13227 a_14010_12170# a_14010_11166# 0.843f
C13228 VDD a_9994_3134# 0.483f
C13229 m2_8760_18014# a_2275_18218# 0.28f
C13230 col[12] a_15014_9158# 0.367f
C13231 a_7894_16186# a_8290_16226# 0.0313f
C13232 a_2275_16210# a_14922_16186# 0.136f
C13233 VDD a_33486_13536# 0.0779f
C13234 rowon_n[3] a_3970_5142# 0.248f
C13235 col_n[5] a_2275_11190# 0.113f
C13236 a_24050_1126# m2_23820_946# 0.0249f
C13237 col[19] a_21950_11166# 0.0682f
C13238 ctop a_14010_17190# 4.06f
C13239 rowoff_n[7] a_27062_9158# 0.294f
C13240 a_2475_4162# a_28978_4138# 0.264f
C13241 col_n[27] a_30074_5142# 0.251f
C13242 a_2275_4162# a_26362_4178# 0.144f
C13243 m3_32988_1078# ctop 0.21f
C13244 a_26058_9158# a_26362_9198# 0.0931f
C13245 a_26970_9158# a_27462_9520# 0.0658f
C13246 rowoff_n[13] a_34090_15182# 0.294f
C13247 rowon_n[3] col[9] 0.0323f
C13248 rowon_n[7] col[17] 0.0323f
C13249 rowon_n[5] col[13] 0.0323f
C13250 row_n[10] col[22] 0.0342f
C13251 row_n[13] col[28] 0.0342f
C13252 rowon_n[11] col[25] 0.0323f
C13253 rowon_n[4] col[11] 0.0323f
C13254 row_n[9] col[20] 0.0342f
C13255 col_n[25] a_2475_10186# 0.0531f
C13256 row_n[5] col[12] 0.0342f
C13257 rowon_n[8] col[19] 0.0323f
C13258 row_n[15] sample_n 0.0596f
C13259 rowon_n[12] col[27] 0.0323f
C13260 row_n[12] col[26] 0.0342f
C13261 rowon_n[2] col[7] 0.0323f
C13262 row_n[0] col[2] 0.0342f
C13263 row_n[1] col[4] 0.0342f
C13264 rowon_n[6] col[15] 0.0323f
C13265 rowon_n[0] col[3] 0.0323f
C13266 row_n[8] col[18] 0.0342f
C13267 row_n[3] col[8] 0.0342f
C13268 row_n[4] col[10] 0.0342f
C13269 row_n[6] col[14] 0.0342f
C13270 row_n[7] col[16] 0.0342f
C13271 rowon_n[9] col[21] 0.0323f
C13272 rowon_n[14] col[31] 0.0323f
C13273 row_n[14] col[30] 0.0342f
C13274 rowon_n[15] rowoff_n[15] 20.2f
C13275 rowon_n[1] col[5] 0.0323f
C13276 row_n[2] col[6] 0.0342f
C13277 row_n[11] col[24] 0.0342f
C13278 rowon_n[13] col[29] 0.0323f
C13279 rowon_n[10] col[23] 0.0323f
C13280 ctop analog_in 0.885f
C13281 col_n[7] a_10298_9198# 0.084f
C13282 vcm a_28978_17190# 0.1f
C13283 a_2475_13198# a_6982_13174# 0.316f
C13284 a_3970_13174# a_4974_13174# 0.843f
C13285 VDD a_25054_7150# 0.483f
C13286 m2_4744_18014# a_2475_18218# 0.286f
C13287 a_2275_18218# a_29982_18194# 0.136f
C13288 VDD a_14410_16548# 0.0779f
C13289 a_2275_1150# a_19942_1126# 0.106f
C13290 row_n[12] a_15014_14178# 0.282f
C13291 col_n[18] a_21438_3496# 0.0283f
C13292 vcm a_31078_2130# 0.56f
C13293 a_22954_6146# a_23046_6146# 0.326f
C13294 col[15] a_2475_7174# 0.136f
C13295 col_n[28] a_31478_15544# 0.0283f
C13296 m2_20808_946# m2_21236_1374# 0.165f
C13297 m2_1732_8978# a_2275_9182# 0.191f
C13298 row_n[2] a_25054_4138# 0.282f
C13299 VDD a_15318_1166# 0.0149f
C13300 row_n[14] a_3878_16186# 0.0437f
C13301 m2_31852_18014# a_32082_17190# 0.843f
C13302 rowon_n[6] a_24962_8154# 0.118f
C13303 a_29070_16186# a_29070_15182# 0.843f
C13304 a_2475_15206# a_22042_15182# 0.316f
C13305 VDD a_5978_10162# 0.483f
C13306 col[1] a_3970_7150# 0.367f
C13307 row_n[4] a_12306_6186# 0.0117f
C13308 col_n[22] a_2275_13198# 0.113f
C13309 a_2275_3158# a_35002_3134# 0.136f
C13310 a_2475_18218# a_27974_18194# 0.264f
C13311 a_17934_3134# a_18330_3174# 0.0313f
C13312 col_n[27] a_2275_2154# 0.113f
C13313 col[8] a_10906_9158# 0.0682f
C13314 vcm a_12002_5142# 0.56f
C13315 rowoff_n[10] a_5978_12170# 0.294f
C13316 col_n[16] a_19030_3134# 0.251f
C13317 a_25966_1126# vcm 0.0989f
C13318 row_n[6] a_2161_8178# 0.0221f
C13319 col_n[26] a_29070_15182# 0.251f
C13320 m2_1732_3958# rowon_n[2] 0.236f
C13321 a_7894_12170# a_8386_12532# 0.0658f
C13322 a_6982_12170# a_7286_12210# 0.0931f
C13323 a_2275_12194# a_13006_12170# 0.399f
C13324 col_n[23] a_25966_5142# 0.0765f
C13325 rowon_n[10] a_2475_12194# 0.31f
C13326 m2_21812_18014# VDD 1f
C13327 col[12] a_2275_10186# 0.0899f
C13328 col[19] rowoff_n[12] 0.0901f
C13329 row_n[15] a_34394_17230# 0.0117f
C13330 a_19030_17190# a_20034_17190# 0.843f
C13331 VDD a_21038_14178# 0.483f
C13332 a_35398_2170# m2_34864_1950# 0.087f
C13333 rowon_n[0] a_12002_2130# 0.248f
C13334 vcm a_27062_9158# 0.56f
C13335 col_n[7] a_10394_1488# 0.0283f
C13336 a_2275_9182# a_3270_9198# 0.144f
C13337 a_2475_9182# a_5886_9158# 0.264f
C13338 rowoff_n[14] a_22042_16186# 0.294f
C13339 col_n[17] a_20434_13536# 0.0283f
C13340 m2_10192_17438# rowon_n[15] 0.0322f
C13341 a_2275_14202# a_28066_14178# 0.399f
C13342 m2_16216_13422# rowon_n[11] 0.0322f
C13343 m2_22240_9406# rowon_n[7] 0.0322f
C13344 m2_28264_5390# rowon_n[3] 0.0322f
C13345 VDD a_2475_17214# 26.1f
C13346 col_n[2] a_2475_6170# 0.0531f
C13347 row_n[9] a_23046_11166# 0.282f
C13348 vcm a_17326_3174# 0.155f
C13349 a_32994_7150# a_33390_7190# 0.0313f
C13350 col[0] a_2874_17190# 0.0682f
C13351 m2_34864_10986# a_34090_11166# 0.843f
C13352 rowon_n[13] a_22954_15182# 0.118f
C13353 vcm a_7986_12170# 0.56f
C13354 a_2275_11190# a_18330_11206# 0.144f
C13355 a_2475_11190# a_20946_11166# 0.264f
C13356 col[3] rowoff_n[13] 0.0901f
C13357 VDD a_4882_2130# 0.181f
C13358 col_n[15] a_18026_13174# 0.251f
C13359 row_n[11] a_10298_13214# 0.0117f
C13360 a_22042_16186# a_22346_16226# 0.0931f
C13361 a_22954_16186# a_23446_16548# 0.0658f
C13362 rowon_n[3] a_32994_5142# 0.118f
C13363 col[29] a_2275_12194# 0.0899f
C13364 col_n[12] a_14922_3134# 0.0765f
C13365 m2_16792_18014# m3_16924_18146# 3.79f
C13366 col_n[22] a_24962_15182# 0.0765f
C13367 a_29070_4138# a_30074_4138# 0.843f
C13368 row_n[1] a_20338_3174# 0.0117f
C13369 vcm a_32386_7190# 0.155f
C13370 rowoff_n[12] a_28466_14540# 0.0133f
C13371 a_2275_8178# a_11910_8154# 0.136f
C13372 col_n[0] a_2275_9182# 0.113f
C13373 vcm a_23046_16186# 0.56f
C13374 a_2275_13198# a_33390_13214# 0.144f
C13375 a_18938_13174# a_19030_13174# 0.326f
C13376 VDD a_19942_6146# 0.181f
C13377 row_n[3] a_10906_5142# 0.0437f
C13378 col_n[6] a_9390_11528# 0.0283f
C13379 rowon_n[7] a_9994_9158# 0.248f
C13380 col_n[19] a_2475_8178# 0.0531f
C13381 a_2475_5166# a_3970_5142# 0.316f
C13382 a_20034_6146# a_20034_5142# 0.843f
C13383 a_2275_5166# a_2966_5142# 0.399f
C13384 m3_28972_18146# m3_29976_18146# 0.202f
C13385 m2_20808_946# m3_19936_1078# 0.0341f
C13386 vcm a_13310_10202# 0.155f
C13387 rowoff_n[15] a_9994_17190# 0.294f
C13388 a_2275_10186# a_26970_10162# 0.136f
C13389 a_13918_10162# a_14314_10202# 0.0313f
C13390 rowoff_n[4] a_8898_6146# 0.202f
C13391 ctop a_26058_5142# 4.11f
C13392 VDD a_35002_10162# 0.258f
C13393 col[4] a_2475_16210# 0.136f
C13394 col[9] a_2475_5166# 0.136f
C13395 col_n[30] a_33390_12210# 0.084f
C13396 col_n[4] a_6982_11166# 0.251f
C13397 a_32994_3134# a_33486_3496# 0.0658f
C13398 a_32082_3134# a_32386_3174# 0.0931f
C13399 col_n[11] a_13918_13174# 0.0765f
C13400 vcm a_6890_4138# 0.1f
C13401 rowoff_n[2] a_17934_4138# 0.202f
C13402 a_9994_7150# a_10998_7150# 0.843f
C13403 rowoff_n[10] a_35002_12170# 0.202f
C13404 a_2475_7174# a_19030_7150# 0.316f
C13405 row_n[6] a_31078_8154# 0.282f
C13406 vcm a_28370_14218# 0.155f
C13407 col_n[16] a_2275_11190# 0.113f
C13408 rowon_n[10] a_30986_12170# 0.118f
C13409 VDD a_26458_4500# 0.0779f
C13410 ctop a_6982_8154# 4.11f
C13411 a_33998_17190# a_34090_17190# 0.326f
C13412 VDD a_15926_13174# 0.181f
C13413 row_n[8] a_18330_10202# 0.0117f
C13414 rowoff_n[7] a_9390_9520# 0.0133f
C13415 rowoff_n[0] a_26970_2130# 0.202f
C13416 a_2275_4162# a_9994_4138# 0.399f
C13417 m3_28972_18146# ctop 0.209f
C13418 rowon_n[5] col[24] 0.0323f
C13419 rowon_n[6] col[26] 0.0323f
C13420 rowon_n[2] col[18] 0.0323f
C13421 row_n[7] col[27] 0.0342f
C13422 row_n[6] col[25] 0.0342f
C13423 row_n[4] col[21] 0.0342f
C13424 row_n[5] col[23] 0.0342f
C13425 row_n[2] col[17] 0.0342f
C13426 rowon_n[7] col[28] 0.0323f
C13427 row_n[9] col[31] 0.0342f
C13428 row_n[0] col[13] 0.0342f
C13429 row_n[3] col[19] 0.0342f
C13430 rowon_n[3] col[20] 0.0323f
C13431 row_n[1] col[15] 0.0342f
C13432 rowon_n[0] col[14] 0.0323f
C13433 rowon_n[9] sample_n 0.0692f
C13434 ctop col[10] 0.123f
C13435 rowon_n[1] col[16] 0.0323f
C13436 row_n[8] col[29] 0.0342f
C13437 rowon_n[4] col[22] 0.0323f
C13438 rowon_n[8] col[30] 0.0323f
C13439 m2_9188_16434# row_n[14] 0.0128f
C13440 col[24] a_27062_10162# 0.367f
C13441 vcm a_21950_8154# 0.1f
C13442 col[6] a_2275_8178# 0.0899f
C13443 m2_15212_12418# row_n[10] 0.0128f
C13444 a_2475_9182# a_34090_9158# 0.316f
C13445 rowoff_n[13] a_16418_15544# 0.0133f
C13446 m2_21236_8402# row_n[6] 0.0128f
C13447 m2_27260_4386# row_n[2] 0.0128f
C13448 row_n[10] a_8898_12170# 0.0437f
C13449 col[31] a_33998_12170# 0.0682f
C13450 vcm a_9294_17230# 0.155f
C13451 rowon_n[14] a_7986_16186# 0.248f
C13452 a_28978_14178# a_29374_14218# 0.0313f
C13453 VDD a_7382_7512# 0.0779f
C13454 rowoff_n[5] a_18426_7512# 0.0133f
C13455 ctop a_22042_12170# 4.11f
C13456 a_2275_18218# a_10298_18234# 0.145f
C13457 row_n[0] a_18938_2130# 0.0437f
C13458 VDD a_30986_17190# 0.181f
C13459 col[26] a_2475_7174# 0.136f
C13460 rowon_n[4] a_18026_6146# 0.248f
C13461 col_n[19] a_22346_10202# 0.084f
C13462 a_13006_6146# a_13310_6186# 0.0931f
C13463 a_2275_6170# a_25054_6146# 0.399f
C13464 a_13918_6146# a_14410_6508# 0.0658f
C13465 rowoff_n[3] a_27462_5504# 0.0133f
C13466 vcm a_2161_11190# 0.0169f
C13467 a_25054_11166# a_26058_11166# 0.843f
C13468 m2_35292_17438# row_n[15] 0.0128f
C13469 VDD a_33086_2130# 0.483f
C13470 m2_10192_17438# a_9994_17190# 0.165f
C13471 a_2874_15182# a_2966_15182# 0.326f
C13472 col_n[30] a_33486_4500# 0.0283f
C13473 VDD a_22442_11528# 0.0779f
C13474 a_2275_3158# a_15318_3174# 0.144f
C13475 a_9902_3134# a_9994_3134# 0.326f
C13476 a_2475_3158# a_17934_3134# 0.264f
C13477 rowoff_n[8] a_19030_10162# 0.294f
C13478 a_31078_1126# a_2475_1150# 0.0299f
C13479 row_n[13] a_29070_15182# 0.282f
C13480 rowoff_n[11] a_22954_13174# 0.202f
C13481 col[23] a_2275_10186# 0.0899f
C13482 col[30] rowoff_n[12] 0.0901f
C13483 m2_29268_13422# a_29070_13174# 0.165f
C13484 col[13] a_16018_8154# 0.367f
C13485 vcm a_17934_15182# 0.1f
C13486 a_16018_13174# a_16018_12170# 0.843f
C13487 VDD a_14010_5142# 0.483f
C13488 a_27974_1126# VDD 0.405f
C13489 row_n[15] a_16322_17230# 0.0117f
C13490 col[20] a_22954_10162# 0.0682f
C13491 a_2275_17214# a_18938_17190# 0.136f
C13492 a_9902_17190# a_10298_17230# 0.0313f
C13493 rowoff_n[6] a_28066_8154# 0.294f
C13494 VDD a_2966_14178# 0.485f
C13495 col_n[28] a_31078_4138# 0.251f
C13496 a_2475_5166# a_32994_5142# 0.264f
C13497 row_n[5] a_26362_7190# 0.0117f
C13498 a_2275_5166# a_30378_5182# 0.144f
C13499 m3_18932_1078# m3_19936_1078# 0.116f
C13500 a_30986_1126# a_31078_1126# 0.0991f
C13501 col_n[8] a_11302_8194# 0.084f
C13502 rowoff_n[14] a_4370_16548# 0.0133f
C13503 a_28978_10162# a_29470_10524# 0.0658f
C13504 a_28066_10162# a_28370_10202# 0.0931f
C13505 m2_30848_946# a_2275_1150# 0.28f
C13506 col_n[8] a_2475_17214# 0.0531f
C13507 m2_11772_946# a_11910_1126# 0.225f
C13508 a_2475_14202# a_10998_14178# 0.316f
C13509 a_5978_14178# a_6982_14178# 0.843f
C13510 VDD a_29070_9158# 0.483f
C13511 row_n[7] a_16930_9158# 0.0437f
C13512 col_n[13] a_2475_6170# 0.0531f
C13513 rowon_n[11] a_16018_13174# 0.248f
C13514 VDD a_18426_18556# 0.0858f
C13515 col_n[19] a_22442_2492# 0.0283f
C13516 a_2275_2154# a_23958_2130# 0.136f
C13517 col_n[29] a_32482_14540# 0.0283f
C13518 m2_25252_1374# VDD 0.0194f
C13519 vcm a_35094_4138# 0.165f
C13520 a_24962_7150# a_25054_7150# 0.326f
C13521 col[14] rowoff_n[13] 0.0901f
C13522 rowon_n[1] a_26058_3134# 0.248f
C13523 m2_20232_11414# a_20034_11166# 0.165f
C13524 a_1957_11190# a_2161_11190# 0.115f
C13525 a_2475_11190# a_2275_11190# 2.76f
C13526 col[3] a_2475_3158# 0.136f
C13527 VDD rowoff_n[9] 1.51f
C13528 m2_11772_18014# a_12002_18194# 0.0249f
C13529 col[2] a_4974_6146# 0.367f
C13530 a_2475_16210# a_26058_16186# 0.316f
C13531 a_31078_17190# a_31078_16186# 0.843f
C13532 VDD a_9994_12170# 0.483f
C13533 a_30378_1166# m2_29844_946# 0.087f
C13534 a_33390_1166# col_n[30] 0.084f
C13535 col[9] a_11910_8154# 0.0682f
C13536 a_19942_4138# a_20338_4178# 0.0313f
C13537 row_n[1] a_3970_3134# 0.282f
C13538 col_n[10] a_2275_9182# 0.113f
C13539 col_n[17] a_20034_2130# 0.25f
C13540 vcm a_16018_7150# 0.56f
C13541 col_n[27] a_30074_14178# 0.251f
C13542 rowoff_n[12] a_10906_14178# 0.202f
C13543 col_n[24] a_26970_4138# 0.0765f
C13544 a_8990_13174# a_9294_13214# 0.0931f
C13545 a_2275_13198# a_17022_13174# 0.399f
C13546 a_9902_13174# a_10394_13536# 0.0658f
C13547 VDD a_35398_7190# 0.0882f
C13548 col_n[7] a_10298_18234# 0.084f
C13549 col_n[30] a_2475_8178# 0.0531f
C13550 VDD a_25054_16186# 0.483f
C13551 col[0] a_2275_6170# 0.099f
C13552 row_n[12] a_24354_14218# 0.0117f
C13553 vcm a_6282_1166# 0.16f
C13554 m2_5172_11414# rowon_n[9] 0.0322f
C13555 m2_11196_7398# rowon_n[5] 0.0322f
C13556 m2_11196_9406# a_10998_9158# 0.165f
C13557 m2_17220_3382# rowon_n[1] 0.0322f
C13558 m2_12776_946# col[10] 0.425f
C13559 col_n[18] a_21438_12532# 0.0283f
C13560 row_n[2] a_35398_4178# 0.0117f
C13561 vcm a_31078_11166# 0.56f
C13562 a_2475_10186# a_9902_10162# 0.264f
C13563 a_5886_10162# a_5978_10162# 0.326f
C13564 a_2275_10186# a_7286_10202# 0.144f
C13565 col[15] a_2475_16210# 0.136f
C13566 row_n[14] a_14922_16186# 0.0437f
C13567 col[20] a_2475_5166# 0.136f
C13568 a_2275_15206# a_32082_15182# 0.399f
C13569 row_n[4] a_24962_6146# 0.0437f
C13570 rowon_n[8] a_24050_10162# 0.248f
C13571 a_6982_3134# a_6982_2130# 0.843f
C13572 col[1] a_3970_16186# 0.367f
C13573 m2_30272_5390# a_30074_5142# 0.165f
C13574 vcm a_21342_5182# 0.155f
C13575 col_n[27] a_2275_11190# 0.113f
C13576 col[8] a_10906_18194# 0.0682f
C13577 m2_3740_18014# vcm 0.353f
C13578 m2_26256_16434# rowon_n[14] 0.0322f
C13579 m2_32280_12418# rowon_n[10] 0.0322f
C13580 vcm a_12002_14178# 0.56f
C13581 a_2275_12194# a_22346_12210# 0.144f
C13582 a_2475_12194# a_24962_12170# 0.264f
C13583 col_n[16] a_19030_12170# 0.251f
C13584 VDD a_8898_4138# 0.181f
C13585 col_n[13] a_15926_2130# 0.0765f
C13586 m2_5748_18014# col[3] 0.347f
C13587 a_24962_17190# a_25454_17552# 0.0658f
C13588 a_24050_17190# a_24354_17230# 0.0931f
C13589 col_n[23] a_25966_14178# 0.0765f
C13590 VDD sample 4.82f
C13591 row_n[4] sample_n 0.0596f
C13592 row_n[8] a_2475_10186# 0.405f
C13593 rowon_n[1] col[27] 0.0323f
C13594 row_n[1] col[26] 0.0342f
C13595 rowon_n[0] col[25] 0.0323f
C13596 row_n[3] col[30] 0.0342f
C13597 row_n[0] col[24] 0.0342f
C13598 en_bit_n[0] col[17] 0.142f
C13599 ctop col[21] 0.123f
C13600 rowon_n[2] col[29] 0.0323f
C13601 row_n[2] col[28] 0.0342f
C13602 rowon_n[3] col[31] 0.0323f
C13603 col[7] col[8] 0.0355f
C13604 col[17] a_2275_8178# 0.0899f
C13605 a_31078_5142# a_32082_5142# 0.843f
C13606 m2_1732_6970# a_1957_7174# 0.245f
C13607 m2_20808_18014# m2_21812_18014# 0.843f
C13608 vcm a_3878_8154# 0.1f
C13609 a_2275_9182# a_15926_9158# 0.136f
C13610 rowon_n[2] a_11910_4138# 0.118f
C13611 col_n[7] a_10394_10524# 0.0283f
C13612 ctop a_15014_3134# 4.11f
C13613 vcm a_27062_18194# 0.165f
C13614 a_20946_14178# a_21038_14178# 0.326f
C13615 VDD a_23958_8154# 0.181f
C13616 m2_21236_3382# a_21038_3134# 0.165f
C13617 m3_27968_1078# VDD 0.0157f
C13618 vcm a_29982_3134# 0.1f
C13619 row_n[9] a_32386_11206# 0.0117f
C13620 a_2475_6170# a_7986_6146# 0.316f
C13621 a_22042_7150# a_22042_6146# 0.843f
C13622 col_n[2] a_2475_15206# 0.0531f
C13623 col_n[7] a_2475_4162# 0.0531f
C13624 rowoff_n[3] a_9902_5142# 0.202f
C13625 vcm a_17326_12210# 0.155f
C13626 a_2275_11190# a_30986_11166# 0.136f
C13627 a_15926_11166# a_16322_11206# 0.0313f
C13628 VDD a_15414_2492# 0.0779f
C13629 m2_30848_18014# a_31078_18194# 0.0249f
C13630 ctop a_30074_7150# 4.11f
C13631 row_n[11] a_22954_13174# 0.0437f
C13632 VDD a_4882_11166# 0.181f
C13633 m2_30848_18014# m3_31984_18146# 0.0341f
C13634 col_n[5] a_7986_10162# 0.251f
C13635 rowon_n[15] a_22042_17190# 0.248f
C13636 col_n[12] a_14922_12170# 0.0765f
C13637 a_35002_4138# a_35494_4500# 0.0658f
C13638 rowoff_n[1] a_18938_3134# 0.202f
C13639 row_n[1] a_32994_3134# 0.0437f
C13640 m2_21812_18014# col_n[19] 0.243f
C13641 en_bit_n[2] a_2475_1150# 0.0162f
C13642 vcm a_10906_6146# 0.1f
C13643 rowon_n[5] a_32082_7150# 0.248f
C13644 a_12002_8154# a_13006_8154# 0.843f
C13645 a_2475_8178# a_23046_8154# 0.316f
C13646 vcm a_32386_16226# 0.155f
C13647 VDD a_30474_6508# 0.0779f
C13648 col_n[0] a_2275_18218# 0.113f
C13649 ctop a_10998_10162# 4.11f
C13650 VDD a_19942_15182# 0.181f
C13651 col_n[4] a_2275_7174# 0.113f
C13652 rowoff_n[6] a_10394_8516# 0.0133f
C13653 m2_4168_10410# row_n[8] 0.0128f
C13654 m2_10192_6394# row_n[4] 0.0128f
C13655 m2_15212_2378# row_n[0] 0.0128f
C13656 col[25] a_28066_9158# 0.367f
C13657 a_2275_5166# a_14010_5142# 0.399f
C13658 row_n[5] a_9994_7150# 0.282f
C13659 m2_34864_946# m3_34996_1078# 3.79f
C13660 m3_1864_10114# m3_1864_9110# 0.202f
C13661 rowon_n[9] a_9902_11166# 0.118f
C13662 vcm a_25966_10162# 0.1f
C13663 col_n[19] a_2475_17214# 0.0531f
C13664 col_n[24] a_2475_6170# 0.0531f
C13665 rowoff_n[4] a_19430_6508# 0.0133f
C13666 ctop a_2275_4162# 0.0683f
C13667 m2_22816_946# a_23046_2130# 0.843f
C13668 a_30986_15182# a_31382_15222# 0.0313f
C13669 VDD a_11398_9520# 0.0779f
C13670 m2_31852_18014# ctop 0.0422f
C13671 ctop a_26058_14178# 4.11f
C13672 col[25] rowoff_n[13] 0.0901f
C13673 a_2275_2154# a_4274_2170# 0.144f
C13674 a_2475_2154# a_6890_2130# 0.264f
C13675 col_n[20] a_23350_9198# 0.084f
C13676 m2_25252_15430# row_n[13] 0.0128f
C13677 m2_31276_11414# row_n[9] 0.0128f
C13678 col[9] a_2475_14202# 0.136f
C13679 m2_1732_9982# m2_1732_8978# 0.843f
C13680 col[14] a_2475_3158# 0.136f
C13681 rowoff_n[2] a_28466_4500# 0.0133f
C13682 a_15014_7150# a_15318_7190# 0.0931f
C13683 col_n[4] rowoff_n[5] 0.0471f
C13684 col_n[7] rowoff_n[8] 0.0471f
C13685 col_n[5] rowoff_n[6] 0.0471f
C13686 rowoff_n[9] a_10998_11166# 0.294f
C13687 a_2275_7174# a_29070_7150# 0.399f
C13688 a_15926_7150# a_16418_7512# 0.0658f
C13689 vcm rowoff_n[1] 0.533f
C13690 col_n[3] rowoff_n[4] 0.0471f
C13691 col_n[8] rowoff_n[9] 0.0471f
C13692 col_n[6] rowoff_n[7] 0.0471f
C13693 col_n[1] rowoff_n[2] 0.0471f
C13694 col_n[2] rowoff_n[3] 0.0471f
C13695 col_n[0] rowoff_n[0] 0.0471f
C13696 vcm a_6890_13174# 0.1f
C13697 a_27062_12170# a_28066_12170# 0.843f
C13698 VDD a_2874_3134# 0.182f
C13699 col_n[31] a_34490_3496# 0.0283f
C13700 a_2275_16210# a_7894_16186# 0.136f
C13701 VDD a_26458_13536# 0.0779f
C13702 col_n[21] a_2275_9182# 0.113f
C13703 ctop a_6982_17190# 4.06f
C13704 row_n[8] a_30986_10162# 0.0437f
C13705 rowoff_n[7] a_20034_9158# 0.294f
C13706 m2_1732_9982# rowoff_n[8] 0.415f
C13707 rowon_n[12] a_30074_14178# 0.248f
C13708 a_2275_4162# a_19334_4178# 0.144f
C13709 a_2475_4162# a_21950_4138# 0.264f
C13710 a_11910_4138# a_12002_4138# 0.326f
C13711 m3_4876_1078# ctop 0.21f
C13712 col[14] a_17022_7150# 0.367f
C13713 rowoff_n[13] a_27062_15182# 0.294f
C13714 vcm a_21950_17190# 0.1f
C13715 col[6] a_2275_17214# 0.0899f
C13716 col[21] a_23958_9158# 0.0682f
C13717 a_18026_14178# a_18026_13174# 0.843f
C13718 VDD a_18026_7150# 0.483f
C13719 rowoff_n[5] a_29070_7150# 0.294f
C13720 col[11] a_2275_6170# 0.0899f
C13721 col_n[29] a_32082_3134# 0.251f
C13722 col[9] rowoff_n[14] 0.0901f
C13723 a_2275_18218# a_22954_18194# 0.136f
C13724 a_11910_18194# a_12306_18234# 0.0313f
C13725 VDD a_7382_16548# 0.0779f
C13726 row_n[12] a_7986_14178# 0.282f
C13727 a_2275_1150# a_12914_1126# 0.136f
C13728 a_6890_1126# a_7286_1166# 0.0313f
C13729 vcm a_24050_2130# 0.56f
C13730 col[26] a_2475_16210# 0.136f
C13731 a_2275_6170# a_35398_6186# 0.145f
C13732 col_n[9] a_12306_7190# 0.084f
C13733 col[31] a_2475_5166# 0.136f
C13734 row_n[2] a_18026_4138# 0.282f
C13735 a_30986_11166# a_31478_11528# 0.0658f
C13736 a_30074_11166# a_30378_11206# 0.0931f
C13737 VDD a_8290_1166# 0.0149f
C13738 rowon_n[6] a_17934_8154# 0.118f
C13739 a_2475_15206# a_15014_15182# 0.316f
C13740 a_7986_15182# a_8990_15182# 0.843f
C13741 VDD a_33086_11166# 0.483f
C13742 col_n[20] a_23446_1488# 0.0283f
C13743 rowon_n[0] m2_22240_2378# 0.0322f
C13744 m2_1732_4962# col[0] 0.0137f
C13745 row_n[4] a_5278_6186# 0.0117f
C13746 col_n[30] a_33486_13536# 0.0283f
C13747 col_n[1] a_2475_2154# 0.0531f
C13748 a_2275_3158# a_27974_3134# 0.136f
C13749 a_2475_18218# a_20946_18194# 0.264f
C13750 vcm a_4974_5142# 0.56f
C13751 rowoff_n[11] a_33486_13536# 0.0133f
C13752 a_26970_8154# a_27062_8154# 0.326f
C13753 m2_3164_12418# a_2966_12170# 0.165f
C13754 a_2275_12194# a_5978_12170# 0.399f
C13755 col[3] a_5978_5142# 0.367f
C13756 VDD col_n[9] 5.17f
C13757 vcm col_n[6] 1.94f
C13758 m2_7756_18014# VDD 1.07f
C13759 row_n[15] a_28978_17190# 0.0437f
C13760 col[13] a_16018_17190# 0.367f
C13761 col[28] a_2275_8178# 0.0899f
C13762 a_2475_17214# a_30074_17190# 0.316f
C13763 col[10] a_12914_7150# 0.0682f
C13764 VDD a_14010_14178# 0.483f
C13765 a_30074_2130# m2_30272_2378# 0.165f
C13766 rowon_n[0] a_4974_2130# 0.248f
C13767 a_21950_5142# a_22346_5182# 0.0313f
C13768 col_n[28] a_31078_13174# 0.251f
C13769 col_n[25] a_27974_3134# 0.0765f
C13770 vcm a_20034_9158# 0.56f
C13771 rowoff_n[14] a_15014_16186# 0.294f
C13772 m3_22948_1078# a_23046_2130# 0.0302f
C13773 col_n[8] a_11302_17230# 0.084f
C13774 m2_19228_1374# a_19030_1126# 0.165f
C13775 a_11910_14178# a_12402_14540# 0.0658f
C13776 a_10998_14178# a_11302_14218# 0.0931f
C13777 a_2275_14202# a_21038_14178# 0.399f
C13778 m2_34864_15002# ctop 0.0422f
C13779 m2_5748_946# vcm 0.353f
C13780 col[1] a_3878_5142# 0.0682f
C13781 VDD a_29070_18194# 0.0356f
C13782 a_2475_2154# a_35094_2130# 0.0299f
C13783 a_18026_2130# a_19030_2130# 0.843f
C13784 col_n[13] a_2475_15206# 0.0531f
C13785 m3_23952_18146# VDD 0.0656f
C13786 col_n[18] a_2475_4162# 0.0531f
C13787 row_n[9] a_16018_11166# 0.282f
C13788 col_n[19] a_22442_11528# 0.0283f
C13789 vcm a_10298_3174# 0.155f
C13790 rowon_n[13] a_15926_15182# 0.118f
C13791 vcm a_35094_13174# 0.165f
C13792 a_2475_11190# a_13918_11166# 0.264f
C13793 a_2275_11190# a_11302_11206# 0.144f
C13794 a_7894_11166# a_7986_11166# 0.326f
C13795 VDD a_31990_3134# 0.181f
C13796 m2_17796_18014# a_18330_18234# 0.087f
C13797 row_n[11] a_3270_13214# 0.0117f
C13798 rowon_n[3] a_25966_5142# 0.118f
C13799 col[3] a_2475_12194# 0.136f
C13800 m2_7756_18014# m3_6884_18146# 0.0341f
C13801 m2_15212_14426# rowon_n[12] 0.0322f
C13802 col[8] a_2475_1150# 0.136f
C13803 col[2] a_4974_15182# 0.367f
C13804 m2_21236_10410# rowon_n[8] 0.0322f
C13805 m2_27260_6394# rowon_n[4] 0.0322f
C13806 a_8990_4138# a_8990_3134# 0.843f
C13807 row_n[1] a_13310_3174# 0.0117f
C13808 col[9] a_11910_17190# 0.0682f
C13809 vcm a_25358_7190# 0.155f
C13810 a_2275_8178# a_4882_8154# 0.136f
C13811 rowoff_n[12] a_21438_14540# 0.0133f
C13812 a_2966_8154# a_3970_8154# 0.843f
C13813 col_n[17] a_20034_11166# 0.251f
C13814 m2_34864_13998# a_35094_14178# 0.0249f
C13815 col_n[10] a_2275_18218# 0.113f
C13816 col_n[14] a_16930_1126# 0.0765f
C13817 ctop a_3970_1126# 0.544f
C13818 vcm a_16018_16186# 0.56f
C13819 a_2475_13198# a_28978_13174# 0.264f
C13820 col_n[15] a_2275_7174# 0.113f
C13821 a_2275_13198# a_26362_13214# 0.144f
C13822 VDD a_12914_6146# 0.181f
C13823 col_n[24] a_26970_13174# 0.0765f
C13824 rowon_n[7] a_2874_9158# 0.118f
C13825 a_26970_18194# a_27462_18556# 0.0658f
C13826 VDD a_35398_16226# 0.0882f
C13827 a_21950_1126# a_22442_1488# 0.0658f
C13828 col_n[30] a_2475_17214# 0.0531f
C13829 vcm a_18938_1126# 0.0983f
C13830 a_33086_6146# a_34090_6146# 0.843f
C13831 col[0] a_2275_15206# 0.099f
C13832 m2_9764_946# m3_10900_1078# 0.0341f
C13833 m3_14916_18146# m3_15920_18146# 0.202f
C13834 col[5] a_2275_4162# 0.0899f
C13835 vcm a_6282_10202# 0.155f
C13836 a_2275_10186# a_19942_10162# 0.136f
C13837 col_n[8] a_11398_9520# 0.0283f
C13838 rowoff_n[15] a_2874_17190# 0.202f
C13839 m2_7180_16434# a_6982_16186# 0.165f
C13840 m2_2736_1950# VDD 0.476f
C13841 ctop a_19030_5142# 4.11f
C13842 a_22954_15182# a_23046_15182# 0.326f
C13843 VDD a_27974_10162# 0.181f
C13844 col[20] a_2475_14202# 0.136f
C13845 col_n[14] rowoff_n[4] 0.0471f
C13846 col_n[19] rowoff_n[9] 0.0471f
C13847 col[25] a_2475_3158# 0.136f
C13848 col_n[18] rowoff_n[8] 0.0471f
C13849 col_n[11] rowoff_n[1] 0.0471f
C13850 col_n[15] rowoff_n[5] 0.0471f
C13851 col_n[12] rowoff_n[2] 0.0471f
C13852 col_n[16] rowoff_n[6] 0.0471f
C13853 col_n[13] rowoff_n[3] 0.0471f
C13854 col_n[17] rowoff_n[7] 0.0471f
C13855 col_n[10] rowoff_n[0] 0.0471f
C13856 vcm a_33998_5142# 0.1f
C13857 a_24050_8154# a_24050_7150# 0.843f
C13858 a_2475_7174# a_12002_7150# 0.316f
C13859 rowoff_n[2] a_10906_4138# 0.202f
C13860 rowoff_n[10] a_27974_12170# 0.202f
C13861 m2_26256_12418# a_26058_12170# 0.165f
C13862 row_n[6] a_24050_8154# 0.282f
C13863 vcm a_21342_14218# 0.155f
C13864 a_2275_12194# a_35002_12170# 0.136f
C13865 a_17934_12170# a_18330_12210# 0.0313f
C13866 rowon_n[10] a_23958_12170# 0.118f
C13867 VDD a_19430_4500# 0.0779f
C13868 col_n[6] a_8990_9158# 0.251f
C13869 ctop a_34090_9158# 4.06f
C13870 m3_34996_7102# a_34090_7150# 0.0303f
C13871 VDD a_8898_13174# 0.181f
C13872 col_n[13] a_15926_11166# 0.0765f
C13873 row_n[8] a_11302_10202# 0.0117f
C13874 rowoff_n[0] a_19942_2130# 0.202f
C13875 rowon_n[0] a_33998_2130# 0.118f
C13876 rowoff_n[7] a_1957_9182# 0.0219f
C13877 a_2275_4162# a_2874_4138# 0.136f
C13878 a_2475_4162# a_3878_4138# 0.264f
C13879 m2_22816_946# col[20] 0.425f
C13880 col[17] a_2275_17214# 0.0899f
C13881 m2_31852_18014# m2_32280_18442# 0.165f
C13882 vcm a_14922_8154# 0.1f
C13883 rowoff_n[13] a_9390_15544# 0.0133f
C13884 a_2475_9182# a_27062_9158# 0.316f
C13885 a_14010_9158# a_15014_9158# 0.843f
C13886 col[22] a_2275_6170# 0.0899f
C13887 col[20] rowoff_n[14] 0.0901f
C13888 vcm a_3878_17190# 0.1f
C13889 VDD a_34490_8516# 0.0779f
C13890 rowoff_n[5] a_11398_7512# 0.0133f
C13891 ctop a_15014_12170# 4.11f
C13892 col_n[3] rowoff_n[10] 0.0471f
C13893 a_2275_18218# a_3270_18234# 0.145f
C13894 row_n[0] a_11910_2130# 0.0437f
C13895 VDD a_23958_17190# 0.181f
C13896 col[26] a_29070_8154# 0.367f
C13897 a_32994_2130# a_33086_2130# 0.326f
C13898 rowon_n[4] a_10998_6146# 0.248f
C13899 a_2275_6170# a_18026_6146# 0.399f
C13900 m2_17220_10410# a_17022_10162# 0.165f
C13901 rowoff_n[3] a_20434_5504# 0.0133f
C13902 vcm a_29982_12170# 0.1f
C13903 a_4974_11166# a_4974_10162# 0.843f
C13904 VDD a_26058_2130# 0.483f
C13905 m2_8184_17438# row_n[15] 0.0128f
C13906 m2_14208_13422# row_n[11] 0.0128f
C13907 m2_20232_9406# row_n[7] 0.0128f
C13908 col_n[7] a_2475_13198# 0.0531f
C13909 m2_26256_5390# row_n[3] 0.0128f
C13910 a_32994_16186# a_33390_16226# 0.0313f
C13911 VDD a_15414_11528# 0.0779f
C13912 col_n[12] a_2475_2154# 0.0531f
C13913 col_n[21] a_24354_8194# 0.084f
C13914 ctop a_30074_16186# 4.11f
C13915 a_2475_18218# a_2275_18218# 2.77f
C13916 a_2475_3158# a_10906_3134# 0.264f
C13917 a_2275_3158# a_8290_3174# 0.144f
C13918 rowoff_n[1] a_29470_3496# 0.0133f
C13919 rowoff_n[8] a_12002_10162# 0.294f
C13920 col_n[2] a_4882_9158# 0.0765f
C13921 a_24050_1126# a_2475_1150# 0.0299f
C13922 row_n[13] a_22042_15182# 0.282f
C13923 a_17934_8154# a_18426_8516# 0.0658f
C13924 rowoff_n[11] a_15926_13174# 0.202f
C13925 a_17022_8154# a_17326_8194# 0.0931f
C13926 a_2275_8178# a_33086_8154# 0.399f
C13927 vcm col_n[17] 1.93f
C13928 VDD col_n[20] 5.17f
C13929 col_n[8] col_n[9] 0.0101f
C13930 col[18] col[19] 0.0355f
C13931 col[4] rowoff_n[15] 0.0901f
C13932 vcm a_10906_15182# 0.1f
C13933 a_29070_13174# a_30074_13174# 0.843f
C13934 VDD a_6982_5142# 0.483f
C13935 row_n[3] a_32082_5142# 0.282f
C13936 row_n[15] a_9294_17230# 0.0117f
C13937 a_2275_17214# a_11910_17190# 0.136f
C13938 rowon_n[7] a_31990_9158# 0.118f
C13939 rowoff_n[6] a_21038_8154# 0.294f
C13940 VDD a_30474_15544# 0.0779f
C13941 col_n[4] a_2275_16210# 0.113f
C13942 row_n[5] a_19334_7190# 0.0117f
C13943 a_13918_5142# a_14010_5142# 0.326f
C13944 a_2275_5166# a_23350_5182# 0.144f
C13945 a_2475_5166# a_25966_5142# 0.264f
C13946 col[15] a_18026_6146# 0.367f
C13947 col_n[9] a_2275_5166# 0.113f
C13948 m2_8184_8402# a_7986_8154# 0.165f
C13949 m3_4876_1078# m3_5880_1078# 0.202f
C13950 vcm a_1957_9182# 0.139f
C13951 rowoff_n[15] a_31990_17190# 0.202f
C13952 col[22] a_24962_8154# 0.0682f
C13953 rowoff_n[4] a_30074_6146# 0.294f
C13954 m2_16792_946# a_2475_1150# 0.286f
C13955 a_2475_14202# a_3970_14178# 0.316f
C13956 a_2275_14202# a_2966_14178# 0.399f
C13957 m2_6752_946# a_6982_1126# 0.0249f
C13958 a_20034_15182# a_20034_14178# 0.843f
C13959 col_n[30] a_33086_2130# 0.251f
C13960 row_n[7] a_9902_9158# 0.0437f
C13961 VDD a_22042_9158# 0.483f
C13962 col_n[24] a_2475_15206# 0.0531f
C13963 ctop a_2275_13198# 0.0683f
C13964 rowon_n[11] a_8990_13174# 0.248f
C13965 col_n[29] a_2475_4162# 0.0531f
C13966 VDD a_11398_18556# 0.0858f
C13967 a_2275_2154# a_16930_2130# 0.136f
C13968 a_8898_2130# a_9294_2170# 0.0313f
C13969 col_n[10] a_13310_6186# 0.084f
C13970 m2_27260_4386# a_27062_4138# 0.165f
C13971 m2_9764_946# VDD 1f
C13972 vcm a_28066_4138# 0.56f
C13973 rowon_n[1] a_19030_3134# 0.248f
C13974 col_n[20] a_23350_18234# 0.084f
C13975 a_32994_12170# a_33486_12532# 0.0658f
C13976 col[14] a_2475_12194# 0.136f
C13977 a_32082_12170# a_32386_12210# 0.0931f
C13978 col[19] a_2475_1150# 0.136f
C13979 a_2475_16210# a_19030_16186# 0.316f
C13980 a_9994_16186# a_10998_16186# 0.843f
C13981 VDD a_2874_12170# 0.182f
C13982 col_n[31] a_34490_12532# 0.0283f
C13983 a_2275_4162# a_31990_4138# 0.136f
C13984 col_n[21] a_2275_18218# 0.113f
C13985 vcm a_8990_7150# 0.56f
C13986 col_n[26] a_2275_7174# 0.113f
C13987 rowoff_n[12] a_3366_14540# 0.0133f
C13988 a_28978_9158# a_29070_9158# 0.326f
C13989 row_n[10] a_30074_12170# 0.282f
C13990 col[4] a_6982_4138# 0.367f
C13991 rowon_n[14] a_29982_16186# 0.118f
C13992 col[14] a_17022_16186# 0.367f
C13993 a_2275_13198# a_9994_13174# 0.399f
C13994 col[11] a_13918_6146# 0.0682f
C13995 col[21] a_23958_18194# 0.0682f
C13996 VDD a_18026_16186# 0.483f
C13997 col[11] a_2275_15206# 0.0899f
C13998 row_n[12] a_17326_14218# 0.0117f
C13999 col_n[29] a_32082_12170# 0.251f
C14000 col[16] a_2275_4162# 0.0899f
C14001 col_n[26] a_28978_2130# 0.0765f
C14002 vcm a_33390_2170# 0.155f
C14003 a_23958_6146# a_24354_6186# 0.0313f
C14004 row_n[2] a_27366_4178# 0.0117f
C14005 vcm a_24050_11166# 0.56f
C14006 row_n[14] a_7894_16186# 0.0437f
C14007 VDD a_20946_1126# 0.405f
C14008 col_n[9] a_12306_16226# 0.084f
C14009 col[31] a_2475_14202# 0.136f
C14010 a_2275_15206# a_25054_15182# 0.399f
C14011 a_13918_15182# a_14410_15544# 0.0658f
C14012 a_13006_15182# a_13310_15222# 0.0931f
C14013 col_n[23] rowoff_n[2] 0.0471f
C14014 col_n[25] rowoff_n[4] 0.0471f
C14015 col_n[27] rowoff_n[6] 0.0471f
C14016 col_n[30] rowoff_n[9] 0.0471f
C14017 col_n[28] rowoff_n[7] 0.0471f
C14018 col_n[24] rowoff_n[3] 0.0471f
C14019 col_n[22] rowoff_n[1] 0.0471f
C14020 col_n[29] rowoff_n[8] 0.0471f
C14021 col_n[26] rowoff_n[5] 0.0471f
C14022 col_n[21] rowoff_n[0] 0.0471f
C14023 row_n[4] a_17934_6146# 0.0437f
C14024 col_n[7] a_2475_18218# 0.0529f
C14025 rowon_n[8] a_17022_10162# 0.248f
C14026 col_n[20] a_23446_10524# 0.0283f
C14027 a_20034_3134# a_21038_3134# 0.843f
C14028 vcm a_14314_5182# 0.155f
C14029 col_n[1] a_2475_11190# 0.0531f
C14030 m2_4168_12418# rowon_n[10] 0.0322f
C14031 m2_10192_8402# rowon_n[6] 0.0322f
C14032 vcm a_4974_14178# 0.56f
C14033 a_2275_12194# a_15318_12210# 0.144f
C14034 a_9902_12170# a_9994_12170# 0.326f
C14035 a_2475_12194# a_17934_12170# 0.264f
C14036 m2_16216_4386# rowon_n[2] 0.0322f
C14037 m2_29268_18442# VDD 0.0456f
C14038 col[3] a_5978_14178# 0.367f
C14039 col[28] a_2275_17214# 0.0899f
C14040 col[10] a_12914_16186# 0.0682f
C14041 a_10998_5142# a_10998_4138# 0.843f
C14042 col_n[18] a_21038_10162# 0.251f
C14043 col[31] rowoff_n[14] 0.0901f
C14044 vcm a_29374_9198# 0.155f
C14045 m2_13780_18014# m2_14784_18014# 0.843f
C14046 a_2275_9182# a_8898_9158# 0.136f
C14047 a_4882_9158# a_5278_9198# 0.0313f
C14048 VDD m2_34864_1950# 0.785f
C14049 col_n[25] a_27974_12170# 0.0765f
C14050 rowon_n[2] a_4882_4138# 0.118f
C14051 vcm a_20034_18194# 0.165f
C14052 col_n[14] rowoff_n[10] 0.0471f
C14053 ctop a_7986_3134# 4.11f
C14054 m2_25252_17438# rowon_n[15] 0.0322f
C14055 a_2475_14202# a_32994_14178# 0.264f
C14056 a_2275_14202# a_30378_14218# 0.144f
C14057 VDD a_16930_8154# 0.181f
C14058 m2_31276_13422# rowon_n[11] 0.0322f
C14059 col[0] m2_2736_946# 0.425f
C14060 m2_28840_946# vcm 0.353f
C14061 col_n[3] a_2275_3158# 0.113f
C14062 a_23046_2130# a_23350_2170# 0.0931f
C14063 a_23958_2130# a_24450_2492# 0.0658f
C14064 col[1] a_3878_14178# 0.0682f
C14065 vcm a_22954_3134# 0.1f
C14066 row_n[9] a_25358_11206# 0.0117f
C14067 col_n[9] a_12402_8516# 0.0283f
C14068 m2_1732_9982# a_2966_10162# 0.843f
C14069 col_n[18] a_2475_13198# 0.0531f
C14070 rowoff_n[3] a_2161_5166# 0.0226f
C14071 vcm a_10298_12210# 0.155f
C14072 a_2275_11190# a_23958_11166# 0.136f
C14073 col_n[23] a_2475_2154# 0.0531f
C14074 VDD a_8386_2492# 0.0779f
C14075 m2_34864_9982# VDD 0.784f
C14076 ctop a_23046_7150# 4.11f
C14077 row_n[11] a_15926_13174# 0.0437f
C14078 a_24962_16186# a_25054_16186# 0.326f
C14079 VDD a_31990_12170# 0.181f
C14080 m2_21812_18014# m3_21944_18146# 3.79f
C14081 rowon_n[15] a_15014_17190# 0.248f
C14082 vcm col_n[28] 1.94f
C14083 VDD col_n[31] 5.04f
C14084 row_n[1] a_25966_3134# 0.0437f
C14085 rowoff_n[1] a_11910_3134# 0.202f
C14086 col[15] rowoff_n[15] 0.0901f
C14087 col[8] a_2475_10186# 0.136f
C14088 m2_34864_15002# m2_35292_15430# 0.165f
C14089 rowon_n[5] a_25054_7150# 0.248f
C14090 rowoff_n[12] a_32082_14178# 0.294f
C14091 a_26058_9158# a_26058_8154# 0.843f
C14092 a_2475_8178# a_16018_8154# 0.316f
C14093 sample rowoff_n[11] 0.0775f
C14094 m2_34864_12994# a_2275_13198# 0.278f
C14095 col_n[7] a_9994_8154# 0.251f
C14096 vcm a_25358_16226# 0.155f
C14097 a_19942_13174# a_20338_13214# 0.0313f
C14098 VDD a_23446_6508# 0.0779f
C14099 col_n[14] a_16930_10162# 0.0765f
C14100 ctop a_3970_10162# 4.11f
C14101 col_n[15] a_2275_16210# 0.113f
C14102 VDD a_12914_15182# 0.181f
C14103 rowoff_n[6] a_2966_8154# 0.294f
C14104 col_n[20] a_2275_5166# 0.113f
C14105 m3_5880_18146# a_5978_17190# 0.0303f
C14106 a_2275_5166# a_6982_5142# 0.399f
C14107 a_4882_5142# a_5374_5504# 0.0658f
C14108 a_3970_5142# a_4274_5182# 0.0931f
C14109 row_n[5] a_2874_7150# 0.0436f
C14110 m3_1864_17142# m3_1864_16138# 0.202f
C14111 m2_25828_946# m3_24956_1078# 0.0341f
C14112 rowon_n[9] a_2161_11190# 0.0177f
C14113 vcm a_18938_10162# 0.1f
C14114 a_2475_10186# a_31078_10162# 0.316f
C14115 a_16018_10162# a_17022_10162# 0.843f
C14116 col[5] a_2275_13198# 0.0899f
C14117 rowoff_n[4] a_12402_6508# 0.0133f
C14118 col_n[8] a_11398_18556# 0.0283f
C14119 VDD a_4370_9520# 0.0779f
C14120 col[10] a_2275_2154# 0.0899f
C14121 m2_17796_18014# ctop 0.0422f
C14122 col_n[31] a_34394_9198# 0.084f
C14123 col[27] a_30074_7150# 0.367f
C14124 ctop a_19030_14178# 4.11f
C14125 a_35002_3134# a_35094_3134# 0.0991f
C14126 a_34090_3134# a_34394_3174# 0.0931f
C14127 m2_3164_11414# row_n[9] 0.0128f
C14128 m2_9188_7398# row_n[5] 0.0128f
C14129 m2_15212_3382# row_n[1] 0.0128f
C14130 col[25] a_2475_12194# 0.136f
C14131 a_2275_7174# a_22042_7150# 0.399f
C14132 rowoff_n[2] a_21438_4500# 0.0133f
C14133 rowoff_n[9] a_3970_11166# 0.294f
C14134 m2_34864_11990# a_35002_12170# 0.225f
C14135 col[30] a_2475_1150# 0.136f
C14136 row_n[6] a_33390_8194# 0.0117f
C14137 vcm a_33998_14178# 0.1f
C14138 a_6982_12170# a_6982_11166# 0.843f
C14139 VDD a_30074_4138# 0.483f
C14140 col_n[22] a_25358_7190# 0.084f
C14141 VDD a_19430_13536# 0.0779f
C14142 row_n[8] a_23958_10162# 0.0437f
C14143 rowoff_n[0] a_30474_2492# 0.0133f
C14144 col_n[3] a_5886_8154# 0.0765f
C14145 rowoff_n[7] a_13006_9158# 0.294f
C14146 rowon_n[12] a_23046_14178# 0.248f
C14147 a_2275_4162# a_12306_4178# 0.144f
C14148 a_2475_4162# a_14922_4138# 0.264f
C14149 m3_1864_13126# ctop 0.21f
C14150 a_29982_1126# col_n[27] 0.0774f
C14151 m2_24248_16434# row_n[14] 0.0128f
C14152 m2_30272_12418# row_n[10] 0.0128f
C14153 a_19942_9158# a_20434_9520# 0.0658f
C14154 m2_35292_8402# row_n[6] 0.0128f
C14155 rowoff_n[13] a_20034_15182# 0.294f
C14156 a_19030_9158# a_19334_9198# 0.0931f
C14157 rowon_n[2] a_33086_4138# 0.248f
C14158 vcm a_14922_17190# 0.1f
C14159 a_31078_14178# a_32082_14178# 0.843f
C14160 VDD a_10998_7150# 0.483f
C14161 col[22] a_2275_15206# 0.0899f
C14162 rowoff_n[5] a_22042_7150# 0.294f
C14163 col[27] a_2275_4162# 0.0899f
C14164 a_2275_18218# a_15926_18194# 0.136f
C14165 VDD a_34490_17552# 0.0779f
C14166 a_2275_1150# a_5886_1126# 0.136f
C14167 m2_2736_1950# a_3970_2130# 0.843f
C14168 col[16] a_19030_5142# 0.367f
C14169 vcm a_17022_2130# 0.56f
C14170 a_2475_6170# a_29982_6146# 0.264f
C14171 col[26] a_29070_17190# 0.367f
C14172 a_15926_6146# a_16018_6146# 0.326f
C14173 a_2275_6170# a_27366_6186# 0.144f
C14174 col[23] a_25966_7150# 0.0682f
C14175 rowoff_n[3] a_31078_5142# 0.294f
C14176 row_n[2] a_10998_4138# 0.282f
C14177 VDD a_2275_1150# 21f
C14178 m2_13204_17438# a_13006_17190# 0.165f
C14179 rowon_n[6] a_10906_8154# 0.118f
C14180 a_2475_15206# a_7986_15182# 0.316f
C14181 a_22042_16186# a_22042_15182# 0.843f
C14182 col_n[18] a_2475_18218# 0.0529f
C14183 VDD a_26058_11166# 0.483f
C14184 col_n[11] a_14314_5182# 0.084f
C14185 col_n[12] a_2475_11190# 0.0531f
C14186 a_10906_3134# a_11302_3174# 0.0313f
C14187 a_2275_3158# a_20946_3134# 0.136f
C14188 a_2475_18218# a_13918_18194# 0.264f
C14189 col_n[21] a_24354_17230# 0.084f
C14190 a_35094_1126# a_2275_1150# 0.0924f
C14191 row_n[13] a_31382_15222# 0.0117f
C14192 vcm a_32082_6146# 0.56f
C14193 rowoff_n[11] a_26458_13536# 0.0133f
C14194 col_n[2] a_4882_18194# 0.0762f
C14195 m2_32280_13422# a_32082_13174# 0.165f
C14196 a_35002_13174# a_35494_13536# 0.0658f
C14197 a_31478_1488# VDD 0.0977f
C14198 row_n[15] a_21950_17190# 0.0437f
C14199 a_12002_17190# a_13006_17190# 0.843f
C14200 col[2] a_2475_8178# 0.136f
C14201 a_2475_17214# a_23046_17190# 0.316f
C14202 VDD a_6982_14178# 0.483f
C14203 row_n[5] a_31990_7150# 0.0437f
C14204 a_2275_5166# a_34394_5182# 0.144f
C14205 col[5] a_7986_3134# 0.367f
C14206 col_n[25] rowoff_n[10] 0.0471f
C14207 rowon_n[9] a_31078_11166# 0.248f
C14208 a_31990_1126# a_32386_1166# 0.0313f
C14209 vcm a_13006_9158# 0.56f
C14210 rowoff_n[14] a_7986_16186# 0.294f
C14211 a_30986_10162# a_31078_10162# 0.326f
C14212 col_n[9] a_2275_14202# 0.113f
C14213 col[15] a_18026_15182# 0.367f
C14214 m2_4168_15430# a_3970_15182# 0.165f
C14215 col[12] a_14922_5142# 0.0682f
C14216 col_n[14] a_2275_3158# 0.113f
C14217 vcm a_1957_18218# 0.139f
C14218 m2_12776_946# a_13310_1166# 0.087f
C14219 a_2275_14202# a_14010_14178# 0.399f
C14220 col[22] a_24962_17190# 0.0682f
C14221 col_n[30] a_33086_11166# 0.251f
C14222 VDD a_22042_18194# 0.0356f
C14223 a_2475_2154# a_28066_2130# 0.316f
C14224 a_32082_3134# a_32082_2130# 0.843f
C14225 col_n[29] a_2475_13198# 0.0531f
C14226 m2_34864_3958# a_35398_4178# 0.087f
C14227 m2_32856_946# VDD 1.01f
C14228 vcm a_3270_3174# 0.155f
C14229 row_n[9] a_8990_11166# 0.282f
C14230 rowoff_n[9] a_32994_11166# 0.202f
C14231 a_25966_7150# a_26362_7190# 0.0313f
C14232 m2_1732_16006# sample_n 0.0522f
C14233 m2_23244_11414# a_23046_11166# 0.165f
C14234 rowon_n[13] a_8898_15182# 0.118f
C14235 col_n[10] a_13310_15222# 0.084f
C14236 vcm a_28066_13174# 0.56f
C14237 a_2475_11190# a_6890_11166# 0.264f
C14238 a_2275_11190# a_4274_11206# 0.144f
C14239 VDD a_24962_3134# 0.181f
C14240 a_15926_16186# a_16418_16548# 0.0658f
C14241 a_15014_16186# a_15318_16226# 0.0931f
C14242 a_2275_16210# a_29070_16186# 0.399f
C14243 rowon_n[3] a_18938_5142# 0.118f
C14244 col_n[2] row_n[13] 0.298f
C14245 vcm row_n[12] 0.616f
C14246 col_n[19] col_n[20] 0.0101f
C14247 col_n[3] rowon_n[13] 0.111f
C14248 col_n[1] rowon_n[12] 0.111f
C14249 col_n[7] rowon_n[15] 0.111f
C14250 VDD rowon_n[10] 3.04f
C14251 col_n[6] row_n[15] 0.298f
C14252 sample row_n[11] 0.423f
C14253 col_n[4] row_n[14] 0.298f
C14254 col_n[0] rowon_n[11] 0.111f
C14255 col_n[5] rowon_n[14] 0.111f
C14256 col[29] col[30] 0.0355f
C14257 col[26] rowoff_n[15] 0.0901f
C14258 col[19] a_2475_10186# 0.136f
C14259 col_n[21] a_24450_9520# 0.0283f
C14260 m2_4168_2378# rowon_n[0] 0.0322f
C14261 a_22042_4138# a_23046_4138# 0.843f
C14262 col_n[9] rowoff_n[11] 0.0471f
C14263 row_n[1] a_6282_3174# 0.0117f
C14264 vcm a_18330_7190# 0.155f
C14265 rowoff_n[12] a_14410_14540# 0.0133f
C14266 sample a_2161_3158# 0.0858f
C14267 ctop a_31078_2130# 4.06f
C14268 col_n[26] a_2275_16210# 0.113f
C14269 vcm a_8990_16186# 0.56f
C14270 a_2475_13198# a_21950_13174# 0.264f
C14271 a_2275_13198# a_19334_13214# 0.144f
C14272 a_11910_13174# a_12002_13174# 0.326f
C14273 VDD a_5886_6146# 0.181f
C14274 col[4] a_6982_13174# 0.367f
C14275 col_n[31] a_2275_5166# 0.113f
C14276 m2_33860_18014# a_2475_18218# 0.286f
C14277 col[11] a_13918_15182# 0.0682f
C14278 row_n[12] a_29982_14178# 0.0437f
C14279 col_n[19] a_22042_9158# 0.251f
C14280 m2_14208_15430# rowon_n[13] 0.0322f
C14281 vcm a_11910_1126# 0.0989f
C14282 a_13006_6146# a_13006_5142# 0.843f
C14283 m2_20232_11414# rowon_n[9] 0.0322f
C14284 m2_26256_7398# rowon_n[5] 0.0322f
C14285 m2_14208_9406# a_14010_9158# 0.165f
C14286 col[16] a_2275_13198# 0.0899f
C14287 m2_32280_3382# rowon_n[1] 0.0322f
C14288 col_n[26] a_28978_11166# 0.0765f
C14289 vcm a_33390_11206# 0.155f
C14290 col[21] a_2275_2154# 0.0899f
C14291 a_6890_10162# a_7286_10202# 0.0313f
C14292 a_2275_10186# a_12914_10162# 0.136f
C14293 ctop a_12002_5142# 4.11f
C14294 a_2275_15206# a_35398_15222# 0.145f
C14295 m2_5748_946# a_5978_2130# 0.843f
C14296 VDD a_20946_10162# 0.181f
C14297 a_25054_3134# a_25358_3174# 0.0931f
C14298 a_25966_3134# a_26458_3496# 0.0658f
C14299 col_n[10] a_13406_7512# 0.0283f
C14300 m2_33284_5390# a_33086_5142# 0.165f
C14301 vcm a_26970_5142# 0.1f
C14302 rowoff_n[2] a_3366_4500# 0.0133f
C14303 rowoff_n[10] a_20946_12170# 0.202f
C14304 a_2475_7174# a_4974_7150# 0.316f
C14305 row_n[6] a_17022_8154# 0.282f
C14306 vcm a_14314_14218# 0.155f
C14307 a_2275_12194# a_27974_12170# 0.136f
C14308 VDD a_12402_4500# 0.0779f
C14309 rowon_n[10] a_16930_12170# 0.118f
C14310 col_n[6] a_2475_9182# 0.0531f
C14311 ctop a_27062_9158# 4.11f
C14312 a_26970_17190# a_27062_17190# 0.326f
C14313 row_n[8] a_4274_10202# 0.0117f
C14314 rowon_n[0] a_26970_2130# 0.118f
C14315 rowoff_n[0] a_12914_2130# 0.202f
C14316 m2_5172_7398# a_4974_7150# 0.165f
C14317 m2_24824_18014# m2_25252_18442# 0.165f
C14318 vcm a_7894_8154# 0.1f
C14319 a_28066_10162# a_28066_9158# 0.843f
C14320 col_n[8] a_10998_7150# 0.251f
C14321 a_2475_9182# a_20034_9158# 0.316f
C14322 rowoff_n[13] a_1957_15206# 0.0219f
C14323 vcm a_29374_18234# 0.16f
C14324 col_n[15] a_17934_9158# 0.0765f
C14325 a_21950_14178# a_22346_14218# 0.0313f
C14326 VDD a_27462_8516# 0.0779f
C14327 rowoff_n[5] a_4370_7512# 0.0133f
C14328 ctop a_7986_12170# 4.11f
C14329 VDD a_16930_17190# 0.181f
C14330 row_n[0] a_4882_2130# 0.0437f
C14331 rowon_n[4] a_3970_6146# 0.248f
C14332 m2_24248_3382# a_24050_3134# 0.165f
C14333 col_n[3] a_2275_12194# 0.113f
C14334 row_n[7] rowoff_n[6] 0.085f
C14335 a_5978_6146# a_6282_6186# 0.0931f
C14336 col_n[8] a_2275_1150# 0.113f
C14337 a_6890_6146# a_7382_6508# 0.0658f
C14338 a_2275_6170# a_10998_6146# 0.399f
C14339 m2_34864_10986# vcm 0.408f
C14340 vcm a_22954_12170# 0.1f
C14341 rowoff_n[3] a_13406_5504# 0.0133f
C14342 col_n[29] a_2475_18218# 0.0529f
C14343 a_2475_11190# a_35094_11166# 0.0299f
C14344 a_18026_11166# a_19030_11166# 0.843f
C14345 col_n[9] a_12402_17552# 0.0283f
C14346 VDD a_19030_2130# 0.483f
C14347 col[28] a_31078_6146# 0.367f
C14348 VDD a_8386_11528# 0.0779f
C14349 col_n[23] a_2475_11190# 0.0531f
C14350 ctop a_23046_16186# 4.11f
C14351 m2_6752_946# col[4] 0.425f
C14352 rowoff_n[1] a_22442_3496# 0.0133f
C14353 rowoff_n[8] a_4974_10162# 0.294f
C14354 row_n[13] a_15014_15182# 0.282f
C14355 a_2275_8178# a_26058_8154# 0.399f
C14356 rowoff_n[11] a_8898_13174# 0.202f
C14357 col[13] a_2475_8178# 0.136f
C14358 a_8990_13174# a_8990_12170# 0.843f
C14359 VDD a_34090_6146# 0.483f
C14360 col_n[23] a_26362_6186# 0.084f
C14361 row_n[3] a_25054_5142# 0.282f
C14362 row_n[15] a_3878_17190# 0.0437f
C14363 col_n[7] a_9994_17190# 0.251f
C14364 rowon_n[7] a_24962_9158# 0.118f
C14365 m2_13204_14426# row_n[12] 0.0128f
C14366 a_2966_17190# a_3970_17190# 0.843f
C14367 a_2275_17214# a_4882_17190# 0.136f
C14368 m2_19228_10410# row_n[8] 0.0128f
C14369 col_n[4] a_6890_7150# 0.0765f
C14370 rowoff_n[6] a_14010_8154# 0.294f
C14371 VDD a_23446_15544# 0.0779f
C14372 m2_25252_6394# row_n[4] 0.0128f
C14373 row_n[5] a_12306_7190# 0.0117f
C14374 col_n[20] a_2275_14202# 0.113f
C14375 a_2275_5166# a_16322_5182# 0.144f
C14376 a_2475_5166# a_18938_5142# 0.264f
C14377 m2_1732_7974# a_2275_8178# 0.191f
C14378 col_n[25] a_2275_3158# 0.113f
C14379 a_21038_10162# a_21342_10202# 0.0931f
C14380 a_21950_10162# a_22442_10524# 0.0658f
C14381 rowoff_n[15] a_24962_17190# 0.202f
C14382 rowoff_n[4] a_23046_6146# 0.294f
C14383 m3_2868_2082# a_3970_2130# 0.0303f
C14384 a_33086_15182# a_34090_15182# 0.843f
C14385 VDD a_15014_9158# 0.483f
C14386 row_n[7] a_2161_9182# 0.0221f
C14387 rowon_n[11] a_2475_13198# 0.31f
C14388 col[17] a_20034_4138# 0.367f
C14389 col[10] a_2275_11190# 0.0899f
C14390 VDD a_4370_18556# 0.0858f
C14391 col_n[31] a_34394_18234# 0.084f
C14392 a_2275_2154# a_9902_2130# 0.136f
C14393 col[27] a_30074_16186# 0.367f
C14394 col[24] a_26970_6146# 0.0682f
C14395 vcm a_21038_4138# 0.56f
C14396 a_2275_7174# a_31382_7190# 0.144f
C14397 rowon_n[1] a_12002_3134# 0.248f
C14398 a_17934_7150# a_18026_7150# 0.326f
C14399 rowoff_n[2] a_32082_4138# 0.294f
C14400 a_2475_7174# a_33998_7150# 0.264f
C14401 m2_1732_1950# sample 0.2f
C14402 col_n[18] rowon_n[15] 0.111f
C14403 col_n[7] row_n[10] 0.298f
C14404 col_n[13] row_n[13] 0.298f
C14405 col_n[16] rowon_n[14] 0.111f
C14406 col_n[3] row_n[8] 0.298f
C14407 col_n[2] rowon_n[7] 0.111f
C14408 col_n[5] row_n[9] 0.298f
C14409 col_n[0] row_n[6] 0.298f
C14410 col_n[8] rowon_n[10] 0.111f
C14411 col_n[17] row_n[15] 0.298f
C14412 col_n[10] rowon_n[11] 0.111f
C14413 vcm rowon_n[6] 0.65f
C14414 VDD row_n[5] 3.29f
C14415 col_n[6] rowon_n[9] 0.111f
C14416 col_n[4] rowon_n[8] 0.111f
C14417 col_n[1] row_n[7] 0.298f
C14418 col_n[11] row_n[12] 0.298f
C14419 sample rowon_n[5] 0.0935f
C14420 col_n[9] row_n[11] 0.298f
C14421 col_n[15] row_n[14] 0.298f
C14422 col_n[12] rowon_n[12] 0.111f
C14423 col_n[14] rowon_n[13] 0.111f
C14424 col[30] a_2475_10186# 0.136f
C14425 m2_1732_12994# VDD 0.856f
C14426 a_2475_16210# a_12002_16186# 0.316f
C14427 a_24050_17190# a_24050_16186# 0.843f
C14428 VDD a_30074_13174# 0.483f
C14429 col_n[12] a_15318_4178# 0.084f
C14430 col_n[20] rowoff_n[11] 0.0471f
C14431 col_n[22] a_25358_16226# 0.084f
C14432 a_2275_4162# a_24962_4138# 0.136f
C14433 a_12914_4138# a_13310_4178# 0.0313f
C14434 m3_19936_1078# ctop 0.317f
C14435 col_n[3] a_5886_17190# 0.0765f
C14436 vcm a_2475_7174# 1.08f
C14437 row_n[10] a_23046_12170# 0.282f
C14438 a_2475_13198# a_3878_13174# 0.264f
C14439 rowon_n[14] a_22954_16186# 0.118f
C14440 a_2275_13198# a_2874_13174# 0.136f
C14441 m2_15788_18014# col_n[13] 0.243f
C14442 row_n[0] a_33086_2130# 0.282f
C14443 VDD a_10998_16186# 0.483f
C14444 a_2475_1150# a_17022_1126# 0.0299f
C14445 row_n[12] a_10298_14218# 0.0117f
C14446 rowon_n[4] a_32994_6146# 0.118f
C14447 col[27] a_2275_13198# 0.0899f
C14448 col[6] a_8990_2130# 0.367f
C14449 vcm a_26362_2170# 0.155f
C14450 m2_15788_946# m2_16792_946# 0.843f
C14451 m2_34864_9982# a_34090_10162# 0.843f
C14452 col[16] a_19030_14178# 0.367f
C14453 col[13] a_15926_4138# 0.0682f
C14454 row_n[2] a_20338_4178# 0.0117f
C14455 vcm a_17022_11166# 0.56f
C14456 a_32994_11166# a_33086_11166# 0.326f
C14457 VDD a_13918_1126# 0.405f
C14458 col[23] a_25966_16186# 0.0682f
C14459 a_2275_15206# a_18026_15182# 0.399f
C14460 col_n[4] rowoff_n[12] 0.0471f
C14461 VDD a_2275_10186# 1.96f
C14462 col_n[31] a_34090_10162# 0.251f
C14463 row_n[4] a_10906_6146# 0.0437f
C14464 col_n[1] a_4274_2170# 0.0839f
C14465 a_2475_3158# a_32082_3134# 0.316f
C14466 a_34090_4138# a_34090_3134# 0.843f
C14467 rowon_n[8] a_9994_10162# 0.248f
C14468 rowoff_n[8] a_33998_10162# 0.202f
C14469 a_24050_1126# a_23958_1126# 0.0991f
C14470 col_n[11] a_14314_14218# 0.084f
C14471 vcm a_7286_5182# 0.155f
C14472 a_27974_8154# a_28370_8194# 0.0313f
C14473 rowoff_n[10] a_2275_12194# 0.151f
C14474 col_n[17] a_2475_9182# 0.0531f
C14475 vcm a_32082_15182# 0.56f
C14476 a_2475_12194# a_10906_12170# 0.264f
C14477 a_2275_12194# a_8290_12210# 0.144f
C14478 VDD a_28978_5142# 0.181f
C14479 m2_15212_18442# VDD 0.0456f
C14480 a_17934_17190# a_18426_17552# 0.0658f
C14481 col_n[22] a_25454_8516# 0.0283f
C14482 a_2275_17214# a_33086_17190# 0.399f
C14483 a_17022_17190# a_17326_17230# 0.0931f
C14484 a_33086_2130# m2_33284_2378# 0.165f
C14485 col[2] a_2475_17214# 0.136f
C14486 m3_1864_16138# a_2966_16186# 0.0302f
C14487 col[7] a_2475_6170# 0.136f
C14488 a_24050_5142# a_25054_5142# 0.843f
C14489 col_n[0] a_3366_2492# 0.0283f
C14490 m2_6752_18014# m2_7756_18014# 0.843f
C14491 vcm a_22346_9198# 0.155f
C14492 a_2475_9182# a_1957_9182# 0.0734f
C14493 col[5] a_7986_12170# 0.367f
C14494 vcm a_13006_18194# 0.165f
C14495 a_13918_14178# a_14010_14178# 0.326f
C14496 col[2] a_4882_2130# 0.0682f
C14497 m3_25960_1078# a_26058_2130# 0.0302f
C14498 a_2475_14202# a_25966_14178# 0.264f
C14499 a_2275_14202# a_23350_14218# 0.144f
C14500 VDD a_9902_8154# 0.181f
C14501 row_n[7] a_31078_9158# 0.282f
C14502 m2_3164_13422# rowon_n[11] 0.0322f
C14503 m2_9188_9406# rowon_n[7] 0.0322f
C14504 m2_15212_5390# rowon_n[3] 0.0322f
C14505 col[12] a_14922_14178# 0.0682f
C14506 col_n[14] a_2275_12194# 0.113f
C14507 rowon_n[11] a_30986_13174# 0.118f
C14508 row_n[3] rowoff_n[3] 0.209f
C14509 VDD a_31382_18234# 0.019f
C14510 col_n[19] a_2275_1150# 0.113f
C14511 col_n[20] a_23046_8154# 0.251f
C14512 vcm a_15926_3134# 0.1f
C14513 row_n[9] a_18330_11206# 0.0117f
C14514 a_15014_7150# a_15014_6146# 0.843f
C14515 col_n[27] a_29982_10162# 0.0765f
C14516 vcm a_3270_12210# 0.155f
C14517 a_8898_11166# a_9294_11206# 0.0313f
C14518 a_2275_11190# a_16930_11166# 0.136f
C14519 VDD a_35494_3496# 0.106f
C14520 m2_21812_18014# a_21950_18194# 0.225f
C14521 col[4] a_2275_9182# 0.0899f
C14522 ctop a_16018_7150# 4.11f
C14523 row_n[11] a_8898_13174# 0.0437f
C14524 VDD a_24962_12170# 0.181f
C14525 m2_12776_18014# m3_11904_18146# 0.0341f
C14526 rowon_n[15] a_7986_17190# 0.248f
C14527 m2_30272_14426# rowon_n[12] 0.0322f
C14528 m2_35292_10410# rowon_n[8] 0.0322f
C14529 col_n[11] a_14410_6508# 0.0283f
C14530 a_27974_4138# a_28466_4500# 0.0658f
C14531 a_27062_4138# a_27366_4178# 0.0931f
C14532 row_n[1] a_18938_3134# 0.0437f
C14533 col_n[21] a_24450_18556# 0.0283f
C14534 rowoff_n[1] a_4882_3134# 0.202f
C14535 col[24] a_2475_8178# 0.136f
C14536 vcm a_30986_7150# 0.1f
C14537 rowon_n[5] a_18026_7150# 0.248f
C14538 rowoff_n[12] a_25054_14178# 0.294f
C14539 a_4974_8154# a_5978_8154# 0.843f
C14540 a_2475_8178# a_8990_8154# 0.316f
C14541 vcm a_18330_16226# 0.155f
C14542 a_2275_13198# a_31990_13174# 0.136f
C14543 VDD a_16418_6508# 0.0779f
C14544 sample a_2161_12194# 0.0858f
C14545 ctop a_31078_11166# 4.11f
C14546 a_28978_18194# a_29070_18194# 0.0991f
C14547 VDD a_5886_15182# 0.181f
C14548 col_n[31] a_2275_14202# 0.113f
C14549 m2_34864_4962# m2_34864_3958# 0.843f
C14550 col_n[9] a_12002_6146# 0.251f
C14551 m2_14784_946# m3_15920_1078# 0.0341f
C14552 vcm a_11910_10162# 0.1f
C14553 a_30074_11166# a_30074_10162# 0.843f
C14554 a_2475_10186# a_24050_10162# 0.316f
C14555 col_n[16] a_18938_8154# 0.0765f
C14556 row_n[14] a_29070_16186# 0.282f
C14557 m2_10192_16434# a_9994_16186# 0.165f
C14558 rowoff_n[4] a_5374_6508# 0.0133f
C14559 col[21] a_2275_11190# 0.0899f
C14560 a_23958_15182# a_24354_15222# 0.0313f
C14561 VDD a_31478_10524# 0.0779f
C14562 m2_3740_18014# ctop 0.0422f
C14563 ctop a_12002_14178# 4.11f
C14564 vcm a_2966_4138# 0.56f
C14565 rowoff_n[2] a_14410_4500# 0.0133f
C14566 col_n[9] rowon_n[5] 0.111f
C14567 col_n[6] row_n[4] 0.298f
C14568 col_n[22] row_n[12] 0.298f
C14569 col_n[28] row_n[15] 0.298f
C14570 col_n[15] rowon_n[8] 0.111f
C14571 col_n[19] rowon_n[10] 0.111f
C14572 col_n[18] row_n[10] 0.298f
C14573 sample row_n[0] 0.425f
C14574 col_n[27] rowon_n[14] 0.111f
C14575 a_7986_7150# a_8290_7190# 0.0931f
C14576 col_n[23] rowon_n[12] 0.111f
C14577 a_8898_7150# a_9390_7512# 0.0658f
C14578 col_n[26] row_n[14] 0.298f
C14579 rowoff_n[10] a_31478_12532# 0.0133f
C14580 col_n[13] rowon_n[7] 0.111f
C14581 col_n[11] rowon_n[6] 0.111f
C14582 col_n[0] rowon_n[0] 0.111f
C14583 col_n[2] row_n[2] 0.298f
C14584 col_n[10] row_n[6] 0.298f
C14585 col_n[30] col_n[31] 0.0125f
C14586 col_n[12] row_n[7] 0.298f
C14587 a_2275_7174# a_15014_7150# 0.399f
C14588 VDD sw 0.276f
C14589 col_n[21] rowon_n[11] 0.111f
C14590 col_n[7] rowon_n[4] 0.111f
C14591 vcm row_n[1] 0.616f
C14592 col_n[3] rowon_n[2] 0.111f
C14593 col_n[4] row_n[3] 0.298f
C14594 col_n[24] row_n[13] 0.298f
C14595 col_n[29] rowon_n[15] 0.111f
C14596 col_n[5] rowon_n[3] 0.111f
C14597 col_n[8] row_n[5] 0.298f
C14598 col_n[20] row_n[11] 0.298f
C14599 col_n[1] rowon_n[1] 0.111f
C14600 col_n[17] rowon_n[9] 0.111f
C14601 col_n[25] rowon_n[13] 0.111f
C14602 col_n[14] row_n[8] 0.298f
C14603 col_n[16] row_n[9] 0.298f
C14604 m2_32856_18014# vcm 0.353f
C14605 m2_29268_12418# a_29070_12170# 0.165f
C14606 col_n[10] a_13406_16548# 0.0283f
C14607 row_n[6] a_26362_8194# 0.0117f
C14608 vcm a_26970_14178# 0.1f
C14609 a_20034_12170# a_21038_12170# 0.843f
C14610 col[29] a_32082_5142# 0.367f
C14611 VDD a_23046_4138# 0.483f
C14612 col_n[31] rowoff_n[11] 0.0471f
C14613 VDD a_12402_13536# 0.0779f
C14614 row_n[8] a_16930_10162# 0.0437f
C14615 rowoff_n[0] a_23446_2492# 0.0133f
C14616 rowoff_n[7] a_5978_9158# 0.294f
C14617 col_n[11] a_2475_7174# 0.0531f
C14618 rowon_n[12] a_16018_14178# 0.248f
C14619 a_3878_4138# a_4274_4178# 0.0313f
C14620 a_4882_4138# a_4974_4138# 0.326f
C14621 a_2275_4162# a_5278_4178# 0.144f
C14622 a_2475_4162# a_7894_4138# 0.264f
C14623 m3_15920_18146# ctop 0.209f
C14624 m2_2160_12418# row_n[10] 0.0194f
C14625 rowoff_n[13] a_13006_15182# 0.294f
C14626 a_2275_9182# a_30074_9158# 0.399f
C14627 m2_8184_8402# row_n[6] 0.0128f
C14628 m2_14208_4386# row_n[2] 0.0128f
C14629 col_n[24] a_27366_5182# 0.084f
C14630 rowon_n[2] a_26058_4138# 0.248f
C14631 vcm a_7894_17190# 0.1f
C14632 col_n[8] a_10998_16186# 0.251f
C14633 a_10998_14178# a_10998_13174# 0.843f
C14634 VDD a_3970_7150# 0.483f
C14635 rowoff_n[5] a_15014_7150# 0.294f
C14636 col_n[5] a_7894_6146# 0.0765f
C14637 col[1] a_2475_4162# 0.136f
C14638 a_2275_18218# a_8898_18194# 0.136f
C14639 a_4882_18194# a_5278_18234# 0.0313f
C14640 col_n[15] a_17934_18194# 0.0762f
C14641 VDD a_27462_17552# 0.0779f
C14642 vcm a_9994_2130# 0.56f
C14643 a_2275_6170# a_20338_6186# 0.144f
C14644 a_2475_6170# a_22954_6146# 0.264f
C14645 m2_20232_10410# a_20034_10162# 0.165f
C14646 rowoff_n[3] a_24050_5142# 0.294f
C14647 row_n[2] a_3970_4138# 0.282f
C14648 col_n[15] rowoff_n[12] 0.0471f
C14649 col_n[8] a_2275_10186# 0.113f
C14650 a_23046_11166# a_23350_11206# 0.0931f
C14651 a_23958_11166# a_24450_11528# 0.0658f
C14652 m2_23244_17438# row_n[15] 0.0128f
C14653 m2_29268_13422# row_n[11] 0.0128f
C14654 m2_17796_18014# a_18026_17190# 0.843f
C14655 m2_34864_8978# row_n[7] 0.267f
C14656 VDD a_19030_11166# 0.483f
C14657 col[18] a_21038_3134# 0.367f
C14658 col[28] a_31078_15182# 0.367f
C14659 col[25] a_27974_5142# 0.0682f
C14660 a_2275_3158# a_13918_3134# 0.136f
C14661 a_2475_18218# a_6890_18194# 0.264f
C14662 rowoff_n[1] a_33086_3134# 0.294f
C14663 col_n[28] a_2475_9182# 0.0531f
C14664 a_27062_1126# a_2275_1150# 0.0924f
C14665 row_n[13] a_24354_15222# 0.0117f
C14666 vcm a_25054_6146# 0.56f
C14667 a_2275_8178# a_2275_7174# 0.0715f
C14668 a_19942_8154# a_20034_8154# 0.326f
C14669 rowoff_n[11] a_19430_13536# 0.0133f
C14670 row_n[3] a_35398_5182# 0.0117f
C14671 a_24450_1488# VDD 0.0977f
C14672 col_n[13] a_16322_3174# 0.084f
C14673 col[13] a_2475_17214# 0.136f
C14674 row_n[15] a_14922_17190# 0.0437f
C14675 a_2475_17214# a_16018_17190# 0.316f
C14676 VDD a_34090_15182# 0.483f
C14677 col_n[23] a_26362_15222# 0.084f
C14678 col[18] a_2475_6170# 0.136f
C14679 col_n[4] a_6890_16186# 0.0765f
C14680 m2_1732_1950# m2_2736_1950# 0.843f
C14681 row_n[5] a_24962_7150# 0.0437f
C14682 a_2275_5166# a_28978_5142# 0.136f
C14683 a_14922_5142# a_15318_5182# 0.0313f
C14684 m2_11196_8402# a_10998_8154# 0.165f
C14685 rowon_n[9] a_24050_11166# 0.248f
C14686 col_n[0] rowoff_n[13] 0.0471f
C14687 vcm a_5978_9158# 0.56f
C14688 rowoff_n[15] a_35494_17552# 0.0133f
C14689 col_n[25] a_2275_12194# 0.113f
C14690 col[1] rowoff_n[8] 0.0901f
C14691 col[0] rowoff_n[7] 0.0901f
C14692 col[2] rowoff_n[9] 0.0901f
C14693 ctop rowoff_n[1] 0.177f
C14694 m2_25828_946# a_2475_1150# 0.286f
C14695 a_4882_14178# a_5374_14540# 0.0658f
C14696 a_2275_14202# a_6982_14178# 0.399f
C14697 a_3970_14178# a_4274_14218# 0.0931f
C14698 col_n[30] a_2275_1150# 0.127f
C14699 VDD a_15014_18194# 0.0356f
C14700 a_10998_2130# a_12002_2130# 0.843f
C14701 a_2475_2154# a_21038_2130# 0.316f
C14702 m2_30272_4386# a_30074_4138# 0.165f
C14703 col[17] a_20034_13174# 0.367f
C14704 m2_17220_1374# VDD 0.0194f
C14705 row_n[9] a_2475_11190# 0.405f
C14706 vcm a_30378_4178# 0.155f
C14707 rowoff_n[9] a_25966_11166# 0.202f
C14708 col[14] a_16930_3134# 0.0682f
C14709 m2_1732_13998# vcm 0.316f
C14710 col[15] a_2275_9182# 0.0899f
C14711 col[24] a_26970_15182# 0.0682f
C14712 vcm a_21038_13174# 0.56f
C14713 a_34090_12170# a_34394_12210# 0.0931f
C14714 a_35002_12170# a_35094_12170# 0.0991f
C14715 VDD a_17934_3134# 0.181f
C14716 m2_23820_18014# a_2275_18218# 0.28f
C14717 a_2275_16210# a_22042_16186# 0.399f
C14718 rowon_n[3] a_11910_5142# 0.118f
C14719 a_29070_1126# m2_28840_946# 0.0249f
C14720 col_n[2] a_5278_1166# 0.0839f
C14721 rowoff_n[7] a_35002_9158# 0.202f
C14722 col_n[12] a_15318_13214# 0.084f
C14723 a_2475_4162# a_2475_3158# 0.0666f
C14724 m2_1732_5966# a_1957_6170# 0.245f
C14725 vcm a_11302_7190# 0.155f
C14726 a_29982_9158# a_30378_9198# 0.0313f
C14727 rowoff_n[12] a_7382_14540# 0.0133f
C14728 row_n[10] a_32386_12210# 0.0117f
C14729 ctop a_24050_2130# 4.06f
C14730 vcm a_2475_16210# 1.08f
C14731 a_2475_13198# a_14922_13174# 0.264f
C14732 a_2275_13198# a_12306_13214# 0.144f
C14733 col_n[23] a_26458_7512# 0.0283f
C14734 VDD a_32994_7150# 0.181f
C14735 col_n[5] a_2475_5166# 0.0531f
C14736 m2_19804_18014# a_2475_18218# 0.286f
C14737 a_19942_18194# a_20434_18556# 0.0658f
C14738 a_14922_1126# a_15414_1488# 0.0658f
C14739 row_n[12] a_22954_14178# 0.0437f
C14740 vcm a_4882_1126# 0.0989f
C14741 a_26058_6146# a_27062_6146# 0.843f
C14742 m2_4168_3382# rowon_n[1] 0.0322f
C14743 m2_32856_946# col_n[30] 0.369f
C14744 row_n[2] a_32994_4138# 0.0437f
C14745 vcm a_26362_11206# 0.155f
C14746 col[6] a_8990_11166# 0.367f
C14747 a_2275_10186# a_5886_10162# 0.136f
C14748 col[3] a_5886_1126# 0.0682f
C14749 rowon_n[6] a_32082_8154# 0.248f
C14750 col[13] a_15926_13174# 0.0682f
C14751 ctop a_4974_5142# 4.11f
C14752 m3_1864_3086# a_2966_3134# 0.0302f
C14753 a_2275_15206# a_27366_15222# 0.144f
C14754 a_2475_15206# a_29982_15182# 0.264f
C14755 a_15926_15182# a_16018_15182# 0.326f
C14756 VDD a_13918_10162# 0.181f
C14757 m2_30848_18014# col[28] 0.347f
C14758 col_n[21] a_24050_7150# 0.251f
C14759 col_n[6] ctop 0.0594f
C14760 col_n[30] rowon_n[10] 0.111f
C14761 col_n[20] rowon_n[5] 0.111f
C14762 col_n[15] row_n[3] 0.298f
C14763 col_n[0] col[1] 7.13f
C14764 col_n[16] rowon_n[3] 0.111f
C14765 col_n[28] rowon_n[9] 0.111f
C14766 col_n[9] row_n[0] 0.298f
C14767 col_n[13] row_n[2] 0.298f
C14768 col_n[11] row_n[1] 0.298f
C14769 col_n[19] row_n[5] 0.298f
C14770 col_n[14] rowon_n[2] 0.111f
C14771 col_n[31] row_n[11] 0.298f
C14772 col_n[17] row_n[4] 0.298f
C14773 vcm col[0] 5.46f
C14774 col_n[10] rowon_n[0] 0.111f
C14775 col_n[21] row_n[6] 0.298f
C14776 VDD col[3] 3.83f
C14777 col_n[26] rowon_n[8] 0.111f
C14778 col_n[12] rowon_n[1] 0.111f
C14779 col_n[18] rowon_n[4] 0.111f
C14780 col_n[27] row_n[9] 0.298f
C14781 col_n[29] row_n[10] 0.298f
C14782 col_n[22] rowon_n[6] 0.111f
C14783 col_n[25] row_n[8] 0.298f
C14784 col_n[24] rowon_n[7] 0.111f
C14785 col_n[23] row_n[7] 0.298f
C14786 a_2475_18218# a_35094_18194# 0.0299f
C14787 col_n[28] a_30986_9158# 0.0765f
C14788 col_n[2] a_2275_8178# 0.113f
C14789 m2_34864_11990# rowoff_n[10] 0.278f
C14790 vcm a_19942_5142# 0.1f
C14791 col_n[1] a_4274_11206# 0.084f
C14792 a_17022_8154# a_17022_7150# 0.843f
C14793 rowoff_n[10] a_13918_12170# 0.202f
C14794 a_33086_1126# vcm 0.165f
C14795 sample a_1957_1150# 0.345f
C14796 m2_13204_16434# rowon_n[14] 0.0322f
C14797 row_n[6] a_9994_8154# 0.282f
C14798 m2_19228_12418# rowon_n[10] 0.0322f
C14799 vcm a_7286_14218# 0.155f
C14800 m2_25252_8402# rowon_n[6] 0.0322f
C14801 m2_31276_4386# rowon_n[2] 0.0322f
C14802 a_10906_12170# a_11302_12210# 0.0313f
C14803 a_2275_12194# a_20946_12170# 0.136f
C14804 rowon_n[10] a_9902_12170# 0.118f
C14805 VDD a_5374_4500# 0.0779f
C14806 ctop a_20034_9158# 4.11f
C14807 col_n[22] a_2475_7174# 0.0531f
C14808 VDD a_28978_14178# 0.181f
C14809 col_n[12] a_15414_5504# 0.0283f
C14810 rowon_n[0] a_19942_2130# 0.118f
C14811 col_n[22] a_25454_17552# 0.0283f
C14812 rowoff_n[0] a_5886_2130# 0.202f
C14813 a_29070_5142# a_29374_5182# 0.0931f
C14814 a_29982_5142# a_30474_5504# 0.0658f
C14815 m2_5748_946# ctop 0.0428f
C14816 vcm a_35002_9158# 0.101f
C14817 m2_17796_18014# m2_18224_18442# 0.165f
C14818 rowoff_n[14] a_29982_16186# 0.202f
C14819 a_2475_9182# a_13006_9158# 0.316f
C14820 a_6982_9158# a_7986_9158# 0.843f
C14821 col[7] a_2475_15206# 0.136f
C14822 col_n[0] a_3366_11528# 0.0283f
C14823 col[12] a_2475_4162# 0.136f
C14824 vcm a_22346_18234# 0.16f
C14825 a_2275_14202# a_34394_14218# 0.144f
C14826 VDD a_20434_8516# 0.0779f
C14827 col[2] a_4882_11166# 0.0682f
C14828 VDD a_9902_17190# 0.181f
C14829 a_25966_2130# a_26058_2130# 0.326f
C14830 col_n[10] a_13006_5142# 0.251f
C14831 m3_14916_1078# VDD 0.0157f
C14832 row_n[9] a_30986_11166# 0.0437f
C14833 col_n[19] a_2275_10186# 0.113f
C14834 col_n[26] rowoff_n[12] 0.0471f
C14835 a_2275_6170# a_3970_6146# 0.399f
C14836 col_n[20] a_23046_17190# 0.251f
C14837 rowon_n[13] a_30074_15182# 0.248f
C14838 col_n[17] a_19942_7150# 0.0765f
C14839 rowoff_n[3] a_6378_5504# 0.0133f
C14840 vcm a_15926_12170# 0.1f
C14841 a_32082_12170# a_32082_11166# 0.843f
C14842 a_2475_11190# a_28066_11166# 0.316f
C14843 VDD a_12002_2130# 0.483f
C14844 a_25966_16186# a_26362_16226# 0.0313f
C14845 VDD a_35494_12532# 0.106f
C14846 col[4] a_2275_18218# 0.0899f
C14847 m2_26832_18014# m3_26964_18146# 3.79f
C14848 ctop a_16018_16186# 4.11f
C14849 col[9] a_2275_7174# 0.0899f
C14850 col_n[1] a_4370_3496# 0.0283f
C14851 rowoff_n[1] a_15414_3496# 0.0133f
C14852 m2_34864_17010# rowoff_n[15] 0.278f
C14853 col_n[11] a_14410_15544# 0.0283f
C14854 row_n[13] a_7986_15182# 0.282f
C14855 a_2275_8178# a_19030_8154# 0.399f
C14856 a_9994_8154# a_10298_8194# 0.0931f
C14857 a_10906_8154# a_11398_8516# 0.0658f
C14858 col[30] a_33086_4138# 0.367f
C14859 col[24] a_2475_17214# 0.136f
C14860 vcm a_30986_16186# 0.1f
C14861 a_22042_13174# a_23046_13174# 0.843f
C14862 col[29] a_2475_6170# 0.136f
C14863 VDD a_27062_6146# 0.483f
C14864 row_n[3] a_18026_5142# 0.282f
C14865 rowon_n[7] a_17934_9158# 0.118f
C14866 VDD a_16418_15544# 0.0779f
C14867 rowoff_n[6] a_6982_8154# 0.294f
C14868 m2_2736_1950# row_n[0] 0.269f
C14869 m3_8892_18146# a_8990_17190# 0.0303f
C14870 col_n[10] rowoff_n[13] 0.0471f
C14871 row_n[5] a_5278_7190# 0.0117f
C14872 a_2475_5166# a_11910_5142# 0.264f
C14873 a_2275_5166# a_9294_5182# 0.144f
C14874 a_6890_5142# a_6982_5142# 0.326f
C14875 m2_30848_946# m3_29976_1078# 0.0341f
C14876 col_n[25] a_28370_4178# 0.084f
C14877 col_n[0] a_2475_3158# 0.0532f
C14878 col[13] rowoff_n[9] 0.0901f
C14879 col[5] rowoff_n[1] 0.0901f
C14880 col[6] rowoff_n[2] 0.0901f
C14881 col[11] rowoff_n[7] 0.0901f
C14882 col[4] rowoff_n[0] 0.0901f
C14883 col[7] rowoff_n[3] 0.0901f
C14884 col[12] rowoff_n[8] 0.0901f
C14885 col[8] rowoff_n[4] 0.0901f
C14886 col[9] rowoff_n[5] 0.0901f
C14887 col[10] rowoff_n[6] 0.0901f
C14888 a_2275_10186# a_34090_10162# 0.399f
C14889 rowoff_n[15] a_17934_17190# 0.202f
C14890 col_n[9] a_12002_15182# 0.251f
C14891 col_n[6] a_8898_5142# 0.0765f
C14892 rowoff_n[4] a_16018_6146# 0.294f
C14893 a_13006_15182# a_13006_14178# 0.843f
C14894 VDD a_7986_9158# 0.483f
C14895 col_n[16] a_18938_17190# 0.0765f
C14896 m2_12200_15430# row_n[13] 0.0128f
C14897 col[26] a_2275_9182# 0.0899f
C14898 a_2161_2154# a_2275_2154# 0.183f
C14899 a_2475_2154# a_2966_2130# 0.0299f
C14900 m2_18224_11414# row_n[9] 0.0128f
C14901 m2_24248_7398# row_n[5] 0.0128f
C14902 m2_30272_3382# row_n[1] 0.0128f
C14903 vcm a_14010_4138# 0.56f
C14904 rowoff_n[2] a_25054_4138# 0.294f
C14905 rowon_n[1] a_4974_3134# 0.248f
C14906 a_2275_7174# a_24354_7190# 0.144f
C14907 a_2475_7174# a_26970_7150# 0.264f
C14908 m2_3164_11414# a_2966_11166# 0.165f
C14909 vcm a_2966_13174# 0.56f
C14910 a_25054_12170# a_25358_12210# 0.0931f
C14911 a_25966_12170# a_26458_12532# 0.0658f
C14912 col[19] a_22042_2130# 0.367f
C14913 a_2475_16210# a_4974_16186# 0.316f
C14914 VDD a_23046_13174# 0.483f
C14915 col[29] a_32082_14178# 0.367f
C14916 col[26] a_28978_4138# 0.0682f
C14917 rowoff_n[0] a_34090_2130# 0.294f
C14918 a_2275_4162# a_17934_4138# 0.136f
C14919 m3_34996_6098# ctop 0.209f
C14920 col_n[11] a_2475_16210# 0.0531f
C14921 vcm a_29070_8154# 0.56f
C14922 a_21950_9158# a_22042_9158# 0.326f
C14923 col_n[16] a_2475_5166# 0.0531f
C14924 row_n[10] a_16018_12170# 0.282f
C14925 col_n[14] a_17326_2170# 0.084f
C14926 rowon_n[14] a_15926_16186# 0.118f
C14927 m2_1732_1950# m3_2868_2082# 0.0341f
C14928 col_n[24] a_27366_14218# 0.084f
C14929 row_n[0] a_26058_2130# 0.282f
C14930 VDD a_3970_16186# 0.483f
C14931 col_n[5] a_7894_15182# 0.0765f
C14932 a_2475_1150# a_9994_1126# 0.0299f
C14933 row_n[12] a_3270_14218# 0.0117f
C14934 col[1] a_2475_13198# 0.136f
C14935 rowon_n[4] a_25966_6146# 0.118f
C14936 vcm a_19334_2170# 0.155f
C14937 col[6] a_2475_2154# 0.136f
C14938 a_16930_6146# a_17326_6186# 0.0313f
C14939 a_2275_6170# a_32994_6146# 0.136f
C14940 m2_8760_946# m2_9764_946# 0.843f
C14941 row_n[2] a_13310_4178# 0.0117f
C14942 vcm a_9994_11166# 0.56f
C14943 VDD a_6890_1126# 0.405f
C14944 m2_16216_17438# a_16018_17190# 0.165f
C14945 a_6890_15182# a_7382_15544# 0.0658f
C14946 a_2275_15206# a_10998_15182# 0.399f
C14947 a_5978_15182# a_6282_15222# 0.0931f
C14948 col_n[29] rowon_n[4] 0.111f
C14949 col_n[25] rowon_n[2] 0.111f
C14950 col_n[24] row_n[2] 0.298f
C14951 col_n[5] col[6] 7.13f
C14952 col_n[27] rowon_n[3] 0.111f
C14953 col_n[30] row_n[5] 0.298f
C14954 col_n[21] rowon_n[0] 0.111f
C14955 col_n[20] row_n[0] 0.298f
C14956 col_n[17] ctop 0.0596f
C14957 col_n[15] en_bit_n[1] 0.187f
C14958 VDD col[14] 3.83f
C14959 col_n[31] rowon_n[5] 0.111f
C14960 col_n[26] row_n[3] 0.298f
C14961 vcm col[11] 5.46f
C14962 col_n[22] row_n[1] 0.298f
C14963 col_n[28] row_n[4] 0.298f
C14964 col_n[23] rowon_n[1] 0.111f
C14965 col_n[13] a_2275_8178# 0.113f
C14966 col[18] a_21038_12170# 0.367f
C14967 a_13006_3134# a_14010_3134# 0.843f
C14968 a_2475_3158# a_25054_3134# 0.316f
C14969 rowon_n[8] a_2874_10162# 0.118f
C14970 col[15] a_17934_2130# 0.0682f
C14971 rowoff_n[8] a_26970_10162# 0.202f
C14972 m2_1732_12994# rowoff_n[11] 0.415f
C14973 col[25] a_27974_14178# 0.0682f
C14974 vcm a_35398_6186# 0.161f
C14975 rowoff_n[11] a_30074_13174# 0.294f
C14976 m2_34864_12994# a_35094_13174# 0.0249f
C14977 col_n[0] a_3270_8194# 0.084f
C14978 vcm a_25054_15182# 0.56f
C14979 col[3] a_2275_5166# 0.0899f
C14980 VDD a_21950_5142# 0.181f
C14981 m2_1046_19620# VDD 0.635f
C14982 a_2275_17214# a_26058_17190# 0.399f
C14983 col_n[13] a_16322_12210# 0.084f
C14984 col[18] a_2475_15206# 0.136f
C14985 a_3970_5142# a_3970_4138# 0.843f
C14986 m3_33992_1078# m3_34568_1078# 0.0133f
C14987 col[23] a_2475_4162# 0.136f
C14988 vcm a_15318_9198# 0.155f
C14989 a_31990_10162# a_32386_10202# 0.0313f
C14990 m2_7180_15430# a_6982_15182# 0.165f
C14991 col_n[24] a_27462_6508# 0.0283f
C14992 ctop a_28066_4138# 4.11f
C14993 vcm a_5978_18194# 0.165f
C14994 m2_16792_946# a_16930_1126# 0.225f
C14995 a_2475_14202# a_18938_14178# 0.264f
C14996 a_2275_14202# a_16322_14218# 0.144f
C14997 VDD a_2161_8178# 0.187f
C14998 row_n[7] a_24050_9158# 0.282f
C14999 rowon_n[11] a_23958_13174# 0.118f
C15000 VDD a_24354_18234# 0.019f
C15001 row_n[13] rowoff_n[12] 0.085f
C15002 col_n[30] a_2275_10186# 0.113f
C15003 a_16018_2130# a_16322_2170# 0.0931f
C15004 a_2275_2154# a_31078_2130# 0.399f
C15005 a_16930_2130# a_17422_2492# 0.0658f
C15006 m3_10900_18146# VDD 0.0868f
C15007 vcm a_8898_3134# 0.1f
C15008 row_n[9] a_11302_11206# 0.0117f
C15009 a_28066_7150# a_29070_7150# 0.843f
C15010 col[7] a_9994_10162# 0.367f
C15011 rowon_n[1] a_33998_3134# 0.118f
C15012 m2_26256_11414# a_26058_11166# 0.165f
C15013 vcm a_30378_13214# 0.155f
C15014 col[14] a_16930_12170# 0.0682f
C15015 a_2275_11190# a_9902_11166# 0.136f
C15016 col[15] a_2275_18218# 0.0899f
C15017 VDD a_28466_3496# 0.0779f
C15018 m2_16792_18014# a_17022_18194# 0.0249f
C15019 col[20] a_2275_7174# 0.0899f
C15020 ctop a_8990_7150# 4.11f
C15021 col_n[22] a_25054_6146# 0.251f
C15022 a_2275_16210# a_31382_16226# 0.144f
C15023 a_2475_16210# a_33998_16186# 0.264f
C15024 a_17934_16186# a_18026_16186# 0.326f
C15025 VDD a_17934_12170# 0.181f
C15026 m2_2736_18014# m3_3872_18146# 0.0341f
C15027 m2_2160_14426# rowon_n[12] 0.0219f
C15028 m2_8184_10410# rowon_n[8] 0.0322f
C15029 col_n[29] a_31990_8154# 0.0765f
C15030 m2_14208_6394# rowon_n[4] 0.0322f
C15031 m2_19228_2378# rowon_n[0] 0.0322f
C15032 row_n[1] a_11910_3134# 0.0437f
C15033 col_n[2] a_5278_10202# 0.084f
C15034 rowon_n[5] a_10998_7150# 0.248f
C15035 vcm a_23958_7150# 0.1f
C15036 rowoff_n[12] a_18026_14178# 0.294f
C15037 a_19030_9158# a_19030_8154# 0.843f
C15038 vcm a_11302_16226# 0.155f
C15039 a_12914_13174# a_13310_13214# 0.0313f
C15040 a_2275_13198# a_24962_13174# 0.136f
C15041 VDD a_9390_6508# 0.0779f
C15042 col_n[13] a_16418_4500# 0.0283f
C15043 ctop a_24050_11166# 4.11f
C15044 col_n[21] rowoff_n[13] 0.0471f
C15045 col_n[23] a_26458_16548# 0.0283f
C15046 VDD a_32994_16186# 0.181f
C15047 col_n[5] a_2475_14202# 0.0531f
C15048 col_n[10] a_2475_3158# 0.0531f
C15049 col[22] rowoff_n[7] 0.0901f
C15050 col[21] rowoff_n[6] 0.0901f
C15051 col[20] rowoff_n[5] 0.0901f
C15052 col[16] rowoff_n[1] 0.0901f
C15053 col[18] rowoff_n[3] 0.0901f
C15054 col[24] rowoff_n[9] 0.0901f
C15055 col[15] rowoff_n[0] 0.0901f
C15056 col[23] rowoff_n[8] 0.0901f
C15057 col[19] rowoff_n[4] 0.0901f
C15058 col[17] rowoff_n[2] 0.0901f
C15059 m2_29268_15430# rowon_n[13] 0.0322f
C15060 m2_34864_10986# rowon_n[9] 0.231f
C15061 a_31078_6146# a_31382_6186# 0.0931f
C15062 a_31990_6146# a_32482_6508# 0.0658f
C15063 m2_5748_946# m3_5880_1078# 3.79f
C15064 m2_17220_9406# a_17022_9158# 0.165f
C15065 vcm a_4882_10162# 0.1f
C15066 col[1] a_2475_18218# 0.136f
C15067 a_2475_10186# a_17022_10162# 0.316f
C15068 a_8990_10162# a_9994_10162# 0.843f
C15069 row_n[14] a_22042_16186# 0.282f
C15070 col[3] a_5886_10162# 0.0682f
C15071 VDD a_24450_10524# 0.0779f
C15072 ctop a_4974_14178# 4.11f
C15073 row_n[4] a_32082_6146# 0.282f
C15074 col_n[11] a_14010_4138# 0.251f
C15075 a_27974_3134# a_28066_3134# 0.326f
C15076 rowon_n[8] a_31990_10162# 0.118f
C15077 col_n[21] a_24050_16186# 0.251f
C15078 col_n[18] a_20946_6146# 0.0765f
C15079 rowoff_n[10] a_24450_12532# 0.0133f
C15080 a_2275_7174# a_7986_7150# 0.399f
C15081 rowoff_n[2] a_7382_4500# 0.0133f
C15082 col_n[28] a_30986_18194# 0.0762f
C15083 col_n[2] a_2275_17214# 0.113f
C15084 m2_18800_18014# vcm 0.353f
C15085 row_n[6] a_19334_8194# 0.0117f
C15086 vcm a_19942_14178# 0.1f
C15087 col_n[7] a_2275_6170# 0.113f
C15088 a_2475_12194# a_32082_12170# 0.316f
C15089 a_34090_13174# a_34090_12170# 0.843f
C15090 VDD a_16018_4138# 0.483f
C15091 sample a_1957_10186# 0.345f
C15092 col_n[5] rowoff_n[14] 0.0471f
C15093 a_27974_17190# a_28370_17230# 0.0313f
C15094 row_n[0] m2_34864_1950# 0.267f
C15095 VDD a_5374_13536# 0.0779f
C15096 col[8] rowoff_n[10] 0.0901f
C15097 row_n[8] a_9902_10162# 0.0437f
C15098 col_n[2] a_5374_2492# 0.0283f
C15099 rowoff_n[0] a_16418_2492# 0.0133f
C15100 col_n[22] a_2475_16210# 0.0531f
C15101 col_n[12] a_15414_14540# 0.0283f
C15102 rowon_n[12] a_8990_14178# 0.248f
C15103 col_n[27] a_2475_5166# 0.0531f
C15104 m2_28840_946# ctop 0.0428f
C15105 m2_8184_7398# a_7986_7150# 0.165f
C15106 col[31] a_34090_3134# 0.367f
C15107 a_2275_9182# a_23046_9158# 0.399f
C15108 a_12002_9158# a_12306_9198# 0.0931f
C15109 a_12914_9158# a_13406_9520# 0.0658f
C15110 rowoff_n[13] a_5978_15182# 0.294f
C15111 rowon_n[2] a_19030_4138# 0.248f
C15112 vcm a_35002_18194# 0.101f
C15113 a_24050_14178# a_25054_14178# 0.843f
C15114 VDD a_31078_8154# 0.483f
C15115 rowoff_n[5] a_7986_7150# 0.294f
C15116 col[12] a_2475_13198# 0.136f
C15117 col[17] a_2475_2154# 0.136f
C15118 VDD a_20434_17552# 0.0779f
C15119 m2_27260_3382# a_27062_3134# 0.165f
C15120 vcm a_2874_2130# 0.101f
C15121 col_n[26] a_29374_3174# 0.084f
C15122 a_8898_6146# a_8990_6146# 0.326f
C15123 a_2475_6170# a_15926_6146# 0.264f
C15124 a_2275_6170# a_13310_6186# 0.144f
C15125 col_n[10] a_13006_14178# 0.251f
C15126 rowoff_n[3] a_17022_5142# 0.294f
C15127 col_n[7] a_9902_4138# 0.0765f
C15128 vcm col[22] 5.46f
C15129 col_n[11] col[11] 0.489f
C15130 col_n[31] row_n[0] 0.297f
C15131 VDD col[25] 3.83f
C15132 col_n[28] ctop 0.0596f
C15133 rowon_n[8] rowon_n[7] 0.0632f
C15134 m2_1732_17010# a_2475_17214# 0.139f
C15135 m2_1732_12994# row_n[11] 0.292f
C15136 col_n[17] a_19942_16186# 0.0765f
C15137 col_n[24] a_2275_8178# 0.113f
C15138 m2_7180_9406# row_n[7] 0.0128f
C15139 m2_13204_5390# row_n[3] 0.0128f
C15140 row_n[11] a_30074_13174# 0.282f
C15141 a_15014_16186# a_15014_15182# 0.843f
C15142 VDD a_12002_11166# 0.483f
C15143 rowon_n[15] a_29982_17190# 0.118f
C15144 a_2275_3158# a_6890_3134# 0.136f
C15145 rowoff_n[1] a_26058_3134# 0.294f
C15146 col[9] a_2275_16210# 0.0899f
C15147 row_n[13] a_17326_15222# 0.0117f
C15148 vcm a_18026_6146# 0.56f
C15149 rowoff_n[11] a_12402_13536# 0.0133f
C15150 a_2275_8178# a_28370_8194# 0.144f
C15151 col[14] a_2275_5166# 0.0899f
C15152 col_n[1] a_4370_12532# 0.0283f
C15153 a_2475_8178# a_30986_8154# 0.264f
C15154 m3_34996_3086# m2_34864_1950# 0.0341f
C15155 a_27974_13174# a_28466_13536# 0.0658f
C15156 a_27062_13174# a_27366_13214# 0.0931f
C15157 VDD a_3878_5142# 0.181f
C15158 col[30] a_33086_13174# 0.367f
C15159 row_n[3] a_27366_5182# 0.0117f
C15160 row_n[15] a_7894_17190# 0.0437f
C15161 col[27] a_29982_3134# 0.0682f
C15162 m2_28264_14426# row_n[12] 0.0128f
C15163 a_2475_17214# a_8990_17190# 0.316f
C15164 a_4974_17190# a_5978_17190# 0.843f
C15165 m2_34288_10410# row_n[8] 0.0128f
C15166 col[29] a_2475_15206# 0.136f
C15167 VDD a_27062_15182# 0.483f
C15168 a_2275_5166# a_21950_5142# 0.136f
C15169 row_n[5] a_17934_7150# 0.0437f
C15170 rowon_n[9] a_17022_11166# 0.248f
C15171 a_24962_1126# a_25358_1166# 0.0313f
C15172 vcm a_33086_10162# 0.56f
C15173 col_n[15] a_18330_1166# 0.0572f
C15174 rowoff_n[15] a_28466_17552# 0.0133f
C15175 a_23958_10162# a_24050_10162# 0.326f
C15176 col_n[25] a_28370_13214# 0.084f
C15177 col_n[0] a_2475_12194# 0.0532f
C15178 m2_27836_946# a_28066_2130# 0.843f
C15179 m2_8760_946# a_2275_1150# 0.28f
C15180 col_n[4] a_2475_1150# 0.0531f
C15181 col_n[6] a_8898_14178# 0.0765f
C15182 VDD a_7986_18194# 0.0356f
C15183 a_25054_3134# a_25054_2130# 0.843f
C15184 a_2475_2154# a_14010_2130# 0.316f
C15185 vcm a_23350_4178# 0.155f
C15186 a_18938_7150# a_19334_7190# 0.0313f
C15187 rowoff_n[9] a_18938_11166# 0.202f
C15188 col[26] a_2275_18218# 0.0899f
C15189 col[31] a_2275_7174# 0.0899f
C15190 vcm a_14010_13174# 0.56f
C15191 VDD a_10906_3134# 0.181f
C15192 m2_9764_18014# a_2275_18218# 0.28f
C15193 m2_3740_18014# a_4274_18234# 0.087f
C15194 a_7986_16186# a_8290_16226# 0.0931f
C15195 a_8898_16186# a_9390_16548# 0.0658f
C15196 a_2275_16210# a_15014_16186# 0.399f
C15197 rowon_n[3] a_4882_5142# 0.118f
C15198 col[19] a_22042_11166# 0.367f
C15199 col[16] a_18938_1126# 0.0699f
C15200 rowoff_n[7] a_27974_9158# 0.202f
C15201 a_15014_4138# a_16018_4138# 0.843f
C15202 a_2475_4162# a_29070_4138# 0.316f
C15203 col[26] a_28978_13174# 0.0682f
C15204 col_n[1] a_2275_4162# 0.113f
C15205 m3_34568_1078# ctop 0.358f
C15206 vcm a_4274_7190# 0.155f
C15207 rowoff_n[13] a_35002_15182# 0.202f
C15208 row_n[10] a_25358_12210# 0.0117f
C15209 ctop a_17022_2130# 4.06f
C15210 vcm a_29070_17190# 0.56f
C15211 a_2275_13198# a_5278_13214# 0.144f
C15212 a_3878_13174# a_4274_13214# 0.0313f
C15213 a_2475_13198# a_7894_13174# 0.264f
C15214 a_4882_13174# a_4974_13174# 0.326f
C15215 VDD a_25966_7150# 0.181f
C15216 col_n[16] a_2475_14202# 0.0531f
C15217 col_n[21] a_2475_3158# 0.0531f
C15218 col_n[14] a_17326_11206# 0.084f
C15219 col[28] rowoff_n[2] 0.0901f
C15220 col[30] rowoff_n[4] 0.0901f
C15221 col[26] rowoff_n[0] 0.0901f
C15222 sample_n rowoff_n[6] 0.14f
C15223 col[29] rowoff_n[3] 0.0901f
C15224 col[31] rowoff_n[5] 0.0901f
C15225 col[27] rowoff_n[1] 0.0901f
C15226 a_2275_18218# a_30074_18194# 0.0924f
C15227 m2_5748_18014# a_2475_18218# 0.286f
C15228 row_n[12] a_15926_14178# 0.0437f
C15229 a_2275_1150# a_20034_1126# 0.399f
C15230 col[12] a_2475_18218# 0.136f
C15231 vcm a_31990_2130# 0.1f
C15232 a_5978_6146# a_5978_5142# 0.843f
C15233 m2_1732_8978# a_2966_9158# 0.843f
C15234 col_n[25] a_28466_5504# 0.0283f
C15235 col[6] a_2475_11190# 0.136f
C15236 row_n[2] a_25966_4138# 0.0437f
C15237 vcm a_19334_11206# 0.155f
C15238 VDD a_17422_1488# 0.0977f
C15239 rowon_n[6] a_25054_8154# 0.248f
C15240 ctop a_32082_6146# 4.11f
C15241 a_2475_15206# a_22954_15182# 0.264f
C15242 a_2275_15206# a_20338_15222# 0.144f
C15243 VDD a_6890_10162# 0.181f
C15244 a_18026_3134# a_18330_3174# 0.0931f
C15245 a_2275_3158# a_35094_3134# 0.0924f
C15246 a_18938_3134# a_19430_3496# 0.0658f
C15247 a_2475_18218# a_28066_18194# 0.0299f
C15248 col_n[13] a_2275_17214# 0.113f
C15249 col[8] a_10998_9158# 0.367f
C15250 col_n[18] a_2275_6170# 0.113f
C15251 vcm a_12914_5142# 0.1f
C15252 a_30074_8154# a_31078_8154# 0.843f
C15253 rowoff_n[10] a_6890_12170# 0.202f
C15254 col[15] a_17934_11166# 0.0682f
C15255 col_n[16] rowoff_n[14] 0.0471f
C15256 a_26058_1126# vcm 0.165f
C15257 m2_34864_11990# a_2275_12194# 0.278f
C15258 row_n[6] a_2874_8154# 0.0436f
C15259 vcm a_35398_15222# 0.161f
C15260 m2_3164_4386# rowon_n[2] 0.0322f
C15261 a_2275_12194# a_13918_12170# 0.136f
C15262 col_n[23] a_26058_5142# 0.251f
C15263 VDD a_32482_5504# 0.0779f
C15264 rowon_n[10] a_2161_12194# 0.0177f
C15265 m2_22816_18014# VDD 1.1f
C15266 col_n[0] a_3270_17230# 0.084f
C15267 col[19] rowoff_n[10] 0.0901f
C15268 ctop a_13006_9158# 4.11f
C15269 a_2275_17214# a_2275_16210# 0.0715f
C15270 a_19942_17190# a_20034_17190# 0.326f
C15271 col_n[30] a_32994_7150# 0.0765f
C15272 col[3] a_2275_14202# 0.0899f
C15273 VDD a_21950_14178# 0.181f
C15274 col[8] a_2275_3158# 0.0899f
C15275 rowon_n[0] a_12914_2130# 0.118f
C15276 col_n[3] a_6282_9198# 0.084f
C15277 m2_16792_946# col_n[14] 0.331f
C15278 m2_10768_18014# m2_11196_18442# 0.165f
C15279 vcm a_27974_9158# 0.1f
C15280 a_21038_10162# a_21038_9158# 0.843f
C15281 a_2966_9158# a_3270_9198# 0.0931f
C15282 a_3878_9158# a_4370_9520# 0.0658f
C15283 rowoff_n[14] a_22954_16186# 0.202f
C15284 a_2475_9182# a_5978_9158# 0.316f
C15285 col[23] a_2475_13198# 0.136f
C15286 col_n[14] a_17422_3496# 0.0283f
C15287 vcm a_15318_18234# 0.16f
C15288 m3_28972_1078# a_29070_2130# 0.0302f
C15289 m2_12200_17438# rowon_n[15] 0.0322f
C15290 col[28] a_2475_2154# 0.136f
C15291 a_14922_14178# a_15318_14218# 0.0313f
C15292 a_2275_14202# a_28978_14178# 0.136f
C15293 row_n[7] a_33390_9198# 0.0117f
C15294 VDD a_13406_8516# 0.0779f
C15295 m2_18224_13422# rowon_n[11] 0.0322f
C15296 col_n[24] a_27462_15544# 0.0283f
C15297 m2_24248_9406# rowon_n[7] 0.0322f
C15298 m2_30272_5390# rowon_n[3] 0.0322f
C15299 ctop a_28066_13174# 4.11f
C15300 VDD a_2161_17214# 0.187f
C15301 rowon_n[15] col[1] 0.0323f
C15302 row_n[12] ctop 0.186f
C15303 rowon_n[5] row_n[5] 18.9f
C15304 vcm rowoff_n[15] 0.535f
C15305 row_n[9] a_23958_11166# 0.0437f
C15306 row_n[15] col[0] 0.0322f
C15307 col_n[16] col[17] 7.13f
C15308 m2_1732_7974# m2_1732_6970# 0.843f
C15309 a_33998_7150# a_34490_7512# 0.0658f
C15310 a_33086_7150# a_33390_7190# 0.0931f
C15311 rowon_n[13] a_23046_15182# 0.248f
C15312 m2_34864_10986# a_35002_11166# 0.225f
C15313 vcm a_8898_12170# 0.1f
C15314 a_10998_11166# a_12002_11166# 0.843f
C15315 a_2475_11190# a_21038_11166# 0.316f
C15316 col[3] rowoff_n[11] 0.0901f
C15317 VDD a_4974_2130# 0.483f
C15318 m2_9764_18014# col_n[7] 0.243f
C15319 col[4] a_6890_9158# 0.0682f
C15320 m2_22816_18014# a_23350_18234# 0.087f
C15321 rowon_n[3] a_33086_5142# 0.248f
C15322 VDD a_28466_12532# 0.0779f
C15323 col_n[12] a_15014_3134# 0.251f
C15324 m2_17796_18014# m3_16924_18146# 0.0341f
C15325 ctop a_8990_16186# 4.11f
C15326 col[20] a_2275_16210# 0.0899f
C15327 col_n[22] a_25054_15182# 0.251f
C15328 col_n[19] a_21950_5142# 0.0765f
C15329 col[25] a_2275_5166# 0.0899f
C15330 a_29982_4138# a_30074_4138# 0.326f
C15331 rowoff_n[1] a_8386_3496# 0.0133f
C15332 col_n[29] a_31990_17190# 0.0765f
C15333 a_2275_8178# a_12002_8154# 0.399f
C15334 col_n[0] a_2966_9158# 0.251f
C15335 vcm a_23958_16186# 0.1f
C15336 a_2475_13198# a_2475_12194# 0.0666f
C15337 VDD a_20034_6146# 0.483f
C15338 row_n[3] a_10998_5142# 0.282f
C15339 rowon_n[7] a_10906_9158# 0.118f
C15340 col_n[3] a_6378_1488# 0.0283f
C15341 a_29982_18194# a_30378_18234# 0.0313f
C15342 VDD a_9390_15544# 0.0779f
C15343 col_n[13] a_16418_13536# 0.0283f
C15344 a_2475_5166# a_4882_5142# 0.264f
C15345 a_2275_5166# a_3878_5142# 0.136f
C15346 a_2874_5142# a_3366_5504# 0.0658f
C15347 col_n[10] a_2475_12194# 0.0531f
C15348 m2_20808_946# m3_21944_1078# 0.0341f
C15349 m3_29976_18146# m3_30980_18146# 0.202f
C15350 a_2275_10186# a_27062_10162# 0.399f
C15351 a_14922_10162# a_15414_10524# 0.0658f
C15352 rowoff_n[15] a_10906_17190# 0.202f
C15353 a_14010_10162# a_14314_10202# 0.0931f
C15354 col_n[15] a_2475_1150# 0.0486f
C15355 row_n[14] a_31382_16226# 0.0117f
C15356 m2_13204_16434# a_13006_16186# 0.165f
C15357 rowoff_n[4] a_8990_6146# 0.294f
C15358 a_26058_15182# a_27062_15182# 0.843f
C15359 col_n[1] a_3970_1126# 0.303f
C15360 col_n[27] a_30378_2170# 0.084f
C15361 col[0] a_2475_9182# 0.148f
C15362 m2_2160_3382# row_n[1] 0.0194f
C15363 col_n[11] a_14010_13174# 0.251f
C15364 vcm a_6982_4138# 0.56f
C15365 a_2475_7174# a_19942_7150# 0.264f
C15366 rowoff_n[10] a_35094_12170# 0.0135f
C15367 a_10906_7150# a_10998_7150# 0.326f
C15368 col_n[8] a_10906_3134# 0.0765f
C15369 a_2275_7174# a_17326_7190# 0.144f
C15370 rowoff_n[2] a_18026_4138# 0.294f
C15371 m2_32280_12418# a_32082_12170# 0.165f
C15372 row_n[6] a_31990_8154# 0.0437f
C15373 col_n[18] a_20946_15182# 0.0765f
C15374 rowon_n[10] a_31078_12170# 0.248f
C15375 col_n[7] a_2275_15206# 0.113f
C15376 a_17022_17190# a_17022_16186# 0.843f
C15377 VDD a_16018_13174# 0.483f
C15378 col_n[12] a_2275_4162# 0.113f
C15379 rowoff_n[0] a_27062_2130# 0.294f
C15380 a_2275_4162# a_10906_4138# 0.136f
C15381 a_5886_4138# a_6282_4178# 0.0313f
C15382 m3_30980_18146# ctop 0.209f
C15383 col_n[2] a_5374_11528# 0.0283f
C15384 m2_11196_16434# row_n[14] 0.0128f
C15385 m2_17220_12418# row_n[10] 0.0128f
C15386 vcm a_22042_8154# 0.56f
C15387 a_2275_9182# a_32386_9198# 0.144f
C15388 col_n[27] a_2475_14202# 0.0531f
C15389 a_2475_9182# a_35002_9158# 0.264f
C15390 m2_23244_8402# row_n[6] 0.0128f
C15391 m2_29268_4386# row_n[2] 0.0128f
C15392 row_n[10] a_8990_12170# 0.282f
C15393 m2_4168_14426# a_3970_14178# 0.165f
C15394 col[31] a_34090_12170# 0.367f
C15395 m2_1732_17010# sample 0.2f
C15396 col[28] a_30986_2130# 0.0682f
C15397 a_29982_14178# a_30474_14540# 0.0658f
C15398 rowon_n[14] a_8898_16186# 0.118f
C15399 col[2] a_2275_1150# 0.0896f
C15400 a_29070_14178# a_29374_14218# 0.0931f
C15401 m2_34864_10986# ctop 0.0422f
C15402 col[23] a_2475_18218# 0.136f
C15403 row_n[0] a_19030_2130# 0.282f
C15404 VDD a_31078_17190# 0.484f
C15405 a_1957_1150# a_2275_1150# 0.158f
C15406 a_2475_1150# a_2874_1126# 0.264f
C15407 rowon_n[4] a_18938_6146# 0.118f
C15408 m2_34864_2954# a_35398_3174# 0.087f
C15409 col[17] a_2475_11190# 0.136f
C15410 vcm a_12306_2170# 0.155f
C15411 a_2275_6170# a_25966_6146# 0.136f
C15412 m2_23244_10410# a_23046_10162# 0.165f
C15413 row_n[2] a_6282_4178# 0.0117f
C15414 col_n[26] a_29374_12210# 0.084f
C15415 vcm a_2874_11166# 0.1f
C15416 a_25966_11166# a_26058_11166# 0.326f
C15417 VDD a_33998_2130# 0.163f
C15418 col_n[7] a_9902_13174# 0.0765f
C15419 a_2275_15206# a_3970_15182# 0.399f
C15420 col_n[24] a_2275_17214# 0.113f
C15421 col_n[29] a_2275_6170# 0.113f
C15422 col_n[27] rowoff_n[14] 0.0471f
C15423 a_27062_4138# a_27062_3134# 0.843f
C15424 a_2475_3158# a_18026_3134# 0.316f
C15425 rowoff_n[8] a_19942_10162# 0.202f
C15426 a_31990_1126# a_2475_1150# 0.264f
C15427 a_29374_1166# a_2275_1150# 0.145f
C15428 row_n[13] a_29982_15182# 0.0437f
C15429 vcm a_27366_6186# 0.155f
C15430 rowoff_n[11] a_23046_13174# 0.294f
C15431 a_20946_8154# a_21342_8194# 0.0313f
C15432 col[30] rowoff_n[10] 0.0901f
C15433 vcm a_18026_15182# 0.56f
C15434 col[14] a_2275_14202# 0.0899f
C15435 VDD a_14922_5142# 0.181f
C15436 a_28066_1126# VDD 0.035f
C15437 col[19] a_2275_3158# 0.0899f
C15438 col[20] a_23046_10162# 0.367f
C15439 a_2275_17214# a_19030_17190# 0.399f
C15440 a_9994_17190# a_10298_17230# 0.0931f
C15441 a_10906_17190# a_11398_17552# 0.0658f
C15442 VDD a_3878_14178# 0.181f
C15443 rowoff_n[6] a_28978_8154# 0.202f
C15444 col[27] a_29982_12170# 0.0682f
C15445 a_17022_5142# a_18026_5142# 0.843f
C15446 a_2475_5166# a_33086_5142# 0.316f
C15447 m2_14208_8402# a_14010_8154# 0.165f
C15448 m3_19936_1078# m3_20940_1078# 0.202f
C15449 vcm a_8290_9198# 0.155f
C15450 ctop a_21038_4138# 4.11f
C15451 m2_31852_946# a_2275_1150# 0.28f
C15452 m2_11772_946# a_12002_1126# 0.0249f
C15453 col_n[15] a_18330_10202# 0.084f
C15454 a_2475_14202# a_11910_14178# 0.264f
C15455 a_6890_14178# a_6982_14178# 0.326f
C15456 a_2275_14202# a_9294_14218# 0.144f
C15457 VDD a_29982_9158# 0.181f
C15458 row_n[7] a_17022_9158# 0.282f
C15459 rowon_n[11] a_16930_13174# 0.118f
C15460 rowon_n[10] col[2] 0.0323f
C15461 col_n[22] col[22] 0.489f
C15462 row_n[15] col[11] 0.0342f
C15463 rowon_n[11] col[4] 0.0323f
C15464 rowon_n[9] col[0] 0.0318f
C15465 col_n[11] rowoff_n[15] 0.0471f
C15466 row_n[14] col[9] 0.0342f
C15467 rowon_n[13] col[8] 0.0323f
C15468 rowon_n[14] col[10] 0.0323f
C15469 rowon_n[12] col[6] 0.0323f
C15470 rowon_n[15] col[12] 0.0323f
C15471 row_n[11] col[3] 0.0342f
C15472 row_n[12] col[5] 0.0342f
C15473 row_n[10] col[1] 0.0342f
C15474 rowon_n[6] ctop 0.203f
C15475 row_n[13] col[7] 0.0342f
C15476 col_n[4] a_2475_10186# 0.0531f
C15477 VDD a_17326_18234# 0.019f
C15478 a_2275_2154# a_24050_2130# 0.399f
C15479 m2_33284_4386# a_33086_4138# 0.165f
C15480 m2_26256_1374# VDD 0.0194f
C15481 vcm a_34394_4178# 0.155f
C15482 row_n[9] a_4274_11206# 0.0117f
C15483 col_n[26] a_29470_4500# 0.0283f
C15484 rowon_n[1] a_26970_3134# 0.118f
C15485 col[14] rowoff_n[11] 0.0901f
C15486 a_7986_7150# a_7986_6146# 0.843f
C15487 rowoff_n[9] a_29470_11528# 0.0133f
C15488 vcm a_23350_13214# 0.155f
C15489 a_2161_11190# a_2275_11190# 0.183f
C15490 a_2475_11190# a_2966_11166# 0.317f
C15491 VDD a_21438_3496# 0.0779f
C15492 col[31] a_2275_16210# 0.0899f
C15493 ctop a_2475_7174# 0.0488f
C15494 a_2275_16210# a_24354_16226# 0.144f
C15495 a_2475_16210# a_26970_16186# 0.264f
C15496 VDD a_10906_12170# 0.181f
C15497 col[9] a_12002_8154# 0.367f
C15498 a_20946_4138# a_21438_4500# 0.0658f
C15499 a_20034_4138# a_20338_4178# 0.0931f
C15500 row_n[1] a_4882_3134# 0.0437f
C15501 m2_5172_6394# a_4974_6146# 0.165f
C15502 col[16] a_18938_10162# 0.0682f
C15503 rowon_n[5] a_3970_7150# 0.248f
C15504 vcm a_16930_7150# 0.1f
C15505 a_32082_9158# a_33086_9158# 0.843f
C15506 rowoff_n[12] a_10998_14178# 0.294f
C15507 col_n[1] a_2275_13198# 0.113f
C15508 col_n[24] a_27062_4138# 0.251f
C15509 col_n[6] a_2275_2154# 0.113f
C15510 vcm a_4274_16226# 0.155f
C15511 a_2275_13198# a_17934_13174# 0.136f
C15512 VDD a_1957_6170# 0.196f
C15513 col_n[31] a_33998_6146# 0.0765f
C15514 ctop a_17022_11166# 4.11f
C15515 a_21950_18194# a_22042_18194# 0.0991f
C15516 VDD a_25966_16186# 0.181f
C15517 col_n[4] a_7286_8194# 0.084f
C15518 col[0] a_2966_6146# 0.367f
C15519 a_16930_1126# a_17022_1126# 0.0991f
C15520 col_n[21] a_2475_12194# 0.0531f
C15521 a_31382_1166# col_n[28] 0.0839f
C15522 col_n[26] a_2475_1150# 0.0531f
C15523 m2_1732_15002# rowon_n[13] 0.236f
C15524 m2_7180_11414# rowon_n[9] 0.0322f
C15525 m2_13204_7398# rowon_n[5] 0.0322f
C15526 m2_19228_3382# rowon_n[1] 0.0322f
C15527 m2_31852_946# m2_32856_946# 0.843f
C15528 vcm a_31990_11166# 0.1f
C15529 col_n[15] a_18426_2492# 0.0283f
C15530 a_23046_11166# a_23046_10162# 0.843f
C15531 a_2475_10186# a_9994_10162# 0.316f
C15532 row_n[14] a_15014_16186# 0.282f
C15533 col_n[25] a_28466_14540# 0.0283f
C15534 a_16930_15182# a_17326_15222# 0.0313f
C15535 a_2275_15206# a_32994_15182# 0.136f
C15536 VDD a_17422_10524# 0.0779f
C15537 col[11] a_2475_9182# 0.136f
C15538 ctop a_32082_15182# 4.11f
C15539 row_n[4] a_25054_6146# 0.282f
C15540 rowon_n[8] a_24962_10162# 0.118f
C15541 rowoff_n[10] a_17422_12532# 0.0133f
C15542 m2_4744_18014# vcm 0.353f
C15543 m2_28264_16434# rowon_n[14] 0.0322f
C15544 col_n[18] a_2275_15206# 0.113f
C15545 m2_34288_12418# rowon_n[10] 0.0322f
C15546 col[5] a_7894_8154# 0.0682f
C15547 row_n[6] a_12306_8194# 0.0117f
C15548 vcm a_12914_14178# 0.1f
C15549 a_13006_12170# a_14010_12170# 0.843f
C15550 a_2475_12194# a_25054_12170# 0.316f
C15551 VDD a_8990_4138# 0.483f
C15552 col_n[23] a_2275_4162# 0.113f
C15553 a_31990_1126# col[29] 0.0682f
C15554 col_n[13] a_16018_2130# 0.251f
C15555 col_n[23] a_26058_14178# 0.251f
C15556 VDD a_32482_14540# 0.0779f
C15557 col_n[20] a_22954_4138# 0.0765f
C15558 row_n[8] a_2161_10186# 0.0221f
C15559 rowoff_n[0] a_9390_2492# 0.0133f
C15560 col_n[30] a_32994_16186# 0.0765f
C15561 rowon_n[12] a_2475_14202# 0.31f
C15562 a_31990_5142# a_32082_5142# 0.326f
C15563 col[8] a_2275_12194# 0.0899f
C15564 col_n[3] a_6282_18234# 0.084f
C15565 m2_1732_6970# a_2275_7174# 0.191f
C15566 col[13] a_2275_1150# 0.0899f
C15567 a_2275_9182# a_16018_9158# 0.399f
C15568 rowoff_n[14] a_33486_16548# 0.0133f
C15569 rowon_n[2] a_12002_4138# 0.248f
C15570 vcm a_27974_18194# 0.101f
C15571 a_3970_14178# a_3970_13174# 0.843f
C15572 VDD a_24050_8154# 0.483f
C15573 col_n[14] a_17422_12532# 0.0283f
C15574 col[28] a_2475_11190# 0.136f
C15575 VDD a_13406_17552# 0.0779f
C15576 a_26970_2130# a_27366_2170# 0.0313f
C15577 m3_29976_1078# VDD 0.0157f
C15578 vcm a_30074_3134# 0.56f
C15579 a_2475_6170# a_8898_6146# 0.264f
C15580 a_2275_6170# a_6282_6186# 0.144f
C15581 rowoff_n[3] a_9994_5142# 0.294f
C15582 a_16018_11166# a_16322_11206# 0.0931f
C15583 a_2275_11190# a_31078_11166# 0.399f
C15584 a_16930_11166# a_17422_11528# 0.0658f
C15585 m2_1732_6970# rowoff_n[5] 0.415f
C15586 row_n[11] a_23046_13174# 0.282f
C15587 a_28066_16186# a_29070_16186# 0.843f
C15588 VDD a_4974_11166# 0.483f
C15589 m2_31852_18014# m3_31984_18146# 3.79f
C15590 col[4] a_6890_18194# 0.0682f
C15591 rowon_n[15] a_22954_17190# 0.118f
C15592 col_n[12] a_15014_12170# 0.251f
C15593 m2_26832_946# col_n[24] 0.331f
C15594 a_35002_4138# a_35398_4178# 0.0313f
C15595 col_n[9] a_11910_2130# 0.0765f
C15596 rowoff_n[1] a_19030_3134# 0.294f
C15597 row_n[1] a_33086_3134# 0.282f
C15598 row_n[13] a_10298_15222# 0.0117f
C15599 col[25] a_2275_14202# 0.0899f
C15600 rowon_n[5] a_32994_7150# 0.118f
C15601 col_n[19] a_21950_14178# 0.0765f
C15602 vcm a_10998_6146# 0.56f
C15603 a_2275_8178# a_21342_8194# 0.144f
C15604 rowoff_n[11] a_5374_13536# 0.0133f
C15605 a_12914_8154# a_13006_8154# 0.326f
C15606 a_2475_8178# a_23958_8154# 0.264f
C15607 col[30] a_2275_3158# 0.0899f
C15608 m2_24824_18014# col[22] 0.347f
C15609 row_n[3] a_20338_5182# 0.0117f
C15610 m2_6176_10410# row_n[8] 0.0128f
C15611 VDD a_20034_15182# 0.483f
C15612 m2_12200_6394# row_n[4] 0.0128f
C15613 m2_17220_2378# row_n[0] 0.0128f
C15614 col_n[3] a_6378_10524# 0.0283f
C15615 m3_11904_18146# a_12002_17190# 0.0303f
C15616 a_7894_5142# a_8290_5182# 0.0313f
C15617 row_n[5] a_10906_7150# 0.0437f
C15618 a_2275_5166# a_14922_5142# 0.136f
C15619 m3_34996_10114# m3_34996_9110# 0.202f
C15620 m2_34864_8978# a_34090_9158# 0.843f
C15621 rowon_n[9] a_9994_11166# 0.248f
C15622 vcm a_26058_10162# 0.56f
C15623 a_2966_10162# a_2966_9158# 0.843f
C15624 rowoff_n[15] a_21438_17552# 0.0133f
C15625 ctop a_2966_4138# 4.06f
C15626 row_n[9] col[10] 0.0342f
C15627 rowon_n[5] col[3] 0.0323f
C15628 rowon_n[7] col[7] 0.0323f
C15629 rowon_n[12] col[17] 0.0323f
C15630 row_n[6] col[4] 0.0342f
C15631 rowon_n[10] col[13] 0.0323f
C15632 row_n[7] col[6] 0.0342f
C15633 rowon_n[9] col[11] 0.0323f
C15634 rowon_n[11] col[15] 0.0323f
C15635 rowon_n[13] col[19] 0.0323f
C15636 col_n[15] a_2475_10186# 0.0531f
C15637 rowon_n[6] col[5] 0.0323f
C15638 row_n[5] col[2] 0.0342f
C15639 rowon_n[4] col[1] 0.0323f
C15640 row_n[8] col[8] 0.0342f
C15641 row_n[13] col[18] 0.0342f
C15642 col_n[22] rowoff_n[15] 0.0471f
C15643 rowon_n[8] col[9] 0.0323f
C15644 rowon_n[15] col[23] 0.0323f
C15645 row_n[4] col[0] 0.0322f
C15646 row_n[15] col[22] 0.0342f
C15647 row_n[10] col[12] 0.0342f
C15648 row_n[12] col[16] 0.0342f
C15649 row_n[11] col[14] 0.0342f
C15650 row_n[14] col[20] 0.0342f
C15651 row_n[1] ctop 0.186f
C15652 col_n[27] col[28] 7.08f
C15653 rowon_n[14] col[21] 0.0323f
C15654 a_31078_15182# a_31382_15222# 0.0931f
C15655 a_31990_15182# a_32482_15544# 0.0658f
C15656 m2_32856_18014# ctop 0.0422f
C15657 col[25] rowoff_n[11] 0.0901f
C15658 a_3970_2130# a_4974_2130# 0.843f
C15659 a_2475_2154# a_6982_2130# 0.316f
C15660 m2_27260_15430# row_n[13] 0.0128f
C15661 m2_33284_11414# row_n[9] 0.0128f
C15662 vcm a_16322_4178# 0.155f
C15663 col_n[27] a_30378_11206# 0.084f
C15664 rowoff_n[9] a_11910_11166# 0.202f
C15665 a_2275_7174# a_29982_7150# 0.136f
C15666 col_n[1] a_3970_10162# 0.251f
C15667 col[5] a_2475_7174# 0.136f
C15668 vcm a_6982_13174# 0.56f
C15669 col_n[8] a_10906_12170# 0.0765f
C15670 a_27974_12170# a_28066_12170# 0.326f
C15671 VDD a_3366_3496# 0.0779f
C15672 a_2275_16210# a_7986_16186# 0.399f
C15673 row_n[8] a_31078_10162# 0.282f
C15674 rowoff_n[7] a_20946_9158# 0.202f
C15675 rowon_n[12] a_30986_14178# 0.118f
C15676 col_n[12] a_2275_13198# 0.113f
C15677 a_29070_5142# a_29070_4138# 0.843f
C15678 a_2475_4162# a_22042_4138# 0.316f
C15679 m3_6884_1078# ctop 0.21f
C15680 col_n[17] a_2275_2154# 0.113f
C15681 vcm a_31382_8194# 0.155f
C15682 rowoff_n[13] a_27974_15182# 0.202f
C15683 a_22954_9158# a_23350_9198# 0.0313f
C15684 row_n[10] a_18330_12210# 0.0117f
C15685 ctop a_9994_2130# 4.06f
C15686 vcm a_22042_17190# 0.56f
C15687 col[21] a_24050_9158# 0.367f
C15688 VDD a_18938_7150# 0.181f
C15689 rowoff_n[5] a_29982_7150# 0.202f
C15690 col[2] a_2275_10186# 0.0899f
C15691 col[28] a_30986_11166# 0.0682f
C15692 col[9] rowoff_n[12] 0.0901f
C15693 a_2275_18218# a_23046_18194# 0.0924f
C15694 a_12914_18194# a_13406_18556# 0.0658f
C15695 row_n[0] a_28370_2170# 0.0117f
C15696 a_7894_1126# a_8386_1488# 0.0658f
C15697 a_2275_1150# a_13006_1126# 0.0924f
C15698 row_n[12] a_8898_14178# 0.0437f
C15699 vcm a_24962_2130# 0.1f
C15700 a_19030_6146# a_20034_6146# 0.843f
C15701 m2_12776_946# m2_13204_1374# 0.165f
C15702 row_n[2] a_18938_4138# 0.0437f
C15703 vcm a_12306_11206# 0.155f
C15704 col_n[16] a_19334_9198# 0.084f
C15705 col[22] a_2475_9182# 0.136f
C15706 VDD a_10394_1488# 0.0977f
C15707 m2_19228_17438# a_19030_17190# 0.165f
C15708 rowon_n[6] a_18026_8154# 0.248f
C15709 m2_34864_5966# VDD 0.784f
C15710 ctop a_25054_6146# 4.11f
C15711 a_2475_15206# a_15926_15182# 0.264f
C15712 a_2275_15206# a_13310_15222# 0.144f
C15713 a_8898_15182# a_8990_15182# 0.326f
C15714 VDD a_33998_11166# 0.181f
C15715 rowon_n[0] m2_24248_2378# 0.0322f
C15716 a_2475_18218# a_21038_18194# 0.0299f
C15717 col_n[27] a_30474_3496# 0.0283f
C15718 a_2275_3158# a_28066_3134# 0.399f
C15719 rowoff_n[8] a_30474_10524# 0.0133f
C15720 col_n[29] a_2275_15206# 0.113f
C15721 vcm a_5886_5142# 0.1f
C15722 m2_34864_12994# m2_35292_13422# 0.165f
C15723 a_9994_8154# a_9994_7150# 0.843f
C15724 vcm a_27366_15222# 0.155f
C15725 a_2275_12194# a_6890_12170# 0.136f
C15726 VDD a_25454_5504# 0.0779f
C15727 m2_8760_18014# VDD 0.993f
C15728 row_n[15] a_29070_17190# 0.282f
C15729 ctop a_5978_9158# 4.11f
C15730 a_2475_17214# a_30986_17190# 0.264f
C15731 a_2275_17214# a_28370_17230# 0.144f
C15732 VDD a_14922_14178# 0.181f
C15733 col[10] a_13006_7150# 0.367f
C15734 col[19] a_2275_12194# 0.0899f
C15735 rowon_n[0] a_5886_2130# 0.118f
C15736 col[24] a_2275_1150# 0.0899f
C15737 col[17] a_19942_9158# 0.0682f
C15738 a_22954_5142# a_23446_5504# 0.0658f
C15739 a_22042_5142# a_22346_5182# 0.0931f
C15740 col_n[25] a_28066_3134# 0.251f
C15741 m2_3740_18014# m2_4168_18442# 0.165f
C15742 vcm a_20946_9158# 0.1f
C15743 rowoff_n[14] a_15926_16186# 0.202f
C15744 a_33998_10162# a_34394_10202# 0.0313f
C15745 m2_10192_15430# a_9994_15182# 0.165f
C15746 vcm a_8290_18234# 0.16f
C15747 a_2275_14202# a_21950_14178# 0.136f
C15748 VDD a_6378_8516# 0.0779f
C15749 row_n[7] a_26362_9198# 0.0117f
C15750 m2_1732_13998# ctop 0.0428f
C15751 col_n[5] a_8290_7190# 0.084f
C15752 m2_2160_5390# rowon_n[3] 0.0219f
C15753 m2_6752_946# vcm 0.353f
C15754 ctop a_21038_13174# 4.11f
C15755 VDD a_29982_18194# 0.343f
C15756 a_2275_2154# a_33390_2170# 0.144f
C15757 a_18938_2130# a_19030_2130# 0.326f
C15758 m3_25960_18146# VDD 0.0313f
C15759 row_n[9] a_16930_11166# 0.0437f
C15760 col_n[9] a_2475_8178# 0.0531f
C15761 rowon_n[13] a_16018_15182# 0.248f
C15762 m2_29268_11414# a_29070_11166# 0.165f
C15763 vcm a_34394_13214# 0.155f
C15764 col_n[26] a_29470_13536# 0.0283f
C15765 a_2475_11190# a_14010_11166# 0.316f
C15766 a_25054_12170# a_25054_11166# 0.843f
C15767 VDD a_32082_3134# 0.483f
C15768 a_18938_16186# a_19334_16226# 0.0313f
C15769 VDD a_21438_12532# 0.0779f
C15770 rowon_n[3] a_26058_5142# 0.248f
C15771 m2_7756_18014# m3_8892_18146# 0.0341f
C15772 m2_17220_14426# rowon_n[12] 0.0322f
C15773 ctop a_2475_16210# 0.0488f
C15774 m2_23244_10410# rowon_n[8] 0.0322f
C15775 m2_29268_6394# rowon_n[4] 0.0322f
C15776 col[9] a_12002_17190# 0.367f
C15777 col[6] a_8898_7150# 0.0682f
C15778 a_2275_8178# a_4974_8154# 0.399f
C15779 a_2874_8154# a_3270_8194# 0.0313f
C15780 a_3878_8154# a_3970_8154# 0.326f
C15781 vcm a_16930_16186# 0.1f
C15782 a_2475_13198# a_29070_13174# 0.316f
C15783 a_15014_13174# a_16018_13174# 0.843f
C15784 VDD a_13006_6146# 0.483f
C15785 row_n[3] a_3970_5142# 0.282f
C15786 col_n[24] a_27062_13174# 0.251f
C15787 col_n[6] a_2275_11190# 0.113f
C15788 col_n[21] a_23958_3134# 0.0765f
C15789 VDD a_1957_15206# 0.196f
C15790 col_n[31] a_33998_15182# 0.0765f
C15791 col_n[4] a_7286_17230# 0.084f
C15792 vcm a_19030_1126# 0.557f
C15793 a_33998_6146# a_34090_6146# 0.326f
C15794 col[0] a_2966_15182# 0.367f
C15795 m2_20232_9406# a_20034_9158# 0.165f
C15796 m2_10768_946# m3_10900_1078# 3.79f
C15797 m3_15920_18146# m3_16924_18146# 0.202f
C15798 rowon_n[5] col[14] 0.0323f
C15799 row_n[11] col[25] 0.0342f
C15800 row_n[14] col[31] 0.0342f
C15801 row_n[12] col[27] 0.0342f
C15802 row_n[6] col[15] 0.0342f
C15803 row_n[15] rowoff_n[15] 0.209f
C15804 rowon_n[0] col[4] 0.0323f
C15805 rowon_n[8] col[20] 0.0323f
C15806 rowon_n[6] col[16] 0.0323f
C15807 row_n[1] col[5] 0.0342f
C15808 row_n[0] col[3] 0.0342f
C15809 row_n[5] col[13] 0.0342f
C15810 rowon_n[1] col[6] 0.0323f
C15811 row_n[2] col[7] 0.0342f
C15812 rowon_n[4] col[12] 0.0323f
C15813 row_n[8] col[19] 0.0342f
C15814 rowon_n[12] col[28] 0.0323f
C15815 row_n[10] col[23] 0.0342f
C15816 rowon_n[3] col[10] 0.0323f
C15817 row_n[3] col[9] 0.0342f
C15818 row_n[9] col[21] 0.0342f
C15819 row_n[13] col[29] 0.0342f
C15820 col_n[26] a_2475_10186# 0.0531f
C15821 ctop col[0] 0.0915f
C15822 rowon_n[7] col[18] 0.0323f
C15823 row_n[7] col[17] 0.0342f
C15824 row_n[4] col[11] 0.0342f
C15825 rowon_n[11] col[26] 0.0323f
C15826 rowon_n[13] col[30] 0.0323f
C15827 rowon_n[2] col[8] 0.0323f
C15828 rowon_n[9] col[22] 0.0323f
C15829 rowon_n[14] sample_n 0.0692f
C15830 rowon_n[10] col[24] 0.0323f
C15831 a_2275_10186# a_20034_10162# 0.399f
C15832 rowoff_n[15] a_3366_17552# 0.0133f
C15833 row_n[14] a_24354_16226# 0.0117f
C15834 rowoff_n[4] a_2475_6170# 3.9f
C15835 m2_10768_946# a_10998_2130# 0.843f
C15836 a_5978_15182# a_5978_14178# 0.843f
C15837 col_n[15] a_18426_11528# 0.0283f
C15838 VDD a_28066_10162# 0.483f
C15839 row_n[4] a_35398_6186# 0.0117f
C15840 a_28978_3134# a_29374_3174# 0.0313f
C15841 col[16] a_2475_7174# 0.136f
C15842 vcm a_34090_5142# 0.56f
C15843 a_2275_7174# a_10298_7190# 0.144f
C15844 rowoff_n[10] a_28066_12170# 0.294f
C15845 rowoff_n[2] a_10998_4138# 0.294f
C15846 a_2475_7174# a_12914_7150# 0.264f
C15847 col_n[0] a_2874_7150# 0.0765f
C15848 row_n[6] a_24962_8154# 0.0437f
C15849 a_18026_12170# a_18330_12210# 0.0931f
C15850 a_18938_12170# a_19430_12532# 0.0658f
C15851 a_2275_12194# a_35094_12170# 0.0924f
C15852 rowon_n[10] a_24050_12170# 0.248f
C15853 col[5] a_7894_17190# 0.0682f
C15854 a_30074_17190# a_31078_17190# 0.843f
C15855 VDD a_8990_13174# 0.483f
C15856 col_n[23] a_2275_13198# 0.113f
C15857 col_n[13] a_16018_11166# 0.251f
C15858 col_n[28] a_2275_2154# 0.113f
C15859 rowoff_n[0] a_20034_2130# 0.294f
C15860 col_n[10] a_12914_1126# 0.0765f
C15861 rowon_n[0] a_34090_2130# 0.248f
C15862 rowoff_n[7] a_2275_9182# 0.151f
C15863 a_2874_4138# a_2966_4138# 0.326f
C15864 col_n[20] a_22954_13174# 0.0765f
C15865 m3_2868_18146# ctop 0.209f
C15866 m2_11196_7398# a_10998_7150# 0.165f
C15867 vcm a_15014_8154# 0.56f
C15868 a_2475_9182# a_27974_9158# 0.264f
C15869 a_14922_9158# a_15014_9158# 0.326f
C15870 a_2275_9182# a_25358_9198# 0.144f
C15871 m2_1732_3958# row_n[2] 0.292f
C15872 row_n[10] a_2475_12194# 0.405f
C15873 col[13] a_2275_10186# 0.0899f
C15874 col[20] rowoff_n[12] 0.0901f
C15875 m3_18932_1078# a_19030_1126# 1.82f
C15876 a_3878_18194# a_4370_18556# 0.0658f
C15877 col_n[4] a_7382_9520# 0.0283f
C15878 row_n[0] a_12002_2130# 0.282f
C15879 VDD a_24050_17190# 0.484f
C15880 rowon_n[4] a_11910_6146# 0.118f
C15881 m2_30272_3382# a_30074_3134# 0.165f
C15882 vcm a_5278_2170# 0.155f
C15883 a_2275_6170# a_18938_6146# 0.136f
C15884 a_9902_6146# a_10298_6186# 0.0313f
C15885 m2_1732_11990# sample_n 0.0522f
C15886 vcm a_30074_12170# 0.56f
C15887 VDD a_26970_2130# 0.181f
C15888 m2_10192_17438# row_n[15] 0.0128f
C15889 m2_16216_13422# row_n[11] 0.0128f
C15890 m2_22240_9406# row_n[7] 0.0128f
C15891 m2_28264_5390# row_n[3] 0.0128f
C15892 a_33998_16186# a_34490_16548# 0.0658f
C15893 a_33086_16186# a_33390_16226# 0.0931f
C15894 row_n[11] a_32386_13214# 0.0117f
C15895 m3_34996_14130# a_34090_14178# 0.0303f
C15896 col_n[3] a_2475_6170# 0.0531f
C15897 a_5978_3134# a_6982_3134# 0.843f
C15898 a_2475_3158# a_10998_3134# 0.316f
C15899 a_2475_18218# a_2966_18194# 0.0299f
C15900 col_n[2] a_4974_9158# 0.251f
C15901 rowoff_n[8] a_12914_10162# 0.202f
C15902 col_n[28] a_31382_10202# 0.084f
C15903 a_24962_1126# a_2475_1150# 0.264f
C15904 a_22346_1166# a_2275_1150# 0.145f
C15905 m2_1732_4962# a_1957_5166# 0.245f
C15906 row_n[13] a_22954_15182# 0.0437f
C15907 vcm a_20338_6186# 0.155f
C15908 a_2275_8178# a_33998_8154# 0.136f
C15909 rowoff_n[11] a_16018_13174# 0.294f
C15910 col_n[9] a_11910_11166# 0.0765f
C15911 col[4] rowoff_n[13] 0.0901f
C15912 vcm a_10998_15182# 0.56f
C15913 a_29982_13174# a_30074_13174# 0.326f
C15914 VDD a_7894_5142# 0.181f
C15915 col[30] a_2275_12194# 0.0899f
C15916 row_n[3] a_32994_5142# 0.0437f
C15917 rowon_n[7] a_32082_9158# 0.248f
C15918 a_2275_17214# a_12002_17190# 0.399f
C15919 rowoff_n[6] a_21950_8154# 0.202f
C15920 a_2475_5166# a_26058_5142# 0.316f
C15921 a_31078_6146# a_31078_5142# 0.843f
C15922 m3_5880_1078# m3_6884_1078# 0.202f
C15923 vcm a_2275_9182# 6.49f
C15924 a_24962_10162# a_25358_10202# 0.0313f
C15925 rowoff_n[15] a_32082_17190# 0.294f
C15926 col[22] a_25054_8154# 0.367f
C15927 rowoff_n[4] a_30986_6146# 0.202f
C15928 ctop a_14010_4138# 4.11f
C15929 a_2475_14202# a_4882_14178# 0.264f
C15930 a_2874_14178# a_3366_14540# 0.0658f
C15931 a_2275_14202# a_3878_14178# 0.136f
C15932 col[29] a_31990_10162# 0.0682f
C15933 VDD a_22954_9158# 0.181f
C15934 row_n[7] a_9994_9158# 0.282f
C15935 rowon_n[11] a_9902_13174# 0.118f
C15936 ctop a_2966_13174# 4.06f
C15937 VDD a_10298_18234# 0.019f
C15938 a_9902_2130# a_10394_2492# 0.0658f
C15939 a_2275_2154# a_17022_2130# 0.399f
C15940 a_8990_2130# a_9294_2170# 0.0931f
C15941 col_n[20] a_2475_8178# 0.0531f
C15942 m2_10768_946# VDD 1f
C15943 vcm a_28978_4138# 0.1f
C15944 rowoff_n[9] a_22442_11528# 0.0133f
C15945 a_21038_7150# a_22042_7150# 0.843f
C15946 rowon_n[1] a_19942_3134# 0.118f
C15947 col_n[17] a_20338_8194# 0.084f
C15948 vcm a_16322_13214# 0.155f
C15949 VDD a_14410_3496# 0.0779f
C15950 m2_7756_18014# a_7894_18194# 0.225f
C15951 col[5] a_2475_16210# 0.136f
C15952 ctop a_29070_8154# 4.11f
C15953 a_2275_16210# a_17326_16226# 0.144f
C15954 a_10906_16186# a_10998_16186# 0.326f
C15955 a_2475_16210# a_19942_16186# 0.264f
C15956 VDD a_3366_12532# 0.0779f
C15957 col[10] a_2475_5166# 0.136f
C15958 col_n[28] a_31478_2492# 0.0283f
C15959 rowoff_n[7] a_31478_9520# 0.0133f
C15960 a_2275_4162# a_32082_4138# 0.399f
C15961 vcm a_9902_7150# 0.1f
C15962 a_12002_9158# a_12002_8154# 0.843f
C15963 rowoff_n[12] a_3970_14178# 0.294f
C15964 col_n[17] a_2275_11190# 0.113f
C15965 row_n[10] a_30986_12170# 0.0437f
C15966 vcm a_31382_17230# 0.155f
C15967 rowon_n[14] a_30074_16186# 0.248f
C15968 a_5886_13174# a_6282_13214# 0.0313f
C15969 a_2275_13198# a_10906_13174# 0.136f
C15970 VDD a_29470_7512# 0.0779f
C15971 col[11] a_14010_6146# 0.367f
C15972 ctop a_9994_11166# 4.11f
C15973 a_2275_18218# a_32386_18234# 0.145f
C15974 VDD a_18938_16186# 0.181f
C15975 col[18] a_20946_8154# 0.0682f
C15976 col[2] col[3] 0.0355f
C15977 row_n[7] col[28] 0.0342f
C15978 row_n[3] col[20] 0.0342f
C15979 rowon_n[4] col[23] 0.0323f
C15980 row_n[0] col[14] 0.0342f
C15981 row_n[1] col[16] 0.0342f
C15982 row_n[4] col[22] 0.0342f
C15983 rowon_n[8] col[31] 0.0323f
C15984 row_n[5] col[24] 0.0342f
C15985 rowon_n[5] col[25] 0.0323f
C15986 row_n[9] sample_n 0.0596f
C15987 row_n[6] col[26] 0.0342f
C15988 rowon_n[2] col[19] 0.0323f
C15989 rowon_n[6] col[27] 0.0323f
C15990 rowon_n[1] col[17] 0.0323f
C15991 row_n[8] col[30] 0.0342f
C15992 rowon_n[7] col[29] 0.0323f
C15993 ctop col[11] 0.123f
C15994 row_n[2] col[18] 0.0342f
C15995 rowon_n[3] col[21] 0.0323f
C15996 rowon_n[0] col[15] 0.0323f
C15997 col_n[26] a_29070_2130# 0.251f
C15998 a_24962_6146# a_25454_6508# 0.0658f
C15999 col[7] a_2275_8178# 0.0899f
C16000 a_24050_6146# a_24354_6186# 0.0931f
C16001 m2_34864_6970# vcm 0.408f
C16002 m2_24824_946# m2_25828_946# 0.843f
C16003 vcm a_24962_11166# 0.1f
C16004 a_1957_10186# a_2275_10186# 0.158f
C16005 a_2475_10186# a_2874_10162# 0.264f
C16006 VDD a_21038_1126# 0.0349f
C16007 row_n[14] a_7986_16186# 0.282f
C16008 col_n[6] a_9294_6186# 0.084f
C16009 a_2275_15206# a_25966_15182# 0.136f
C16010 col_n[16] a_19334_18234# 0.084f
C16011 VDD a_10394_10524# 0.0779f
C16012 col[27] a_2475_7174# 0.136f
C16013 ctop a_25054_15182# 4.11f
C16014 row_n[4] a_18026_6146# 0.282f
C16015 rowon_n[8] a_17934_10162# 0.118f
C16016 a_20946_3134# a_21038_3134# 0.326f
C16017 col_n[27] a_30474_12532# 0.0283f
C16018 rowoff_n[10] a_10394_12532# 0.0133f
C16019 a_28370_1166# vcm 0.16f
C16020 row_n[6] a_5278_8194# 0.0117f
C16021 m2_6176_12418# rowon_n[10] 0.0322f
C16022 m2_12200_8402# rowon_n[6] 0.0322f
C16023 vcm a_5886_14178# 0.1f
C16024 m2_18224_4386# rowon_n[2] 0.0322f
C16025 a_2475_12194# a_18026_12170# 0.316f
C16026 a_27062_13174# a_27062_12170# 0.843f
C16027 VDD a_2475_4162# 26.1f
C16028 m2_30272_18442# VDD 0.0456f
C16029 a_20946_17190# a_21342_17230# 0.0313f
C16030 VDD a_25454_14540# 0.0779f
C16031 col[0] a_2874_4138# 0.0682f
C16032 rowoff_n[0] a_1957_2154# 0.0219f
C16033 col[10] a_13006_16186# 0.367f
C16034 col[7] a_9902_6146# 0.0682f
C16035 col[17] a_19942_18194# 0.0682f
C16036 col[24] a_2275_10186# 0.0899f
C16037 col[31] rowoff_n[12] 0.0901f
C16038 VDD m2_1732_946# 1.56f
C16039 rowoff_n[14] a_26458_16548# 0.0133f
C16040 a_2275_9182# a_8990_9158# 0.399f
C16041 a_4974_9158# a_5278_9198# 0.0931f
C16042 a_5886_9158# a_6378_9520# 0.0658f
C16043 rowon_n[2] a_4974_4138# 0.248f
C16044 col_n[25] a_28066_12170# 0.251f
C16045 vcm a_20946_18194# 0.101f
C16046 a_2475_14202# a_33086_14178# 0.316f
C16047 a_17022_14178# a_18026_14178# 0.843f
C16048 m3_31984_1078# a_32082_2130# 0.0302f
C16049 m2_27260_17438# rowon_n[15] 0.0322f
C16050 col_n[22] a_24962_2130# 0.0765f
C16051 m2_33284_13422# rowon_n[11] 0.0322f
C16052 VDD a_17022_8154# 0.483f
C16053 m2_29844_946# vcm 0.353f
C16054 VDD a_6378_17552# 0.0779f
C16055 col_n[5] a_8290_16226# 0.084f
C16056 m3_1864_1078# VDD 0.0281f
C16057 vcm a_23046_3134# 0.56f
C16058 en_bit_n[1] a_17934_1126# 0.0724f
C16059 m2_3164_10410# a_2966_10162# 0.165f
C16060 rowoff_n[3] a_2874_5142# 0.202f
C16061 a_2275_11190# a_24050_11166# 0.399f
C16062 col_n[16] a_19430_10524# 0.0283f
C16063 col_n[9] a_2475_17214# 0.0531f
C16064 m2_26832_18014# a_26970_18194# 0.225f
C16065 m2_3740_18014# a_3970_17190# 0.843f
C16066 m2_1732_8978# VDD 0.856f
C16067 col_n[14] a_2475_6170# 0.0531f
C16068 row_n[11] a_16018_13174# 0.282f
C16069 a_7986_16186# a_7986_15182# 0.843f
C16070 VDD a_32082_12170# 0.483f
C16071 m2_22816_18014# m3_21944_18146# 0.0341f
C16072 rowon_n[15] a_15926_17190# 0.118f
C16073 a_30986_4138# a_31382_4178# 0.0313f
C16074 col[15] rowoff_n[13] 0.0901f
C16075 row_n[1] a_26058_3134# 0.282f
C16076 rowoff_n[1] a_12002_3134# 0.294f
C16077 row_n[13] a_3270_15222# 0.0117f
C16078 rowon_n[5] a_25966_7150# 0.118f
C16079 vcm a_3970_6146# 0.56f
C16080 a_2275_8178# a_14314_8194# 0.144f
C16081 rowoff_n[12] a_32994_14178# 0.202f
C16082 a_2475_8178# a_16930_8154# 0.264f
C16083 VDD rowoff_n[8] 1.51f
C16084 col[4] a_2475_3158# 0.136f
C16085 sample rowoff_n[9] 0.0775f
C16086 col[6] a_8898_16186# 0.0682f
C16087 a_20034_13174# a_20338_13214# 0.0931f
C16088 a_20946_13174# a_21438_13536# 0.0658f
C16089 row_n[3] a_13310_5182# 0.0117f
C16090 col_n[14] a_17022_10162# 0.251f
C16091 VDD a_13006_15182# 0.483f
C16092 rowoff_n[6] a_3878_8154# 0.202f
C16093 col_n[21] a_23958_12170# 0.0765f
C16094 col_n[11] a_2275_9182# 0.113f
C16095 a_2275_5166# a_7894_5142# 0.136f
C16096 m3_34996_17142# m3_34996_16138# 0.202f
C16097 m2_25828_946# m3_26964_1078# 0.0341f
C16098 rowon_n[9] a_2874_11166# 0.118f
C16099 vcm a_19030_10162# 0.56f
C16100 a_16930_10162# a_17022_10162# 0.326f
C16101 rowoff_n[15] a_14410_17552# 0.0133f
C16102 a_2275_10186# a_29374_10202# 0.144f
C16103 a_2475_10186# a_31990_10162# 0.264f
C16104 m2_16216_16434# a_16018_16186# 0.165f
C16105 m2_18800_18014# ctop 0.0422f
C16106 col_n[31] a_2475_8178# 0.0531f
C16107 col_n[5] a_8386_8516# 0.0283f
C16108 col[1] a_2275_6170# 0.0899f
C16109 m2_10768_946# col_n[8] 0.331f
C16110 a_32482_1488# col_n[29] 0.0283f
C16111 a_18026_3134# a_18026_2130# 0.843f
C16112 m2_5172_11414# row_n[9] 0.0128f
C16113 m2_11196_7398# row_n[5] 0.0128f
C16114 m2_17220_3382# row_n[1] 0.0128f
C16115 vcm a_9294_4178# 0.155f
C16116 rowoff_n[9] a_4882_11166# 0.202f
C16117 a_11910_7150# a_12306_7190# 0.0313f
C16118 a_2275_7174# a_22954_7150# 0.136f
C16119 m2_34864_11990# a_35094_12170# 0.0249f
C16120 col[16] a_2475_16210# 0.136f
C16121 vcm a_34090_14178# 0.56f
C16122 col[21] a_2475_5166# 0.136f
C16123 VDD a_30986_4138# 0.181f
C16124 col_n[0] a_2874_16186# 0.0765f
C16125 row_n[8] a_24050_10162# 0.282f
C16126 rowoff_n[7] a_13918_9158# 0.202f
C16127 col_n[3] a_5978_8154# 0.251f
C16128 col_n[29] a_32386_9198# 0.084f
C16129 rowon_n[12] a_23958_14178# 0.118f
C16130 a_2475_4162# a_15014_4138# 0.316f
C16131 a_7986_4138# a_8990_4138# 0.843f
C16132 col_n[28] a_2275_11190# 0.113f
C16133 m3_1864_12122# ctop 0.21f
C16134 col_n[10] a_12914_10162# 0.0765f
C16135 m2_3740_18014# col_n[1] 0.243f
C16136 m2_26256_16434# row_n[14] 0.0128f
C16137 vcm a_24354_8194# 0.155f
C16138 m2_32280_12418# row_n[10] 0.0128f
C16139 rowoff_n[13] a_20946_15182# 0.202f
C16140 row_n[10] a_11302_12210# 0.0117f
C16141 m2_7180_14426# a_6982_14178# 0.165f
C16142 rowon_n[2] a_33998_4138# 0.118f
C16143 vcm a_15014_17190# 0.56f
C16144 a_31990_14178# a_32082_14178# 0.326f
C16145 VDD a_11910_7150# 0.181f
C16146 rowoff_n[5] a_22954_7150# 0.202f
C16147 VDD col_n[0] 5.18f
C16148 rowon_n[2] col[30] 0.0323f
C16149 rowon_n[1] col[28] 0.0323f
C16150 ctop col[22] 0.123f
C16151 row_n[3] col[31] 0.0342f
C16152 rowon_n[0] col[26] 0.0323f
C16153 row_n[1] col[27] 0.0342f
C16154 row_n[0] col[25] 0.0342f
C16155 row_n[2] col[29] 0.0342f
C16156 rowon_n[3] sample_n 0.0692f
C16157 a_2275_18218# a_16018_18194# 0.0924f
C16158 row_n[0] a_21342_2170# 0.0117f
C16159 col[18] a_2275_8178# 0.0899f
C16160 a_2275_1150# a_5978_1126# 0.0924f
C16161 m2_4168_2378# a_3970_2130# 0.165f
C16162 col_n[4] a_7382_18556# 0.0283f
C16163 vcm a_17934_2130# 0.1f
C16164 col_n[1] a_3878_8154# 0.0765f
C16165 a_2475_6170# a_30074_6146# 0.316f
C16166 a_33086_7150# a_33086_6146# 0.843f
C16167 m2_5748_946# m2_6176_1374# 0.165f
C16168 col[23] a_26058_7150# 0.367f
C16169 m2_26256_10410# a_26058_10162# 0.165f
C16170 rowoff_n[3] a_31990_5142# 0.202f
C16171 row_n[2] a_11910_4138# 0.0437f
C16172 vcm a_5278_11206# 0.155f
C16173 a_26970_11166# a_27366_11206# 0.0313f
C16174 VDD a_2966_1126# 0.0351f
C16175 col[30] a_32994_9158# 0.0682f
C16176 rowon_n[6] a_10998_8154# 0.248f
C16177 m2_22816_18014# a_23046_17190# 0.843f
C16178 ctop a_18026_6146# 4.11f
C16179 a_2275_15206# a_6282_15222# 0.144f
C16180 a_2475_15206# a_8898_15182# 0.264f
C16181 VDD a_26970_11166# 0.181f
C16182 m2_1732_15002# m3_1864_16138# 0.0341f
C16183 a_2275_3158# a_21038_3134# 0.399f
C16184 a_11910_3134# a_12402_3496# 0.0658f
C16185 a_10998_3134# a_11302_3174# 0.0931f
C16186 a_2475_18218# a_14010_18194# 0.0299f
C16187 rowoff_n[8] a_23446_10524# 0.0133f
C16188 a_33390_1166# a_2275_1150# 0.145f
C16189 col_n[3] a_2475_15206# 0.0531f
C16190 col_n[18] a_21342_7190# 0.084f
C16191 vcm a_32994_6146# 0.1f
C16192 a_23046_8154# a_24050_8154# 0.843f
C16193 col_n[8] a_2475_4162# 0.0531f
C16194 vcm a_20338_15222# 0.155f
C16195 a_35002_13174# a_35398_13214# 0.0313f
C16196 VDD a_18426_5504# 0.0779f
C16197 a_30378_1166# VDD 0.0149f
C16198 a_25966_1126# col_n[23] 0.0765f
C16199 ctop a_33086_10162# 4.11f
C16200 row_n[15] a_22042_17190# 0.282f
C16201 a_2275_17214# a_21342_17230# 0.144f
C16202 a_2475_17214# a_23958_17190# 0.264f
C16203 a_12914_17190# a_13006_17190# 0.326f
C16204 rowoff_n[6] a_32482_8516# 0.0133f
C16205 VDD a_7894_14178# 0.181f
C16206 en_bit_n[0] a_2475_1150# 0.0162f
C16207 row_n[5] a_32082_7150# 0.282f
C16208 m2_17220_8402# a_17022_8154# 0.165f
C16209 rowon_n[9] a_31990_11166# 0.118f
C16210 a_32994_1126# a_33486_1488# 0.0658f
C16211 vcm a_13918_9158# 0.1f
C16212 a_14010_10162# a_14010_9158# 0.843f
C16213 rowoff_n[14] a_8898_16186# 0.202f
C16214 col[12] a_15014_5142# 0.367f
C16215 vcm a_2275_18218# 7.11f
C16216 a_2275_14202# a_14922_14178# 0.136f
C16217 a_7894_14178# a_8290_14218# 0.0313f
C16218 VDD a_33486_9520# 0.0779f
C16219 row_n[7] a_19334_9198# 0.0117f
C16220 col[22] a_25054_17190# 0.367f
C16221 col_n[5] a_2275_7174# 0.113f
C16222 col[19] a_21950_7150# 0.0682f
C16223 ctop a_14010_13174# 4.11f
C16224 VDD a_22954_18194# 0.343f
C16225 a_2475_2154# a_28978_2130# 0.264f
C16226 a_2275_2154# a_26362_2170# 0.144f
C16227 m2_33860_946# VDD 0.791f
C16228 row_n[9] a_9902_11166# 0.0437f
C16229 rowoff_n[9] a_33086_11166# 0.294f
C16230 a_26970_7150# a_27462_7512# 0.0658f
C16231 col_n[20] a_2475_17214# 0.0531f
C16232 a_26058_7150# a_26362_7190# 0.0931f
C16233 rowon_n[13] a_8990_15182# 0.248f
C16234 col_n[25] a_2475_6170# 0.0531f
C16235 vcm a_28978_13174# 0.1f
C16236 col_n[7] a_10298_5182# 0.084f
C16237 a_3970_11166# a_4974_11166# 0.843f
C16238 a_2475_11190# a_6982_11166# 0.316f
C16239 VDD a_25054_3134# 0.483f
C16240 col_n[17] a_20338_17230# 0.084f
C16241 a_2275_16210# a_29982_16186# 0.136f
C16242 VDD a_14410_12532# 0.0779f
C16243 rowon_n[3] a_19030_5142# 0.248f
C16244 a_33390_1166# m2_32856_946# 0.087f
C16245 col[26] rowoff_n[13] 0.0901f
C16246 ctop a_29070_17190# 4.06f
C16247 m2_1732_5966# rowon_n[4] 0.236f
C16248 col[10] a_2475_14202# 0.136f
C16249 m2_6176_2378# rowon_n[0] 0.0322f
C16250 a_22954_4138# a_23046_4138# 0.326f
C16251 col_n[2] rowoff_n[2] 0.0471f
C16252 col_n[1] rowoff_n[1] 0.0471f
C16253 col[15] a_2475_3158# 0.136f
C16254 col_n[6] rowoff_n[6] 0.0471f
C16255 col_n[8] rowoff_n[8] 0.0471f
C16256 col_n[28] a_31478_11528# 0.0283f
C16257 col_n[9] rowoff_n[9] 0.0471f
C16258 col_n[5] rowoff_n[5] 0.0471f
C16259 vcm rowoff_n[0] 0.533f
C16260 col_n[7] rowoff_n[7] 0.0471f
C16261 col_n[3] rowoff_n[3] 0.0471f
C16262 col_n[4] rowoff_n[4] 0.0471f
C16263 m2_8184_6394# a_7986_6146# 0.165f
C16264 vcm a_9902_16186# 0.1f
C16265 a_29070_14178# a_29070_13174# 0.843f
C16266 a_2475_13198# a_22042_13174# 0.316f
C16267 VDD a_5978_6146# 0.483f
C16268 col[1] a_3970_3134# 0.367f
C16269 m2_34864_18014# a_2475_18218# 0.282f
C16270 col_n[22] a_2275_9182# 0.113f
C16271 a_22954_18194# a_23350_18234# 0.0313f
C16272 VDD a_29470_16548# 0.0779f
C16273 col[11] a_14010_15182# 0.367f
C16274 a_17934_1126# a_18330_1166# 0.0346f
C16275 row_n[12] a_30074_14178# 0.282f
C16276 col[8] a_10906_5142# 0.0682f
C16277 vcm a_12002_1126# 0.165f
C16278 col[18] a_20946_17190# 0.0682f
C16279 m2_16216_15430# rowon_n[13] 0.0322f
C16280 m2_22240_11414# rowon_n[9] 0.0322f
C16281 m2_28264_7398# rowon_n[5] 0.0322f
C16282 m3_1864_18146# m3_2868_18146# 0.202f
C16283 m2_34288_3382# rowon_n[1] 0.0322f
C16284 col_n[26] a_29070_11166# 0.251f
C16285 col[7] a_2275_17214# 0.0899f
C16286 a_7894_10162# a_8386_10524# 0.0658f
C16287 a_6982_10162# a_7286_10202# 0.0931f
C16288 a_2275_10186# a_13006_10162# 0.399f
C16289 row_n[14] a_17326_16226# 0.0117f
C16290 m2_1732_16006# a_2475_16210# 0.139f
C16291 col[12] a_2275_6170# 0.0899f
C16292 a_19030_15182# a_20034_15182# 0.843f
C16293 VDD a_21038_10162# 0.483f
C16294 col[10] rowoff_n[14] 0.0901f
C16295 m2_1732_11990# m3_1864_13126# 0.0341f
C16296 col_n[6] a_9294_15222# 0.084f
C16297 row_n[4] a_27366_6186# 0.0117f
C16298 col[27] a_2475_16210# 0.136f
C16299 vcm a_27062_5142# 0.56f
C16300 a_2475_7174# a_5886_7150# 0.264f
C16301 rowoff_n[10] a_21038_12170# 0.294f
C16302 a_2275_7174# a_3270_7190# 0.144f
C16303 rowoff_n[2] a_3970_4138# 0.294f
C16304 col_n[17] a_20434_9520# 0.0283f
C16305 row_n[6] a_17934_8154# 0.0437f
C16306 a_2275_12194# a_28066_12170# 0.399f
C16307 rowon_n[10] a_17022_12170# 0.248f
C16308 row_n[0] m2_22240_2378# 0.0128f
C16309 a_9994_17190# a_9994_16186# 0.843f
C16310 VDD a_2475_13198# 26.1f
C16311 col_n[2] a_2475_2154# 0.0531f
C16312 m2_1732_16006# col[0] 0.0137f
C16313 rowon_n[0] a_27062_2130# 0.248f
C16314 rowoff_n[0] a_13006_2130# 0.294f
C16315 col[0] a_2874_13174# 0.0682f
C16316 a_32994_5142# a_33390_5182# 0.0313f
C16317 vcm a_7986_8154# 0.56f
C16318 a_2475_9182# a_20946_9158# 0.264f
C16319 a_2275_9182# a_18330_9198# 0.144f
C16320 col[7] a_9902_15182# 0.0682f
C16321 rowoff_n[13] a_2275_15206# 0.151f
C16322 VDD col_n[10] 5.17f
C16323 vcm col_n[7] 1.94f
C16324 col_n[3] col_n[4] 0.0101f
C16325 col[13] col[14] 0.0355f
C16326 ctop rowoff_n[15] 0.177f
C16327 a_22042_14178# a_22346_14218# 0.0931f
C16328 col_n[15] a_18026_9158# 0.251f
C16329 a_22954_14178# a_23446_14540# 0.0658f
C16330 col[29] a_2275_8178# 0.0899f
C16331 col_n[22] a_24962_11166# 0.0765f
C16332 row_n[0] a_4974_2130# 0.282f
C16333 VDD a_17022_17190# 0.484f
C16334 a_29070_2130# a_30074_2130# 0.843f
C16335 rowon_n[4] a_4882_6146# 0.118f
C16336 vcm a_32386_3174# 0.155f
C16337 a_2275_6170# a_11910_6146# 0.136f
C16338 m2_1732_9982# vcm 0.316f
C16339 col_n[0] a_2275_5166# 0.113f
C16340 vcm a_23046_12170# 0.56f
C16341 a_18938_11166# a_19030_11166# 0.326f
C16342 a_2275_11190# a_33390_11206# 0.144f
C16343 VDD a_19942_2130# 0.181f
C16344 col_n[6] a_9390_7512# 0.0283f
C16345 row_n[11] a_25358_13214# 0.0117f
C16346 col_n[14] a_2475_15206# 0.0531f
C16347 col_n[19] a_2475_4162# 0.0531f
C16348 a_2475_3158# a_3970_3134# 0.316f
C16349 a_2275_3158# a_2966_3134# 0.399f
C16350 a_20034_4138# a_20034_3134# 0.843f
C16351 rowoff_n[8] a_5886_10162# 0.202f
C16352 row_n[13] a_15926_15182# 0.0437f
C16353 vcm a_13310_6186# 0.155f
C16354 a_13918_8154# a_14314_8194# 0.0313f
C16355 rowoff_n[11] a_8990_13174# 0.294f
C16356 a_2275_8178# a_26970_8154# 0.136f
C16357 vcm a_3970_15182# 0.56f
C16358 VDD a_35002_6146# 0.258f
C16359 col[4] a_2475_12194# 0.136f
C16360 row_n[3] a_25966_5142# 0.0437f
C16361 col[9] a_2475_1150# 0.136f
C16362 a_3878_17190# a_3970_17190# 0.326f
C16363 rowon_n[7] a_25054_9158# 0.248f
C16364 a_2874_17190# a_3270_17230# 0.0313f
C16365 m2_15212_14426# row_n[12] 0.0128f
C16366 a_2275_17214# a_4974_17190# 0.399f
C16367 rowoff_n[6] a_14922_8154# 0.202f
C16368 col_n[30] a_33390_8194# 0.084f
C16369 col_n[4] a_6982_7150# 0.251f
C16370 m2_21236_10410# row_n[8] 0.0128f
C16371 m2_27260_6394# row_n[4] 0.0128f
C16372 m3_14916_18146# a_15014_17190# 0.0303f
C16373 col_n[11] a_13918_9158# 0.0765f
C16374 a_9994_5142# a_10998_5142# 0.843f
C16375 a_2475_5166# a_19030_5142# 0.316f
C16376 m2_1732_7974# a_2966_8154# 0.843f
C16377 col_n[11] a_2275_18218# 0.113f
C16378 vcm a_28370_10202# 0.155f
C16379 en_C0_n a_3970_1126# 0.208f
C16380 rowoff_n[15] a_25054_17190# 0.294f
C16381 col_n[16] a_2275_7174# 0.113f
C16382 rowoff_n[4] a_23958_6146# 0.202f
C16383 ctop a_6982_4138# 4.11f
C16384 a_33998_15182# a_34090_15182# 0.326f
C16385 row_n[7] a_2874_9158# 0.0436f
C16386 VDD a_15926_9158# 0.181f
C16387 m2_1732_8978# m3_1864_10114# 0.0341f
C16388 rowon_n[11] a_2161_13198# 0.0177f
C16389 VDD a_3270_18234# 0.019f
C16390 col_n[31] a_2475_17214# 0.0531f
C16391 col_n[5] a_8386_17552# 0.0283f
C16392 a_2275_2154# a_9994_2130# 0.399f
C16393 col[1] a_2275_15206# 0.0899f
C16394 col[24] a_27062_6146# 0.367f
C16395 col[6] a_2275_4162# 0.0899f
C16396 vcm a_21950_4138# 0.1f
C16397 rowoff_n[2] a_32994_4138# 0.202f
C16398 rowoff_n[9] a_15414_11528# 0.0133f
C16399 a_2475_7174# a_34090_7150# 0.316f
C16400 rowon_n[1] a_12914_3134# 0.118f
C16401 m2_34864_10986# a_2275_11190# 0.278f
C16402 col[31] a_33998_8154# 0.0682f
C16403 vcm a_9294_13214# 0.155f
C16404 a_28978_12170# a_29374_12210# 0.0313f
C16405 VDD a_7382_3496# 0.0779f
C16406 m2_2736_18014# a_2874_18194# 0.225f
C16407 ctop a_22042_8154# 4.11f
C16408 col[21] a_2475_14202# 0.136f
C16409 a_2275_16210# a_10298_16226# 0.144f
C16410 a_2475_16210# a_12914_16186# 0.264f
C16411 VDD a_30986_13174# 0.181f
C16412 col_n[16] rowoff_n[5] 0.0471f
C16413 col_n[12] rowoff_n[1] 0.0471f
C16414 col_n[17] rowoff_n[6] 0.0471f
C16415 col_n[11] rowoff_n[0] 0.0471f
C16416 col_n[20] rowoff_n[9] 0.0471f
C16417 col_n[15] rowoff_n[4] 0.0471f
C16418 col_n[14] rowoff_n[3] 0.0471f
C16419 col_n[19] rowoff_n[8] 0.0471f
C16420 col_n[18] rowoff_n[7] 0.0471f
C16421 col[26] a_2475_3158# 0.136f
C16422 col_n[13] rowoff_n[2] 0.0471f
C16423 row_n[8] a_33390_10202# 0.0117f
C16424 rowoff_n[7] a_24450_9520# 0.0133f
C16425 col_n[19] a_22346_6186# 0.084f
C16426 a_13006_4138# a_13310_4178# 0.0931f
C16427 a_2275_4162# a_25054_4138# 0.399f
C16428 a_13918_4138# a_14410_4500# 0.0658f
C16429 m3_21944_1078# ctop 0.21f
C16430 VDD a_2475_18218# 26.8f
C16431 col_n[3] a_5978_17190# 0.251f
C16432 col_n[29] a_32386_18234# 0.084f
C16433 vcm a_2161_7174# 0.0169f
C16434 m2_1732_16006# m2_2160_16434# 0.165f
C16435 rowoff_n[13] a_31478_15544# 0.0133f
C16436 a_25054_9158# a_26058_9158# 0.843f
C16437 row_n[10] a_23958_12170# 0.0437f
C16438 vcm a_24354_17230# 0.155f
C16439 rowon_n[14] a_23046_16186# 0.248f
C16440 a_2874_13174# a_2966_13174# 0.326f
C16441 VDD a_22442_7512# 0.0779f
C16442 rowoff_n[5] a_33486_7512# 0.0133f
C16443 m2_20808_946# col_n[18] 0.331f
C16444 a_14922_18194# a_15014_18194# 0.0991f
C16445 a_2275_18218# a_25358_18234# 0.145f
C16446 VDD a_11910_16186# 0.181f
C16447 row_n[0] a_33998_2130# 0.0437f
C16448 a_9902_1126# a_9994_1126# 0.0991f
C16449 a_2275_1150# a_15318_1166# 0.145f
C16450 a_2475_1150# a_17934_1126# 0.285f
C16451 rowon_n[4] a_33086_6146# 0.248f
C16452 m2_18800_18014# col[16] 0.347f
C16453 col[18] a_2275_17214# 0.0899f
C16454 m2_34864_9982# a_35002_10162# 0.225f
C16455 col[23] a_2275_6170# 0.0899f
C16456 vcm a_17934_11166# 0.1f
C16457 col[13] a_16018_4138# 0.367f
C16458 col[21] rowoff_n[14] 0.0901f
C16459 col_n[1] a_3878_17190# 0.0765f
C16460 a_16018_11166# a_16018_10162# 0.843f
C16461 VDD a_14010_1126# 0.035f
C16462 m2_22240_17438# a_22042_17190# 0.165f
C16463 col[23] a_26058_16186# 0.367f
C16464 col[20] a_22954_6146# 0.0682f
C16465 a_9902_15182# a_10298_15222# 0.0313f
C16466 a_2275_15206# a_18938_15182# 0.136f
C16467 VDD a_2966_10162# 0.485f
C16468 col_n[4] rowoff_n[10] 0.0471f
C16469 col[30] a_32994_18194# 0.0682f
C16470 ctop a_18026_15182# 4.11f
C16471 row_n[4] a_10998_6146# 0.282f
C16472 rowon_n[8] a_10906_10162# 0.118f
C16473 a_2475_3158# a_32994_3134# 0.264f
C16474 a_2275_3158# a_30378_3174# 0.144f
C16475 rowoff_n[8] a_34090_10162# 0.294f
C16476 col_n[8] a_11302_4178# 0.084f
C16477 rowoff_n[10] a_2966_12170# 0.294f
C16478 a_28066_8154# a_28370_8194# 0.0931f
C16479 a_28978_8154# a_29470_8516# 0.0658f
C16480 col_n[18] a_21342_16226# 0.084f
C16481 vcm a_32994_15182# 0.1f
C16482 a_5978_12170# a_6982_12170# 0.843f
C16483 a_2475_12194# a_10998_12170# 0.316f
C16484 col_n[8] a_2475_13198# 0.0531f
C16485 VDD a_29070_5142# 0.483f
C16486 m2_16216_18442# VDD 0.0456f
C16487 col_n[13] a_2475_2154# 0.0531f
C16488 row_n[15] a_31382_17230# 0.0117f
C16489 a_2275_17214# a_33998_17190# 0.136f
C16490 VDD a_18426_14540# 0.0779f
C16491 col_n[29] a_32482_10524# 0.0283f
C16492 a_24962_5142# a_25054_5142# 0.326f
C16493 VDD col_n[21] 5.17f
C16494 vcm col_n[18] 1.94f
C16495 col[5] rowoff_n[15] 0.0901f
C16496 a_1957_9182# a_2161_9182# 0.115f
C16497 a_2475_9182# a_2275_9182# 2.76f
C16498 rowoff_n[14] a_19430_16548# 0.0133f
C16499 m2_13204_15430# a_13006_15182# 0.165f
C16500 vcm a_13918_18194# 0.101f
C16501 m2_20808_946# a_21342_1166# 0.087f
C16502 col[2] a_4974_2130# 0.367f
C16503 a_2475_14202# a_26058_14178# 0.316f
C16504 a_31078_15182# a_31078_14178# 0.843f
C16505 row_n[7] a_31990_9158# 0.0437f
C16506 VDD a_9994_8154# 0.483f
C16507 m2_5172_13422# rowon_n[11] 0.0322f
C16508 m2_11196_9406# rowon_n[7] 0.0322f
C16509 m2_1732_5966# m3_1864_7102# 0.0341f
C16510 col[12] a_15014_14178# 0.367f
C16511 m2_17220_5390# rowon_n[3] 0.0322f
C16512 rowon_n[11] a_31078_13174# 0.248f
C16513 col[9] a_11910_4138# 0.0682f
C16514 VDD a_33486_18556# 0.0858f
C16515 col_n[5] a_2275_16210# 0.113f
C16516 a_19942_2130# a_20338_2170# 0.0313f
C16517 col[19] a_21950_16186# 0.0682f
C16518 col_n[10] a_2275_5166# 0.113f
C16519 vcm a_16018_3134# 0.56f
C16520 col_n[27] a_30074_10162# 0.251f
C16521 m2_32280_11414# a_32082_11166# 0.165f
C16522 a_8990_11166# a_9294_11206# 0.0931f
C16523 a_9902_11166# a_10394_11528# 0.0658f
C16524 a_2275_11190# a_17022_11166# 0.399f
C16525 VDD a_35398_3174# 0.0882f
C16526 m2_21812_18014# a_22042_18194# 0.0249f
C16527 col_n[25] a_2475_15206# 0.0531f
C16528 col_n[7] a_10298_14218# 0.084f
C16529 row_n[11] a_8990_13174# 0.282f
C16530 a_21038_16186# a_22042_16186# 0.843f
C16531 col_n[30] a_2475_4162# 0.0531f
C16532 VDD a_25054_12170# 0.483f
C16533 m2_12776_18014# m3_13912_18146# 0.0341f
C16534 m2_1732_18014# m3_1864_17142# 0.0341f
C16535 col[0] a_2275_2154# 0.099f
C16536 rowon_n[15] a_8898_17190# 0.118f
C16537 m2_32280_14426# rowon_n[12] 0.0322f
C16538 row_n[1] a_19030_3134# 0.282f
C16539 rowoff_n[1] a_4974_3134# 0.294f
C16540 col_n[18] a_21438_8516# 0.0283f
C16541 rowon_n[5] a_18938_7150# 0.118f
C16542 vcm a_31078_7150# 0.56f
C16543 rowoff_n[12] a_25966_14178# 0.202f
C16544 a_2275_8178# a_7286_8194# 0.144f
C16545 a_5886_8154# a_5978_8154# 0.326f
C16546 a_2475_8178# a_9902_8154# 0.264f
C16547 col[15] a_2475_12194# 0.136f
C16548 m2_4168_13422# a_3970_13174# 0.165f
C16549 col[20] a_2475_1150# 0.136f
C16550 a_2275_13198# a_32082_13174# 0.399f
C16551 row_n[3] a_6282_5182# 0.0117f
C16552 VDD a_5978_15182# 0.483f
C16553 col[1] a_3970_12170# 0.367f
C16554 col_n[22] a_2275_18218# 0.113f
C16555 vcm a_21342_1166# 0.16f
C16556 col_n[27] a_2275_7174# 0.113f
C16557 col[8] a_10906_14178# 0.0682f
C16558 m2_23244_9406# a_23046_9158# 0.165f
C16559 m2_15788_946# m3_15920_1078# 3.79f
C16560 vcm a_12002_10162# 0.56f
C16561 a_2275_10186# a_22346_10202# 0.144f
C16562 rowoff_n[15] a_7382_17552# 0.0133f
C16563 a_2475_10186# a_24962_10162# 0.264f
C16564 col_n[16] a_19030_8154# 0.251f
C16565 row_n[14] a_29982_16186# 0.0437f
C16566 a_24962_15182# a_25454_15544# 0.0658f
C16567 a_24050_15182# a_24354_15222# 0.0931f
C16568 m2_4744_18014# ctop 0.0422f
C16569 col_n[23] a_25966_10162# 0.0765f
C16570 col[12] a_2275_15206# 0.0899f
C16571 col[17] a_2275_4162# 0.0899f
C16572 a_31078_3134# a_32082_3134# 0.843f
C16573 vcm a_3878_4138# 0.1f
C16574 a_2275_7174# a_15926_7150# 0.136f
C16575 m2_33860_18014# vcm 0.353f
C16576 vcm a_27062_14178# 0.56f
C16577 col_n[7] a_10394_6508# 0.0283f
C16578 a_20946_12170# a_21038_12170# 0.326f
C16579 VDD a_23958_4138# 0.181f
C16580 col_n[29] rowoff_n[7] 0.0471f
C16581 col_n[25] rowoff_n[3] 0.0471f
C16582 col_n[23] rowoff_n[1] 0.0471f
C16583 col_n[31] rowoff_n[9] 0.0471f
C16584 col_n[22] rowoff_n[0] 0.0471f
C16585 col_n[24] rowoff_n[2] 0.0471f
C16586 col_n[26] rowoff_n[4] 0.0471f
C16587 col_n[27] rowoff_n[5] 0.0471f
C16588 col_n[30] rowoff_n[8] 0.0471f
C16589 col_n[28] rowoff_n[6] 0.0471f
C16590 col_n[17] a_20434_18556# 0.0283f
C16591 col_n[8] a_2475_18218# 0.0529f
C16592 row_n[8] a_17022_10162# 0.282f
C16593 rowoff_n[7] a_6890_9158# 0.202f
C16594 rowon_n[12] a_16930_14178# 0.118f
C16595 a_22042_5142# a_22042_4138# 0.843f
C16596 a_2475_4162# a_7986_4138# 0.316f
C16597 m3_17928_18146# ctop 0.209f
C16598 col_n[2] a_2475_11190# 0.0531f
C16599 m2_14208_7398# a_14010_7150# 0.165f
C16600 m2_4168_12418# row_n[10] 0.0128f
C16601 vcm a_17326_8194# 0.155f
C16602 m2_10192_8402# row_n[6] 0.0128f
C16603 a_2275_9182# a_30986_9158# 0.136f
C16604 rowoff_n[13] a_13918_15182# 0.202f
C16605 a_15926_9158# a_16322_9198# 0.0313f
C16606 m2_16216_4386# row_n[2] 0.0128f
C16607 row_n[10] a_4274_12210# 0.0117f
C16608 rowon_n[2] a_26970_4138# 0.118f
C16609 ctop a_30074_3134# 4.11f
C16610 vcm a_7986_17190# 0.56f
C16611 VDD a_4882_7150# 0.181f
C16612 m2_1732_2954# m3_1864_4090# 0.0341f
C16613 col_n[5] a_7986_6146# 0.251f
C16614 rowoff_n[5] a_15926_7150# 0.202f
C16615 a_2275_18218# a_8990_18194# 0.0924f
C16616 a_5886_18194# a_6378_18556# 0.0658f
C16617 row_n[0] a_14314_2170# 0.0117f
C16618 col[29] a_2275_17214# 0.0899f
C16619 col_n[12] a_14922_8154# 0.0765f
C16620 a_35002_2130# a_35494_2492# 0.0658f
C16621 m2_33284_3382# a_33086_3134# 0.165f
C16622 vcm a_10906_2130# 0.1f
C16623 sample_n rowoff_n[14] 0.14f
C16624 a_12002_6146# a_13006_6146# 0.843f
C16625 a_2475_6170# a_23046_6146# 0.316f
C16626 rowoff_n[3] a_24962_5142# 0.202f
C16627 row_n[2] a_4882_4138# 0.0437f
C16628 vcm a_32386_12210# 0.155f
C16629 col_n[15] rowoff_n[10] 0.0471f
C16630 VDD a_30474_2492# 0.0779f
C16631 m2_25252_17438# row_n[15] 0.0128f
C16632 rowon_n[6] a_3970_8154# 0.248f
C16633 m2_31276_13422# row_n[11] 0.0128f
C16634 col_n[0] a_2275_14202# 0.113f
C16635 ctop a_10998_6146# 4.11f
C16636 VDD a_19942_11166# 0.181f
C16637 col_n[4] a_2275_3158# 0.113f
C16638 col_n[6] a_9390_16548# 0.0283f
C16639 col[25] a_28066_5142# 0.367f
C16640 a_2275_3158# a_14010_3134# 0.399f
C16641 a_2475_18218# a_6982_18194# 0.0299f
C16642 rowoff_n[1] a_33998_3134# 0.202f
C16643 rowoff_n[8] a_16418_10524# 0.0133f
C16644 a_27974_1126# a_2275_1150# 0.136f
C16645 m2_5172_5390# a_4974_5142# 0.165f
C16646 col_n[19] a_2475_13198# 0.0531f
C16647 vcm a_25966_6146# 0.1f
C16648 col_n[24] a_2475_2154# 0.0531f
C16649 vcm a_13310_15222# 0.155f
C16650 a_30986_13174# a_31382_13214# 0.0313f
C16651 VDD a_11398_5504# 0.0779f
C16652 a_23350_1166# VDD 0.0149f
C16653 row_n[15] a_15014_17190# 0.282f
C16654 ctop a_26058_10162# 4.11f
C16655 a_2475_17214# a_16930_17190# 0.264f
C16656 a_2275_17214# a_14314_17230# 0.144f
C16657 VDD a_35002_15182# 0.258f
C16658 rowoff_n[6] a_25454_8516# 0.0133f
C16659 col_n[20] a_23350_5182# 0.084f
C16660 VDD rowon_n[15] 3.1f
C16661 vcm col_n[29] 1.94f
C16662 col[24] col[25] 0.0355f
C16663 col[16] rowoff_n[15] 0.0901f
C16664 col[9] a_2475_10186# 0.136f
C16665 col_n[4] a_6982_16186# 0.251f
C16666 col_n[30] a_33390_17230# 0.084f
C16667 a_2275_5166# a_29070_5142# 0.399f
C16668 a_15014_5142# a_15318_5182# 0.0931f
C16669 a_15926_5142# a_16418_5504# 0.0658f
C16670 row_n[5] a_25054_7150# 0.282f
C16671 col_n[11] a_13918_18194# 0.0762f
C16672 col_n[0] rowoff_n[11] 0.0471f
C16673 rowon_n[9] a_24962_11166# 0.118f
C16674 vcm a_6890_9158# 0.1f
C16675 a_27062_10162# a_28066_10162# 0.843f
C16676 rowoff_n[4] a_34490_6508# 0.0133f
C16677 m2_26832_946# a_2475_1150# 0.286f
C16678 a_2275_14202# a_7894_14178# 0.136f
C16679 m2_32856_946# a_33086_2130# 0.843f
C16680 VDD a_26458_9520# 0.0779f
C16681 row_n[7] a_12306_9198# 0.0117f
C16682 col_n[16] a_2275_16210# 0.113f
C16683 col_n[21] a_2275_5166# 0.113f
C16684 ctop a_6982_13174# 4.11f
C16685 VDD a_15926_18194# 0.343f
C16686 a_11910_2130# a_12002_2130# 0.326f
C16687 a_2475_2154# a_21950_2130# 0.264f
C16688 a_2275_2154# a_19334_2170# 0.144f
C16689 m2_19228_1374# VDD 0.0209f
C16690 row_n[9] a_2161_11190# 0.0221f
C16691 rowoff_n[9] a_26058_11166# 0.294f
C16692 col[14] a_17022_3134# 0.367f
C16693 rowon_n[13] a_2475_15206# 0.31f
C16694 col[24] a_27062_15182# 0.367f
C16695 col[6] a_2275_13198# 0.0899f
C16696 vcm a_21950_13174# 0.1f
C16697 col[21] a_23958_5142# 0.0682f
C16698 a_18026_12170# a_18026_11166# 0.843f
C16699 VDD a_18026_3134# 0.483f
C16700 col[11] a_2275_2154# 0.0899f
C16701 m2_8760_18014# a_9294_18234# 0.087f
C16702 m2_24824_18014# a_2275_18218# 0.28f
C16703 col[31] a_33998_17190# 0.0682f
C16704 a_11910_16186# a_12306_16226# 0.0313f
C16705 a_2275_16210# a_22954_16186# 0.136f
C16706 rowon_n[3] a_12002_5142# 0.248f
C16707 VDD a_7382_12532# 0.0779f
C16708 ctop a_22042_17190# 4.06f
C16709 rowoff_n[7] a_35094_9158# 0.0135f
C16710 col[26] a_2475_12194# 0.136f
C16711 a_2275_4162# a_35398_4178# 0.145f
C16712 col_n[9] a_12306_3174# 0.084f
C16713 m2_1732_5966# a_2275_6170# 0.191f
C16714 col[31] a_2475_1150# 0.0298f
C16715 col_n[19] a_22346_15222# 0.084f
C16716 a_30074_9158# a_30378_9198# 0.0931f
C16717 a_30986_9158# a_31478_9520# 0.0658f
C16718 vcm a_2161_16210# 0.0169f
C16719 a_2475_13198# a_15014_13174# 0.316f
C16720 a_7986_13174# a_8990_13174# 0.843f
C16721 VDD a_33086_7150# 0.483f
C16722 m2_20808_18014# a_2475_18218# 0.286f
C16723 col_n[30] a_33486_9520# 0.0283f
C16724 VDD a_22442_16548# 0.0779f
C16725 row_n[12] a_23046_14178# 0.282f
C16726 vcm a_4974_1126# 0.165f
C16727 a_26970_6146# a_27062_6146# 0.326f
C16728 m2_6176_3382# rowon_n[1] 0.0322f
C16729 m2_28840_946# m2_29268_1374# 0.165f
C16730 row_n[2] a_33086_4138# 0.282f
C16731 a_2275_10186# a_5978_10162# 0.399f
C16732 row_n[14] a_10298_16226# 0.0117f
C16733 rowon_n[6] a_32994_8154# 0.118f
C16734 col[23] a_2275_15206# 0.0899f
C16735 col[13] a_16018_13174# 0.367f
C16736 col[28] a_2275_4162# 0.0899f
C16737 a_2475_15206# a_30074_15182# 0.316f
C16738 a_33086_16186# a_33086_15182# 0.843f
C16739 col[10] a_12914_3134# 0.0682f
C16740 VDD a_14010_10162# 0.483f
C16741 col[20] a_22954_15182# 0.0682f
C16742 row_n[4] a_20338_6186# 0.0117f
C16743 a_21950_3134# a_22346_3174# 0.0313f
C16744 col_n[28] a_31078_9158# 0.251f
C16745 vcm a_20034_5142# 0.56f
C16746 rowoff_n[10] a_14010_12170# 0.294f
C16747 a_35002_1126# vcm 0.0989f
C16748 m2_15212_16434# rowon_n[14] 0.0322f
C16749 row_n[6] a_10906_8154# 0.0437f
C16750 m2_21236_12418# rowon_n[10] 0.0322f
C16751 m2_27260_8402# rowon_n[6] 0.0322f
C16752 a_2275_12194# a_21038_12170# 0.399f
C16753 a_11910_12170# a_12402_12532# 0.0658f
C16754 col_n[8] a_11302_13214# 0.084f
C16755 a_10998_12170# a_11302_12210# 0.0931f
C16756 m2_33284_4386# rowon_n[2] 0.0322f
C16757 rowon_n[10] a_9994_12170# 0.248f
C16758 col_n[19] a_2475_18218# 0.0529f
C16759 col[1] a_3878_1126# 0.0703f
C16760 a_23046_17190# a_24050_17190# 0.843f
C16761 VDD a_29070_14178# 0.483f
C16762 col_n[13] a_2475_11190# 0.0531f
C16763 rowoff_n[0] a_5978_2130# 0.294f
C16764 rowon_n[0] a_20034_2130# 0.248f
C16765 col_n[19] a_22442_7512# 0.0283f
C16766 m2_6752_946# ctop 0.0428f
C16767 m2_34864_7974# a_34090_8154# 0.843f
C16768 vcm a_35094_9158# 0.165f
C16769 rowoff_n[14] a_30074_16186# 0.294f
C16770 a_2275_9182# a_11302_9198# 0.144f
C16771 a_7894_9158# a_7986_9158# 0.326f
C16772 a_2475_9182# a_13918_9158# 0.264f
C16773 col[3] a_2475_8178# 0.136f
C16774 col[2] a_4974_11166# 0.367f
C16775 m3_1864_10114# a_2966_10162# 0.0302f
C16776 VDD a_9994_17190# 0.484f
C16777 col[9] a_11910_13174# 0.0682f
C16778 m3_16924_1078# VDD 0.0157f
C16779 row_n[9] a_31078_11166# 0.282f
C16780 vcm a_25358_3174# 0.155f
C16781 col_n[26] rowoff_n[10] 0.0471f
C16782 a_2966_6146# a_3970_6146# 0.843f
C16783 a_2275_6170# a_4882_6146# 0.136f
C16784 col_n[17] a_20034_7150# 0.251f
C16785 rowon_n[13] a_30986_15182# 0.118f
C16786 col_n[10] a_2275_14202# 0.113f
C16787 vcm a_16018_12170# 0.56f
C16788 col_n[15] a_2275_3158# 0.113f
C16789 a_2275_11190# a_26362_11206# 0.144f
C16790 a_2475_11190# a_28978_11166# 0.264f
C16791 VDD a_12914_2130# 0.181f
C16792 col_n[24] a_26970_9158# 0.0765f
C16793 m2_27836_18014# a_28370_18234# 0.087f
C16794 a_26058_16186# a_26362_16226# 0.0931f
C16795 a_26970_16186# a_27462_16548# 0.0658f
C16796 row_n[11] a_18330_13214# 0.0117f
C16797 VDD a_35398_12210# 0.0882f
C16798 m2_27836_18014# m3_26964_18146# 0.0341f
C16799 col_n[30] a_2475_13198# 0.0531f
C16800 a_33086_4138# a_34090_4138# 0.843f
C16801 col[0] a_2275_11190# 0.099f
C16802 row_n[1] a_28370_3174# 0.0117f
C16803 row_n[13] a_8898_15182# 0.0437f
C16804 vcm a_6282_6186# 0.155f
C16805 rowoff_n[11] a_2475_13198# 3.9f
C16806 a_2275_8178# a_19942_8154# 0.136f
C16807 col_n[8] a_11398_5504# 0.0283f
C16808 col_n[18] a_21438_17552# 0.0283f
C16809 ctop a_19030_1126# 2.06f
C16810 vcm a_31078_16186# 0.56f
C16811 a_22954_13174# a_23046_13174# 0.326f
C16812 VDD a_27974_6146# 0.181f
C16813 row_n[3] a_18938_5142# 0.0437f
C16814 col_n[8] rowon_n[15] 0.111f
C16815 col_n[3] row_n[13] 0.298f
C16816 col_n[5] row_n[14] 0.298f
C16817 col_n[2] rowon_n[12] 0.111f
C16818 vcm rowon_n[11] 0.65f
C16819 col_n[7] row_n[15] 0.298f
C16820 col_n[4] rowon_n[13] 0.111f
C16821 col_n[0] row_n[11] 0.298f
C16822 sample rowon_n[10] 0.0935f
C16823 col_n[1] row_n[12] 0.298f
C16824 col_n[6] rowon_n[14] 0.111f
C16825 VDD row_n[10] 3.29f
C16826 col[20] a_2475_10186# 0.136f
C16827 col[27] rowoff_n[15] 0.0901f
C16828 rowon_n[7] a_18026_9158# 0.248f
C16829 rowoff_n[6] a_7894_8154# 0.202f
C16830 m2_4168_2378# row_n[0] 0.0128f
C16831 col_n[10] rowoff_n[11] 0.0471f
C16832 a_24050_6146# a_24050_5142# 0.843f
C16833 a_2475_5166# a_12002_5142# 0.316f
C16834 m2_30848_946# m3_31984_1078# 0.0341f
C16835 vcm a_21342_10202# 0.155f
C16836 a_2275_10186# a_35002_10162# 0.136f
C16837 col_n[27] a_2275_16210# 0.113f
C16838 rowoff_n[15] a_18026_17190# 0.294f
C16839 a_17934_10162# a_18330_10202# 0.0313f
C16840 m2_19228_16434# a_19030_16186# 0.165f
C16841 rowoff_n[4] a_16930_6146# 0.202f
C16842 col_n[6] a_8990_5142# 0.251f
C16843 ctop a_34090_5142# 4.06f
C16844 VDD a_8898_9158# 0.181f
C16845 col_n[16] a_19030_17190# 0.251f
C16846 col_n[13] a_15926_7150# 0.0765f
C16847 a_2275_2154# a_2874_2130# 0.136f
C16848 m2_14208_15430# row_n[13] 0.0128f
C16849 a_2475_2154# a_3878_2130# 0.264f
C16850 m2_20232_11414# row_n[9] 0.0128f
C16851 m2_26256_7398# row_n[5] 0.0128f
C16852 m2_32280_3382# row_n[1] 0.0128f
C16853 col[17] a_2275_13198# 0.0899f
C16854 vcm a_14922_4138# 0.1f
C16855 a_14010_7150# a_15014_7150# 0.843f
C16856 a_2475_7174# a_27062_7150# 0.316f
C16857 rowoff_n[2] a_25966_4138# 0.202f
C16858 rowoff_n[9] a_8386_11528# 0.0133f
C16859 rowon_n[1] a_5886_3134# 0.118f
C16860 col[22] a_2275_2154# 0.0899f
C16861 vcm a_3878_13174# 0.1f
C16862 VDD a_34490_4500# 0.0779f
C16863 col_n[7] a_10394_15544# 0.0283f
C16864 ctop a_15014_8154# 4.11f
C16865 a_2275_16210# a_3270_16226# 0.144f
C16866 a_2475_16210# a_5886_16186# 0.264f
C16867 VDD a_23958_13174# 0.181f
C16868 col[26] a_29070_4138# 0.367f
C16869 m2_1732_1950# m2_1732_946# 0.843f
C16870 row_n[8] a_26362_10202# 0.0117f
C16871 rowoff_n[7] a_17422_9520# 0.0133f
C16872 rowoff_n[0] a_35002_2130# 0.202f
C16873 a_2275_4162# a_18026_4138# 0.399f
C16874 m3_34996_5094# ctop 0.209f
C16875 vcm a_29982_8154# 0.1f
C16876 a_4974_9158# a_4974_8154# 0.843f
C16877 rowoff_n[13] a_24450_15544# 0.0133f
C16878 row_n[10] a_16930_12170# 0.0437f
C16879 m2_10192_14426# a_9994_14178# 0.165f
C16880 col_n[7] a_2475_9182# 0.0531f
C16881 vcm a_17326_17230# 0.155f
C16882 a_32994_14178# a_33390_14218# 0.0313f
C16883 rowon_n[14] a_16018_16186# 0.248f
C16884 VDD a_15414_7512# 0.0779f
C16885 m2_1732_1950# m3_1864_1078# 0.0341f
C16886 m2_2736_1950# m3_2868_2082# 3.79f
C16887 rowoff_n[5] a_26458_7512# 0.0133f
C16888 ctop a_30074_12170# 4.11f
C16889 col_n[21] a_24354_4178# 0.084f
C16890 a_2275_18218# a_18330_18234# 0.145f
C16891 row_n[0] a_26970_2130# 0.0437f
C16892 VDD a_4882_16186# 0.181f
C16893 col_n[5] a_7986_15182# 0.251f
C16894 a_2475_1150# a_10906_1126# 0.264f
C16895 a_2275_1150# a_8290_1166# 0.145f
C16896 rowon_n[4] a_26058_6146# 0.248f
C16897 col_n[2] a_4882_5142# 0.0765f
C16898 m2_7180_2378# a_6982_2130# 0.165f
C16899 m2_1732_5966# m2_1732_4962# 0.843f
C16900 col_n[12] a_14922_17190# 0.0765f
C16901 a_2275_6170# a_33086_6146# 0.399f
C16902 a_17934_6146# a_18426_6508# 0.0658f
C16903 a_17022_6146# a_17326_6186# 0.0931f
C16904 m2_29268_10410# a_29070_10162# 0.165f
C16905 rowoff_n[3] a_35494_5504# 0.0133f
C16906 vcm a_10906_11166# 0.1f
C16907 a_29070_11166# a_30074_11166# 0.843f
C16908 VDD a_6982_1126# 0.035f
C16909 a_2275_15206# a_11910_15182# 0.136f
C16910 VDD a_30474_11528# 0.0779f
C16911 ctop a_10998_15182# 4.11f
C16912 row_n[4] a_3970_6146# 0.282f
C16913 col_n[4] a_2275_12194# 0.113f
C16914 rowon_n[6] rowoff_n[6] 20.2f
C16915 a_2275_3158# a_23350_3174# 0.144f
C16916 a_13918_3134# a_14010_3134# 0.326f
C16917 a_2475_3158# a_25966_3134# 0.264f
C16918 col[15] a_18026_2130# 0.367f
C16919 rowoff_n[8] a_27062_10162# 0.294f
C16920 col_n[9] a_2275_1150# 0.113f
C16921 vcm a_1957_5166# 0.139f
C16922 col[25] a_28066_14178# 0.367f
C16923 rowoff_n[11] a_30986_13174# 0.202f
C16924 col[22] a_24962_4138# 0.0682f
C16925 col_n[30] a_2475_18218# 0.0529f
C16926 vcm a_25966_15182# 0.1f
C16927 a_20034_13174# a_20034_12170# 0.843f
C16928 a_2475_12194# a_3970_12170# 0.316f
C16929 a_2275_12194# a_2966_12170# 0.399f
C16930 VDD a_22042_5142# 0.483f
C16931 m2_4744_946# col_n[2] 0.331f
C16932 col_n[24] a_2475_11190# 0.0531f
C16933 m2_2160_18442# VDD 0.0428f
C16934 row_n[15] a_24354_17230# 0.0117f
C16935 ctop a_2275_9182# 0.0683f
C16936 a_13918_17190# a_14314_17230# 0.0313f
C16937 a_2275_17214# a_26970_17190# 0.136f
C16938 VDD a_11398_14540# 0.0779f
C16939 col_n[10] a_13310_2170# 0.084f
C16940 rowon_n[0] a_1957_2154# 0.0172f
C16941 row_n[5] a_35398_7190# 0.0117f
C16942 col_n[20] a_23350_14218# 0.084f
C16943 m2_20232_8402# a_20034_8154# 0.165f
C16944 m3_34568_1078# m3_34996_1078# 0.202f
C16945 col[14] a_2475_8178# 0.136f
C16946 a_32994_10162# a_33486_10524# 0.0658f
C16947 rowoff_n[14] a_12402_16548# 0.0133f
C16948 a_32082_10162# a_32386_10202# 0.0931f
C16949 vcm a_6890_18194# 0.101f
C16950 a_9994_14178# a_10998_14178# 0.843f
C16951 a_2475_14202# a_19030_14178# 0.316f
C16952 m2_16792_946# a_17022_1126# 0.0249f
C16953 VDD a_2874_8154# 0.182f
C16954 row_n[7] a_24962_9158# 0.0437f
C16955 col_n[31] a_34490_8516# 0.0283f
C16956 rowon_n[11] a_24050_13174# 0.248f
C16957 VDD a_26458_18556# 0.0858f
C16958 a_2275_2154# a_31990_2130# 0.136f
C16959 col_n[21] a_2275_14202# 0.113f
C16960 m3_12908_18146# VDD 0.0277f
C16961 vcm a_8990_3134# 0.56f
C16962 col_n[26] a_2275_3158# 0.113f
C16963 a_28978_7150# a_29070_7150# 0.326f
C16964 rowon_n[1] a_34090_3134# 0.248f
C16965 a_2275_11190# a_9994_11166# 0.399f
C16966 col[14] a_17022_12170# 0.367f
C16967 col[11] a_13918_2130# 0.0682f
C16968 row_n[11] a_2475_13198# 0.405f
C16969 col[21] a_23958_14178# 0.0682f
C16970 a_2475_16210# a_34090_16186# 0.316f
C16971 VDD a_18026_12170# 0.483f
C16972 col[11] a_2275_11190# 0.0899f
C16973 m2_3740_18014# m3_3872_18146# 3.79f
C16974 m2_4168_14426# rowon_n[12] 0.0322f
C16975 col_n[29] a_32082_8154# 0.251f
C16976 m2_10192_10410# rowon_n[8] 0.0322f
C16977 m2_16216_6394# rowon_n[4] 0.0322f
C16978 a_23958_4138# a_24354_4178# 0.0313f
C16979 row_n[1] a_12002_3134# 0.282f
C16980 m2_11196_6394# a_10998_6146# 0.165f
C16981 rowon_n[5] a_11910_7150# 0.118f
C16982 vcm a_24050_7150# 0.56f
C16983 rowoff_n[12] a_18938_14178# 0.202f
C16984 col_n[9] a_12306_12210# 0.084f
C16985 vcm row_n[6] 0.616f
C16986 col_n[8] row_n[10] 0.298f
C16987 col_n[18] row_n[15] 0.298f
C16988 col_n[1] rowon_n[6] 0.111f
C16989 col_n[25] col_n[26] 0.0102f
C16990 col_n[3] rowon_n[7] 0.111f
C16991 col_n[13] rowon_n[12] 0.111f
C16992 col_n[5] rowon_n[8] 0.111f
C16993 col_n[4] row_n[8] 0.298f
C16994 col_n[6] row_n[9] 0.298f
C16995 VDD rowon_n[4] 3.04f
C16996 col_n[10] row_n[11] 0.298f
C16997 col_n[12] row_n[12] 0.298f
C16998 col_n[16] row_n[14] 0.298f
C16999 col_n[7] rowon_n[9] 0.111f
C17000 col_n[14] row_n[13] 0.298f
C17001 col_n[19] rowon_n[15] 0.111f
C17002 col_n[15] rowon_n[13] 0.111f
C17003 col_n[0] rowon_n[5] 0.111f
C17004 sample row_n[5] 0.423f
C17005 col_n[2] row_n[7] 0.298f
C17006 col_n[9] rowon_n[10] 0.111f
C17007 col_n[17] rowon_n[14] 0.111f
C17008 col_n[11] rowon_n[11] 0.111f
C17009 col[31] a_2475_10186# 0.136f
C17010 m2_1732_12994# sample 0.2f
C17011 a_13006_13174# a_13310_13214# 0.0931f
C17012 a_13918_13174# a_14410_13536# 0.0658f
C17013 a_2275_13198# a_25054_13174# 0.399f
C17014 m2_34864_6970# ctop 0.0422f
C17015 col_n[21] rowoff_n[11] 0.0471f
C17016 VDD a_33086_16186# 0.483f
C17017 row_n[12] a_32386_14218# 0.0117f
C17018 col_n[20] a_23446_6508# 0.0283f
C17019 col_n[30] a_33486_18556# 0.0283f
C17020 m2_31276_15430# rowon_n[13] 0.0322f
C17021 vcm a_14314_1166# 0.16f
C17022 col_n[1] a_2475_7174# 0.0531f
C17023 m2_6752_946# m3_5880_1078# 0.0341f
C17024 vcm a_4974_10162# 0.56f
C17025 a_9902_10162# a_9994_10162# 0.326f
C17026 a_2275_10186# a_15318_10202# 0.144f
C17027 a_2475_10186# a_17934_10162# 0.264f
C17028 row_n[14] a_22954_16186# 0.0437f
C17029 col[3] a_5978_10162# 0.367f
C17030 row_n[4] a_32994_6146# 0.0437f
C17031 col[28] a_2275_13198# 0.0899f
C17032 col[10] a_12914_12170# 0.0682f
C17033 a_10998_3134# a_10998_2130# 0.843f
C17034 rowon_n[8] a_32082_10162# 0.248f
C17035 m2_1732_3958# a_1957_4162# 0.245f
C17036 col_n[18] a_21038_6146# 0.251f
C17037 vcm a_29374_5182# 0.155f
C17038 a_2275_7174# a_8898_7150# 0.136f
C17039 a_4882_7150# a_5278_7190# 0.0313f
C17040 m2_19804_18014# vcm 0.353f
C17041 col_n[25] a_27974_8154# 0.0765f
C17042 vcm a_20034_14178# 0.56f
C17043 a_2275_12194# a_30378_12210# 0.144f
C17044 a_2475_12194# a_32994_12170# 0.264f
C17045 VDD a_16930_4138# 0.181f
C17046 col_n[5] rowoff_n[12] 0.0471f
C17047 a_28066_17190# a_28370_17230# 0.0931f
C17048 a_28978_17190# a_29470_17552# 0.0658f
C17049 row_n[8] a_9994_10162# 0.282f
C17050 col[1] a_3878_10162# 0.0682f
C17051 rowon_n[12] a_9902_14178# 0.118f
C17052 col_n[9] a_12402_4500# 0.0283f
C17053 m2_29844_946# ctop 0.0428f
C17054 col_n[18] a_2475_9182# 0.0531f
C17055 m2_28840_18014# m2_29844_18014# 0.843f
C17056 vcm a_10298_8194# 0.155f
C17057 col_n[19] a_22442_16548# 0.0283f
C17058 rowoff_n[13] a_6890_15182# 0.202f
C17059 a_2275_9182# a_23958_9158# 0.136f
C17060 rowon_n[2] a_19942_4138# 0.118f
C17061 ctop a_23046_3134# 4.11f
C17062 vcm a_35094_18194# 0.165f
C17063 a_24962_14178# a_25054_14178# 0.326f
C17064 VDD a_31990_8154# 0.181f
C17065 rowoff_n[5] a_8898_7150# 0.202f
C17066 a_1957_18218# a_2161_18218# 0.115f
C17067 col[3] a_2475_17214# 0.136f
C17068 row_n[0] a_7286_2170# 0.0117f
C17069 col[8] a_2475_6170# 0.136f
C17070 a_2475_6170# a_16018_6146# 0.316f
C17071 a_26058_7150# a_26058_6146# 0.843f
C17072 col_n[7] a_9994_4138# 0.251f
C17073 vcm a_25358_12210# 0.155f
C17074 rowoff_n[3] a_17934_5142# 0.202f
C17075 a_19942_11166# a_20338_11206# 0.0313f
C17076 VDD a_23446_2492# 0.0779f
C17077 m2_3164_13422# row_n[11] 0.0128f
C17078 col_n[17] a_20034_16186# 0.251f
C17079 m2_1732_17010# a_2161_17214# 0.0454f
C17080 m2_9188_9406# row_n[7] 0.0128f
C17081 m2_15212_5390# row_n[3] 0.0128f
C17082 ctop a_3970_6146# 4.11f
C17083 col_n[14] a_16930_6146# 0.0765f
C17084 col_n[15] a_2275_12194# 0.113f
C17085 row_n[11] a_30986_13174# 0.0437f
C17086 VDD a_12914_11166# 0.181f
C17087 col_n[24] a_26970_18194# 0.0762f
C17088 row_n[3] rowoff_n[2] 0.085f
C17089 rowon_n[15] a_30074_17190# 0.248f
C17090 col_n[20] a_2275_1150# 0.113f
C17091 a_2275_3158# a_6982_3134# 0.399f
C17092 a_4882_3134# a_5374_3496# 0.0658f
C17093 a_3970_3134# a_4274_3174# 0.0931f
C17094 rowoff_n[8] a_9390_10524# 0.0133f
C17095 rowoff_n[1] a_26970_3134# 0.202f
C17096 vcm a_18938_6146# 0.1f
C17097 a_16018_8154# a_17022_8154# 0.843f
C17098 a_2475_8178# a_31078_8154# 0.316f
C17099 col[5] a_2275_9182# 0.0899f
C17100 vcm a_6282_15222# 0.155f
C17101 col_n[8] a_11398_14540# 0.0283f
C17102 VDD a_4370_5504# 0.0779f
C17103 col_n[31] a_34394_5182# 0.084f
C17104 ctop a_19030_10162# 4.11f
C17105 col[27] a_30074_3134# 0.367f
C17106 row_n[15] a_7986_17190# 0.282f
C17107 m2_30272_14426# row_n[12] 0.0128f
C17108 a_2475_17214# a_9902_17190# 0.264f
C17109 a_5886_17190# a_5978_17190# 0.326f
C17110 a_2275_17214# a_7286_17230# 0.144f
C17111 rowoff_n[6] a_18426_8516# 0.0133f
C17112 VDD a_27974_15182# 0.181f
C17113 m2_35292_10410# row_n[8] 0.0128f
C17114 m3_17928_18146# a_18026_17190# 0.0303f
C17115 col[25] a_2475_8178# 0.136f
C17116 a_2275_5166# a_22042_5142# 0.399f
C17117 row_n[5] a_18026_7150# 0.282f
C17118 rowon_n[9] a_17934_11166# 0.118f
C17119 vcm a_33998_10162# 0.1f
C17120 a_25966_1126# a_26458_1488# 0.0658f
C17121 a_6982_10162# a_6982_9158# 0.843f
C17122 rowoff_n[4] a_27462_6508# 0.0133f
C17123 m2_9764_946# a_2275_1150# 0.28f
C17124 col_n[22] a_25358_3174# 0.084f
C17125 row_n[7] a_5278_9198# 0.0117f
C17126 VDD a_19430_9520# 0.0779f
C17127 col_n[6] a_8990_14178# 0.251f
C17128 ctop a_34090_14178# 4.06f
C17129 col_n[3] a_5886_4138# 0.0765f
C17130 VDD a_8898_18194# 0.343f
C17131 a_2275_2154# a_12306_2170# 0.144f
C17132 a_2475_2154# a_14922_2130# 0.264f
C17133 col_n[13] a_15926_16186# 0.0765f
C17134 m2_4168_1374# VDD 0.0208f
C17135 rowoff_n[9] a_19030_11166# 0.294f
C17136 a_19030_7150# a_19334_7190# 0.0931f
C17137 a_19942_7150# a_20434_7512# 0.0658f
C17138 vcm a_14922_13174# 0.1f
C17139 a_31078_12170# a_32082_12170# 0.843f
C17140 col[22] a_2275_11190# 0.0899f
C17141 VDD a_10998_3134# 0.483f
C17142 m2_10768_18014# a_2275_18218# 0.28f
C17143 a_2275_16210# a_15926_16186# 0.136f
C17144 VDD a_34490_13536# 0.0779f
C17145 rowon_n[3] a_4974_5142# 0.248f
C17146 a_24962_1126# m2_24824_946# 0.225f
C17147 ctop a_15014_17190# 4.06f
C17148 col[16] a_19030_1126# 0.428f
C17149 rowoff_n[7] a_28066_9158# 0.294f
C17150 col[26] a_29070_13174# 0.367f
C17151 a_2475_4162# a_29982_4138# 0.264f
C17152 a_15926_4138# a_16018_4138# 0.326f
C17153 a_2275_4162# a_27366_4178# 0.144f
C17154 col_n[12] rowon_n[6] 0.111f
C17155 col_n[7] row_n[4] 0.298f
C17156 col_n[0] row_n[0] 0.298f
C17157 vcm rowon_n[0] 0.65f
C17158 col_n[3] row_n[2] 0.298f
C17159 VDD sw_n 0.326f
C17160 col_n[1] row_n[1] 0.298f
C17161 col_n[22] rowon_n[11] 0.111f
C17162 col_n[27] row_n[14] 0.298f
C17163 col_n[26] rowon_n[13] 0.111f
C17164 col_n[5] row_n[3] 0.298f
C17165 col_n[9] row_n[5] 0.298f
C17166 col_n[21] row_n[11] 0.298f
C17167 col_n[28] rowon_n[14] 0.111f
C17168 col_n[19] row_n[10] 0.298f
C17169 col_n[25] row_n[13] 0.298f
C17170 col_n[17] row_n[9] 0.298f
C17171 col_n[8] rowon_n[4] 0.111f
C17172 col_n[18] rowon_n[9] 0.111f
C17173 col_n[15] row_n[8] 0.298f
C17174 col_n[30] rowon_n[15] 0.111f
C17175 col_n[11] row_n[6] 0.298f
C17176 col_n[4] rowon_n[2] 0.111f
C17177 col_n[14] rowon_n[7] 0.111f
C17178 col_n[13] row_n[7] 0.298f
C17179 col_n[16] rowon_n[8] 0.111f
C17180 col_n[10] rowon_n[5] 0.111f
C17181 col_n[20] rowon_n[10] 0.111f
C17182 col_n[6] rowon_n[3] 0.111f
C17183 col_n[24] rowon_n[12] 0.111f
C17184 col_n[2] rowon_n[1] 0.111f
C17185 col_n[23] row_n[12] 0.298f
C17186 col_n[29] row_n[15] 0.298f
C17187 col[23] a_25966_3134# 0.0682f
C17188 rowoff_n[13] a_35094_15182# 0.0135f
C17189 vcm a_29982_17190# 0.1f
C17190 a_22042_14178# a_22042_13174# 0.843f
C17191 a_2475_13198# a_7986_13174# 0.316f
C17192 VDD a_26058_7150# 0.483f
C17193 m2_6752_18014# a_2475_18218# 0.286f
C17194 a_2275_18218# a_30986_18194# 0.136f
C17195 a_15926_18194# a_16322_18234# 0.0313f
C17196 col_n[11] a_14314_1166# 0.0839f
C17197 VDD a_15414_16548# 0.0779f
C17198 col_n[12] a_2475_7174# 0.0531f
C17199 a_10906_1126# a_11302_1166# 0.0313f
C17200 a_2275_1150# a_20946_1126# 0.136f
C17201 row_n[12] a_16018_14178# 0.282f
C17202 col_n[21] a_24354_13214# 0.084f
C17203 vcm a_32082_2130# 0.56f
C17204 col_n[2] a_4882_14178# 0.0765f
C17205 m2_3164_9406# a_2966_9158# 0.165f
C17206 m2_21812_946# m2_22240_1374# 0.165f
C17207 row_n[2] a_26058_4138# 0.282f
C17208 a_35002_11166# a_35494_11528# 0.0658f
C17209 VDD a_16322_1166# 0.0149f
C17210 row_n[14] a_3270_16226# 0.0117f
C17211 m2_25252_17438# a_25054_17190# 0.165f
C17212 rowon_n[6] a_25966_8154# 0.118f
C17213 col[2] a_2475_4162# 0.136f
C17214 a_12002_15182# a_13006_15182# 0.843f
C17215 a_2475_15206# a_23046_15182# 0.316f
C17216 VDD a_6982_10162# 0.483f
C17217 row_n[4] a_13310_6186# 0.0117f
C17218 a_2475_18218# a_28978_18194# 0.264f
C17219 a_2275_3158# a_34394_3174# 0.144f
C17220 vcm a_13006_5142# 0.56f
C17221 rowoff_n[10] a_6982_12170# 0.294f
C17222 a_30986_8154# a_31078_8154# 0.326f
C17223 col_n[16] rowoff_n[12] 0.0471f
C17224 a_26970_1126# vcm 0.0989f
C17225 col[15] a_18026_11166# 0.367f
C17226 col_n[9] a_2275_10186# 0.113f
C17227 col[12] a_14922_1126# 0.0682f
C17228 vcm a_1957_14202# 0.139f
C17229 m2_5172_4386# rowon_n[2] 0.0322f
C17230 a_2275_12194# a_14010_12170# 0.399f
C17231 col[22] a_24962_13174# 0.0682f
C17232 rowon_n[10] a_2874_12170# 0.118f
C17233 m2_23820_18014# VDD 1.06f
C17234 VDD a_22042_14178# 0.483f
C17235 col_n[30] a_33086_7150# 0.251f
C17236 a_1957_1150# m2_1732_946# 0.245f
C17237 rowon_n[0] a_13006_2130# 0.248f
C17238 col_n[29] a_2475_9182# 0.0531f
C17239 a_25966_5142# a_26362_5182# 0.0313f
C17240 col_n[10] a_13310_11206# 0.084f
C17241 vcm a_28066_9158# 0.56f
C17242 a_2475_9182# a_6890_9158# 0.264f
C17243 rowoff_n[14] a_23046_16186# 0.294f
C17244 a_2275_9182# a_4274_9198# 0.144f
C17245 m2_16216_15430# a_16018_15182# 0.165f
C17246 m2_14208_17438# rowon_n[15] 0.0322f
C17247 a_15014_14178# a_15318_14218# 0.0931f
C17248 a_2275_14202# a_29070_14178# 0.399f
C17249 col[14] a_2475_17214# 0.136f
C17250 a_15926_14178# a_16418_14540# 0.0658f
C17251 m2_20232_13422# rowon_n[11] 0.0322f
C17252 m2_26256_9406# rowon_n[7] 0.0322f
C17253 m2_32280_5390# rowon_n[3] 0.0322f
C17254 col[19] a_2475_6170# 0.136f
C17255 col_n[21] a_24450_5504# 0.0283f
C17256 VDD a_2874_17190# 0.182f
C17257 col_n[31] a_34490_17552# 0.0283f
C17258 a_22042_2130# a_23046_2130# 0.843f
C17259 vcm rowoff_n[13] 0.533f
C17260 vcm a_18330_3174# 0.155f
C17261 row_n[9] a_24050_11166# 0.282f
C17262 m2_34864_10986# a_35094_11166# 0.0249f
C17263 rowon_n[13] a_23958_15182# 0.118f
C17264 col_n[26] a_2275_12194# 0.113f
C17265 vcm a_8990_12170# 0.56f
C17266 a_11910_11166# a_12002_11166# 0.326f
C17267 a_2475_11190# a_21950_11166# 0.264f
C17268 a_2275_11190# a_19334_11206# 0.144f
C17269 VDD a_5886_2130# 0.181f
C17270 col[3] rowoff_n[9] 0.0901f
C17271 col[1] rowoff_n[7] 0.0901f
C17272 col[0] rowoff_n[6] 0.0901f
C17273 ctop rowoff_n[0] 0.172f
C17274 col[2] rowoff_n[8] 0.0901f
C17275 col[4] a_6982_9158# 0.367f
C17276 col_n[31] a_2275_1150# 0.118f
C17277 row_n[11] a_11302_13214# 0.0117f
C17278 rowon_n[3] a_33998_5142# 0.118f
C17279 m2_17796_18014# m3_18932_18146# 0.0341f
C17280 col[11] a_13918_11166# 0.0682f
C17281 m2_12776_18014# col[10] 0.347f
C17282 col_n[19] a_22042_5142# 0.251f
C17283 a_13006_4138# a_13006_3134# 0.843f
C17284 row_n[1] a_21342_3174# 0.0117f
C17285 col[16] a_2275_9182# 0.0899f
C17286 col_n[29] a_32082_17190# 0.251f
C17287 col_n[26] a_28978_7150# 0.0765f
C17288 vcm a_33390_7190# 0.155f
C17289 a_2275_8178# a_12914_8154# 0.136f
C17290 a_6890_8154# a_7286_8194# 0.0313f
C17291 rowoff_n[12] a_29470_14540# 0.0133f
C17292 m2_7180_13422# a_6982_13174# 0.165f
C17293 vcm a_24050_16186# 0.56f
C17294 a_2275_13198# a_35398_13214# 0.145f
C17295 VDD a_20946_6146# 0.181f
C17296 row_n[3] a_11910_5142# 0.0437f
C17297 rowon_n[7] a_10998_9158# 0.248f
C17298 a_30986_18194# a_31478_18556# 0.0658f
C17299 col_n[10] a_13406_3496# 0.0283f
C17300 a_2475_5166# a_4974_5142# 0.316f
C17301 col_n[20] a_23446_15544# 0.0283f
C17302 m2_21812_946# m3_21944_1078# 3.79f
C17303 m3_30980_18146# m3_31984_18146# 0.202f
C17304 m2_26256_9406# a_26058_9158# 0.165f
C17305 vcm a_14314_10202# 0.155f
C17306 a_2275_10186# a_27974_10162# 0.136f
C17307 rowoff_n[15] a_10998_17190# 0.294f
C17308 col_n[1] a_2475_16210# 0.0531f
C17309 rowoff_n[4] a_9902_6146# 0.202f
C17310 col_n[6] a_2475_5166# 0.0531f
C17311 ctop a_27062_5142# 4.11f
C17312 a_26970_15182# a_27062_15182# 0.326f
C17313 m2_15788_946# a_16018_2130# 0.843f
C17314 m2_4168_3382# row_n[1] 0.0128f
C17315 vcm a_7894_4138# 0.1f
C17316 m2_34864_10986# m2_35292_11414# 0.165f
C17317 a_2475_7174# a_20034_7150# 0.316f
C17318 a_28066_8154# a_28066_7150# 0.843f
C17319 rowoff_n[2] a_18938_4138# 0.202f
C17320 col_n[8] a_10998_3134# 0.251f
C17321 m2_28840_18014# col_n[26] 0.243f
C17322 row_n[6] a_32082_8154# 0.282f
C17323 col_n[18] a_21038_15182# 0.251f
C17324 vcm a_29374_14218# 0.155f
C17325 a_21950_12170# a_22346_12210# 0.0313f
C17326 col_n[15] a_17934_5142# 0.0765f
C17327 rowon_n[10] a_31990_12170# 0.118f
C17328 VDD a_27462_4500# 0.0779f
C17329 col_n[25] a_27974_17190# 0.0765f
C17330 ctop a_7986_8154# 4.11f
C17331 VDD a_16930_13174# 0.181f
C17332 col_n[28] row_n[9] 0.298f
C17333 col_n[15] rowon_n[2] 0.111f
C17334 col_n[20] row_n[5] 0.298f
C17335 col_n[19] rowon_n[4] 0.111f
C17336 col_n[22] row_n[6] 0.298f
C17337 col_n[7] ctop 0.0594f
C17338 col_n[18] row_n[4] 0.298f
C17339 col_n[10] row_n[0] 0.298f
C17340 col_n[12] row_n[1] 0.298f
C17341 col_n[31] rowon_n[10] 0.111f
C17342 col_n[26] row_n[8] 0.298f
C17343 col_n[29] rowon_n[9] 0.111f
C17344 col_n[27] rowon_n[8] 0.111f
C17345 col_n[24] row_n[7] 0.298f
C17346 col_n[23] rowon_n[6] 0.111f
C17347 rowon_n[13] row_n[13] 18.9f
C17348 col_n[30] row_n[10] 0.298f
C17349 vcm col[1] 5.46f
C17350 col_n[25] rowon_n[7] 0.111f
C17351 col_n[11] rowon_n[0] 0.111f
C17352 VDD col[4] 3.83f
C17353 col_n[21] rowon_n[5] 0.111f
C17354 col_n[13] rowon_n[1] 0.111f
C17355 col_n[16] row_n[3] 0.298f
C17356 col_n[14] row_n[2] 0.298f
C17357 col_n[17] rowon_n[3] 0.111f
C17358 row_n[8] a_19334_10202# 0.0117f
C17359 rowoff_n[0] a_27974_2130# 0.202f
C17360 col_n[3] a_2275_8178# 0.113f
C17361 rowoff_n[7] a_10394_9520# 0.0133f
C17362 a_5978_4138# a_6282_4178# 0.0931f
C17363 a_2275_4162# a_10998_4138# 0.399f
C17364 a_6890_4138# a_7382_4500# 0.0658f
C17365 m3_32988_18146# ctop 0.209f
C17366 m2_17220_7398# a_17022_7150# 0.165f
C17367 m2_13204_16434# row_n[14] 0.0128f
C17368 m2_19228_12418# row_n[10] 0.0128f
C17369 vcm a_22954_8154# 0.1f
C17370 a_18026_9158# a_19030_9158# 0.843f
C17371 a_2475_9182# a_35094_9158# 0.0299f
C17372 rowoff_n[13] a_17422_15544# 0.0133f
C17373 m2_25252_8402# row_n[6] 0.0128f
C17374 m2_31276_4386# row_n[2] 0.0128f
C17375 col_n[9] a_12402_13536# 0.0283f
C17376 row_n[10] a_9902_12170# 0.0437f
C17377 vcm a_10298_17230# 0.155f
C17378 col[28] a_31078_2130# 0.367f
C17379 rowon_n[14] a_8990_16186# 0.248f
C17380 VDD a_8386_7512# 0.0779f
C17381 m2_1732_9982# ctop 0.0428f
C17382 col_n[23] a_2475_7174# 0.0531f
C17383 rowoff_n[5] a_19430_7512# 0.0133f
C17384 ctop a_23046_12170# 4.11f
C17385 a_2275_18218# a_11302_18234# 0.145f
C17386 a_7894_18194# a_7986_18194# 0.0991f
C17387 row_n[0] a_19942_2130# 0.0437f
C17388 VDD a_31990_17190# 0.181f
C17389 rowon_n[4] a_19030_6146# 0.248f
C17390 a_2275_6170# a_26058_6146# 0.399f
C17391 col[8] a_2475_15206# 0.136f
C17392 col[13] a_2475_4162# 0.136f
C17393 rowoff_n[3] a_28466_5504# 0.0133f
C17394 a_8990_11166# a_8990_10162# 0.843f
C17395 VDD a_34090_2130# 0.474f
C17396 col_n[23] a_26362_2170# 0.084f
C17397 col_n[7] a_9994_13174# 0.251f
C17398 a_2275_15206# a_4882_15182# 0.136f
C17399 a_2966_15182# a_3970_15182# 0.843f
C17400 VDD a_23446_11528# 0.0779f
C17401 col_n[4] a_6890_3134# 0.0765f
C17402 ctop a_3970_15182# 4.11f
C17403 col_n[14] a_16930_15182# 0.0765f
C17404 a_2275_3158# a_16322_3174# 0.144f
C17405 col_n[20] a_2275_10186# 0.113f
C17406 a_2475_3158# a_18938_3134# 0.264f
C17407 col_n[27] rowoff_n[12] 0.0471f
C17408 rowoff_n[8] a_20034_10162# 0.294f
C17409 a_32082_1126# a_2475_1150# 0.0299f
C17410 en_bit_n[2] a_19334_1166# 0.0266f
C17411 m2_8184_5390# a_7986_5142# 0.165f
C17412 row_n[13] a_30074_15182# 0.282f
C17413 rowoff_n[11] a_23958_13174# 0.202f
C17414 a_21038_8154# a_21342_8194# 0.0931f
C17415 a_21950_8154# a_22442_8516# 0.0658f
C17416 vcm a_18938_15182# 0.1f
C17417 a_33086_13174# a_34090_13174# 0.843f
C17418 VDD a_15014_5142# 0.483f
C17419 a_28978_1126# VDD 0.405f
C17420 col[5] a_2275_18218# 0.0899f
C17421 row_n[15] a_17326_17230# 0.0117f
C17422 a_2275_17214# a_19942_17190# 0.136f
C17423 col[10] a_2275_7174# 0.0899f
C17424 VDD a_4370_14540# 0.0779f
C17425 rowoff_n[6] a_29070_8154# 0.294f
C17426 col_n[31] a_34394_14218# 0.084f
C17427 col[27] a_30074_12170# 0.367f
C17428 col[24] a_26970_2130# 0.0682f
C17429 row_n[5] a_27366_7190# 0.0117f
C17430 a_17934_5142# a_18026_5142# 0.326f
C17431 a_2475_5166# a_33998_5142# 0.264f
C17432 a_2275_5166# a_31382_5182# 0.144f
C17433 m3_20940_1078# m3_21944_1078# 0.202f
C17434 col[25] a_2475_17214# 0.136f
C17435 rowoff_n[14] a_5374_16548# 0.0133f
C17436 m2_1732_15002# a_2475_15206# 0.139f
C17437 col[30] a_2475_6170# 0.136f
C17438 m2_32856_946# a_2275_1150# 0.283f
C17439 m2_34864_946# a_2475_1150# 0.282f
C17440 a_24050_15182# a_24050_14178# 0.843f
C17441 a_2475_14202# a_12002_14178# 0.316f
C17442 VDD a_30074_9158# 0.483f
C17443 row_n[7] a_17934_9158# 0.0437f
C17444 rowon_n[11] a_17022_13174# 0.248f
C17445 col_n[22] a_25358_12210# 0.084f
C17446 col_n[11] rowoff_n[13] 0.0471f
C17447 VDD a_19430_18556# 0.0858f
C17448 a_2275_2154# a_24962_2130# 0.136f
C17449 a_12914_2130# a_13310_2170# 0.0313f
C17450 a_20034_2130# m2_20232_2378# 0.165f
C17451 col_n[3] a_5886_13174# 0.0765f
C17452 m2_27260_1374# VDD 0.0194f
C17453 vcm a_2475_3158# 1.08f
C17454 col[8] rowoff_n[3] 0.0901f
C17455 col[10] rowoff_n[5] 0.0901f
C17456 col[5] rowoff_n[0] 0.0901f
C17457 col[14] rowoff_n[9] 0.0901f
C17458 col[12] rowoff_n[7] 0.0901f
C17459 rowon_n[1] a_27062_3134# 0.248f
C17460 col[9] rowoff_n[4] 0.0901f
C17461 col[13] rowoff_n[8] 0.0901f
C17462 col[11] rowoff_n[6] 0.0901f
C17463 col[6] rowoff_n[1] 0.0901f
C17464 col[7] rowoff_n[2] 0.0901f
C17465 a_2475_11190# a_3878_11166# 0.264f
C17466 a_2275_11190# a_2874_11166# 0.136f
C17467 m2_12776_18014# a_12914_18194# 0.225f
C17468 a_14010_16186# a_15014_16186# 0.843f
C17469 a_2475_16210# a_27062_16186# 0.316f
C17470 VDD a_10998_12170# 0.483f
C17471 col[27] a_2275_9182# 0.0899f
C17472 row_n[1] a_4974_3134# 0.282f
C17473 col[16] a_19030_10162# 0.367f
C17474 vcm a_17022_7150# 0.56f
C17475 rowon_n[5] a_4882_7150# 0.118f
C17476 rowoff_n[12] a_11910_14178# 0.202f
C17477 a_32994_9158# a_33086_9158# 0.326f
C17478 col[23] a_25966_12170# 0.0682f
C17479 a_2275_13198# a_18026_13174# 0.399f
C17480 VDD a_2275_6170# 1.96f
C17481 col_n[31] a_34090_6146# 0.251f
C17482 VDD a_26058_16186# 0.483f
C17483 row_n[12] a_25358_14218# 0.0117f
C17484 col_n[11] a_14314_10202# 0.084f
C17485 m2_3164_15430# rowon_n[13] 0.0322f
C17486 col_n[12] a_2475_16210# 0.0531f
C17487 vcm a_7286_1166# 0.16f
C17488 m2_9188_11414# rowon_n[9] 0.0322f
C17489 a_27974_6146# a_28370_6186# 0.0313f
C17490 m2_15212_7398# rowon_n[5] 0.0322f
C17491 m2_1732_7974# sample_n 0.0522f
C17492 col_n[17] a_2475_5166# 0.0531f
C17493 m2_21236_3382# rowon_n[1] 0.0322f
C17494 m2_1732_3958# rowoff_n[2] 0.415f
C17495 vcm a_32082_11166# 0.56f
C17496 a_2275_10186# a_8290_10202# 0.144f
C17497 a_2475_10186# a_10906_10162# 0.264f
C17498 row_n[14] a_15926_16186# 0.0437f
C17499 col_n[22] a_25454_4500# 0.0283f
C17500 a_17022_15182# a_17326_15222# 0.0931f
C17501 a_17934_15182# a_18426_15544# 0.0658f
C17502 a_2275_15206# a_33086_15182# 0.399f
C17503 row_n[4] a_25966_6146# 0.0437f
C17504 col[2] a_2475_13198# 0.136f
C17505 a_24050_3134# a_25054_3134# 0.843f
C17506 col[7] a_2475_2154# 0.136f
C17507 rowon_n[8] a_25054_10162# 0.248f
C17508 vcm a_22346_5182# 0.155f
C17509 a_2475_7174# a_1957_7174# 0.0734f
C17510 m2_5748_18014# vcm 0.353f
C17511 m2_30272_16434# rowon_n[14] 0.0322f
C17512 col[5] a_7986_8154# 0.367f
C17513 m2_35292_12418# rowon_n[10] 0.0322f
C17514 vcm a_13006_14178# 0.56f
C17515 a_13918_12170# a_14010_12170# 0.326f
C17516 a_2275_12194# a_23350_12210# 0.144f
C17517 a_2475_12194# a_25966_12170# 0.264f
C17518 VDD a_9902_4138# 0.181f
C17519 col_n[6] col[6] 0.489f
C17520 col_n[18] ctop 0.0594f
C17521 col_n[22] rowon_n[0] 0.111f
C17522 col_n[30] rowon_n[4] 0.111f
C17523 col_n[27] row_n[3] 0.298f
C17524 col_n[23] row_n[1] 0.298f
C17525 vcm col[12] 5.46f
C17526 col_n[24] rowon_n[1] 0.111f
C17527 col_n[31] row_n[5] 0.298f
C17528 col_n[28] rowon_n[3] 0.111f
C17529 col_n[26] rowon_n[2] 0.111f
C17530 col_n[29] row_n[4] 0.298f
C17531 VDD col[15] 3.83f
C17532 col_n[25] row_n[2] 0.298f
C17533 col_n[21] row_n[0] 0.298f
C17534 col[12] a_14922_10162# 0.0682f
C17535 col_n[14] a_2275_8178# 0.113f
C17536 col_n[20] a_23046_4138# 0.251f
C17537 row_n[8] a_2874_10162# 0.0436f
C17538 col_n[30] a_33086_16186# 0.251f
C17539 rowon_n[12] a_2161_14202# 0.0177f
C17540 a_15014_5142# a_15014_4138# 0.843f
C17541 col_n[27] a_29982_6146# 0.0765f
C17542 m2_1732_6970# a_2966_7150# 0.843f
C17543 vcm a_3270_8194# 0.155f
C17544 m2_21812_18014# m2_22816_18014# 0.843f
C17545 a_2275_9182# a_16930_9158# 0.136f
C17546 a_8898_9158# a_9294_9198# 0.0313f
C17547 col[4] a_2275_5166# 0.0899f
C17548 rowon_n[2] a_12914_4138# 0.118f
C17549 ctop a_16018_3134# 4.11f
C17550 a_27366_1166# col_n[24] 0.0839f
C17551 vcm a_28066_18194# 0.165f
C17552 VDD a_24962_8154# 0.181f
C17553 col_n[11] a_14410_2492# 0.0283f
C17554 a_27062_2130# a_27366_2170# 0.0931f
C17555 a_27974_2130# a_28466_2492# 0.0658f
C17556 col[19] a_2475_15206# 0.136f
C17557 col_n[21] a_24450_14540# 0.0283f
C17558 m3_31984_1078# VDD 0.0157f
C17559 col[24] a_2475_4162# 0.136f
C17560 row_n[9] a_33390_11206# 0.0117f
C17561 vcm a_30986_3134# 0.1f
C17562 a_4974_6146# a_5978_6146# 0.843f
C17563 a_2475_6170# a_8990_6146# 0.316f
C17564 m2_34864_9982# a_2275_10186# 0.278f
C17565 rowoff_n[3] a_10906_5142# 0.202f
C17566 vcm a_18330_12210# 0.155f
C17567 a_2275_11190# a_31990_11166# 0.136f
C17568 VDD a_16418_2492# 0.0779f
C17569 m2_31852_18014# a_31990_18194# 0.225f
C17570 m2_8760_18014# a_8990_17190# 0.843f
C17571 sample a_2161_8178# 0.0858f
C17572 ctop a_31078_7150# 4.11f
C17573 row_n[11] a_23958_13174# 0.0437f
C17574 a_28978_16186# a_29070_16186# 0.326f
C17575 VDD a_5886_11166# 0.181f
C17576 rowon_n[12] rowoff_n[12] 20.2f
C17577 m2_32856_18014# m3_31984_18146# 0.0341f
C17578 col_n[31] a_2275_10186# 0.113f
C17579 rowon_n[15] a_23046_17190# 0.248f
C17580 col_n[9] a_12002_2130# 0.251f
C17581 a_27974_1126# col[25] 0.0682f
C17582 row_n[1] a_33998_3134# 0.0437f
C17583 rowoff_n[1] a_19942_3134# 0.202f
C17584 rowoff_n[8] a_1957_10186# 0.0219f
C17585 rowon_n[5] a_33086_7150# 0.248f
C17586 col_n[19] a_22042_14178# 0.251f
C17587 vcm a_11910_6146# 0.1f
C17588 a_2475_8178# a_24050_8154# 0.316f
C17589 a_30074_9158# a_30074_8154# 0.843f
C17590 m2_29844_946# col[27] 0.425f
C17591 col_n[16] a_18938_4138# 0.0765f
C17592 col[16] a_2275_18218# 0.0899f
C17593 vcm a_33390_16226# 0.155f
C17594 col_n[26] a_28978_16186# 0.0765f
C17595 col[21] a_2275_7174# 0.0899f
C17596 a_23958_13174# a_24354_13214# 0.0313f
C17597 VDD a_31478_6508# 0.0779f
C17598 ctop a_12002_10162# 4.11f
C17599 m2_2160_14426# row_n[12] 0.0194f
C17600 rowoff_n[6] a_11398_8516# 0.0133f
C17601 m2_8184_10410# row_n[8] 0.0128f
C17602 VDD a_20946_15182# 0.181f
C17603 m2_14208_6394# row_n[4] 0.0128f
C17604 m2_19228_2378# row_n[0] 0.0128f
C17605 row_n[5] a_10998_7150# 0.282f
C17606 a_7986_5142# a_8290_5182# 0.0931f
C17607 a_8898_5142# a_9390_5504# 0.0658f
C17608 a_2275_5166# a_15014_5142# 0.399f
C17609 m2_34864_2954# vcm 0.395f
C17610 m3_1864_9110# m3_1864_8106# 0.202f
C17611 m2_34864_8978# a_35002_9158# 0.225f
C17612 col_n[10] a_13406_12532# 0.0283f
C17613 rowon_n[9] a_10906_11166# 0.118f
C17614 vcm a_26970_10162# 0.1f
C17615 a_20034_10162# a_21038_10162# 0.843f
C17616 m2_22240_16434# a_22042_16186# 0.165f
C17617 rowoff_n[4] a_20434_6508# 0.0133f
C17618 col_n[22] rowoff_n[13] 0.0471f
C17619 m2_33860_18014# ctop 0.0418f
C17620 VDD a_12402_9520# 0.0779f
C17621 col_n[6] a_2475_14202# 0.0531f
C17622 ctop a_27062_14178# 4.11f
C17623 col_n[11] a_2475_3158# 0.0531f
C17624 col[20] rowoff_n[4] 0.0901f
C17625 col[16] rowoff_n[0] 0.0901f
C17626 col[17] rowoff_n[1] 0.0901f
C17627 col[23] rowoff_n[7] 0.0901f
C17628 col[18] rowoff_n[2] 0.0901f
C17629 col[22] rowoff_n[6] 0.0901f
C17630 col[25] rowoff_n[9] 0.0901f
C17631 col[24] rowoff_n[8] 0.0901f
C17632 col[19] rowoff_n[3] 0.0901f
C17633 col[21] rowoff_n[5] 0.0901f
C17634 a_4882_2130# a_4974_2130# 0.326f
C17635 a_3878_2130# a_4274_2170# 0.0313f
C17636 m2_29268_15430# row_n[13] 0.0128f
C17637 a_2475_2154# a_7894_2130# 0.264f
C17638 a_2275_2154# a_5278_2170# 0.144f
C17639 m2_34864_10986# row_n[9] 0.267f
C17640 rowoff_n[2] a_29470_4500# 0.0133f
C17641 col[2] a_2475_18218# 0.136f
C17642 rowoff_n[9] a_12002_11166# 0.294f
C17643 a_2275_7174# a_30074_7150# 0.399f
C17644 vcm a_7894_13174# 0.1f
C17645 col_n[8] a_10998_12170# 0.251f
C17646 a_10998_12170# a_10998_11166# 0.843f
C17647 VDD a_3970_3134# 0.483f
C17648 col_n[5] a_7894_2130# 0.0765f
C17649 col_n[15] a_17934_14178# 0.0765f
C17650 a_2275_16210# a_8898_16186# 0.136f
C17651 a_4882_16186# a_5278_16226# 0.0313f
C17652 VDD a_27462_13536# 0.0779f
C17653 row_n[8] a_31990_10162# 0.0437f
C17654 ctop a_7986_17190# 4.06f
C17655 rowoff_n[7] a_21038_9158# 0.294f
C17656 rowon_n[12] a_31078_14178# 0.248f
C17657 a_2475_4162# a_22954_4138# 0.264f
C17658 a_2275_4162# a_20338_4178# 0.144f
C17659 m3_8892_1078# ctop 0.21f
C17660 col_n[3] a_2275_17214# 0.113f
C17661 a_23046_9158# a_23350_9198# 0.0931f
C17662 a_23958_9158# a_24450_9520# 0.0658f
C17663 rowoff_n[13] a_28066_15182# 0.294f
C17664 col_n[8] a_2275_6170# 0.113f
C17665 m2_13204_14426# a_13006_14178# 0.165f
C17666 col_n[6] rowoff_n[14] 0.0471f
C17667 vcm a_22954_17190# 0.1f
C17668 VDD a_19030_7150# 0.483f
C17669 rowoff_n[5] a_30074_7150# 0.294f
C17670 col[28] a_31078_11166# 0.367f
C17671 col[9] rowoff_n[10] 0.0901f
C17672 a_2275_18218# a_23958_18194# 0.136f
C17673 col_n[23] a_2475_16210# 0.0531f
C17674 VDD a_8386_16548# 0.0779f
C17675 a_2275_1150# a_13918_1126# 0.136f
C17676 row_n[12] a_8990_14178# 0.282f
C17677 col_n[28] a_2475_5166# 0.0531f
C17678 m2_10192_2378# a_9994_2130# 0.165f
C17679 vcm a_25054_2130# 0.56f
C17680 a_2275_6170# a_2275_5166# 0.0715f
C17681 a_19942_6146# a_20034_6146# 0.326f
C17682 m2_32280_10410# a_32082_10162# 0.165f
C17683 row_n[2] a_19030_4138# 0.282f
C17684 VDD a_9294_1166# 0.0149f
C17685 rowon_n[6] a_18938_8154# 0.118f
C17686 m2_27836_18014# a_28066_17190# 0.843f
C17687 m2_1732_4962# VDD 0.856f
C17688 col[13] a_2475_13198# 0.136f
C17689 a_26058_16186# a_26058_15182# 0.843f
C17690 a_2475_15206# a_16018_15182# 0.316f
C17691 VDD a_34090_11166# 0.483f
C17692 col_n[23] a_26362_11206# 0.084f
C17693 col[18] a_2475_2154# 0.136f
C17694 rowon_n[0] m2_26256_2378# 0.0322f
C17695 row_n[4] a_6282_6186# 0.0117f
C17696 col_n[4] a_6890_12170# 0.0765f
C17697 a_2275_3158# a_28978_3134# 0.136f
C17698 a_14922_3134# a_15318_3174# 0.0313f
C17699 a_2475_18218# a_21950_18194# 0.264f
C17700 vcm a_5978_5142# 0.56f
C17701 rowoff_n[11] a_34490_13536# 0.0133f
C17702 vcm col[23] 5.46f
C17703 col_n[11] col[12] 7.13f
C17704 VDD col[26] 3.83f
C17705 col_n[31] sw 0.0457f
C17706 col_n[29] ctop 0.0602f
C17707 m2_4168_12418# a_3970_12170# 0.165f
C17708 col_n[25] a_2275_8178# 0.113f
C17709 a_4882_12170# a_5374_12532# 0.0658f
C17710 a_3970_12170# a_4274_12210# 0.0931f
C17711 a_2275_12194# a_6982_12170# 0.399f
C17712 m2_9764_18014# VDD 1f
C17713 row_n[15] a_29982_17190# 0.0437f
C17714 a_2475_17214# a_31078_17190# 0.316f
C17715 a_16018_17190# a_17022_17190# 0.843f
C17716 VDD a_15014_14178# 0.483f
C17717 rowon_n[0] a_5978_2130# 0.248f
C17718 col[17] a_20034_9158# 0.367f
C17719 col[10] a_2275_16210# 0.0899f
C17720 col[15] a_2275_5166# 0.0899f
C17721 m2_23244_8402# a_23046_8154# 0.165f
C17722 col[24] a_26970_11166# 0.0682f
C17723 vcm a_21038_9158# 0.56f
C17724 a_34090_10162# a_34394_10202# 0.0931f
C17725 a_35002_10162# a_35094_10162# 0.0991f
C17726 rowoff_n[14] a_16018_16186# 0.294f
C17727 a_2275_14202# a_22042_14178# 0.399f
C17728 col[30] a_2475_15206# 0.136f
C17729 m2_4168_5390# rowon_n[3] 0.0322f
C17730 m2_7756_946# vcm 0.353f
C17731 VDD a_30074_18194# 0.0356f
C17732 col_n[12] a_15318_9198# 0.084f
C17733 a_2475_2154# a_2475_1150# 0.0646f
C17734 m3_27968_18146# VDD 0.0646f
C17735 row_n[9] a_17022_11166# 0.282f
C17736 vcm a_11302_3174# 0.155f
C17737 a_29982_7150# a_30378_7190# 0.0313f
C17738 rowon_n[13] a_16930_15182# 0.118f
C17739 vcm a_2475_12194# 1.08f
C17740 a_2475_11190# a_14922_11166# 0.264f
C17741 a_2275_11190# a_12306_11206# 0.144f
C17742 col_n[23] a_26458_3496# 0.0283f
C17743 VDD a_32994_3134# 0.181f
C17744 col_n[5] a_2475_1150# 0.0531f
C17745 a_19030_16186# a_19334_16226# 0.0931f
C17746 a_19942_16186# a_20434_16548# 0.0658f
C17747 row_n[11] a_4274_13214# 0.0117f
C17748 rowon_n[3] a_26970_5142# 0.118f
C17749 m2_8760_18014# m3_8892_18146# 3.79f
C17750 m2_19228_14426# rowon_n[12] 0.0322f
C17751 m2_25252_10410# rowon_n[8] 0.0322f
C17752 m2_31276_6394# rowon_n[4] 0.0322f
C17753 a_26058_4138# a_27062_4138# 0.843f
C17754 col[27] a_2275_18218# 0.0899f
C17755 row_n[1] a_14314_3174# 0.0117f
C17756 m2_14208_6394# a_14010_6146# 0.165f
C17757 vcm a_26362_7190# 0.155f
C17758 col[6] a_8990_7150# 0.367f
C17759 rowoff_n[12] a_22442_14540# 0.0133f
C17760 a_2275_8178# a_5886_8154# 0.136f
C17761 col[13] a_15926_9158# 0.0682f
C17762 vcm a_17022_16186# 0.56f
C17763 a_2275_13198# a_27366_13214# 0.144f
C17764 a_15926_13174# a_16018_13174# 0.326f
C17765 a_2475_13198# a_29982_13174# 0.264f
C17766 VDD a_13918_6146# 0.181f
C17767 row_n[3] a_4882_5142# 0.0437f
C17768 col_n[21] a_24050_3134# 0.251f
C17769 rowon_n[7] a_3970_9158# 0.248f
C17770 col[17] a_18938_1126# 0.011f
C17771 VDD a_2275_15206# 1.96f
C17772 col_n[31] a_34090_15182# 0.251f
C17773 col_n[28] a_30986_5142# 0.0765f
C17774 col_n[2] a_2275_4162# 0.113f
C17775 vcm a_19942_1126# 0.0951f
C17776 a_17022_6146# a_17022_5142# 0.843f
C17777 col_n[1] a_4274_7190# 0.084f
C17778 m3_16924_18146# m3_17928_18146# 0.202f
C17779 m2_11772_946# m3_10900_1078# 0.0341f
C17780 vcm a_7286_10202# 0.155f
C17781 a_10906_10162# a_11302_10202# 0.0313f
C17782 rowoff_n[15] a_3970_17190# 0.294f
C17783 a_2275_10186# a_20946_10162# 0.136f
C17784 col_n[17] a_2475_14202# 0.0531f
C17785 rowoff_n[4] a_2161_6170# 0.0226f
C17786 ctop a_20034_5142# 4.11f
C17787 col_n[22] a_2475_3158# 0.0531f
C17788 VDD a_28978_10162# 0.181f
C17789 col[30] rowoff_n[3] 0.0901f
C17790 col[31] rowoff_n[4] 0.0901f
C17791 col[29] rowoff_n[2] 0.0901f
C17792 col[27] rowoff_n[0] 0.0901f
C17793 col[28] rowoff_n[1] 0.0901f
C17794 sample_n rowoff_n[5] 0.14f
C17795 col_n[12] a_15414_1488# 0.0283f
C17796 sw a_2275_1150# 0.0408f
C17797 col_n[22] a_25454_13536# 0.0283f
C17798 col[13] a_2475_18218# 0.136f
C17799 a_29070_3134# a_29374_3174# 0.0931f
C17800 a_29982_3134# a_30474_3496# 0.0658f
C17801 m2_5172_4386# a_4974_4138# 0.165f
C17802 vcm a_35002_5142# 0.101f
C17803 col[7] a_2475_11190# 0.136f
C17804 rowoff_n[10] a_28978_12170# 0.202f
C17805 a_2475_7174# a_13006_7150# 0.316f
C17806 rowoff_n[2] a_11910_4138# 0.202f
C17807 a_6982_7150# a_7986_7150# 0.843f
C17808 col_n[0] a_3366_7512# 0.0283f
C17809 row_n[6] a_25054_8154# 0.282f
C17810 vcm a_22346_14218# 0.155f
C17811 a_2275_12194# a_34394_12210# 0.144f
C17812 VDD a_20434_4500# 0.0779f
C17813 rowon_n[10] a_24962_12170# 0.118f
C17814 col[5] a_7986_17190# 0.367f
C17815 col[2] a_4882_7150# 0.0682f
C17816 a_30986_17190# a_31078_17190# 0.326f
C17817 VDD a_9902_13174# 0.181f
C17818 col_n[14] a_2275_17214# 0.113f
C17819 row_n[8] a_12306_10202# 0.0117f
C17820 rowon_n[0] a_35002_2130# 0.118f
C17821 rowoff_n[0] a_20946_2130# 0.202f
C17822 rowoff_n[7] a_2966_9158# 0.294f
C17823 col_n[19] a_2275_6170# 0.113f
C17824 a_2275_4162# a_3970_4138# 0.399f
C17825 col_n[20] a_23046_13174# 0.251f
C17826 m3_4876_18146# ctop 0.209f
C17827 col_n[17] rowoff_n[14] 0.0471f
C17828 col_n[17] a_19942_3134# 0.0765f
C17829 vcm a_15926_8154# 0.1f
C17830 m2_32856_18014# m2_33284_18442# 0.165f
C17831 a_2475_9182# a_28066_9158# 0.316f
C17832 rowoff_n[13] a_10394_15544# 0.0133f
C17833 a_32082_10162# a_32082_9158# 0.843f
C17834 col_n[27] a_29982_15182# 0.0765f
C17835 m2_3164_4386# row_n[2] 0.0128f
C17836 row_n[10] a_2161_12194# 0.0221f
C17837 col[20] rowoff_n[10] 0.0901f
C17838 vcm a_3270_17230# 0.155f
C17839 a_25966_14178# a_26362_14218# 0.0313f
C17840 rowon_n[14] a_2475_16210# 0.31f
C17841 VDD a_35494_8516# 0.106f
C17842 col[4] a_2275_14202# 0.0899f
C17843 rowoff_n[5] a_12402_7512# 0.0133f
C17844 ctop a_16018_12170# 4.11f
C17845 col[9] a_2275_3158# 0.0899f
C17846 a_2275_18218# a_4274_18234# 0.145f
C17847 row_n[0] a_12914_2130# 0.0437f
C17848 VDD a_24962_17190# 0.181f
C17849 rowon_n[4] a_12002_6146# 0.248f
C17850 col_n[11] a_14410_11528# 0.0283f
C17851 a_2275_6170# a_19030_6146# 0.399f
C17852 a_10906_6146# a_11398_6508# 0.0658f
C17853 a_9994_6146# a_10298_6186# 0.0931f
C17854 col[24] a_2475_13198# 0.136f
C17855 rowoff_n[3] a_21438_5504# 0.0133f
C17856 vcm a_30986_12170# 0.1f
C17857 a_22042_11166# a_23046_11166# 0.843f
C17858 m2_12200_17438# row_n[15] 0.0128f
C17859 VDD a_27062_2130# 0.483f
C17860 col[29] a_2475_2154# 0.136f
C17861 m2_18224_13422# row_n[11] 0.0128f
C17862 m2_24248_9406# row_n[7] 0.0128f
C17863 m2_30272_5390# row_n[3] 0.0128f
C17864 VDD a_16418_11528# 0.0779f
C17865 m2_34864_17010# m3_34996_18146# 0.0341f
C17866 sample a_2161_17214# 0.0858f
C17867 ctop a_31078_16186# 4.11f
C17868 a_2475_3158# a_11910_3134# 0.264f
C17869 rowon_n[14] col[0] 0.0318f
C17870 a_2475_18218# a_3878_18194# 0.264f
C17871 col_n[1] rowoff_n[15] 0.0471f
C17872 a_6890_3134# a_6982_3134# 0.326f
C17873 rowon_n[5] rowon_n[4] 0.0632f
C17874 row_n[15] col[1] 0.0342f
C17875 rowon_n[11] ctop 0.203f
C17876 col_n[17] col[17] 0.414f
C17877 a_2275_3158# a_9294_3174# 0.144f
C17878 rowon_n[15] col[2] 0.0323f
C17879 rowoff_n[1] a_30474_3496# 0.0133f
C17880 rowoff_n[8] a_13006_10162# 0.294f
C17881 a_25054_1126# a_2475_1150# 0.0299f
C17882 m2_1732_4962# a_2275_5166# 0.191f
C17883 row_n[13] a_23046_15182# 0.282f
C17884 rowoff_n[11] a_16930_13174# 0.202f
C17885 a_2275_8178# a_34090_8154# 0.399f
C17886 col_n[9] a_12002_11166# 0.251f
C17887 col[4] rowoff_n[11] 0.0901f
C17888 col_n[6] a_8898_1126# 0.0765f
C17889 vcm a_11910_15182# 0.1f
C17890 a_13006_13174# a_13006_12170# 0.843f
C17891 VDD a_7986_5142# 0.483f
C17892 col_n[16] a_18938_13174# 0.0765f
C17893 row_n[3] a_33086_5142# 0.282f
C17894 row_n[15] a_10298_17230# 0.0117f
C17895 col[21] a_2275_16210# 0.0899f
C17896 rowon_n[7] a_32994_9158# 0.118f
C17897 a_6890_17190# a_7286_17230# 0.0313f
C17898 a_2275_17214# a_12914_17190# 0.136f
C17899 VDD a_31478_15544# 0.0779f
C17900 rowoff_n[6] a_22042_8154# 0.294f
C17901 col[26] a_2275_5166# 0.0899f
C17902 m3_20940_18146# a_21038_17190# 0.0303f
C17903 a_2475_5166# a_26970_5142# 0.264f
C17904 a_2275_5166# a_24354_5182# 0.144f
C17905 row_n[5] a_20338_7190# 0.0117f
C17906 m3_6884_1078# m3_7888_1078# 0.202f
C17907 vcm a_2966_9158# 0.56f
C17908 a_27974_1126# a_28066_1126# 0.0991f
C17909 a_25054_10162# a_25358_10202# 0.0931f
C17910 a_25966_10162# a_26458_10524# 0.0658f
C17911 rowoff_n[15] a_32994_17190# 0.202f
C17912 rowoff_n[4] a_31078_6146# 0.294f
C17913 a_2475_14202# a_4974_14178# 0.316f
C17914 m2_7756_946# a_7894_1126# 0.225f
C17915 VDD a_23046_9158# 0.483f
C17916 col[29] a_32082_10162# 0.367f
C17917 row_n[7] a_10906_9158# 0.0437f
C17918 rowon_n[11] a_9994_13174# 0.248f
C17919 VDD a_12402_18556# 0.0858f
C17920 a_2275_2154# a_17934_2130# 0.136f
C17921 col_n[11] a_2475_12194# 0.0531f
C17922 m2_11772_946# VDD 1f
C17923 vcm a_29070_4138# 0.56f
C17924 rowon_n[1] a_20034_3134# 0.248f
C17925 a_21950_7150# a_22042_7150# 0.326f
C17926 col_n[16] a_2475_1150# 0.0486f
C17927 col_n[24] a_27366_10202# 0.084f
C17928 m2_7756_18014# a_7986_18194# 0.0249f
C17929 a_2475_16210# a_20034_16186# 0.316f
C17930 a_28066_17190# a_28066_16186# 0.843f
C17931 VDD a_3970_12170# 0.483f
C17932 col_n[5] a_7894_11166# 0.0765f
C17933 a_26362_1166# m2_25828_946# 0.087f
C17934 col[1] a_2475_9182# 0.136f
C17935 m2_1732_11990# col[0] 0.0137f
C17936 a_16930_4138# a_17326_4178# 0.0313f
C17937 a_2275_4162# a_32994_4138# 0.136f
C17938 m2_34864_6970# a_34090_7150# 0.843f
C17939 vcm a_9994_7150# 0.56f
C17940 rowoff_n[12] a_4882_14178# 0.202f
C17941 row_n[10] a_31078_12170# 0.282f
C17942 col_n[8] a_2275_15206# 0.113f
C17943 a_2275_13198# a_10998_13174# 0.399f
C17944 a_6890_13174# a_7382_13536# 0.0658f
C17945 rowon_n[14] a_30986_16186# 0.118f
C17946 a_5978_13174# a_6282_13214# 0.0931f
C17947 col_n[13] a_2275_4162# 0.113f
C17948 VDD a_19030_16186# 0.483f
C17949 col[18] a_21038_8154# 0.367f
C17950 row_n[12] a_18330_14218# 0.0117f
C17951 vcm a_35398_2170# 0.161f
C17952 col[25] a_27974_10162# 0.0682f
C17953 col_n[28] a_2475_14202# 0.0531f
C17954 m2_1732_5966# vcm 0.316f
C17955 col_n[0] a_3270_4178# 0.084f
C17956 row_n[2] a_28370_4178# 0.0117f
C17957 vcm a_25054_11166# 0.56f
C17958 VDD a_21950_1126# 0.405f
C17959 col[3] a_2275_1150# 0.0899f
C17960 row_n[14] a_8898_16186# 0.0437f
C17961 m2_28264_17438# a_28066_17190# 0.165f
C17962 a_2275_15206# a_26058_15182# 0.399f
C17963 col[24] a_2475_18218# 0.136f
C17964 m2_34864_13998# m3_34996_15134# 0.0341f
C17965 col_n[13] a_16322_8194# 0.084f
C17966 row_n[4] a_18938_6146# 0.0437f
C17967 col[18] a_2475_11190# 0.136f
C17968 rowon_n[8] a_18026_10162# 0.248f
C17969 a_3970_3134# a_3970_2130# 0.843f
C17970 vcm a_15318_5182# 0.155f
C17971 a_31990_8154# a_32386_8194# 0.0313f
C17972 col_n[24] a_27462_2492# 0.0283f
C17973 m2_2160_16434# rowon_n[14] 0.0219f
C17974 m2_8184_12418# rowon_n[10] 0.0322f
C17975 m2_14208_8402# rowon_n[6] 0.0322f
C17976 vcm a_5978_14178# 0.56f
C17977 a_2475_12194# a_18938_12170# 0.264f
C17978 a_2275_12194# a_16322_12210# 0.144f
C17979 m2_20232_4386# rowon_n[2] 0.0322f
C17980 VDD a_2161_4162# 0.187f
C17981 m2_31276_18442# VDD 0.0456f
C17982 col_n[25] a_2275_17214# 0.113f
C17983 a_21950_17190# a_22442_17552# 0.0658f
C17984 a_21038_17190# a_21342_17230# 0.0931f
C17985 col_n[30] a_2275_6170# 0.113f
C17986 col_n[28] rowoff_n[14] 0.0471f
C17987 rowoff_n[0] a_2275_2154# 0.151f
C17988 en_bit_n[0] a_20434_1488# 0.018f
C17989 col[7] a_9994_6146# 0.367f
C17990 a_28066_5142# a_29070_5142# 0.843f
C17991 col[31] rowoff_n[10] 0.0901f
C17992 vcm a_30378_9198# 0.155f
C17993 m2_14784_18014# m2_15788_18014# 0.843f
C17994 VDD m2_2736_946# 1f
C17995 a_2275_9182# a_9902_9158# 0.136f
C17996 col[14] a_16930_8154# 0.0682f
C17997 col[15] a_2275_14202# 0.0899f
C17998 m2_19228_15430# a_19030_15182# 0.165f
C17999 rowon_n[2] a_5886_4138# 0.118f
C18000 col[20] a_2275_3158# 0.0899f
C18001 ctop a_8990_3134# 4.11f
C18002 vcm a_21038_18194# 0.165f
C18003 col_n[22] a_25054_2130# 0.251f
C18004 m2_29268_17438# rowon_n[15] 0.0322f
C18005 a_2275_14202# a_31382_14218# 0.144f
C18006 a_2475_14202# a_33998_14178# 0.264f
C18007 a_17934_14178# a_18026_14178# 0.326f
C18008 m2_34864_12994# rowon_n[11] 0.231f
C18009 VDD a_17934_8154# 0.181f
C18010 m2_30848_946# vcm 0.353f
C18011 col_n[29] a_31990_4138# 0.0765f
C18012 col_n[2] a_5278_6186# 0.084f
C18013 m3_3872_1078# VDD 0.0118f
C18014 col_n[12] a_15318_18234# 0.084f
C18015 vcm a_23958_3134# 0.1f
C18016 row_n[9] a_26362_11206# 0.0117f
C18017 a_19030_7150# a_19030_6146# 0.843f
C18018 en_bit_n[1] a_18026_1126# 0.208f
C18019 vcm a_11302_12210# 0.155f
C18020 rowoff_n[3] a_3366_5504# 0.0133f
C18021 a_12914_11166# a_13310_11206# 0.0313f
C18022 a_2275_11190# a_24962_11166# 0.136f
C18023 VDD a_9390_2492# 0.0779f
C18024 m2_26832_18014# a_27062_18194# 0.0249f
C18025 ctop a_24050_7150# 4.11f
C18026 row_n[11] a_16930_13174# 0.0437f
C18027 VDD a_32994_12170# 0.181f
C18028 col_n[23] a_26458_12532# 0.0283f
C18029 rowon_n[2] row_n[2] 18.9f
C18030 rowon_n[12] col[7] 0.0323f
C18031 row_n[11] col[4] 0.0342f
C18032 row_n[15] col[12] 0.0342f
C18033 col_n[5] a_2475_10186# 0.0531f
C18034 rowon_n[13] col[9] 0.0323f
C18035 row_n[6] ctop 0.186f
C18036 row_n[12] col[6] 0.0342f
C18037 col_n[22] col[23] 7.13f
C18038 row_n[13] col[8] 0.0342f
C18039 rowon_n[9] col[1] 0.0323f
C18040 rowon_n[14] col[11] 0.0323f
C18041 m2_22816_18014# m3_23952_18146# 0.0341f
C18042 row_n[10] col[2] 0.0342f
C18043 rowon_n[15] col[13] 0.0323f
C18044 row_n[14] col[10] 0.0342f
C18045 rowon_n[10] col[3] 0.0323f
C18046 col_n[12] rowoff_n[15] 0.0471f
C18047 row_n[9] col[0] 0.0322f
C18048 rowon_n[11] col[5] 0.0323f
C18049 rowon_n[15] a_16018_17190# 0.248f
C18050 a_31990_4138# a_32482_4500# 0.0658f
C18051 a_31078_4138# a_31382_4178# 0.0931f
C18052 col[15] rowoff_n[11] 0.0901f
C18053 rowoff_n[1] a_12914_3134# 0.202f
C18054 row_n[1] a_26970_3134# 0.0437f
C18055 m2_1732_13998# m2_2160_14426# 0.165f
C18056 rowon_n[5] a_26058_7150# 0.248f
C18057 vcm a_4882_6146# 0.1f
C18058 rowoff_n[12] a_33086_14178# 0.294f
C18059 a_2475_8178# a_17022_8154# 0.316f
C18060 a_8990_8154# a_9994_8154# 0.843f
C18061 m2_10192_13422# a_9994_13174# 0.165f
C18062 col[6] a_8990_16186# 0.367f
C18063 vcm a_26362_16226# 0.155f
C18064 VDD a_24450_6508# 0.0779f
C18065 col[3] a_5886_6146# 0.0682f
C18066 col[13] a_15926_18194# 0.0682f
C18067 ctop a_4974_10162# 4.11f
C18068 a_32994_18194# a_33086_18194# 0.0991f
C18069 VDD a_13918_15182# 0.181f
C18070 rowoff_n[6] a_4370_8516# 0.0133f
C18071 col_n[21] a_24050_12170# 0.251f
C18072 col_n[18] a_20946_2130# 0.0765f
C18073 a_2275_5166# a_7986_5142# 0.399f
C18074 row_n[5] a_3970_7150# 0.282f
C18075 col_n[28] a_30986_14178# 0.0765f
C18076 col_n[2] a_2275_13198# 0.113f
C18077 m2_26832_946# m3_26964_1078# 3.79f
C18078 m3_1864_16138# m3_1864_15134# 0.202f
C18079 m2_29268_9406# a_29070_9158# 0.165f
C18080 col_n[7] a_2275_2154# 0.113f
C18081 vcm a_19942_10162# 0.1f
C18082 a_34090_11166# a_34090_10162# 0.843f
C18083 col_n[1] a_4274_16226# 0.084f
C18084 a_2475_10186# a_32082_10162# 0.316f
C18085 sample a_1957_6170# 0.345f
C18086 rowoff_n[4] a_13406_6508# 0.0133f
C18087 a_27974_15182# a_28370_15222# 0.0313f
C18088 m2_19804_18014# ctop 0.0422f
C18089 VDD a_5374_9520# 0.0779f
C18090 m2_34864_10986# m3_34996_12122# 0.0341f
C18091 ctop a_20034_14178# 4.11f
C18092 col_n[22] a_2475_12194# 0.0531f
C18093 col_n[12] a_15414_10524# 0.0283f
C18094 col_n[27] a_2475_1150# 0.0531f
C18095 m2_1732_15002# row_n[13] 0.292f
C18096 m2_7180_11414# row_n[9] 0.0128f
C18097 m2_13204_7398# row_n[5] 0.0128f
C18098 m2_19228_3382# row_n[1] 0.0128f
C18099 m2_13780_946# col[11] 0.425f
C18100 rowoff_n[9] a_4974_11166# 0.294f
C18101 rowon_n[1] a_1957_3158# 0.0172f
C18102 rowoff_n[2] a_22442_4500# 0.0133f
C18103 a_2275_7174# a_23046_7150# 0.399f
C18104 a_12002_7150# a_12306_7190# 0.0931f
C18105 a_12914_7150# a_13406_7512# 0.0658f
C18106 row_n[6] a_35398_8194# 0.0117f
C18107 vcm a_35002_14178# 0.101f
C18108 a_24050_12170# a_25054_12170# 0.843f
C18109 VDD a_31078_4138# 0.483f
C18110 col_n[0] a_3366_16548# 0.0283f
C18111 col[12] a_2475_9182# 0.136f
C18112 a_2475_16210# a_1957_16210# 0.0734f
C18113 VDD a_20434_13536# 0.0779f
C18114 row_n[8] a_24962_10162# 0.0437f
C18115 rowoff_n[7] a_14010_9158# 0.294f
C18116 rowoff_n[0] a_31478_2492# 0.0133f
C18117 col[2] a_4882_16186# 0.0682f
C18118 rowon_n[12] a_24050_14178# 0.248f
C18119 a_2475_4162# a_15926_4138# 0.264f
C18120 a_2275_4162# a_13310_4178# 0.144f
C18121 a_8898_4138# a_8990_4138# 0.326f
C18122 m3_1864_11118# ctop 0.21f
C18123 col_n[10] a_13006_10162# 0.251f
C18124 m2_20232_7398# a_20034_7150# 0.165f
C18125 m2_28264_16434# row_n[14] 0.0128f
C18126 m2_34864_18014# m2_34864_17010# 0.843f
C18127 m2_34288_12418# row_n[10] 0.0128f
C18128 col_n[19] a_2275_15206# 0.113f
C18129 rowoff_n[13] a_21038_15182# 0.294f
C18130 col_n[24] a_2275_4162# 0.113f
C18131 col_n[17] a_19942_12170# 0.0765f
C18132 rowon_n[2] a_34090_4138# 0.248f
C18133 m2_6752_18014# col[4] 0.347f
C18134 vcm a_15926_17190# 0.1f
C18135 a_15014_14178# a_15014_13174# 0.843f
C18136 VDD a_12002_7150# 0.483f
C18137 rowoff_n[5] a_23046_7150# 0.294f
C18138 a_2275_18218# a_16930_18194# 0.136f
C18139 a_8898_18194# a_9294_18234# 0.0313f
C18140 VDD a_35494_17552# 0.106f
C18141 a_2275_1150# a_6890_1126# 0.136f
C18142 row_n[12] a_2475_14202# 0.405f
C18143 col[9] a_2275_12194# 0.0899f
C18144 vcm a_18026_2130# 0.56f
C18145 a_2275_6170# a_28370_6186# 0.144f
C18146 col_n[1] a_4370_8516# 0.0283f
C18147 col[14] a_2275_1150# 0.0899f
C18148 a_2475_6170# a_30986_6146# 0.264f
C18149 row_n[2] a_12002_4138# 0.282f
C18150 rowoff_n[3] a_32082_5142# 0.294f
C18151 a_28466_1488# col_n[25] 0.0283f
C18152 a_27062_11166# a_27366_11206# 0.0931f
C18153 a_27974_11166# a_28466_11528# 0.0658f
C18154 VDD a_3878_1126# 0.404f
C18155 col[30] a_33086_9158# 0.367f
C18156 rowon_n[6] a_11910_8154# 0.118f
C18157 a_4974_15182# a_5978_15182# 0.843f
C18158 a_2475_15206# a_8990_15182# 0.316f
C18159 col[29] a_2475_11190# 0.136f
C18160 VDD a_27062_11166# 0.483f
C18161 m2_1732_15002# m3_1864_15134# 3.79f
C18162 a_2275_3158# a_21950_3134# 0.136f
C18163 a_2475_18218# a_14922_18194# 0.264f
C18164 m2_11196_5390# a_10998_5142# 0.165f
C18165 row_n[13] a_32386_15222# 0.0117f
C18166 vcm a_33086_6146# 0.56f
C18167 rowoff_n[11] a_27462_13536# 0.0133f
C18168 a_23958_8154# a_24050_8154# 0.326f
C18169 col_n[25] a_28370_9198# 0.084f
C18170 col_n[0] a_2475_8178# 0.0532f
C18171 a_32482_1488# VDD 0.0978f
C18172 col_n[6] a_8898_10162# 0.0765f
C18173 row_n[15] a_22954_17190# 0.0437f
C18174 a_2475_17214# a_24050_17190# 0.316f
C18175 m3_34996_8106# a_34090_8154# 0.0303f
C18176 VDD a_7986_14178# 0.483f
C18177 m2_22816_18014# col_n[20] 0.243f
C18178 row_n[5] a_32994_7150# 0.0437f
C18179 a_18938_5142# a_19334_5182# 0.0313f
C18180 col[26] a_2275_14202# 0.0899f
C18181 col[31] a_2275_3158# 0.0899f
C18182 rowon_n[9] a_32082_11166# 0.248f
C18183 vcm a_14010_9158# 0.56f
C18184 rowoff_n[14] a_8990_16186# 0.294f
C18185 vcm a_2966_18194# 0.165f
C18186 a_7986_14178# a_8290_14218# 0.0931f
C18187 a_8898_14178# a_9390_14540# 0.0658f
C18188 a_2275_14202# a_15014_14178# 0.399f
C18189 m2_34864_7974# m3_34996_9110# 0.0341f
C18190 col[19] a_22042_7150# 0.367f
C18191 VDD a_23046_18194# 0.0356f
C18192 a_15014_2130# a_16018_2130# 0.843f
C18193 col[26] a_28978_9158# 0.0682f
C18194 a_2475_2154# a_29070_2130# 0.316f
C18195 m2_1732_2954# a_1957_3158# 0.245f
C18196 m2_35292_1374# VDD 0.0193f
C18197 vcm a_4274_3174# 0.155f
C18198 row_n[9] a_9994_11166# 0.282f
C18199 rowoff_n[9] a_33998_11166# 0.202f
C18200 rowon_n[13] a_9902_15182# 0.118f
C18201 vcm a_29070_13174# 0.56f
C18202 a_4882_11166# a_4974_11166# 0.326f
C18203 a_2275_11190# a_5278_11206# 0.144f
C18204 a_3878_11166# a_4274_11206# 0.0313f
C18205 a_2475_11190# a_7894_11166# 0.264f
C18206 row_n[5] col[3] 0.0342f
C18207 row_n[11] col[15] 0.0342f
C18208 row_n[9] col[11] 0.0342f
C18209 rowon_n[14] col[22] 0.0323f
C18210 rowon_n[3] col[0] 0.0318f
C18211 col_n[23] rowoff_n[15] 0.0471f
C18212 rowon_n[7] col[8] 0.0323f
C18213 rowon_n[9] col[12] 0.0323f
C18214 row_n[14] col[21] 0.0342f
C18215 VDD a_25966_3134# 0.181f
C18216 rowon_n[0] ctop 0.198f
C18217 row_n[8] col[9] 0.0342f
C18218 rowon_n[4] col[2] 0.0323f
C18219 rowon_n[5] col[4] 0.0323f
C18220 col_n[28] col[28] 0.53f
C18221 row_n[10] col[13] 0.0342f
C18222 rowon_n[15] col[24] 0.0323f
C18223 row_n[12] col[17] 0.0342f
C18224 rowon_n[12] col[18] 0.0323f
C18225 row_n[7] col[7] 0.0342f
C18226 rowon_n[13] col[20] 0.0323f
C18227 row_n[15] col[23] 0.0342f
C18228 row_n[6] col[5] 0.0342f
C18229 rowon_n[6] col[6] 0.0323f
C18230 row_n[4] col[1] 0.0342f
C18231 rowon_n[10] col[14] 0.0323f
C18232 col_n[16] a_2475_10186# 0.0531f
C18233 rowon_n[11] col[16] 0.0323f
C18234 row_n[13] col[19] 0.0342f
C18235 rowon_n[8] col[10] 0.0323f
C18236 m2_13780_18014# a_14314_18234# 0.087f
C18237 col_n[14] a_17326_7190# 0.084f
C18238 a_2275_16210# a_30074_16186# 0.399f
C18239 rowon_n[3] a_19942_5142# 0.118f
C18240 col[26] rowoff_n[11] 0.0901f
C18241 m2_3164_6394# rowon_n[4] 0.0322f
C18242 m2_8184_2378# rowon_n[0] 0.0322f
C18243 a_5978_4138# a_5978_3134# 0.843f
C18244 row_n[1] a_7286_3174# 0.0117f
C18245 col[6] a_2475_7174# 0.136f
C18246 vcm a_19334_7190# 0.155f
C18247 rowoff_n[12] a_15414_14540# 0.0133f
C18248 vcm a_9994_16186# 0.56f
C18249 ctop a_32082_2130# 4.06f
C18250 a_2475_13198# a_22954_13174# 0.264f
C18251 a_2275_13198# a_20338_13214# 0.144f
C18252 VDD a_6890_6146# 0.181f
C18253 a_23958_18194# a_24450_18556# 0.0658f
C18254 a_18026_1126# a_18330_1166# 0.0997f
C18255 col_n[13] a_2275_13198# 0.113f
C18256 a_18938_1126# a_19430_1488# 0.0664f
C18257 row_n[12] a_30986_14178# 0.0437f
C18258 col[8] a_10998_5142# 0.367f
C18259 col_n[18] a_2275_2154# 0.113f
C18260 vcm a_12914_1126# 0.0989f
C18261 col[18] a_21038_17190# 0.367f
C18262 m2_18224_15430# rowon_n[13] 0.0322f
C18263 a_30074_6146# a_31078_6146# 0.843f
C18264 m2_24248_11414# rowon_n[9] 0.0322f
C18265 m2_30272_7398# rowon_n[5] 0.0322f
C18266 col[15] a_17934_7150# 0.0682f
C18267 m2_35292_3382# rowon_n[1] 0.0322f
C18268 m3_2868_18146# m3_3872_18146# 0.202f
C18269 vcm a_35398_11206# 0.161f
C18270 a_2275_10186# a_13918_10162# 0.136f
C18271 m2_1732_16006# a_2161_16210# 0.0454f
C18272 col_n[0] a_3270_13214# 0.084f
C18273 ctop a_13006_5142# 4.11f
C18274 a_19942_15182# a_20034_15182# 0.326f
C18275 a_2275_15206# a_2275_14202# 0.0715f
C18276 VDD a_21950_10162# 0.181f
C18277 col[3] a_2275_10186# 0.0899f
C18278 col_n[30] a_32994_3134# 0.0765f
C18279 col[10] rowoff_n[12] 0.0901f
C18280 m2_1732_11990# m3_1864_12122# 3.79f
C18281 col_n[3] a_6282_5182# 0.084f
C18282 col_n[13] a_16322_17230# 0.084f
C18283 vcm a_27974_5142# 0.1f
C18284 rowoff_n[2] a_4882_4138# 0.202f
C18285 a_2966_7150# a_3270_7190# 0.0931f
C18286 a_21038_8154# a_21038_7150# 0.843f
C18287 rowoff_n[10] a_21950_12170# 0.202f
C18288 a_2475_7174# a_5978_7150# 0.316f
C18289 a_3878_7150# a_4370_7512# 0.0658f
C18290 col[23] a_2475_9182# 0.136f
C18291 row_n[6] a_18026_8154# 0.282f
C18292 vcm a_15318_14218# 0.155f
C18293 a_2275_12194# a_28978_12170# 0.136f
C18294 a_14922_12170# a_15318_12210# 0.0313f
C18295 VDD a_13406_4500# 0.0779f
C18296 rowon_n[10] a_17934_12170# 0.118f
C18297 col_n[24] a_27462_11528# 0.0283f
C18298 m2_34864_17010# VDD 0.773f
C18299 ctop a_28066_9158# 4.11f
C18300 row_n[0] m2_24248_2378# 0.0128f
C18301 VDD a_2161_13198# 0.187f
C18302 row_n[8] a_5278_10202# 0.0117f
C18303 rowoff_n[0] a_13918_2130# 0.202f
C18304 rowon_n[0] a_27974_2130# 0.118f
C18305 col_n[30] a_2275_15206# 0.113f
C18306 a_33086_5142# a_33390_5182# 0.0931f
C18307 a_33998_5142# a_34490_5504# 0.0658f
C18308 m2_25828_18014# m2_26256_18442# 0.165f
C18309 vcm a_8898_8154# 0.1f
C18310 col[7] a_9994_15182# 0.367f
C18311 a_2475_9182# a_21038_9158# 0.316f
C18312 a_10998_9158# a_12002_9158# 0.843f
C18313 rowoff_n[13] a_2966_15182# 0.294f
C18314 col[4] a_6890_5142# 0.0682f
C18315 vcm a_30378_18234# 0.16f
C18316 ctop rowoff_n[13] 0.177f
C18317 col[14] a_16930_17190# 0.0682f
C18318 VDD a_28466_8516# 0.0779f
C18319 m2_34864_4962# m3_34996_6098# 0.0341f
C18320 rowoff_n[5] a_5374_7512# 0.0133f
C18321 ctop a_8990_12170# 4.11f
C18322 col[20] a_2275_12194# 0.0899f
C18323 col_n[22] a_25054_11166# 0.251f
C18324 VDD a_17934_17190# 0.181f
C18325 row_n[0] a_5886_2130# 0.0437f
C18326 col_n[19] a_21950_1126# 0.0765f
C18327 col[25] a_2275_1150# 0.0899f
C18328 a_29982_2130# a_30074_2130# 0.326f
C18329 rowon_n[4] a_4974_6146# 0.248f
C18330 col_n[29] a_31990_13174# 0.0765f
C18331 a_2275_6170# a_12002_6146# 0.399f
C18332 col_n[2] a_5278_15222# 0.084f
C18333 col_n[0] a_2966_5142# 0.251f
C18334 rowoff_n[3] a_14410_5504# 0.0133f
C18335 vcm a_23958_12170# 0.1f
C18336 a_2475_11190# a_2475_10186# 0.0666f
C18337 VDD a_20034_2130# 0.483f
C18338 m2_32856_18014# a_33390_18234# 0.087f
C18339 m2_2160_5390# row_n[3] 0.0194f
C18340 a_29982_16186# a_30378_16226# 0.0313f
C18341 VDD a_9390_11528# 0.0779f
C18342 col_n[13] a_16418_9520# 0.0283f
C18343 ctop a_24050_16186# 4.11f
C18344 a_2275_3158# a_3878_3134# 0.136f
C18345 a_2874_3134# a_3366_3496# 0.0658f
C18346 a_2475_3158# a_4882_3134# 0.264f
C18347 rowoff_n[1] a_23446_3496# 0.0133f
C18348 rowoff_n[8] a_5978_10162# 0.294f
C18349 col_n[10] a_2475_8178# 0.0531f
C18350 row_n[13] a_16018_15182# 0.282f
C18351 a_14010_8154# a_14314_8194# 0.0931f
C18352 a_2275_8178# a_27062_8154# 0.399f
C18353 a_14922_8154# a_15414_8516# 0.0658f
C18354 rowoff_n[11] a_9902_13174# 0.202f
C18355 vcm a_4882_15182# 0.1f
C18356 a_26058_13174# a_27062_13174# 0.843f
C18357 row_n[3] a_26058_5142# 0.282f
C18358 row_n[15] a_3270_17230# 0.0117f
C18359 rowon_n[7] a_25966_9158# 0.118f
C18360 m2_17220_14426# row_n[12] 0.0128f
C18361 a_2275_17214# a_5886_17190# 0.136f
C18362 VDD a_24450_15544# 0.0779f
C18363 col[3] a_5886_15182# 0.0682f
C18364 m2_23244_10410# row_n[8] 0.0128f
C18365 rowoff_n[6] a_15014_8154# 0.294f
C18366 m2_29268_6394# row_n[4] 0.0128f
C18367 col[0] a_2475_5166# 0.148f
C18368 col_n[11] a_14010_9158# 0.251f
C18369 a_2275_5166# a_17326_5182# 0.144f
C18370 row_n[5] a_13310_7190# 0.0117f
C18371 a_10906_5142# a_10998_5142# 0.326f
C18372 a_2475_5166# a_19942_5142# 0.264f
C18373 m2_3164_8402# a_2966_8154# 0.165f
C18374 col_n[18] a_20946_11166# 0.0765f
C18375 rowoff_n[15] a_25966_17190# 0.202f
C18376 m2_25252_16434# a_25054_16186# 0.165f
C18377 rowoff_n[4] a_24050_6146# 0.294f
C18378 col_n[7] a_2275_11190# 0.113f
C18379 m3_3872_1078# a_3970_2130# 0.0176f
C18380 m2_4744_946# a_2475_1150# 0.286f
C18381 a_17022_15182# a_17022_14178# 0.843f
C18382 VDD a_16018_9158# 0.483f
C18383 sample a_1957_15206# 0.345f
C18384 m2_1732_8978# m3_1864_9110# 3.79f
C18385 rowon_n[11] a_2874_13174# 0.118f
C18386 VDD a_5374_18556# 0.0858f
C18387 a_2275_2154# a_10906_2130# 0.136f
C18388 a_5886_2130# a_6282_2170# 0.0313f
C18389 col_n[2] a_5374_7512# 0.0283f
C18390 vcm a_22042_4138# 0.56f
C18391 rowon_n[4] col[13] 0.0323f
C18392 rowon_n[7] col[19] 0.0323f
C18393 rowon_n[9] col[23] 0.0323f
C18394 a_2475_7174# a_35002_7150# 0.264f
C18395 rowon_n[13] col[31] 0.0323f
C18396 a_2275_7174# a_32386_7190# 0.144f
C18397 row_n[12] col[28] 0.0342f
C18398 row_n[7] col[18] 0.0342f
C18399 rowon_n[11] col[27] 0.0323f
C18400 rowoff_n[2] a_33086_4138# 0.294f
C18401 rowon_n[6] col[17] 0.0323f
C18402 row_n[5] col[14] 0.0342f
C18403 row_n[14] sample_n 0.0596f
C18404 rowon_n[10] col[25] 0.0323f
C18405 rowon_n[8] col[21] 0.0323f
C18406 rowon_n[5] col[15] 0.0323f
C18407 row_n[10] col[24] 0.0342f
C18408 row_n[13] col[30] 0.0342f
C18409 rowon_n[3] col[11] 0.0323f
C18410 row_n[2] col[8] 0.0342f
C18411 col_n[27] a_2475_10186# 0.0531f
C18412 row_n[11] col[26] 0.0342f
C18413 rowon_n[2] col[9] 0.0323f
C18414 row_n[0] col[4] 0.0342f
C18415 row_n[9] col[22] 0.0342f
C18416 row_n[4] col[12] 0.0342f
C18417 row_n[8] col[20] 0.0342f
C18418 rowon_n[1] col[7] 0.0323f
C18419 rowon_n[0] col[5] 0.0323f
C18420 rowon_n[12] col[29] 0.0323f
C18421 row_n[6] col[16] 0.0342f
C18422 row_n[1] col[6] 0.0342f
C18423 ctop col[1] 0.125f
C18424 rowon_n[1] a_13006_3134# 0.248f
C18425 row_n[3] col[10] 0.0342f
C18426 col[31] a_34090_8154# 0.367f
C18427 a_29070_12170# a_29374_12210# 0.0931f
C18428 a_29982_12170# a_30474_12532# 0.0658f
C18429 a_2475_16210# a_13006_16186# 0.316f
C18430 a_6982_16186# a_7986_16186# 0.843f
C18431 VDD a_31078_13174# 0.483f
C18432 col[17] a_2475_7174# 0.136f
C18433 a_2275_4162# a_25966_4138# 0.136f
C18434 m3_23952_1078# ctop 0.21f
C18435 col_n[26] a_29374_8194# 0.084f
C18436 vcm a_2874_7150# 0.1f
C18437 a_25966_9158# a_26058_9158# 0.326f
C18438 m2_16216_14426# a_16018_14178# 0.165f
C18439 row_n[10] a_24050_12170# 0.282f
C18440 col_n[7] a_9902_9158# 0.0765f
C18441 a_2275_13198# a_3970_13174# 0.399f
C18442 rowon_n[14] a_23958_16186# 0.118f
C18443 col_n[24] a_2275_13198# 0.113f
C18444 col_n[29] a_2275_2154# 0.113f
C18445 row_n[0] a_34090_2130# 0.282f
C18446 VDD a_12002_16186# 0.483f
C18447 a_2475_1150# a_18026_1126# 0.31f
C18448 row_n[12] a_11302_14218# 0.0117f
C18449 rowon_n[4] a_33998_6146# 0.118f
C18450 m2_23820_946# col[21] 0.425f
C18451 m2_13204_2378# a_13006_2130# 0.165f
C18452 vcm a_27366_2170# 0.155f
C18453 a_20946_6146# a_21342_6186# 0.0313f
C18454 m2_34864_9982# a_35094_10162# 0.0249f
C18455 row_n[2] a_21342_4178# 0.0117f
C18456 vcm a_18026_11166# 0.56f
C18457 col[14] a_2275_10186# 0.0899f
C18458 col_n[1] a_4370_17552# 0.0283f
C18459 col[21] rowoff_n[12] 0.0901f
C18460 VDD a_14922_1126# 0.405f
C18461 col[20] a_23046_6146# 0.367f
C18462 a_9994_15182# a_10298_15222# 0.0931f
C18463 a_10906_15182# a_11398_15544# 0.0658f
C18464 a_2275_15206# a_19030_15182# 0.399f
C18465 VDD a_3878_10162# 0.181f
C18466 col[27] a_29982_8154# 0.0682f
C18467 row_n[4] a_11910_6146# 0.0437f
C18468 a_17022_3134# a_18026_3134# 0.843f
C18469 a_2475_3158# a_33086_3134# 0.316f
C18470 rowon_n[8] a_10998_10162# 0.248f
C18471 rowoff_n[8] a_35002_10162# 0.202f
C18472 vcm a_8290_5182# 0.155f
C18473 rowoff_n[10] a_3878_12170# 0.202f
C18474 m2_7180_12418# a_6982_12170# 0.165f
C18475 vcm a_33086_15182# 0.56f
C18476 col_n[15] a_18330_6186# 0.084f
C18477 a_6890_12170# a_6982_12170# 0.326f
C18478 a_2475_12194# a_11910_12170# 0.264f
C18479 a_2275_12194# a_9294_12210# 0.144f
C18480 VDD a_29982_5142# 0.181f
C18481 col_n[25] a_28370_18234# 0.084f
C18482 col_n[0] a_2475_17214# 0.0532f
C18483 m2_17220_18442# VDD 0.0456f
C18484 a_2275_17214# a_34090_17190# 0.399f
C18485 col_n[4] a_2475_6170# 0.0531f
C18486 a_7986_5142# a_7986_4138# 0.843f
C18487 m2_26256_8402# a_26058_8154# 0.165f
C18488 col[5] rowoff_n[13] 0.0901f
C18489 m2_7756_18014# m2_8760_18014# 0.843f
C18490 vcm a_23350_9198# 0.155f
C18491 a_2475_9182# a_2966_9158# 0.317f
C18492 a_2161_9182# a_2275_9182# 0.183f
C18493 col[31] a_2275_12194# 0.0899f
C18494 ctop a_2475_3158# 0.0487f
C18495 vcm a_14010_18194# 0.165f
C18496 m2_1732_17010# rowon_n[15] 0.236f
C18497 a_2275_14202# a_24354_14218# 0.144f
C18498 a_2475_14202# a_26970_14178# 0.264f
C18499 m2_7180_13422# rowon_n[11] 0.0322f
C18500 VDD a_10906_8154# 0.181f
C18501 row_n[7] a_32082_9158# 0.282f
C18502 m2_1732_5966# m3_1864_6098# 3.79f
C18503 m2_13204_9406# rowon_n[7] 0.0322f
C18504 m2_19228_5390# rowon_n[3] 0.0322f
C18505 rowon_n[11] a_31990_13174# 0.118f
C18506 col[9] a_12002_4138# 0.367f
C18507 VDD a_32386_18234# 0.019f
C18508 a_20034_2130# a_20338_2170# 0.0931f
C18509 a_20946_2130# a_21438_2492# 0.0658f
C18510 col[19] a_22042_16186# 0.367f
C18511 col[16] a_18938_6146# 0.0682f
C18512 row_n[9] a_19334_11206# 0.0117f
C18513 vcm a_16930_3134# 0.1f
C18514 a_32082_7150# a_33086_7150# 0.843f
C18515 col_n[1] a_2275_9182# 0.113f
C18516 col[26] a_28978_18194# 0.0682f
C18517 vcm a_4274_12210# 0.155f
C18518 a_2275_11190# a_17934_11166# 0.136f
C18519 VDD a_1957_2154# 0.196f
C18520 col_n[31] a_33998_2130# 0.0765f
C18521 ctop a_17022_7150# 4.11f
C18522 row_n[11] a_9902_13174# 0.0437f
C18523 a_21950_16186# a_22042_16186# 0.326f
C18524 col_n[4] a_7286_4178# 0.084f
C18525 VDD a_25966_12170# 0.181f
C18526 m2_13780_18014# m3_13912_18146# 3.79f
C18527 rowon_n[15] a_8990_17190# 0.248f
C18528 col_n[14] a_17326_16226# 0.084f
C18529 m2_34288_14426# rowon_n[12] 0.0322f
C18530 col_n[21] a_2475_8178# 0.0531f
C18531 row_n[1] a_19942_3134# 0.0437f
C18532 rowoff_n[1] a_5886_3134# 0.202f
C18533 m2_17220_6394# a_17022_6146# 0.165f
C18534 vcm a_31990_7150# 0.1f
C18535 rowon_n[5] a_19030_7150# 0.248f
C18536 a_23046_9158# a_23046_8154# 0.843f
C18537 rowoff_n[12] a_26058_14178# 0.294f
C18538 a_2475_8178# a_9994_8154# 0.316f
C18539 col_n[25] a_28466_10524# 0.0283f
C18540 vcm a_19334_16226# 0.155f
C18541 col[6] a_2475_16210# 0.136f
C18542 a_16930_13174# a_17326_13214# 0.0313f
C18543 a_2275_13198# a_32994_13174# 0.136f
C18544 VDD a_17422_6508# 0.0779f
C18545 col[11] a_2475_5166# 0.136f
C18546 ctop a_32082_11166# 4.11f
C18547 VDD a_6890_15182# 0.181f
C18548 m2_1732_3958# m2_1732_2954# 0.843f
C18549 col[8] a_10998_14178# 0.367f
C18550 m2_16792_946# m3_15920_1078# 0.0341f
C18551 col[5] a_7894_4138# 0.0682f
C18552 col_n[18] a_2275_11190# 0.113f
C18553 vcm a_12914_10162# 0.1f
C18554 a_2475_10186# a_25054_10162# 0.316f
C18555 a_13006_10162# a_14010_10162# 0.843f
C18556 row_n[14] a_30074_16186# 0.282f
C18557 col[15] a_17934_16186# 0.0682f
C18558 rowoff_n[4] a_6378_6508# 0.0133f
C18559 col_n[23] a_26058_10162# 0.251f
C18560 m2_5748_18014# ctop 0.0422f
C18561 VDD a_32482_10524# 0.0779f
C18562 ctop a_13006_14178# 4.11f
C18563 col_n[30] a_32994_12170# 0.0765f
C18564 rowon_n[2] col[20] 0.0323f
C18565 row_n[6] col[27] 0.0342f
C18566 rowon_n[3] col[22] 0.0323f
C18567 rowon_n[4] col[24] 0.0323f
C18568 rowon_n[8] sample_n 0.0692f
C18569 row_n[7] col[29] 0.0342f
C18570 rowon_n[1] col[18] 0.0323f
C18571 row_n[2] col[19] 0.0342f
C18572 row_n[1] col[17] 0.0342f
C18573 row_n[3] col[21] 0.0342f
C18574 row_n[4] col[23] 0.0342f
C18575 row_n[5] col[25] 0.0342f
C18576 rowon_n[6] col[28] 0.0323f
C18577 rowon_n[7] col[30] 0.0323f
C18578 row_n[0] col[15] 0.0342f
C18579 ctop col[12] 0.123f
C18580 rowon_n[0] col[16] 0.0323f
C18581 rowon_n[5] col[26] 0.0323f
C18582 row_n[8] col[31] 0.0342f
C18583 a_31990_3134# a_32082_3134# 0.326f
C18584 col[8] a_2275_8178# 0.0899f
C18585 col_n[3] a_6282_14218# 0.084f
C18586 m2_8184_4386# a_7986_4138# 0.165f
C18587 rowoff_n[10] a_32482_12532# 0.0133f
C18588 rowoff_n[2] a_15414_4500# 0.0133f
C18589 a_2275_7174# a_16018_7150# 0.399f
C18590 m2_34864_18014# vcm 0.408f
C18591 row_n[6] a_27366_8194# 0.0117f
C18592 vcm a_27974_14178# 0.1f
C18593 a_3970_12170# a_3970_11166# 0.843f
C18594 VDD a_24050_4138# 0.483f
C18595 col_n[14] a_17422_8516# 0.0283f
C18596 col[28] a_2475_7174# 0.136f
C18597 a_31990_17190# a_32386_17230# 0.0313f
C18598 VDD a_13406_13536# 0.0779f
C18599 row_n[8] a_17934_10162# 0.0437f
C18600 rowoff_n[0] a_24450_2492# 0.0133f
C18601 rowoff_n[7] a_6982_9158# 0.294f
C18602 rowon_n[12] a_17022_14178# 0.248f
C18603 a_2475_4162# a_8898_4138# 0.264f
C18604 a_2275_4162# a_6282_4178# 0.144f
C18605 m3_19936_18146# ctop 0.209f
C18606 m2_6176_12418# row_n[10] 0.0128f
C18607 a_2275_9182# a_31078_9158# 0.399f
C18608 a_16930_9158# a_17422_9520# 0.0658f
C18609 rowoff_n[13] a_14010_15182# 0.294f
C18610 m2_12200_8402# row_n[6] 0.0128f
C18611 a_16018_9158# a_16322_9198# 0.0931f
C18612 m2_18224_4386# row_n[2] 0.0128f
C18613 m2_1732_13998# a_2475_14202# 0.139f
C18614 rowon_n[2] a_27062_4138# 0.248f
C18615 vcm a_8898_17190# 0.1f
C18616 a_28066_14178# a_29070_14178# 0.843f
C18617 VDD a_4974_7150# 0.483f
C18618 m2_1732_2954# m3_1864_3086# 3.79f
C18619 col[4] a_6890_14178# 0.0682f
C18620 rowoff_n[5] a_16018_7150# 0.294f
C18621 a_2275_18218# a_9902_18194# 0.136f
C18622 VDD a_28466_17552# 0.0779f
C18623 col_n[12] a_15014_8154# 0.251f
C18624 a_35002_2130# a_35398_2170# 0.0313f
C18625 vcm a_10998_2130# 0.56f
C18626 col[25] a_2275_10186# 0.0899f
C18627 col_n[19] a_21950_10162# 0.0765f
C18628 sample_n rowoff_n[12] 0.14f
C18629 a_2475_6170# a_23958_6146# 0.264f
C18630 a_12914_6146# a_13006_6146# 0.326f
C18631 a_2275_6170# a_21342_6186# 0.144f
C18632 sample m2_1732_946# 0.2f
C18633 rowoff_n[3] a_25054_5142# 0.294f
C18634 row_n[2] a_4974_4138# 0.282f
C18635 m2_27260_17438# row_n[15] 0.0128f
C18636 m2_33284_13422# row_n[11] 0.0128f
C18637 rowon_n[6] a_4882_8154# 0.118f
C18638 col_n[0] a_2966_14178# 0.251f
C18639 a_19030_16186# a_19030_15182# 0.843f
C18640 VDD a_20034_11166# 0.483f
C18641 col_n[3] a_6378_6508# 0.0283f
C18642 a_2275_3158# a_14922_3134# 0.136f
C18643 a_7894_3134# a_8290_3174# 0.0313f
C18644 col_n[13] a_16418_18556# 0.0283f
C18645 a_2475_18218# a_7894_18194# 0.264f
C18646 rowoff_n[1] a_34090_3134# 0.294f
C18647 a_28066_1126# a_2275_1150# 0.0924f
C18648 row_n[13] a_25358_15222# 0.0117f
C18649 vcm a_26058_6146# 0.56f
C18650 a_2966_8154# a_2966_7150# 0.843f
C18651 rowoff_n[11] a_20434_13536# 0.0133f
C18652 col_n[10] a_2475_17214# 0.0531f
C18653 m2_1732_8978# sample 0.2f
C18654 col_n[15] a_2475_6170# 0.0531f
C18655 a_31078_13174# a_31382_13214# 0.0931f
C18656 a_31990_13174# a_32482_13536# 0.0658f
C18657 m2_34864_2954# ctop 0.0422f
C18658 a_25454_1488# VDD 0.0977f
C18659 row_n[15] a_15926_17190# 0.0437f
C18660 a_2475_17214# a_17022_17190# 0.316f
C18661 a_8990_17190# a_9994_17190# 0.843f
C18662 col[16] rowoff_n[13] 0.0901f
C18663 m3_23952_18146# a_24050_17190# 0.0303f
C18664 a_2275_5166# a_29982_5142# 0.136f
C18665 col_n[1] a_3970_6146# 0.251f
C18666 row_n[5] a_25966_7150# 0.0437f
C18667 col_n[27] a_30378_7190# 0.084f
C18668 col[0] a_2475_14202# 0.148f
C18669 col[5] a_2475_3158# 0.136f
C18670 sample rowoff_n[8] 0.0775f
C18671 rowon_n[9] a_25054_11166# 0.248f
C18672 VDD rowoff_n[7] 1.51f
C18673 col_n[0] rowoff_n[9] 0.0471f
C18674 a_28978_1126# a_29374_1166# 0.0313f
C18675 vcm a_6982_9158# 0.56f
C18676 col_n[8] a_10906_8154# 0.0765f
C18677 rowoff_n[14] a_2475_16210# 3.9f
C18678 a_27974_10162# a_28066_10162# 0.326f
C18679 m2_27836_946# a_2475_1150# 0.286f
C18680 m2_8760_946# a_9294_1166# 0.087f
C18681 a_2275_14202# a_7986_14178# 0.399f
C18682 VDD a_16018_18194# 0.0356f
C18683 col_n[12] a_2275_9182# 0.113f
C18684 a_29070_3134# a_29070_2130# 0.843f
C18685 a_2475_2154# a_22042_2130# 0.316f
C18686 m2_20808_946# VDD 0.999f
C18687 row_n[9] a_2874_11166# 0.0436f
C18688 vcm a_31382_4178# 0.155f
C18689 rowoff_n[9] a_26970_11166# 0.202f
C18690 a_22954_7150# a_23350_7190# 0.0313f
C18691 col_n[2] a_5374_16548# 0.0283f
C18692 rowon_n[13] a_2161_15206# 0.0177f
C18693 vcm a_22042_13174# 0.56f
C18694 col[21] a_24050_5142# 0.367f
C18695 VDD a_18938_3134# 0.181f
C18696 m2_25828_18014# a_2275_18218# 0.28f
C18697 col[31] a_34090_17190# 0.367f
C18698 a_12002_16186# a_12306_16226# 0.0931f
C18699 a_2275_16210# a_23046_16186# 0.399f
C18700 col[28] a_30986_7150# 0.0682f
C18701 col[2] a_2275_6170# 0.0899f
C18702 a_12914_16186# a_13406_16548# 0.0658f
C18703 rowon_n[3] a_12914_5142# 0.118f
C18704 a_29982_1126# m2_29844_946# 0.225f
C18705 col[0] rowoff_n[14] 0.0901f
C18706 a_19030_4138# a_20034_4138# 0.843f
C18707 m2_1732_5966# a_2966_6146# 0.843f
C18708 col[17] a_2475_16210# 0.136f
C18709 vcm a_12306_7190# 0.155f
C18710 rowoff_n[12] a_8386_14540# 0.0133f
C18711 col[22] a_2475_5166# 0.136f
C18712 col_n[16] a_19334_5182# 0.084f
C18713 row_n[10] a_33390_12210# 0.0117f
C18714 ctop a_25054_2130# 4.06f
C18715 vcm a_2874_16186# 0.1f
C18716 col_n[26] a_29374_17230# 0.084f
C18717 a_8898_13174# a_8990_13174# 0.326f
C18718 a_2475_13198# a_15926_13174# 0.264f
C18719 a_2275_13198# a_13310_13214# 0.144f
C18720 VDD a_33998_7150# 0.181f
C18721 col_n[7] a_9902_18194# 0.0762f
C18722 m2_21812_18014# a_2475_18218# 0.286f
C18723 row_n[12] a_23958_14178# 0.0437f
C18724 col_n[29] a_2275_11190# 0.113f
C18725 vcm a_5886_1126# 0.0989f
C18726 a_9994_6146# a_9994_5142# 0.843f
C18727 m2_2160_7398# rowon_n[5] 0.0219f
C18728 m2_8184_3382# rowon_n[1] 0.0322f
C18729 m2_34864_8978# a_2275_9182# 0.278f
C18730 row_n[2] a_33998_4138# 0.0437f
C18731 vcm a_27366_11206# 0.155f
C18732 a_2275_10186# a_6890_10162# 0.136f
C18733 m2_31276_17438# a_31078_17190# 0.165f
C18734 rowon_n[6] a_33086_8154# 0.248f
C18735 ctop a_5978_5142# 4.11f
C18736 VDD vcm 24.5f
C18737 a_2275_15206# a_28370_15222# 0.144f
C18738 a_2475_15206# a_30986_15182# 0.264f
C18739 row_n[0] col[26] 0.0342f
C18740 row_n[3] sample_n 0.0596f
C18741 col[10] a_13006_3134# 0.367f
C18742 rowon_n[1] col[29] 0.0323f
C18743 rowon_n[2] col[31] 0.0323f
C18744 ctop col[23] 0.123f
C18745 row_n[1] col[28] 0.0342f
C18746 row_n[2] col[30] 0.0342f
C18747 VDD a_14922_10162# 0.181f
C18748 col[8] col[9] 0.0355f
C18749 rowon_n[0] col[27] 0.0323f
C18750 col[19] a_2275_8178# 0.0899f
C18751 col[20] a_23046_15182# 0.367f
C18752 col[17] a_19942_5142# 0.0682f
C18753 a_22954_3134# a_23446_3496# 0.0658f
C18754 a_2475_18218# a_2475_17214# 0.0666f
C18755 a_22042_3134# a_22346_3174# 0.0931f
C18756 col[27] a_29982_17190# 0.0682f
C18757 vcm a_20946_5142# 0.1f
C18758 rowoff_n[10] a_14922_12170# 0.202f
C18759 a_33998_8154# a_34394_8194# 0.0313f
C18760 a_35094_1126# vcm 0.165f
C18761 m2_17220_16434# rowon_n[14] 0.0322f
C18762 m2_23244_12418# rowon_n[10] 0.0322f
C18763 row_n[6] a_10998_8154# 0.282f
C18764 m2_29268_8402# rowon_n[6] 0.0322f
C18765 vcm a_8290_14218# 0.155f
C18766 m2_34864_3958# rowon_n[2] 0.231f
C18767 a_2275_12194# a_21950_12170# 0.136f
C18768 rowon_n[10] a_10906_12170# 0.118f
C18769 VDD a_6378_4500# 0.0779f
C18770 col_n[5] a_8290_3174# 0.084f
C18771 ctop a_21038_9158# 4.11f
C18772 col_n[15] a_18330_15222# 0.084f
C18773 a_23958_17190# a_24050_17190# 0.326f
C18774 VDD a_29982_14178# 0.181f
C18775 rowon_n[0] a_20946_2130# 0.118f
C18776 rowoff_n[0] a_6890_2130# 0.202f
C18777 col_n[4] a_2475_15206# 0.0531f
C18778 col_n[9] a_2475_4162# 0.0531f
C18779 m2_7756_946# ctop 0.0428f
C18780 m2_34864_7974# a_35002_8154# 0.225f
C18781 vcm a_34394_9198# 0.155f
C18782 col_n[26] a_29470_9520# 0.0283f
C18783 m2_18800_18014# m2_19228_18442# 0.165f
C18784 a_25054_10162# a_25054_9158# 0.843f
C18785 rowoff_n[14] a_30986_16186# 0.202f
C18786 a_2475_9182# a_14010_9158# 0.316f
C18787 m2_22240_15430# a_22042_15182# 0.165f
C18788 vcm a_23350_18234# 0.16f
C18789 a_18938_14178# a_19334_14218# 0.0313f
C18790 VDD a_21438_8516# 0.0779f
C18791 ctop a_2475_12194# 0.0488f
C18792 VDD a_10906_17190# 0.181f
C18793 analog_in a_2475_1150# 0.0422f
C18794 col[9] a_12002_13174# 0.367f
C18795 row_n[9] a_31990_11166# 0.0437f
C18796 col[6] a_8898_3134# 0.0682f
C18797 a_3878_6146# a_3970_6146# 0.326f
C18798 a_2275_6170# a_4974_6146# 0.399f
C18799 a_2874_6146# a_3270_6186# 0.0313f
C18800 rowon_n[13] a_31078_15182# 0.248f
C18801 col[16] a_18938_15182# 0.0682f
C18802 rowoff_n[3] a_7382_5504# 0.0133f
C18803 vcm a_16930_12170# 0.1f
C18804 a_15014_11166# a_16018_11166# 0.843f
C18805 a_2475_11190# a_29070_11166# 0.316f
C18806 col_n[1] a_2275_18218# 0.113f
C18807 VDD a_13006_2130# 0.483f
C18808 col_n[24] a_27062_9158# 0.251f
C18809 col_n[6] a_2275_7174# 0.113f
C18810 VDD a_1957_11190# 0.196f
C18811 m2_27836_18014# m3_28972_18146# 0.0341f
C18812 col_n[31] a_33998_11166# 0.0765f
C18813 ctop a_17022_16186# 4.11f
C18814 col_n[4] a_7286_13214# 0.084f
C18815 a_33998_4138# a_34090_4138# 0.326f
C18816 col[0] a_2966_11166# 0.367f
C18817 rowoff_n[1] a_16418_3496# 0.0133f
C18818 col_n[21] a_2475_17214# 0.0531f
C18819 row_n[13] a_8990_15182# 0.282f
C18820 col_n[26] a_2475_6170# 0.0531f
C18821 rowoff_n[11] a_2161_13198# 0.0226f
C18822 a_2275_8178# a_20034_8154# 0.399f
C18823 m2_13204_13422# a_13006_13174# 0.165f
C18824 vcm a_31990_16186# 0.1f
C18825 col_n[15] a_18426_7512# 0.0283f
C18826 a_5978_13174# a_5978_12170# 0.843f
C18827 VDD a_28066_6146# 0.483f
C18828 row_n[3] a_19030_5142# 0.282f
C18829 col[27] rowoff_n[13] 0.0901f
C18830 rowon_n[7] a_18938_9158# 0.118f
C18831 VDD a_17422_15544# 0.0779f
C18832 rowoff_n[6] a_7986_8154# 0.294f
C18833 m2_1732_5966# row_n[4] 0.292f
C18834 col[11] a_2475_14202# 0.136f
C18835 m2_6176_2378# row_n[0] 0.0128f
C18836 col[16] a_2475_3158# 0.136f
C18837 col_n[5] rowoff_n[4] 0.0471f
C18838 col_n[1] rowoff_n[0] 0.0471f
C18839 col_n[7] rowoff_n[6] 0.0471f
C18840 col_n[2] rowoff_n[1] 0.0471f
C18841 col_n[9] rowoff_n[8] 0.0471f
C18842 m3_1864_17142# a_2966_17190# 0.0302f
C18843 col_n[6] rowoff_n[5] 0.0471f
C18844 col_n[8] rowoff_n[7] 0.0471f
C18845 col_n[10] rowoff_n[9] 0.0471f
C18846 col_n[3] rowoff_n[2] 0.0471f
C18847 col_n[4] rowoff_n[3] 0.0471f
C18848 row_n[5] a_6282_7190# 0.0117f
C18849 a_2475_5166# a_12914_5142# 0.264f
C18850 a_2275_5166# a_10298_5182# 0.144f
C18851 m2_31852_946# m3_31984_1078# 3.79f
C18852 m2_32280_9406# a_32082_9158# 0.165f
C18853 col_n[0] a_2874_3134# 0.0765f
C18854 a_2275_10186# a_35094_10162# 0.0924f
C18855 a_18938_10162# a_19430_10524# 0.0658f
C18856 a_18026_10162# a_18330_10202# 0.0931f
C18857 rowoff_n[15] a_18938_17190# 0.202f
C18858 col[5] a_7894_13174# 0.0682f
C18859 rowoff_n[4] a_17022_6146# 0.294f
C18860 a_30074_15182# a_31078_15182# 0.843f
C18861 VDD a_8990_9158# 0.483f
C18862 col_n[23] a_2275_9182# 0.113f
C18863 col_n[13] a_16018_7150# 0.251f
C18864 col_n[20] a_22954_9158# 0.0765f
C18865 m2_16216_15430# row_n[13] 0.0128f
C18866 a_2874_2130# a_2966_2130# 0.0991f
C18867 m2_22240_11414# row_n[9] 0.0128f
C18868 m2_28264_7398# row_n[5] 0.0128f
C18869 m2_34288_3382# row_n[1] 0.0128f
C18870 vcm a_15014_4138# 0.56f
C18871 a_2275_7174# a_25358_7190# 0.144f
C18872 a_2475_7174# a_27974_7150# 0.264f
C18873 rowoff_n[2] a_26058_4138# 0.294f
C18874 rowon_n[1] a_5978_3134# 0.248f
C18875 a_14922_7150# a_15014_7150# 0.326f
C18876 col[8] a_2275_17214# 0.0899f
C18877 m2_4168_11414# a_3970_11166# 0.165f
C18878 col[13] a_2275_6170# 0.0899f
C18879 col[11] rowoff_n[14] 0.0901f
C18880 a_21038_17190# a_21038_16186# 0.843f
C18881 a_2966_16186# a_3270_16226# 0.0931f
C18882 a_2475_16210# a_5978_16186# 0.316f
C18883 a_3878_16186# a_4370_16548# 0.0658f
C18884 col_n[4] a_7382_5504# 0.0283f
C18885 VDD a_24050_13174# 0.483f
C18886 col_n[14] a_17422_17552# 0.0283f
C18887 rowoff_n[0] a_35094_2130# 0.0135f
C18888 col[28] a_2475_16210# 0.136f
C18889 a_2275_4162# a_18938_4138# 0.136f
C18890 a_9902_4138# a_10298_4178# 0.0313f
C18891 m3_34996_4090# ctop 0.209f
C18892 m2_23244_7398# a_23046_7150# 0.165f
C18893 vcm a_30074_8154# 0.56f
C18894 row_n[10] a_17022_12170# 0.282f
C18895 rowon_n[14] a_16930_16186# 0.118f
C18896 a_33998_14178# a_34490_14540# 0.0658f
C18897 a_33086_14178# a_33390_14218# 0.0931f
C18898 col_n[3] a_2475_2154# 0.0531f
C18899 VDD a_4974_16186# 0.483f
C18900 row_n[0] a_27062_2130# 0.282f
C18901 row_n[12] a_4274_14218# 0.0117f
C18902 a_2475_1150# a_10998_1126# 0.0299f
C18903 col_n[28] a_31382_6186# 0.084f
C18904 rowon_n[4] a_26970_6146# 0.118f
C18905 col_n[2] a_4974_5142# 0.251f
C18906 vcm a_20338_2170# 0.155f
C18907 col_n[12] a_15014_17190# 0.251f
C18908 a_2275_6170# a_33998_6146# 0.136f
C18909 col_n[9] a_11910_7150# 0.0765f
C18910 m2_9764_946# m2_10768_946# 0.843f
C18911 row_n[2] a_14314_4178# 0.0117f
C18912 VDD col_n[11] 5.17f
C18913 vcm a_10998_11166# 0.56f
C18914 vcm col_n[8] 1.94f
C18915 a_29982_11166# a_30074_11166# 0.326f
C18916 VDD a_7894_1126# 0.405f
C18917 col[30] a_2275_8178# 0.0899f
C18918 a_2275_15206# a_12002_15182# 0.399f
C18919 row_n[4] a_4882_6146# 0.0437f
C18920 a_31078_4138# a_31078_3134# 0.843f
C18921 rowon_n[8] a_3970_10162# 0.248f
C18922 a_2475_3158# a_26058_3134# 0.316f
C18923 rowoff_n[8] a_27974_10162# 0.202f
C18924 col_n[3] a_6378_15544# 0.0283f
C18925 m2_14208_5390# a_14010_5142# 0.165f
C18926 vcm a_2275_5166# 6.49f
C18927 rowoff_n[11] a_31078_13174# 0.294f
C18928 a_24962_8154# a_25358_8194# 0.0313f
C18929 col[22] a_25054_4138# 0.367f
C18930 vcm a_26058_15182# 0.56f
C18931 a_2874_12170# a_3366_12532# 0.0658f
C18932 a_2475_12194# a_4882_12170# 0.264f
C18933 a_2275_12194# a_3878_12170# 0.136f
C18934 VDD a_22954_5142# 0.181f
C18935 col[29] a_31990_6146# 0.0682f
C18936 m2_3164_18442# VDD 0.0456f
C18937 ctop a_2966_9158# 4.06f
C18938 col_n[15] a_2475_15206# 0.0531f
C18939 a_14010_17190# a_14314_17230# 0.0931f
C18940 a_2275_17214# a_27062_17190# 0.399f
C18941 a_14922_17190# a_15414_17552# 0.0658f
C18942 m2_7756_946# col[5] 0.425f
C18943 col_n[20] a_2475_4162# 0.0531f
C18944 rowon_n[0] a_2275_2154# 1.79f
C18945 a_21038_5142# a_22042_5142# 0.843f
C18946 col_n[17] a_20338_4178# 0.084f
C18947 vcm a_16322_9198# 0.155f
C18948 col_n[27] a_30378_16226# 0.084f
C18949 col_n[1] a_3970_15182# 0.251f
C18950 col[5] a_2475_12194# 0.136f
C18951 ctop a_29070_4138# 4.11f
C18952 vcm a_6982_18194# 0.165f
C18953 a_2275_14202# a_17326_14218# 0.144f
C18954 col_n[8] a_10906_17190# 0.0765f
C18955 a_10906_14178# a_10998_14178# 0.326f
C18956 a_2475_14202# a_19942_14178# 0.264f
C18957 row_n[7] a_25054_9158# 0.282f
C18958 VDD a_3366_8516# 0.0779f
C18959 col[10] a_2475_1150# 0.136f
C18960 rowon_n[11] a_24962_13174# 0.118f
C18961 VDD a_25358_18234# 0.019f
C18962 a_2275_2154# a_32082_2130# 0.399f
C18963 m2_5172_3382# a_4974_3134# 0.165f
C18964 m3_14916_18146# VDD 0.0873f
C18965 m2_34864_8978# m2_35292_9406# 0.165f
C18966 row_n[9] a_12306_11206# 0.0117f
C18967 col_n[12] a_2275_18218# 0.113f
C18968 vcm a_9902_3134# 0.1f
C18969 a_12002_7150# a_12002_6146# 0.843f
C18970 rowon_n[1] a_35002_3134# 0.118f
C18971 col_n[17] a_2275_7174# 0.113f
C18972 vcm a_31382_13214# 0.155f
C18973 a_2275_11190# a_10906_11166# 0.136f
C18974 a_5886_11166# a_6282_11206# 0.0313f
C18975 VDD a_29470_3496# 0.0779f
C18976 col[11] a_14010_2130# 0.367f
C18977 m2_17796_18014# a_17934_18194# 0.225f
C18978 ctop a_9994_7150# 4.11f
C18979 row_n[11] a_2161_13198# 0.0221f
C18980 a_2275_16210# a_32386_16226# 0.144f
C18981 a_2475_16210# a_35002_16186# 0.264f
C18982 col[21] a_24050_14178# 0.367f
C18983 VDD a_18938_12170# 0.181f
C18984 col[18] a_20946_4138# 0.0682f
C18985 m2_4744_18014# m3_3872_18146# 0.0341f
C18986 rowon_n[15] a_2475_17214# 0.31f
C18987 m2_6176_14426# rowon_n[12] 0.0322f
C18988 col[28] a_30986_16186# 0.0682f
C18989 m2_12200_10410# rowon_n[8] 0.0322f
C18990 col[2] a_2275_15206# 0.0899f
C18991 m2_18224_6394# rowon_n[4] 0.0322f
C18992 a_24962_4138# a_25454_4500# 0.0658f
C18993 a_24050_4138# a_24354_4178# 0.0931f
C18994 col[7] a_2275_4162# 0.0899f
C18995 row_n[1] a_12914_3134# 0.0437f
C18996 vcm a_24962_7150# 0.1f
C18997 rowon_n[5] a_12002_7150# 0.248f
C18998 rowoff_n[12] a_19030_14178# 0.294f
C18999 m2_2736_1950# col_n[0] 0.251f
C19000 a_1957_8178# a_2275_8178# 0.158f
C19001 a_2475_8178# a_2874_8154# 0.264f
C19002 col_n[6] a_9294_2170# 0.084f
C19003 vcm a_12306_16226# 0.155f
C19004 a_2275_13198# a_25966_13174# 0.136f
C19005 col_n[16] a_19334_14218# 0.084f
C19006 col[22] a_2475_14202# 0.136f
C19007 VDD a_10394_6508# 0.0779f
C19008 m2_1732_5966# ctop 0.0428f
C19009 col_n[13] rowoff_n[1] 0.0471f
C19010 col_n[15] rowoff_n[3] 0.0471f
C19011 col_n[19] rowoff_n[7] 0.0471f
C19012 col[27] a_2475_3158# 0.136f
C19013 col_n[18] rowoff_n[6] 0.0471f
C19014 col_n[20] rowoff_n[8] 0.0471f
C19015 col_n[14] rowoff_n[2] 0.0471f
C19016 ctop a_25054_11166# 4.11f
C19017 col_n[17] rowoff_n[5] 0.0471f
C19018 col_n[21] rowoff_n[9] 0.0471f
C19019 col_n[16] rowoff_n[4] 0.0471f
C19020 col_n[12] rowoff_n[0] 0.0471f
C19021 a_25966_18194# a_26058_18194# 0.0991f
C19022 VDD a_33998_16186# 0.181f
C19023 a_20946_1126# a_21038_1126# 0.0991f
C19024 m2_33284_15430# rowon_n[13] 0.0322f
C19025 col_n[27] a_30474_8516# 0.0283f
C19026 m2_6752_946# m3_7888_1078# 0.0341f
C19027 vcm a_5886_10162# 0.1f
C19028 a_27062_11166# a_27062_10162# 0.843f
C19029 a_2475_10186# a_18026_10162# 0.316f
C19030 row_n[14] a_23046_16186# 0.282f
C19031 a_20946_15182# a_21342_15222# 0.0313f
C19032 m2_16792_18014# col_n[14] 0.243f
C19033 VDD a_25454_10524# 0.0779f
C19034 ctop a_5978_14178# 4.11f
C19035 row_n[4] a_33086_6146# 0.282f
C19036 col[10] a_13006_12170# 0.367f
C19037 col[7] a_9902_2130# 0.0682f
C19038 col[19] a_2275_17214# 0.0899f
C19039 rowon_n[8] a_32994_10162# 0.118f
C19040 m2_1732_3958# a_2275_4162# 0.191f
C19041 col[17] a_19942_14178# 0.0682f
C19042 col[24] a_2275_6170# 0.0899f
C19043 a_5886_7150# a_6378_7512# 0.0658f
C19044 a_2275_7174# a_8990_7150# 0.399f
C19045 rowoff_n[10] a_25454_12532# 0.0133f
C19046 rowoff_n[2] a_8386_4500# 0.0133f
C19047 a_4974_7150# a_5278_7190# 0.0931f
C19048 col[22] rowoff_n[14] 0.0901f
C19049 m2_20808_18014# vcm 0.353f
C19050 row_n[6] a_20338_8194# 0.0117f
C19051 col_n[25] a_28066_8154# 0.251f
C19052 vcm a_20946_14178# 0.1f
C19053 a_2475_12194# a_33086_12170# 0.316f
C19054 a_17022_12170# a_18026_12170# 0.843f
C19055 VDD a_17022_4138# 0.483f
C19056 col_n[5] rowoff_n[10] 0.0471f
C19057 VDD a_6378_13536# 0.0779f
C19058 col_n[5] a_8290_12210# 0.084f
C19059 row_n[8] a_10906_10162# 0.0437f
C19060 rowoff_n[0] a_17422_2492# 0.0133f
C19061 rowon_n[12] a_9994_14178# 0.248f
C19062 m2_30848_946# ctop 0.0428f
C19063 a_2275_9182# a_24050_9158# 0.399f
C19064 rowoff_n[13] a_6982_15182# 0.294f
C19065 col_n[9] a_2475_13198# 0.0531f
C19066 col_n[16] a_19430_6508# 0.0283f
C19067 rowon_n[2] a_20034_4138# 0.248f
C19068 col_n[14] a_2475_2154# 0.0531f
C19069 col_n[26] a_29470_18556# 0.0283f
C19070 vcm a_34394_18234# 0.16f
C19071 a_7986_14178# a_7986_13174# 0.843f
C19072 VDD a_32082_8154# 0.483f
C19073 rowoff_n[5] a_8990_7150# 0.294f
C19074 a_2161_18218# a_2275_18218# 0.183f
C19075 VDD a_21438_17552# 0.0779f
C19076 a_30986_2130# a_31382_2170# 0.0313f
C19077 vcm col_n[19] 1.94f
C19078 col_n[9] col_n[10] 0.0101f
C19079 VDD col_n[22] 5.17f
C19080 vcm a_3970_2130# 0.56f
C19081 col[19] col[20] 0.0355f
C19082 col[6] rowoff_n[15] 0.0901f
C19083 a_2275_6170# a_14314_6186# 0.144f
C19084 a_2475_6170# a_16930_6146# 0.264f
C19085 rowoff_n[3] a_18026_5142# 0.294f
C19086 col[6] a_8898_12170# 0.0682f
C19087 a_20946_11166# a_21438_11528# 0.0658f
C19088 a_20034_11166# a_20338_11206# 0.0931f
C19089 m2_13780_18014# a_14010_17190# 0.843f
C19090 m2_5172_13422# row_n[11] 0.0128f
C19091 m2_11196_9406# row_n[7] 0.0128f
C19092 col_n[14] a_17022_6146# 0.251f
C19093 m2_17220_5390# row_n[3] 0.0128f
C19094 m3_1864_4090# a_2966_4138# 0.0302f
C19095 row_n[11] a_31078_13174# 0.282f
C19096 a_32082_16186# a_33086_16186# 0.843f
C19097 VDD a_13006_11166# 0.483f
C19098 rowon_n[15] a_30986_17190# 0.118f
C19099 col_n[6] a_2275_16210# 0.113f
C19100 col_n[21] a_23958_8154# 0.0765f
C19101 col_n[11] a_2275_5166# 0.113f
C19102 a_2275_3158# a_7894_3134# 0.136f
C19103 rowoff_n[1] a_27062_3134# 0.294f
C19104 m2_34864_5966# a_34090_6146# 0.843f
C19105 row_n[13] a_18330_15222# 0.0117f
C19106 vcm a_19030_6146# 0.56f
C19107 rowoff_n[11] a_13406_13536# 0.0133f
C19108 a_2475_8178# a_31990_8154# 0.264f
C19109 a_16930_8154# a_17022_8154# 0.326f
C19110 a_2275_8178# a_29374_8194# 0.144f
C19111 col_n[26] a_2475_15206# 0.0531f
C19112 col_n[5] a_8386_4500# 0.0283f
C19113 row_n[3] a_28370_5182# 0.0117f
C19114 col_n[31] a_2475_4162# 0.0531f
C19115 col[1] a_2275_2154# 0.0899f
C19116 row_n[15] a_8898_17190# 0.0437f
C19117 m2_32280_14426# row_n[12] 0.0128f
C19118 col_n[15] a_18426_16548# 0.0283f
C19119 a_2475_17214# a_9994_17190# 0.316f
C19120 VDD a_28066_15182# 0.483f
C19121 row_n[5] a_18938_7150# 0.0437f
C19122 a_11910_5142# a_12306_5182# 0.0313f
C19123 a_2275_5166# a_22954_5142# 0.136f
C19124 m2_1732_3958# sample_n 0.0522f
C19125 col[16] a_2475_12194# 0.136f
C19126 rowon_n[9] a_18026_11166# 0.248f
C19127 vcm a_34090_10162# 0.56f
C19128 col[21] a_2475_1150# 0.136f
C19129 rowoff_n[15] a_29470_17552# 0.0133f
C19130 m2_28264_16434# a_28066_16186# 0.165f
C19131 col_n[0] a_2874_12170# 0.0765f
C19132 m3_6884_1078# a_6982_2130# 0.0302f
C19133 m2_10768_946# a_2275_1150# 0.28f
C19134 col_n[3] a_5978_4138# 0.251f
C19135 col_n[29] a_32386_5182# 0.084f
C19136 VDD a_8990_18194# 0.0356f
C19137 col_n[23] a_2275_18218# 0.113f
C19138 a_2475_2154# a_15014_2130# 0.316f
C19139 a_7986_2130# a_8990_2130# 0.843f
C19140 col_n[13] a_16018_16186# 0.251f
C19141 col_n[28] a_2275_7174# 0.113f
C19142 col_n[10] a_12914_6146# 0.0765f
C19143 m2_5172_1374# VDD 0.0193f
C19144 vcm a_24354_4178# 0.155f
C19145 rowoff_n[9] a_19942_11166# 0.202f
C19146 col_n[20] a_22954_18194# 0.0762f
C19147 vcm a_15014_13174# 0.56f
C19148 a_31990_12170# a_32082_12170# 0.326f
C19149 VDD a_11910_3134# 0.181f
C19150 m2_11772_18014# a_2275_18218# 0.28f
C19151 col[13] a_2275_15206# 0.0899f
C19152 a_2275_16210# a_16018_16186# 0.399f
C19153 rowon_n[3] a_5886_5142# 0.118f
C19154 col[18] a_2275_4162# 0.0899f
C19155 a_25054_1126# m2_24824_946# 0.0249f
C19156 rowoff_n[7] a_28978_9158# 0.202f
C19157 m2_34864_9982# rowoff_n[8] 0.278f
C19158 col_n[4] a_7382_14540# 0.0283f
C19159 a_33086_5142# a_33086_4138# 0.843f
C19160 col_n[1] a_3878_4138# 0.0765f
C19161 a_2475_4162# a_30074_4138# 0.316f
C19162 col[23] a_26058_3134# 0.367f
C19163 vcm a_5278_7190# 0.155f
C19164 a_26970_9158# a_27366_9198# 0.0313f
C19165 col[30] a_32994_5142# 0.0682f
C19166 row_n[10] a_26362_12210# 0.0117f
C19167 m2_19228_14426# a_19030_14178# 0.165f
C19168 col_n[24] rowoff_n[1] 0.0471f
C19169 col_n[28] rowoff_n[5] 0.0471f
C19170 col_n[30] rowoff_n[7] 0.0471f
C19171 col_n[23] rowoff_n[0] 0.0471f
C19172 col_n[25] rowoff_n[2] 0.0471f
C19173 col_n[27] rowoff_n[4] 0.0471f
C19174 col_n[26] rowoff_n[3] 0.0471f
C19175 col_n[29] rowoff_n[6] 0.0471f
C19176 col_n[31] rowoff_n[8] 0.0471f
C19177 ctop a_18026_2130# 4.09f
C19178 vcm a_30074_17190# 0.56f
C19179 a_2475_13198# a_8898_13174# 0.264f
C19180 a_2275_13198# a_6282_13214# 0.144f
C19181 VDD a_26970_7150# 0.181f
C19182 col_n[9] a_2475_18218# 0.0529f
C19183 a_2275_18218# a_31078_18194# 0.0924f
C19184 m2_7756_18014# a_2475_18218# 0.286f
C19185 a_16930_18194# a_17422_18556# 0.0658f
C19186 a_11910_1126# a_12402_1488# 0.0658f
C19187 a_2275_1150# a_21038_1126# 0.0924f
C19188 row_n[12] a_16930_14178# 0.0437f
C19189 col_n[3] a_2475_11190# 0.0531f
C19190 m2_16216_2378# a_16018_2130# 0.165f
C19191 col_n[18] a_21342_3174# 0.084f
C19192 vcm a_32994_2130# 0.1f
C19193 a_23046_6146# a_24050_6146# 0.843f
C19194 col_n[28] a_31382_15222# 0.084f
C19195 col_n[2] a_4974_14178# 0.251f
C19196 vcm a_20338_11206# 0.155f
C19197 row_n[2] a_26970_4138# 0.0437f
C19198 a_35002_11166# a_35398_11206# 0.0313f
C19199 VDD a_18426_1488# 0.0914f
C19200 col_n[9] a_11910_16186# 0.0765f
C19201 rowon_n[6] a_26058_8154# 0.248f
C19202 m2_32856_18014# a_33086_17190# 0.843f
C19203 ctop a_33086_6146# 4.11f
C19204 a_12914_15182# a_13006_15182# 0.326f
C19205 a_2275_15206# a_21342_15222# 0.144f
C19206 a_2475_15206# a_23958_15182# 0.264f
C19207 VDD a_7894_10162# 0.181f
C19208 col[30] a_2275_17214# 0.0899f
C19209 a_2475_18218# a_29070_18194# 0.0299f
C19210 vcm a_13918_5142# 0.1f
C19211 rowoff_n[10] a_7894_12170# 0.202f
C19212 a_14010_8154# a_14010_7150# 0.843f
C19213 col_n[16] rowoff_n[10] 0.0471f
C19214 a_27062_1126# vcm 0.165f
C19215 m2_10192_12418# a_9994_12170# 0.165f
C19216 row_n[6] a_3970_8154# 0.282f
C19217 m2_1732_7974# rowon_n[6] 0.236f
C19218 vcm a_2275_14202# 6.49f
C19219 a_2275_12194# a_14922_12170# 0.136f
C19220 a_7894_12170# a_8290_12210# 0.0313f
C19221 m2_7180_4386# rowon_n[2] 0.0322f
C19222 VDD a_33486_5504# 0.0779f
C19223 col[22] a_25054_13174# 0.367f
C19224 col_n[5] a_2275_3158# 0.113f
C19225 col[19] a_21950_3134# 0.0682f
C19226 m2_24824_18014# VDD 0.993f
C19227 ctop a_14010_9158# 4.11f
C19228 a_2966_17190# a_2966_16186# 0.843f
C19229 VDD a_22954_14178# 0.181f
C19230 col[29] a_31990_15182# 0.0682f
C19231 a_2275_1150# m2_1732_946# 0.191f
C19232 rowon_n[0] a_13918_2130# 0.118f
C19233 col_n[20] a_2475_13198# 0.0531f
C19234 a_26058_5142# a_26362_5182# 0.0931f
C19235 a_26970_5142# a_27462_5504# 0.0658f
C19236 m2_29268_8402# a_29070_8154# 0.165f
C19237 col_n[25] a_2475_2154# 0.0531f
C19238 col_n[7] a_10298_1166# 0.0839f
C19239 vcm a_28978_9158# 0.1f
C19240 m2_11772_18014# m2_12200_18442# 0.165f
C19241 a_2475_9182# a_6982_9158# 0.316f
C19242 a_3970_9158# a_4974_9158# 0.843f
C19243 rowoff_n[14] a_23958_16186# 0.202f
C19244 col_n[17] a_20338_13214# 0.084f
C19245 rowon_n[2] a_1957_4162# 0.0172f
C19246 vcm a_16322_18234# 0.16f
C19247 m2_16216_17438# rowon_n[15] 0.0322f
C19248 a_2275_14202# a_29982_14178# 0.136f
C19249 row_n[7] a_35398_9198# 0.0117f
C19250 VDD a_14410_8516# 0.0779f
C19251 m2_22240_13422# rowon_n[11] 0.0322f
C19252 m2_28264_9406# rowon_n[7] 0.0322f
C19253 m2_34288_5390# rowon_n[3] 0.0322f
C19254 ctop a_29070_13174# 4.11f
C19255 VDD row_n[15] 3.29f
C19256 sample rowon_n[15] 0.0935f
C19257 vcm col_n[30] 1.94f
C19258 col[10] a_2475_10186# 0.136f
C19259 col[17] rowoff_n[15] 0.0901f
C19260 VDD a_3366_17552# 0.0779f
C19261 a_22954_2130# a_23046_2130# 0.326f
C19262 col_n[28] a_31478_7512# 0.0283f
C19263 vcm rowoff_n[11] 0.533f
C19264 row_n[9] a_24962_11166# 0.0437f
C19265 rowon_n[13] a_24050_15182# 0.248f
C19266 vcm a_9902_12170# 0.1f
C19267 a_29070_12170# a_29070_11166# 0.843f
C19268 a_2475_11190# a_22042_11166# 0.316f
C19269 VDD a_5978_2130# 0.483f
C19270 col_n[17] a_2275_16210# 0.113f
C19271 a_22954_16186# a_23350_16226# 0.0313f
C19272 col_n[22] a_2275_5166# 0.113f
C19273 rowon_n[3] a_34090_5142# 0.248f
C19274 VDD a_29470_12532# 0.0779f
C19275 m2_18800_18014# m3_18932_18146# 3.79f
C19276 col[11] a_14010_11166# 0.367f
C19277 col[8] a_10906_1126# 0.0682f
C19278 ctop a_9994_16186# 4.11f
C19279 col[18] a_20946_13174# 0.0682f
C19280 rowoff_n[1] a_9390_3496# 0.0133f
C19281 m2_20232_6394# a_20034_6146# 0.165f
C19282 row_n[13] a_2475_15206# 0.405f
C19283 col_n[26] a_29070_7150# 0.251f
C19284 a_6982_8154# a_7286_8194# 0.0931f
C19285 col[7] a_2275_13198# 0.0899f
C19286 a_7894_8154# a_8386_8516# 0.0658f
C19287 a_2275_8178# a_13006_8154# 0.399f
C19288 col[12] a_2275_2154# 0.0899f
C19289 vcm a_24962_16186# 0.1f
C19290 a_19030_13174# a_20034_13174# 0.843f
C19291 VDD a_21038_6146# 0.483f
C19292 row_n[3] a_12002_5142# 0.282f
C19293 col_n[6] a_9294_11206# 0.084f
C19294 rowon_n[7] a_11910_9158# 0.118f
C19295 VDD a_10394_15544# 0.0779f
C19296 col[27] a_2475_12194# 0.136f
C19297 a_2275_5166# a_3270_5182# 0.144f
C19298 a_2475_5166# a_5886_5142# 0.264f
C19299 col_n[17] a_20434_5504# 0.0283f
C19300 m3_31984_18146# m3_32988_18146# 0.202f
C19301 m2_22816_946# m3_21944_1078# 0.0341f
C19302 col_n[27] a_30474_17552# 0.0283f
C19303 a_2275_10186# a_28066_10162# 0.399f
C19304 rowoff_n[15] a_11910_17190# 0.202f
C19305 row_n[14] a_32386_16226# 0.0117f
C19306 rowoff_n[4] a_9994_6146# 0.294f
C19307 a_9994_15182# a_9994_14178# 0.843f
C19308 VDD a_2475_9182# 26.1f
C19309 a_32994_3134# a_33390_3174# 0.0313f
C19310 col[0] a_2874_9158# 0.0682f
C19311 m2_11196_4386# a_10998_4138# 0.165f
C19312 m2_6176_3382# row_n[1] 0.0128f
C19313 vcm a_7986_4138# 0.56f
C19314 m2_33860_946# col_n[31] 0.637f
C19315 a_2475_7174# a_20946_7150# 0.264f
C19316 a_2275_7174# a_18330_7190# 0.144f
C19317 col[7] a_9902_11166# 0.0682f
C19318 rowoff_n[2] a_19030_4138# 0.294f
C19319 col[24] a_2275_15206# 0.0899f
C19320 row_n[6] a_32994_8154# 0.0437f
C19321 col_n[15] a_18026_5142# 0.251f
C19322 a_22954_12170# a_23446_12532# 0.0658f
C19323 a_22042_12170# a_22346_12210# 0.0931f
C19324 col[29] a_2275_4162# 0.0899f
C19325 rowon_n[10] a_32082_12170# 0.248f
C19326 col_n[25] a_28066_17190# 0.251f
C19327 m2_31852_18014# col[29] 0.347f
C19328 col_n[22] a_24962_7150# 0.0765f
C19329 a_33998_17190# a_34394_17230# 0.0313f
C19330 VDD a_17022_13174# 0.483f
C19331 rowoff_n[0] a_28066_2130# 0.294f
C19332 a_2275_4162# a_11910_4138# 0.136f
C19333 row_n[10] rowoff_n[9] 0.085f
C19334 m2_15212_16434# row_n[14] 0.0128f
C19335 col_n[0] a_2275_1150# 0.113f
C19336 m2_21236_12418# row_n[10] 0.0128f
C19337 vcm a_23046_8154# 0.56f
C19338 a_2275_9182# a_33390_9198# 0.144f
C19339 a_18938_9158# a_19030_9158# 0.326f
C19340 m2_27260_8402# row_n[6] 0.0128f
C19341 m2_33284_4386# row_n[2] 0.0128f
C19342 row_n[10] a_9994_12170# 0.282f
C19343 col_n[20] a_2475_18218# 0.0529f
C19344 col_n[6] a_9390_3496# 0.0283f
C19345 col[2] a_3878_1126# 0.011f
C19346 rowon_n[14] a_9902_16186# 0.118f
C19347 col_n[16] a_19430_15544# 0.0283f
C19348 col_n[14] a_2475_11190# 0.0531f
C19349 row_n[0] a_20034_2130# 0.282f
C19350 VDD a_32082_17190# 0.484f
C19351 a_2275_1150# a_2966_1126# 0.0924f
C19352 a_2475_1150# a_3970_1126# 0.311f
C19353 a_20034_2130# a_20034_1126# 0.843f
C19354 rowon_n[4] a_19942_6146# 0.118f
C19355 m2_1732_1950# a_1957_2154# 0.245f
C19356 vcm a_13310_2170# 0.155f
C19357 a_13918_6146# a_14314_6186# 0.0313f
C19358 a_2275_6170# a_26970_6146# 0.136f
C19359 row_n[2] a_7286_4178# 0.0117f
C19360 vcm a_3970_11166# 0.56f
C19361 VDD a_35002_2130# 0.258f
C19362 col[4] a_2475_8178# 0.136f
C19363 a_2874_15182# a_3270_15222# 0.0313f
C19364 a_3878_15182# a_3970_15182# 0.326f
C19365 a_2275_15206# a_4974_15182# 0.399f
C19366 col_n[4] a_6982_3134# 0.251f
C19367 col_n[30] a_33390_4178# 0.084f
C19368 col_n[14] a_17022_15182# 0.251f
C19369 col_n[11] a_13918_5142# 0.0765f
C19370 a_9994_3134# a_10998_3134# 0.843f
C19371 col_n[27] rowoff_n[10] 0.0471f
C19372 a_2475_3158# a_19030_3134# 0.316f
C19373 rowoff_n[8] a_20946_10162# 0.202f
C19374 col_n[21] a_23958_17190# 0.0765f
C19375 a_30378_1166# a_2275_1150# 0.145f
C19376 a_32994_1126# a_2475_1150# 0.264f
C19377 col_n[11] a_2275_14202# 0.113f
C19378 row_n[13] a_30986_15182# 0.0437f
C19379 vcm a_28370_6186# 0.155f
C19380 rowoff_n[11] a_24050_13174# 0.294f
C19381 col_n[16] a_2275_3158# 0.113f
C19382 vcm a_19030_15182# 0.56f
C19383 a_33998_13174# a_34090_13174# 0.326f
C19384 VDD a_15926_5142# 0.181f
C19385 a_29070_1126# VDD 0.035f
C19386 a_2275_17214# a_20034_17190# 0.399f
C19387 rowoff_n[6] a_29982_8154# 0.202f
C19388 col_n[5] a_8386_13536# 0.0283f
C19389 col_n[31] a_2475_13198# 0.0531f
C19390 col[1] a_2275_11190# 0.0899f
C19391 m3_26964_18146# a_27062_17190# 0.0303f
C19392 col[24] a_27062_2130# 0.367f
C19393 a_2475_5166# a_34090_5142# 0.316f
C19394 m3_21944_1078# m3_22948_1078# 0.202f
C19395 col[31] a_33998_4138# 0.0682f
C19396 vcm a_9294_9198# 0.155f
C19397 a_28978_10162# a_29374_10202# 0.0313f
C19398 m2_1732_15002# a_2161_15206# 0.0454f
C19399 col_n[6] row_n[14] 0.298f
C19400 vcm row_n[11] 0.616f
C19401 sample row_n[10] 0.423f
C19402 col_n[8] row_n[15] 0.298f
C19403 ctop a_22042_4138# 4.11f
C19404 col_n[4] row_n[13] 0.298f
C19405 col_n[3] rowon_n[12] 0.111f
C19406 col_n[20] col_n[21] 0.0101f
C19407 VDD rowon_n[9] 3.04f
C19408 col_n[9] rowon_n[15] 0.111f
C19409 col_n[0] rowon_n[10] 0.111f
C19410 col_n[7] rowon_n[14] 0.111f
C19411 col_n[2] row_n[12] 0.298f
C19412 col_n[1] rowon_n[11] 0.111f
C19413 col_n[5] rowon_n[13] 0.111f
C19414 col[28] rowoff_n[15] 0.0901f
C19415 a_2275_14202# a_10298_14218# 0.144f
C19416 col[21] a_2475_10186# 0.136f
C19417 m2_33860_946# a_2275_1150# 0.222f
C19418 a_2475_14202# a_12914_14178# 0.264f
C19419 col[30] col[31] 0.0337f
C19420 m2_12776_946# a_12914_1126# 0.225f
C19421 row_n[7] a_18026_9158# 0.282f
C19422 VDD a_30986_9158# 0.181f
C19423 rowon_n[11] a_17934_13174# 0.118f
C19424 col_n[11] rowoff_n[11] 0.0471f
C19425 VDD a_18330_18234# 0.019f
C19426 col_n[19] a_22346_2170# 0.084f
C19427 a_13918_2130# a_14410_2492# 0.0658f
C19428 a_13006_2130# a_13310_2170# 0.0931f
C19429 a_2275_2154# a_25054_2130# 0.399f
C19430 col_n[3] a_5978_13174# 0.251f
C19431 col_n[29] a_32386_14218# 0.084f
C19432 m2_28264_1374# VDD 0.0194f
C19433 row_n[9] a_5278_11206# 0.0117f
C19434 vcm a_2161_3158# 0.0169f
C19435 a_25054_7150# a_26058_7150# 0.843f
C19436 rowoff_n[9] a_30474_11528# 0.0133f
C19437 rowon_n[1] a_27974_3134# 0.118f
C19438 col_n[28] a_2275_16210# 0.113f
C19439 col_n[10] a_12914_15182# 0.0765f
C19440 vcm a_24354_13214# 0.155f
C19441 a_2874_11166# a_2966_11166# 0.326f
C19442 VDD a_22442_3496# 0.0779f
C19443 m2_12776_18014# a_13006_18194# 0.0249f
C19444 a_2475_16210# a_27974_16186# 0.264f
C19445 a_2275_16210# a_25358_16226# 0.144f
C19446 a_14922_16186# a_15014_16186# 0.326f
C19447 VDD a_11910_12170# 0.181f
C19448 a_31382_1166# m2_30848_946# 0.087f
C19449 col[18] a_2275_13198# 0.0899f
C19450 row_n[1] a_5886_3134# 0.0437f
C19451 col[23] a_2275_2154# 0.0899f
C19452 vcm a_17934_7150# 0.1f
C19453 rowon_n[5] a_4974_7150# 0.248f
C19454 col_n[1] a_3878_13174# 0.0765f
C19455 a_16018_9158# a_16018_8154# 0.843f
C19456 rowoff_n[12] a_12002_14178# 0.294f
C19457 col[23] a_26058_12170# 0.367f
C19458 vcm a_5278_16226# 0.155f
C19459 col[20] a_22954_2130# 0.0682f
C19460 a_9902_13174# a_10298_13214# 0.0313f
C19461 a_2275_13198# a_18938_13174# 0.136f
C19462 VDD a_2966_6146# 0.485f
C19463 col[30] a_32994_14178# 0.0682f
C19464 ctop a_18026_11166# 4.11f
C19465 VDD a_26970_16186# 0.181f
C19466 m2_5172_15430# rowon_n[13] 0.0322f
C19467 a_28978_6146# a_29470_6508# 0.0658f
C19468 a_28066_6146# a_28370_6186# 0.0931f
C19469 m2_11196_11414# rowon_n[9] 0.0322f
C19470 m2_17220_7398# rowon_n[5] 0.0322f
C19471 m2_23244_3382# rowon_n[1] 0.0322f
C19472 m2_32856_946# m2_33860_946# 0.843f
C19473 col_n[18] a_21342_12210# 0.084f
C19474 vcm a_32994_11166# 0.1f
C19475 col_n[8] a_2475_9182# 0.0531f
C19476 a_2475_10186# a_10998_10162# 0.316f
C19477 a_5978_10162# a_6982_10162# 0.843f
C19478 row_n[14] a_16018_16186# 0.282f
C19479 m2_34288_17438# a_34090_17190# 0.165f
C19480 a_2275_15206# a_33998_15182# 0.136f
C19481 VDD a_18426_10524# 0.0779f
C19482 ctop a_33086_15182# 4.11f
C19483 col_n[29] a_32482_6508# 0.0283f
C19484 row_n[4] a_26058_6146# 0.282f
C19485 a_24962_3134# a_25054_3134# 0.326f
C19486 rowon_n[8] a_25966_10162# 0.118f
C19487 rowoff_n[10] a_18426_12532# 0.0133f
C19488 a_1957_7174# a_2161_7174# 0.115f
C19489 a_2475_7174# a_2275_7174# 2.76f
C19490 m2_6752_18014# vcm 0.353f
C19491 m2_32280_16434# rowon_n[14] 0.0322f
C19492 row_n[6] a_13310_8194# 0.0117f
C19493 vcm a_13918_14178# 0.1f
C19494 a_2475_12194# a_26058_12170# 0.316f
C19495 a_31078_13174# a_31078_12170# 0.843f
C19496 VDD a_9994_4138# 0.483f
C19497 col[12] a_15014_10162# 0.367f
C19498 a_24962_17190# a_25358_17230# 0.0313f
C19499 VDD a_33486_14540# 0.0779f
C19500 col_n[5] a_2275_12194# 0.113f
C19501 col[19] a_21950_12170# 0.0682f
C19502 row_n[6] rowoff_n[6] 0.209f
C19503 col_n[10] a_2275_1150# 0.113f
C19504 rowoff_n[0] a_10394_2492# 0.0133f
C19505 rowon_n[12] a_2874_14178# 0.118f
C19506 col_n[27] a_30074_6146# 0.251f
C19507 col_n[31] a_2475_18218# 0.0529f
C19508 m2_3164_7398# a_2966_7150# 0.165f
C19509 a_8990_9158# a_9294_9198# 0.0931f
C19510 a_2275_9182# a_17022_9158# 0.399f
C19511 a_9902_9158# a_10394_9520# 0.0658f
C19512 rowoff_n[14] a_34490_16548# 0.0133f
C19513 m2_25252_15430# a_25054_15182# 0.165f
C19514 rowon_n[2] a_13006_4138# 0.248f
C19515 col_n[25] a_2475_11190# 0.0531f
C19516 vcm a_28978_18194# 0.101f
C19517 col_n[7] a_10298_10202# 0.084f
C19518 a_21038_14178# a_22042_14178# 0.843f
C19519 VDD a_25054_8154# 0.483f
C19520 rowoff_n[5] a_2475_7174# 3.9f
C19521 row_n[0] a_1957_2154# 0.187f
C19522 VDD a_14410_17552# 0.0779f
C19523 col_n[18] a_21438_4500# 0.0283f
C19524 vcm a_31078_3134# 0.56f
C19525 a_2475_6170# a_9902_6146# 0.264f
C19526 a_5886_6146# a_5978_6146# 0.326f
C19527 a_2275_6170# a_7286_6186# 0.144f
C19528 col[15] a_2475_8178# 0.136f
C19529 col_n[28] a_31478_16548# 0.0283f
C19530 rowoff_n[3] a_10998_5142# 0.294f
C19531 a_2275_11190# a_32082_11166# 0.399f
C19532 m2_31852_18014# a_32082_18194# 0.0249f
C19533 a_12002_16186# a_12002_15182# 0.843f
C19534 row_n[11] a_24050_13174# 0.282f
C19535 VDD a_5978_11166# 0.483f
C19536 m2_32856_18014# m3_33992_18146# 0.0341f
C19537 rowon_n[15] a_23958_17190# 0.118f
C19538 col[1] a_3970_8154# 0.367f
C19539 col_n[22] a_2275_14202# 0.113f
C19540 m2_1732_7974# col[0] 0.0137f
C19541 col_n[27] a_2275_3158# 0.113f
C19542 col[8] a_10906_10162# 0.0682f
C19543 rowoff_n[1] a_20034_3134# 0.294f
C19544 row_n[1] a_34090_3134# 0.282f
C19545 rowoff_n[8] a_2275_10186# 0.151f
C19546 row_n[13] a_11302_15222# 0.0117f
C19547 rowon_n[5] a_33998_7150# 0.118f
C19548 vcm a_12002_6146# 0.56f
C19549 rowoff_n[11] a_6378_13536# 0.0133f
C19550 a_2475_8178# a_24962_8154# 0.264f
C19551 a_2275_8178# a_22346_8194# 0.144f
C19552 col_n[16] a_19030_4138# 0.251f
C19553 m2_16216_13422# a_16018_13174# 0.165f
C19554 col_n[26] a_29070_16186# 0.251f
C19555 a_24962_13174# a_25454_13536# 0.0658f
C19556 a_24050_13174# a_24354_13214# 0.0931f
C19557 col_n[23] a_25966_6146# 0.0765f
C19558 row_n[3] a_21342_5182# 0.0117f
C19559 col[12] a_2275_11190# 0.0899f
C19560 m2_4168_14426# row_n[12] 0.0128f
C19561 a_1957_17214# a_2275_17214# 0.158f
C19562 a_2475_17214# a_2874_17190# 0.264f
C19563 VDD a_21038_15182# 0.483f
C19564 m2_10192_10410# row_n[8] 0.0128f
C19565 m2_16216_6394# row_n[4] 0.0128f
C19566 a_23350_1166# col_n[20] 0.0839f
C19567 row_n[5] a_11910_7150# 0.0437f
C19568 a_2275_5166# a_15926_5142# 0.136f
C19569 m2_1732_1950# vcm 0.316f
C19570 m3_34996_9110# m3_34996_8106# 0.202f
C19571 m2_34864_8978# a_35094_9158# 0.0249f
C19572 col_n[6] rowon_n[8] 0.111f
C19573 col_n[4] rowon_n[7] 0.111f
C19574 rowon_n[9] a_10998_11166# 0.248f
C19575 col_n[17] row_n[14] 0.298f
C19576 col_n[9] row_n[10] 0.298f
C19577 col_n[7] row_n[9] 0.298f
C19578 vcm rowon_n[5] 0.65f
C19579 col_n[2] rowon_n[6] 0.111f
C19580 col_n[20] rowon_n[15] 0.111f
C19581 col_n[15] row_n[13] 0.298f
C19582 col_n[16] rowon_n[13] 0.111f
C19583 col_n[10] rowon_n[10] 0.111f
C19584 col_n[8] rowon_n[9] 0.111f
C19585 sample rowon_n[4] 0.0935f
C19586 col_n[12] rowon_n[11] 0.111f
C19587 col_n[1] row_n[6] 0.298f
C19588 col_n[13] row_n[12] 0.298f
C19589 col_n[18] rowon_n[14] 0.111f
C19590 col_n[3] row_n[7] 0.298f
C19591 col_n[14] rowon_n[12] 0.111f
C19592 col_n[11] row_n[11] 0.298f
C19593 col_n[0] row_n[5] 0.298f
C19594 col_n[19] row_n[15] 0.298f
C19595 col_n[5] row_n[8] 0.298f
C19596 VDD row_n[4] 3.29f
C19597 col_n[7] a_10394_2492# 0.0283f
C19598 vcm a_27062_10162# 0.56f
C19599 a_20946_10162# a_21038_10162# 0.326f
C19600 rowoff_n[15] a_22442_17552# 0.0133f
C19601 col_n[17] a_20434_14540# 0.0283f
C19602 m2_23820_946# a_24050_2130# 0.843f
C19603 col_n[22] rowoff_n[11] 0.0471f
C19604 a_2475_2154# a_7986_2130# 0.316f
C19605 a_22042_3134# a_22042_2130# 0.843f
C19606 m2_31276_15430# row_n[13] 0.0128f
C19607 col_n[2] a_2475_7174# 0.0531f
C19608 vcm a_17326_4178# 0.155f
C19609 col[0] a_2874_18194# 0.0682f
C19610 a_2275_7174# a_30986_7150# 0.136f
C19611 rowoff_n[9] a_12914_11166# 0.202f
C19612 a_15926_7150# a_16322_7190# 0.0313f
C19613 m2_7180_11414# a_6982_11166# 0.165f
C19614 vcm a_7986_13174# 0.56f
C19615 VDD a_4882_3134# 0.181f
C19616 col_n[5] a_7986_2130# 0.251f
C19617 a_2275_16210# a_8990_16186# 0.399f
C19618 col_n[15] a_18026_14178# 0.251f
C19619 a_5886_16186# a_6378_16548# 0.0658f
C19620 a_4974_16186# a_5278_16226# 0.0931f
C19621 col[29] a_2275_13198# 0.0899f
C19622 col_n[12] a_14922_4138# 0.0765f
C19623 row_n[8] a_32082_10162# 0.282f
C19624 rowoff_n[7] a_21950_9158# 0.202f
C19625 col_n[22] a_24962_16186# 0.0765f
C19626 rowon_n[12] a_31990_14178# 0.118f
C19627 a_2475_4162# a_23046_4138# 0.316f
C19628 a_12002_4138# a_13006_4138# 0.843f
C19629 m3_10900_1078# ctop 0.21f
C19630 m2_26256_7398# a_26058_7150# 0.165f
C19631 vcm a_32386_8194# 0.155f
C19632 rowoff_n[13] a_28978_15182# 0.202f
C19633 row_n[10] a_19334_12210# 0.0117f
C19634 col_n[6] rowoff_n[12] 0.0471f
C19635 col_n[0] a_2275_10186# 0.113f
C19636 ctop a_10998_2130# 4.06f
C19637 vcm a_23046_17190# 0.56f
C19638 VDD a_19942_7150# 0.181f
C19639 rowoff_n[5] a_30986_7150# 0.202f
C19640 col_n[6] a_9390_12532# 0.0283f
C19641 a_2275_18218# a_24050_18194# 0.0924f
C19642 row_n[0] a_29374_2170# 0.0117f
C19643 a_2275_1150# a_14010_1126# 0.0924f
C19644 row_n[12] a_9902_14178# 0.0437f
C19645 vcm a_25966_2130# 0.1f
C19646 col_n[19] a_2475_9182# 0.0531f
C19647 m2_13780_946# m2_14208_1374# 0.165f
C19648 row_n[2] a_19942_4138# 0.0437f
C19649 vcm a_13310_11206# 0.155f
C19650 a_30986_11166# a_31382_11206# 0.0313f
C19651 VDD a_11398_1488# 0.0977f
C19652 rowon_n[6] a_19030_8154# 0.248f
C19653 ctop a_26058_6146# 4.11f
C19654 a_2475_15206# a_16930_15182# 0.264f
C19655 a_2275_15206# a_14314_15222# 0.144f
C19656 VDD a_35002_11166# 0.258f
C19657 col[4] a_2475_17214# 0.136f
C19658 rowon_n[0] m2_28264_2378# 0.0322f
C19659 col[9] a_2475_6170# 0.136f
C19660 col_n[30] a_33390_13214# 0.084f
C19661 col_n[4] a_6982_12170# 0.251f
C19662 a_15926_3134# a_16418_3496# 0.0658f
C19663 a_2275_3158# a_29070_3134# 0.399f
C19664 a_15014_3134# a_15318_3174# 0.0931f
C19665 a_2475_18218# a_22042_18194# 0.0299f
C19666 rowoff_n[8] a_31478_10524# 0.0133f
C19667 m2_17220_5390# a_17022_5142# 0.165f
C19668 a_22346_1166# a_21950_1126# 0.0313f
C19669 col_n[11] a_13918_14178# 0.0765f
C19670 m2_1732_11990# m2_2160_12418# 0.165f
C19671 vcm a_6890_5142# 0.1f
C19672 a_27062_8154# a_28066_8154# 0.843f
C19673 vcm a_28370_15222# 0.155f
C19674 a_2275_12194# a_7894_12170# 0.136f
C19675 VDD a_26458_5504# 0.0779f
C19676 col_n[16] a_2275_12194# 0.113f
C19677 m2_10768_18014# VDD 1.1f
C19678 rowon_n[2] rowoff_n[2] 20.2f
C19679 ctop a_6982_9158# 4.11f
C19680 col_n[21] a_2275_1150# 0.113f
C19681 row_n[15] a_30074_17190# 0.282f
C19682 a_2275_17214# a_29374_17230# 0.144f
C19683 a_16930_17190# a_17022_17190# 0.326f
C19684 a_2475_17214# a_31990_17190# 0.264f
C19685 VDD a_15926_14178# 0.181f
C19686 rowon_n[0] a_6890_2130# 0.118f
C19687 col[24] a_27062_11166# 0.367f
C19688 col[6] a_2275_9182# 0.0899f
C19689 m2_4744_18014# m2_5172_18442# 0.165f
C19690 vcm a_21950_9158# 0.1f
C19691 col[21] a_23958_1126# 0.0682f
C19692 a_18026_10162# a_18026_9158# 0.843f
C19693 rowoff_n[14] a_16930_16186# 0.202f
C19694 col[31] a_33998_13174# 0.0682f
C19695 vcm a_9294_18234# 0.16f
C19696 a_11910_14178# a_12306_14218# 0.0313f
C19697 m2_20808_946# a_20034_1126# 0.843f
C19698 a_2275_14202# a_22954_14178# 0.136f
C19699 row_n[7] a_27366_9198# 0.0117f
C19700 VDD a_7382_8516# 0.0779f
C19701 m2_6176_5390# rowon_n[3] 0.0322f
C19702 m2_8760_946# vcm 0.353f
C19703 ctop a_22042_13174# 4.11f
C19704 VDD a_30986_18194# 0.343f
C19705 a_2275_2154# a_35398_2170# 0.145f
C19706 col[26] a_2475_8178# 0.136f
C19707 m2_8184_3382# a_7986_3134# 0.165f
C19708 m3_29976_18146# VDD 0.0314f
C19709 col_n[19] a_22346_11206# 0.084f
C19710 row_n[9] a_17934_11166# 0.0437f
C19711 a_30986_7150# a_31478_7512# 0.0658f
C19712 a_30074_7150# a_30378_7190# 0.0931f
C19713 rowon_n[13] a_17022_15182# 0.248f
C19714 vcm a_2161_12194# 0.0169f
C19715 a_2475_11190# a_15014_11166# 0.316f
C19716 a_7986_11166# a_8990_11166# 0.843f
C19717 VDD a_33086_3134# 0.483f
C19718 m2_18800_18014# a_19334_18234# 0.087f
C19719 col_n[30] a_33486_5504# 0.0283f
C19720 VDD a_22442_12532# 0.0779f
C19721 rowon_n[3] a_27062_5142# 0.248f
C19722 m2_9764_18014# m3_8892_18146# 0.0341f
C19723 m2_21236_14426# rowon_n[12] 0.0322f
C19724 m2_27260_10410# rowon_n[8] 0.0322f
C19725 m2_33284_6394# rowon_n[4] 0.0322f
C19726 a_26970_4138# a_27062_4138# 0.326f
C19727 rowoff_n[1] a_1957_3158# 0.0219f
C19728 m2_34864_16006# m2_34864_15002# 0.843f
C19729 a_2275_8178# a_5978_8154# 0.399f
C19730 col[23] a_2275_11190# 0.0899f
C19731 m2_1732_12994# a_2475_13198# 0.139f
C19732 col[13] a_16018_9158# 0.367f
C19733 vcm a_17934_16186# 0.1f
C19734 a_33086_14178# a_33086_13174# 0.843f
C19735 a_2475_13198# a_30074_13174# 0.316f
C19736 VDD a_14010_6146# 0.483f
C19737 row_n[3] a_4974_5142# 0.282f
C19738 col[20] a_22954_11166# 0.0682f
C19739 rowon_n[7] a_4882_9158# 0.118f
C19740 a_26970_18194# a_27366_18234# 0.0313f
C19741 VDD a_2966_15182# 0.485f
C19742 col_n[28] a_31078_5142# 0.251f
C19743 col_n[19] rowon_n[9] 0.111f
C19744 col_n[11] rowon_n[5] 0.111f
C19745 col_n[22] row_n[11] 0.298f
C19746 col_n[23] rowon_n[11] 0.111f
C19747 col_n[8] row_n[4] 0.298f
C19748 col_n[29] rowon_n[14] 0.111f
C19749 col_n[13] rowon_n[6] 0.111f
C19750 col_n[6] row_n[3] 0.298f
C19751 col_n[5] rowon_n[2] 0.111f
C19752 col_n[27] rowon_n[13] 0.111f
C19753 col_n[20] row_n[10] 0.298f
C19754 col_n[2] row_n[1] 0.298f
C19755 col_n[18] row_n[9] 0.298f
C19756 col_n[17] rowon_n[8] 0.111f
C19757 col_n[14] row_n[7] 0.298f
C19758 col_n[24] row_n[12] 0.298f
C19759 col_n[4] row_n[2] 0.298f
C19760 col_n[12] row_n[6] 0.298f
C19761 col_n[16] row_n[8] 0.298f
C19762 col_n[21] rowon_n[10] 0.111f
C19763 col_n[15] rowon_n[7] 0.111f
C19764 vcm row_n[0] 0.62f
C19765 col_n[1] rowon_n[0] 0.111f
C19766 col_n[25] rowon_n[12] 0.111f
C19767 col_n[28] row_n[14] 0.298f
C19768 col_n[3] rowon_n[1] 0.111f
C19769 col_n[7] rowon_n[3] 0.111f
C19770 col_n[10] row_n[5] 0.298f
C19771 col_n[31] rowon_n[15] 0.111f
C19772 VDD ctop 5.47f
C19773 col_n[26] row_n[13] 0.298f
C19774 col_n[30] row_n[15] 0.298f
C19775 col_n[9] rowon_n[4] 0.111f
C19776 vcm a_20034_1126# 0.557f
C19777 m3_17928_18146# m3_18932_18146# 0.202f
C19778 m2_11772_946# m3_12908_1078# 0.0341f
C19779 a_10998_10162# a_11302_10202# 0.0931f
C19780 col_n[8] a_11302_9198# 0.084f
C19781 a_11910_10162# a_12402_10524# 0.0658f
C19782 a_2275_10186# a_21038_10162# 0.399f
C19783 rowoff_n[15] a_4882_17190# 0.202f
C19784 row_n[14] a_25358_16226# 0.0117f
C19785 rowoff_n[4] a_2874_6146# 0.202f
C19786 a_23046_15182# a_24050_15182# 0.843f
C19787 VDD a_29070_10162# 0.483f
C19788 col_n[13] a_2475_7174# 0.0531f
C19789 col_n[19] a_22442_3496# 0.0283f
C19790 col_n[29] a_32482_15544# 0.0283f
C19791 vcm a_35094_5142# 0.165f
C19792 a_7894_7150# a_7986_7150# 0.326f
C19793 a_2275_7174# a_11302_7190# 0.144f
C19794 a_2475_7174# a_13918_7150# 0.264f
C19795 rowoff_n[10] a_29070_12170# 0.294f
C19796 rowoff_n[2] a_12002_4138# 0.294f
C19797 row_n[6] a_25966_8154# 0.0437f
C19798 col[3] a_2475_4162# 0.136f
C19799 rowon_n[10] a_25054_12170# 0.248f
C19800 col[2] a_4974_7150# 0.367f
C19801 a_14010_17190# a_14010_16186# 0.843f
C19802 VDD a_9994_13174# 0.483f
C19803 rowoff_n[7] a_3878_9158# 0.202f
C19804 col[9] a_11910_9158# 0.0682f
C19805 rowoff_n[0] a_21038_2130# 0.294f
C19806 rowon_n[0] a_35094_2130# 0.0141f
C19807 a_2275_4162# a_4882_4138# 0.136f
C19808 a_2966_4138# a_3970_4138# 0.843f
C19809 m3_6884_18146# ctop 0.209f
C19810 col_n[17] rowoff_n[12] 0.0471f
C19811 col_n[17] a_20034_3134# 0.251f
C19812 col_n[10] a_2275_10186# 0.113f
C19813 vcm a_16018_8154# 0.56f
C19814 col_n[27] a_30074_15182# 0.251f
C19815 a_2475_9182# a_28978_9158# 0.264f
C19816 a_2275_9182# a_26362_9198# 0.144f
C19817 m2_5172_4386# row_n[2] 0.0128f
C19818 row_n[10] a_2874_12170# 0.0436f
C19819 col_n[24] a_26970_5142# 0.0765f
C19820 m3_18932_1078# a_20034_1126# 0.0188f
C19821 a_26058_14178# a_26362_14218# 0.0931f
C19822 a_26970_14178# a_27462_14540# 0.0658f
C19823 rowon_n[14] a_2161_16210# 0.0177f
C19824 VDD a_35398_8194# 0.0882f
C19825 VDD a_25054_17190# 0.484f
C19826 col_n[30] a_2475_9182# 0.0531f
C19827 row_n[0] a_13006_2130# 0.282f
C19828 col[0] a_2275_7174# 0.099f
C19829 a_33086_2130# a_34090_2130# 0.843f
C19830 rowon_n[4] a_12914_6146# 0.118f
C19831 vcm a_6282_2170# 0.155f
C19832 a_2275_6170# a_19942_6146# 0.136f
C19833 col_n[8] a_11398_1488# 0.0283f
C19834 col_n[18] a_21438_13536# 0.0283f
C19835 m2_33860_946# sw 0.304f
C19836 vcm a_31078_12170# 0.56f
C19837 a_22954_11166# a_23046_11166# 0.326f
C19838 col[15] a_2475_17214# 0.136f
C19839 VDD a_27974_2130# 0.181f
C19840 m2_14208_17438# row_n[15] 0.0128f
C19841 m2_20232_13422# row_n[11] 0.0128f
C19842 m2_26256_9406# row_n[7] 0.0128f
C19843 col[20] a_2475_6170# 0.136f
C19844 m2_32280_5390# row_n[3] 0.0128f
C19845 row_n[11] a_33390_13214# 0.0117f
C19846 m2_34864_17010# m3_34996_17142# 3.79f
C19847 col_n[1] rowoff_n[13] 0.0471f
C19848 a_24050_4138# a_24050_3134# 0.843f
C19849 a_2475_3158# a_12002_3134# 0.316f
C19850 col[1] a_3970_17190# 0.367f
C19851 rowoff_n[8] a_13918_10162# 0.202f
C19852 m2_1732_4962# a_2966_5142# 0.843f
C19853 a_25966_1126# a_2475_1150# 0.264f
C19854 a_23350_1166# a_2275_1150# 0.145f
C19855 row_n[13] a_23958_15182# 0.0437f
C19856 vcm a_21342_6186# 0.155f
C19857 rowoff_n[11] a_17022_13174# 0.294f
C19858 a_2275_8178# a_35002_8154# 0.136f
C19859 col_n[27] a_2275_12194# 0.113f
C19860 a_17934_8154# a_18330_8194# 0.0313f
C19861 col[0] rowoff_n[5] 0.0901f
C19862 col[1] rowoff_n[6] 0.0901f
C19863 col[2] rowoff_n[7] 0.0901f
C19864 col[4] rowoff_n[9] 0.0901f
C19865 col[3] rowoff_n[8] 0.0901f
C19866 m2_10768_18014# col_n[8] 0.243f
C19867 vcm a_12002_15182# 0.56f
C19868 col_n[16] a_19030_13174# 0.251f
C19869 VDD a_8898_5142# 0.181f
C19870 row_n[3] a_33998_5142# 0.0437f
C19871 col_n[13] a_15926_3134# 0.0765f
C19872 rowon_n[7] a_33086_9158# 0.248f
C19873 a_6982_17190# a_7286_17230# 0.0931f
C19874 a_2275_17214# a_13006_17190# 0.399f
C19875 a_7894_17190# a_8386_17552# 0.0658f
C19876 col_n[23] a_25966_15182# 0.0765f
C19877 rowoff_n[6] a_22954_8154# 0.202f
C19878 col[17] a_2275_9182# 0.0899f
C19879 a_2475_5166# a_27062_5142# 0.316f
C19880 a_14010_5142# a_15014_5142# 0.843f
C19881 m2_34864_7974# a_2275_8178# 0.278f
C19882 m3_7888_1078# m3_8892_1078# 0.202f
C19883 vcm a_3878_9158# 0.1f
C19884 rowoff_n[15] a_33086_17190# 0.294f
C19885 m2_31276_16434# a_31078_16186# 0.165f
C19886 rowoff_n[4] a_31990_6146# 0.202f
C19887 col_n[7] a_10394_11528# 0.0283f
C19888 ctop a_15014_4138# 4.11f
C19889 m2_7756_946# a_7986_1126# 0.0249f
C19890 m3_9896_1078# a_9994_2130# 0.0302f
C19891 a_2475_14202# a_5886_14178# 0.264f
C19892 a_2275_14202# a_3270_14218# 0.144f
C19893 VDD a_23958_9158# 0.181f
C19894 row_n[7] a_10998_9158# 0.282f
C19895 rowon_n[11] a_10906_13174# 0.118f
C19896 VDD a_11302_18234# 0.019f
C19897 a_2275_2154# a_18026_2130# 0.399f
C19898 m2_12776_946# VDD 1f
C19899 vcm a_29982_4138# 0.1f
C19900 a_4974_7150# a_4974_6146# 0.843f
C19901 rowoff_n[9] a_23446_11528# 0.0133f
C19902 rowon_n[1] a_20946_3134# 0.118f
C19903 col_n[2] a_2475_16210# 0.0531f
C19904 vcm a_17326_13214# 0.155f
C19905 col_n[7] a_2475_5166# 0.0531f
C19906 a_32994_12170# a_33390_12210# 0.0313f
C19907 VDD a_15414_3496# 0.0779f
C19908 m2_34864_12994# VDD 0.772f
C19909 ctop a_30074_8154# 4.11f
C19910 a_2475_16210# a_20946_16186# 0.264f
C19911 a_2275_16210# a_18330_16226# 0.144f
C19912 VDD a_4882_12170# 0.181f
C19913 col_n[5] a_7986_11166# 0.251f
C19914 col_n[2] a_4882_1126# 0.0765f
C19915 rowoff_n[7] a_32482_9520# 0.0133f
C19916 col_n[12] a_14922_13174# 0.0765f
C19917 a_2275_4162# a_33086_4138# 0.399f
C19918 a_17934_4138# a_18426_4500# 0.0658f
C19919 a_17022_4138# a_17326_4178# 0.0931f
C19920 m2_34864_6970# a_35002_7150# 0.225f
C19921 vcm a_10906_7150# 0.1f
C19922 a_29070_9158# a_30074_9158# 0.843f
C19923 rowoff_n[12] a_4974_14178# 0.294f
C19924 row_n[10] a_31990_12170# 0.0437f
C19925 m2_22240_14426# a_22042_14178# 0.165f
C19926 vcm a_32386_17230# 0.155f
C19927 rowon_n[14] a_31078_16186# 0.248f
C19928 a_2275_13198# a_11910_13174# 0.136f
C19929 VDD a_30474_7512# 0.0779f
C19930 col_n[27] row_n[8] 0.298f
C19931 col_n[26] rowon_n[7] 0.111f
C19932 col_n[8] ctop 0.0594f
C19933 col_n[24] rowon_n[6] 0.111f
C19934 col_n[11] row_n[0] 0.298f
C19935 col_n[1] col[1] 0.414f
C19936 col_n[25] row_n[7] 0.298f
C19937 col_n[13] row_n[1] 0.298f
C19938 col_n[30] rowon_n[9] 0.111f
C19939 col_n[14] rowon_n[1] 0.111f
C19940 col_n[17] row_n[3] 0.298f
C19941 col_n[12] rowon_n[0] 0.111f
C19942 col_n[22] rowon_n[5] 0.111f
C19943 VDD col[5] 3.83f
C19944 vcm col[2] 5.46f
C19945 col_n[19] row_n[4] 0.298f
C19946 ctop a_10998_11166# 4.11f
C19947 rowon_n[13] rowon_n[12] 0.0632f
C19948 col_n[31] row_n[10] 0.298f
C19949 col_n[18] rowon_n[3] 0.111f
C19950 col_n[21] row_n[5] 0.298f
C19951 col_n[15] row_n[2] 0.298f
C19952 col_n[16] rowon_n[2] 0.111f
C19953 col_n[23] row_n[6] 0.298f
C19954 col_n[20] rowon_n[4] 0.111f
C19955 col_n[28] rowon_n[8] 0.111f
C19956 col_n[29] row_n[9] 0.298f
C19957 a_2275_18218# a_33390_18234# 0.145f
C19958 a_18938_18194# a_19030_18194# 0.0991f
C19959 col_n[4] a_2275_8178# 0.113f
C19960 VDD a_19942_16186# 0.181f
C19961 a_13918_1126# a_14010_1126# 0.0991f
C19962 m2_19228_2378# a_19030_2130# 0.165f
C19963 col[25] a_28066_10162# 0.367f
C19964 vcm a_1957_1150# 0.139f
C19965 m2_25828_946# m2_26832_946# 0.843f
C19966 vcm a_25966_11166# 0.1f
C19967 a_2475_10186# a_3970_10162# 0.316f
C19968 a_2275_10186# a_2966_10162# 0.399f
C19969 a_20034_11166# a_20034_10162# 0.843f
C19970 VDD a_22042_1126# 0.035f
C19971 row_n[14] a_8990_16186# 0.282f
C19972 col_n[24] a_2475_7174# 0.0531f
C19973 ctop a_2275_5166# 0.0683f
C19974 a_13918_15182# a_14314_15222# 0.0313f
C19975 a_2275_15206# a_26970_15182# 0.136f
C19976 VDD a_11398_10524# 0.0779f
C19977 m2_34864_13998# m3_34996_14130# 3.79f
C19978 ctop a_26058_15182# 4.11f
C19979 row_n[4] a_19030_6146# 0.282f
C19980 rowon_n[8] a_18938_10162# 0.118f
C19981 col_n[20] a_23350_10202# 0.084f
C19982 col[9] a_2475_15206# 0.136f
C19983 col[14] a_2475_4162# 0.136f
C19984 a_32994_8154# a_33486_8516# 0.0658f
C19985 rowoff_n[10] a_11398_12532# 0.0133f
C19986 a_32082_8154# a_32386_8194# 0.0931f
C19987 a_29374_1166# vcm 0.16f
C19988 m2_13204_12418# a_13006_12170# 0.165f
C19989 m2_4168_16434# rowon_n[14] 0.0322f
C19990 m2_10192_12418# rowon_n[10] 0.0322f
C19991 row_n[6] a_6282_8194# 0.0117f
C19992 vcm a_6890_14178# 0.1f
C19993 m2_16216_8402# rowon_n[6] 0.0322f
C19994 m2_22240_4386# rowon_n[2] 0.0322f
C19995 a_2475_12194# a_19030_12170# 0.316f
C19996 a_9994_12170# a_10998_12170# 0.843f
C19997 VDD a_2874_4138# 0.182f
C19998 col_n[31] a_34490_4500# 0.0283f
C19999 m2_32280_18442# VDD 0.0456f
C20000 VDD a_26458_14540# 0.0779f
C20001 col_n[28] rowoff_n[12] 0.0471f
C20002 col_n[21] a_2275_10186# 0.113f
C20003 rowoff_n[0] a_2966_2130# 0.0136f
C20004 a_28978_5142# a_29070_5142# 0.326f
C20005 m2_32280_8402# a_32082_8154# 0.165f
C20006 a_2275_9182# a_9994_9158# 0.399f
C20007 col[14] a_17022_8154# 0.367f
C20008 rowoff_n[14] a_27462_16548# 0.0133f
C20009 rowon_n[2] a_5978_4138# 0.248f
C20010 vcm a_21950_18194# 0.101f
C20011 col[6] a_2275_18218# 0.0899f
C20012 m2_31276_17438# rowon_n[15] 0.0322f
C20013 col[21] a_23958_10162# 0.0682f
C20014 a_2475_14202# a_34090_14178# 0.316f
C20015 VDD a_18026_8154# 0.483f
C20016 col[11] a_2275_7174# 0.0899f
C20017 m2_31852_946# vcm 0.353f
C20018 col_n[29] a_32082_4138# 0.251f
C20019 VDD a_7382_17552# 0.0779f
C20020 a_23958_2130# a_24354_2170# 0.0313f
C20021 m3_5880_1078# VDD 0.0157f
C20022 vcm a_24050_3134# 0.56f
C20023 col[26] a_2475_17214# 0.136f
C20024 col_n[9] a_12306_8194# 0.084f
C20025 m2_4168_10410# a_3970_10162# 0.165f
C20026 col[31] a_2475_6170# 0.136f
C20027 rowoff_n[3] a_3970_5142# 0.294f
C20028 a_13918_11166# a_14410_11528# 0.0658f
C20029 a_13006_11166# a_13310_11206# 0.0931f
C20030 a_2275_11190# a_25054_11166# 0.399f
C20031 row_n[11] a_17022_13174# 0.282f
C20032 a_25054_16186# a_26058_16186# 0.843f
C20033 VDD a_33086_12170# 0.483f
C20034 m2_23820_18014# m3_23952_18146# 3.79f
C20035 col_n[12] rowoff_n[13] 0.0471f
C20036 col_n[20] a_23446_2492# 0.0283f
C20037 rowon_n[15] a_16930_17190# 0.118f
C20038 col_n[30] a_33486_14540# 0.0283f
C20039 col_n[1] a_2475_3158# 0.0531f
C20040 col[10] rowoff_n[4] 0.0901f
C20041 col[8] rowoff_n[2] 0.0901f
C20042 col[13] rowoff_n[7] 0.0901f
C20043 col[7] rowoff_n[1] 0.0901f
C20044 col[11] rowoff_n[5] 0.0901f
C20045 rowoff_n[1] a_13006_3134# 0.294f
C20046 col[15] rowoff_n[9] 0.0901f
C20047 col[14] rowoff_n[8] 0.0901f
C20048 col[6] rowoff_n[0] 0.0901f
C20049 col[9] rowoff_n[3] 0.0901f
C20050 col[12] rowoff_n[6] 0.0901f
C20051 row_n[1] a_27062_3134# 0.282f
C20052 m2_23244_6394# a_23046_6146# 0.165f
C20053 row_n[13] a_4274_15222# 0.0117f
C20054 vcm a_4974_6146# 0.56f
C20055 rowon_n[5] a_26970_7150# 0.118f
C20056 a_9902_8154# a_9994_8154# 0.326f
C20057 a_2475_8178# a_17934_8154# 0.264f
C20058 a_2275_8178# a_15318_8194# 0.144f
C20059 rowoff_n[12] a_33998_14178# 0.202f
C20060 col[3] a_5978_6146# 0.367f
C20061 row_n[3] a_14314_5182# 0.0117f
C20062 col[28] a_2275_9182# 0.0899f
C20063 VDD a_14010_15182# 0.483f
C20064 col[10] a_12914_8154# 0.0682f
C20065 col_n[18] a_21038_2130# 0.251f
C20066 a_2275_5166# a_8898_5142# 0.136f
C20067 row_n[5] a_4882_7150# 0.0437f
C20068 a_4882_5142# a_5278_5182# 0.0313f
C20069 col_n[28] a_31078_14178# 0.251f
C20070 m2_27836_946# m3_26964_1078# 0.0341f
C20071 m3_34996_16138# m3_34996_15134# 0.202f
C20072 rowon_n[9] a_3970_11166# 0.248f
C20073 col_n[25] a_27974_4138# 0.0765f
C20074 vcm a_20034_10162# 0.56f
C20075 a_2475_10186# a_32994_10162# 0.264f
C20076 rowoff_n[15] a_15414_17552# 0.0133f
C20077 a_2275_10186# a_30378_10202# 0.144f
C20078 a_28066_15182# a_28370_15222# 0.0931f
C20079 col_n[8] a_11302_18234# 0.084f
C20080 a_28978_15182# a_29470_15544# 0.0658f
C20081 m2_20808_18014# ctop 0.0422f
C20082 m2_34864_10986# m3_34996_11118# 3.79f
C20083 col[1] a_3878_6146# 0.0682f
C20084 m2_3164_15430# row_n[13] 0.0128f
C20085 col_n[13] a_2475_16210# 0.0531f
C20086 m2_9188_11414# row_n[9] 0.0128f
C20087 m2_15212_7398# row_n[5] 0.0128f
C20088 m2_14208_4386# a_14010_4138# 0.165f
C20089 col_n[18] a_2475_5166# 0.0531f
C20090 m2_21236_3382# row_n[1] 0.0128f
C20091 col_n[19] a_22442_12532# 0.0283f
C20092 vcm a_10298_4178# 0.155f
C20093 a_2275_7174# a_23958_7150# 0.136f
C20094 rowon_n[1] a_2275_3158# 1.79f
C20095 rowoff_n[9] a_5886_11166# 0.202f
C20096 vcm a_35094_14178# 0.165f
C20097 a_24962_12170# a_25054_12170# 0.326f
C20098 VDD a_31990_4138# 0.181f
C20099 a_1957_16210# a_2161_16210# 0.115f
C20100 a_2475_16210# a_2275_16210# 2.76f
C20101 col[3] a_2475_13198# 0.136f
C20102 col[8] a_2475_2154# 0.136f
C20103 row_n[8] a_25054_10162# 0.282f
C20104 rowoff_n[7] a_14922_9158# 0.202f
C20105 col[2] a_4974_16186# 0.367f
C20106 rowon_n[12] a_24962_14178# 0.118f
C20107 a_2475_4162# a_16018_4138# 0.316f
C20108 a_26058_5142# a_26058_4138# 0.843f
C20109 m3_1864_10114# ctop 0.21f
C20110 col[9] a_11910_18194# 0.0682f
C20111 m2_30272_16434# row_n[14] 0.0128f
C20112 vcm a_25358_8194# 0.155f
C20113 m2_35292_12418# row_n[10] 0.0128f
C20114 a_19942_9158# a_20338_9198# 0.0313f
C20115 rowoff_n[13] a_21950_15182# 0.202f
C20116 row_n[10] a_12306_12210# 0.0117f
C20117 col_n[17] a_20034_12170# 0.251f
C20118 col_n[29] rowon_n[3] 0.111f
C20119 col_n[31] rowon_n[4] 0.111f
C20120 col_n[25] rowon_n[1] 0.111f
C20121 col_n[26] row_n[2] 0.298f
C20122 rowon_n[2] a_35002_4138# 0.118f
C20123 vcm col[13] 5.46f
C20124 rowon_n[10] row_n[10] 18.9f
C20125 col_n[16] en_bit_n[2] 0.187f
C20126 VDD col[16] 3.83f
C20127 col_n[27] rowon_n[2] 0.111f
C20128 col_n[6] col[7] 7.13f
C20129 col_n[19] ctop 0.0594f
C20130 col_n[30] row_n[4] 0.298f
C20131 col_n[22] row_n[0] 0.298f
C20132 col_n[23] rowon_n[0] 0.111f
C20133 col_n[28] row_n[3] 0.298f
C20134 col_n[24] row_n[1] 0.298f
C20135 ctop a_3970_2130# 4.03f
C20136 col_n[14] a_16930_2130# 0.0765f
C20137 vcm a_16018_17190# 0.56f
C20138 col_n[15] a_2275_8178# 0.113f
C20139 VDD a_12914_7150# 0.181f
C20140 rowoff_n[5] a_23958_7150# 0.202f
C20141 col_n[24] a_26970_14178# 0.0765f
C20142 a_2275_18218# a_17022_18194# 0.0924f
C20143 a_9902_18194# a_10394_18556# 0.0658f
C20144 VDD a_35398_17230# 0.0882f
C20145 row_n[0] a_22346_2170# 0.0117f
C20146 a_4882_1126# a_5374_1488# 0.0658f
C20147 row_n[12] a_2161_14202# 0.0221f
C20148 a_3970_1126# a_4274_1166# 0.0997f
C20149 a_2275_1150# a_6982_1126# 0.0924f
C20150 vcm a_18938_2130# 0.1f
C20151 a_2475_6170# a_31078_6146# 0.316f
C20152 a_16018_6146# a_17022_6146# 0.843f
C20153 col[0] a_2275_16210# 0.099f
C20154 m2_6752_946# m2_7180_1374# 0.165f
C20155 col[5] a_2275_5166# 0.0899f
C20156 row_n[2] a_12914_4138# 0.0437f
C20157 rowoff_n[3] a_32994_5142# 0.202f
C20158 vcm a_6282_11206# 0.155f
C20159 col_n[8] a_11398_10524# 0.0283f
C20160 VDD a_4370_1488# 0.0913f
C20161 rowon_n[6] a_12002_8154# 0.248f
C20162 ctop a_19030_6146# 4.11f
C20163 a_5886_15182# a_5978_15182# 0.326f
C20164 a_2475_15206# a_9902_15182# 0.264f
C20165 a_2275_15206# a_7286_15222# 0.144f
C20166 VDD a_27974_11166# 0.181f
C20167 m2_1732_15002# m3_1864_14130# 0.0341f
C20168 col[20] a_2475_15206# 0.136f
C20169 col[25] a_2475_4162# 0.136f
C20170 a_2275_3158# a_22042_3134# 0.399f
C20171 a_2475_18218# a_15014_18194# 0.0299f
C20172 rowoff_n[8] a_24450_10524# 0.0133f
C20173 vcm a_33998_6146# 0.1f
C20174 a_6982_8154# a_6982_7150# 0.843f
C20175 vcm a_21342_15222# 0.155f
C20176 VDD a_19430_5504# 0.0779f
C20177 a_31382_1166# VDD 0.0149f
C20178 col_n[6] a_8990_10162# 0.251f
C20179 row_n[12] rowoff_n[12] 0.209f
C20180 row_n[15] a_23046_17190# 0.282f
C20181 ctop a_34090_10162# 4.06f
C20182 a_2275_17214# a_22346_17230# 0.144f
C20183 a_2475_17214# a_24962_17190# 0.264f
C20184 rowoff_n[6] a_33486_8516# 0.0133f
C20185 VDD a_8898_14178# 0.181f
C20186 m2_27836_946# col_n[25] 0.338f
C20187 col_n[13] a_15926_12170# 0.0765f
C20188 m3_29976_18146# a_30074_17190# 0.0303f
C20189 a_19030_5142# a_19334_5182# 0.0931f
C20190 row_n[5] a_33086_7150# 0.282f
C20191 a_19942_5142# a_20434_5504# 0.0658f
C20192 col[17] a_2275_18218# 0.0899f
C20193 rowon_n[9] a_32994_11166# 0.118f
C20194 vcm a_14922_9158# 0.1f
C20195 m2_25828_18014# col[23] 0.347f
C20196 rowoff_n[14] a_9902_16186# 0.202f
C20197 a_31078_10162# a_32082_10162# 0.843f
C20198 col[22] a_2275_7174# 0.0899f
C20199 vcm a_3878_18194# 0.101f
C20200 m2_13780_946# a_14314_1166# 0.087f
C20201 a_2275_14202# a_15926_14178# 0.136f
C20202 row_n[7] a_20338_9198# 0.0117f
C20203 VDD a_34490_9520# 0.0779f
C20204 m2_34864_7974# m3_34996_8106# 3.79f
C20205 ctop a_15014_13174# 4.11f
C20206 a_24450_1488# col_n[21] 0.0283f
C20207 VDD a_23958_18194# 0.343f
C20208 a_2275_2154# a_27366_2170# 0.144f
C20209 col[26] a_29070_9158# 0.367f
C20210 a_2475_2154# a_29982_2130# 0.264f
C20211 a_15926_2130# a_16018_2130# 0.326f
C20212 m2_1732_2954# a_2275_3158# 0.191f
C20213 m3_1864_18146# VDD 0.0306f
C20214 row_n[9] a_10906_11166# 0.0437f
C20215 rowoff_n[9] a_34090_11166# 0.294f
C20216 m2_34864_13998# vcm 0.408f
C20217 rowon_n[13] a_9994_15182# 0.248f
C20218 vcm a_29982_13174# 0.1f
C20219 a_22042_12170# a_22042_11166# 0.843f
C20220 a_2475_11190# a_7986_11166# 0.316f
C20221 col_n[23] rowoff_n[13] 0.0471f
C20222 VDD a_26058_3134# 0.483f
C20223 col_n[7] a_2475_14202# 0.0531f
C20224 a_2275_16210# a_30986_16186# 0.136f
C20225 a_15926_16186# a_16322_16226# 0.0313f
C20226 VDD a_15414_12532# 0.0779f
C20227 rowon_n[3] a_20034_5142# 0.248f
C20228 col_n[12] a_2475_3158# 0.0531f
C20229 a_35398_1166# m2_34864_946# 0.087f
C20230 col[17] rowoff_n[0] 0.0901f
C20231 col[20] rowoff_n[3] 0.0901f
C20232 col[24] rowoff_n[7] 0.0901f
C20233 col[21] rowoff_n[4] 0.0901f
C20234 col[23] rowoff_n[6] 0.0901f
C20235 col[18] rowoff_n[1] 0.0901f
C20236 col[22] rowoff_n[5] 0.0901f
C20237 col[19] rowoff_n[2] 0.0901f
C20238 col[25] rowoff_n[8] 0.0901f
C20239 col[26] rowoff_n[9] 0.0901f
C20240 ctop a_30074_17190# 4.06f
C20241 col_n[21] a_24354_9198# 0.084f
C20242 m3_34996_15134# a_34090_15182# 0.0303f
C20243 m2_5172_6394# rowon_n[4] 0.0322f
C20244 m2_10192_2378# rowon_n[0] 0.0322f
C20245 col_n[2] a_4882_10162# 0.0765f
C20246 col[3] a_2475_18218# 0.136f
C20247 a_35002_9158# a_35494_9520# 0.0658f
C20248 vcm a_10906_16186# 0.1f
C20249 a_2475_13198# a_23046_13174# 0.316f
C20250 a_12002_13174# a_13006_13174# 0.843f
C20251 VDD a_6982_6146# 0.483f
C20252 VDD a_30474_16548# 0.0779f
C20253 row_n[12] a_31078_14178# 0.282f
C20254 col_n[4] a_2275_17214# 0.113f
C20255 m2_20232_15430# rowon_n[13] 0.0322f
C20256 vcm a_13006_1126# 0.165f
C20257 a_30986_6146# a_31078_6146# 0.326f
C20258 m2_26256_11414# rowon_n[9] 0.0322f
C20259 col_n[9] a_2275_6170# 0.113f
C20260 m2_32280_7398# rowon_n[5] 0.0322f
C20261 col[15] a_18026_7150# 0.367f
C20262 m3_3872_18146# m3_4876_18146# 0.202f
C20263 vcm a_1957_10186# 0.139f
C20264 col_n[7] rowoff_n[14] 0.0471f
C20265 a_2275_10186# a_14010_10162# 0.399f
C20266 col[22] a_24962_9158# 0.0682f
C20267 row_n[14] a_18330_16226# 0.0117f
C20268 m2_6752_946# a_6982_2130# 0.843f
C20269 col[10] rowoff_n[10] 0.0901f
C20270 VDD a_22042_10162# 0.483f
C20271 col_n[30] a_33086_3134# 0.251f
C20272 col_n[24] a_2475_16210# 0.0531f
C20273 m2_1732_11990# m3_1864_11118# 0.0341f
C20274 ctop a_2275_14202# 0.0683f
C20275 row_n[4] a_28370_6186# 0.0117f
C20276 col_n[29] a_2475_5166# 0.0531f
C20277 a_25966_3134# a_26362_3174# 0.0313f
C20278 m2_34864_4962# a_34090_5142# 0.843f
C20279 col_n[10] a_13310_7190# 0.084f
C20280 vcm a_28066_5142# 0.56f
C20281 rowoff_n[2] a_4974_4138# 0.294f
C20282 a_2475_7174# a_6890_7150# 0.264f
C20283 a_2275_7174# a_4274_7190# 0.144f
C20284 rowoff_n[10] a_22042_12170# 0.294f
C20285 row_n[6] a_18938_8154# 0.0437f
C20286 m2_1732_4962# sample 0.2f
C20287 col[14] a_2475_13198# 0.136f
C20288 a_15014_12170# a_15318_12210# 0.0931f
C20289 a_2275_12194# a_29070_12170# 0.399f
C20290 a_15926_12170# a_16418_12532# 0.0658f
C20291 rowon_n[10] a_18026_12170# 0.248f
C20292 col[19] a_2475_2154# 0.136f
C20293 m2_1732_16006# VDD 0.856f
C20294 row_n[0] m2_26256_2378# 0.0128f
C20295 a_27062_17190# a_28066_17190# 0.843f
C20296 VDD a_2874_13174# 0.182f
C20297 col_n[31] a_34490_13536# 0.0283f
C20298 rowon_n[0] a_28066_2130# 0.248f
C20299 rowoff_n[0] a_14010_2130# 0.294f
C20300 col_n[31] sw_n 0.418f
C20301 vcm col[24] 5.46f
C20302 col_n[30] ctop 0.0675f
C20303 VDD col[27] 3.83f
C20304 col_n[12] col[12] 0.489f
C20305 col_n[26] a_2275_8178# 0.113f
C20306 vcm a_8990_8154# 0.56f
C20307 rowoff_n[13] a_3878_15182# 0.202f
C20308 a_2275_9182# a_19334_9198# 0.144f
C20309 a_2475_9182# a_21950_9158# 0.264f
C20310 a_11910_9158# a_12002_9158# 0.326f
C20311 col[4] a_6982_5142# 0.367f
C20312 m2_28264_15430# a_28066_15182# 0.165f
C20313 ctop rowoff_n[11] 0.177f
C20314 col[14] a_17022_17190# 0.367f
C20315 m2_34864_4962# m3_34996_5094# 3.79f
C20316 col[11] a_13918_7150# 0.0682f
C20317 row_n[0] a_5978_2130# 0.282f
C20318 VDD a_18026_17190# 0.484f
C20319 col[11] a_2275_16210# 0.0899f
C20320 rowon_n[4] a_5886_6146# 0.118f
C20321 col_n[29] a_32082_13174# 0.251f
C20322 col[16] a_2275_5166# 0.0899f
C20323 col_n[26] a_28978_3134# 0.0765f
C20324 vcm a_33390_3174# 0.155f
C20325 a_2275_6170# a_12914_6146# 0.136f
C20326 a_6890_6146# a_7286_6186# 0.0313f
C20327 vcm a_24050_12170# 0.56f
C20328 a_2275_11190# a_35398_11206# 0.145f
C20329 VDD a_20946_2130# 0.181f
C20330 col_n[9] a_12306_17230# 0.084f
C20331 col[31] a_2475_15206# 0.136f
C20332 m2_4168_5390# row_n[3] 0.0128f
C20333 row_n[11] a_26362_13214# 0.0117f
C20334 a_30986_16186# a_31478_16548# 0.0658f
C20335 a_30074_16186# a_30378_16226# 0.0931f
C20336 col_n[20] a_23446_11528# 0.0283f
C20337 a_2475_3158# a_4974_3134# 0.316f
C20338 rowoff_n[8] a_6890_10162# 0.202f
C20339 row_n[13] a_16930_15182# 0.0437f
C20340 vcm a_14314_6186# 0.155f
C20341 rowoff_n[11] a_9994_13174# 0.294f
C20342 col_n[1] a_2475_12194# 0.0531f
C20343 a_2275_8178# a_27974_8154# 0.136f
C20344 m2_19228_13422# a_19030_13174# 0.165f
C20345 col_n[6] a_2475_1150# 0.0531f
C20346 vcm a_4974_15182# 0.56f
C20347 a_26970_13174# a_27062_13174# 0.326f
C20348 row_n[3] a_26970_5142# 0.0437f
C20349 rowon_n[7] a_26058_9158# 0.248f
C20350 m2_19228_14426# row_n[12] 0.0128f
C20351 a_2275_17214# a_5978_17190# 0.399f
C20352 col[3] a_5978_15182# 0.367f
C20353 m2_25252_10410# row_n[8] 0.0128f
C20354 rowoff_n[6] a_15926_8154# 0.202f
C20355 m2_31276_6394# row_n[4] 0.0128f
C20356 col[28] a_2275_18218# 0.0899f
C20357 col[10] a_12914_17190# 0.0682f
C20358 a_2475_5166# a_20034_5142# 0.316f
C20359 a_28066_6146# a_28066_5142# 0.843f
C20360 col_n[18] a_21038_11166# 0.251f
C20361 vcm a_29374_10202# 0.155f
C20362 col_n[15] a_17934_1126# 0.0785f
C20363 a_21950_10162# a_22346_10202# 0.0313f
C20364 rowoff_n[15] a_26058_17190# 0.294f
C20365 rowoff_n[4] a_24962_6146# 0.202f
C20366 col_n[25] a_27974_13174# 0.0765f
C20367 ctop a_7986_4138# 4.11f
C20368 m2_5748_946# a_2475_1150# 0.286f
C20369 row_n[7] a_3970_9158# 0.282f
C20370 VDD a_16930_9158# 0.181f
C20371 m2_1732_8978# m3_1864_8106# 0.0341f
C20372 col_n[3] a_2275_4162# 0.113f
C20373 VDD a_4274_18234# 0.019f
C20374 a_2275_2154# a_10998_2130# 0.399f
C20375 a_6890_2130# a_7382_2492# 0.0658f
C20376 a_5978_2130# a_6282_2170# 0.0931f
C20377 col[1] a_3878_15182# 0.0682f
C20378 vcm a_22954_4138# 0.1f
C20379 rowon_n[1] a_13918_3134# 0.118f
C20380 a_2475_7174# a_35094_7150# 0.0299f
C20381 a_18026_7150# a_19030_7150# 0.843f
C20382 rowoff_n[9] a_16418_11528# 0.0133f
C20383 rowoff_n[2] a_33998_4138# 0.202f
C20384 col_n[9] a_12402_9520# 0.0283f
C20385 m2_10192_11414# a_9994_11166# 0.165f
C20386 col_n[18] a_2475_14202# 0.0531f
C20387 vcm a_10298_13214# 0.155f
C20388 col_n[23] a_2475_3158# 0.0531f
C20389 VDD a_8386_3496# 0.0779f
C20390 col[30] rowoff_n[2] 0.0901f
C20391 col[28] rowoff_n[0] 0.0901f
C20392 sample_n rowoff_n[4] 0.14f
C20393 col[31] rowoff_n[3] 0.0901f
C20394 col[29] rowoff_n[1] 0.0901f
C20395 sw_n a_2275_1150# 0.0415f
C20396 ctop a_23046_8154# 4.11f
C20397 a_2275_16210# a_11302_16226# 0.144f
C20398 a_2475_16210# a_13918_16186# 0.264f
C20399 a_7894_16186# a_7986_16186# 0.326f
C20400 VDD a_31990_13174# 0.181f
C20401 rowon_n[3] a_1957_5166# 0.0172f
C20402 col[14] a_2475_18218# 0.136f
C20403 row_n[8] a_35398_10202# 0.0117f
C20404 rowoff_n[7] a_25454_9520# 0.0133f
C20405 a_2275_4162# a_26058_4138# 0.399f
C20406 m3_25960_1078# ctop 0.21f
C20407 col[8] a_2475_11190# 0.136f
C20408 m2_29268_7398# a_29070_7150# 0.165f
C20409 rowoff_n[13] a_32482_15544# 0.0133f
C20410 a_8990_9158# a_8990_8154# 0.843f
C20411 row_n[10] a_24962_12170# 0.0437f
C20412 vcm a_25358_17230# 0.155f
C20413 col_n[7] a_9994_9158# 0.251f
C20414 a_2966_13174# a_3970_13174# 0.843f
C20415 a_2275_13198# a_4882_13174# 0.136f
C20416 rowon_n[14] a_24050_16186# 0.248f
C20417 VDD a_23446_7512# 0.0779f
C20418 rowoff_n[5] a_34490_7512# 0.0133f
C20419 ctop a_3970_11166# 4.11f
C20420 col_n[14] a_16930_11166# 0.0765f
C20421 a_2275_18218# a_26362_18234# 0.145f
C20422 col_n[15] a_2275_17214# 0.113f
C20423 VDD a_12914_16186# 0.181f
C20424 row_n[0] a_35002_2130# 0.0437f
C20425 col_n[20] a_2275_6170# 0.113f
C20426 a_2475_1150# a_18938_1126# 0.285f
C20427 a_2275_1150# a_16322_1166# 0.145f
C20428 rowon_n[4] a_34090_6146# 0.248f
C20429 col_n[18] rowoff_n[14] 0.0471f
C20430 a_21950_6146# a_22442_6508# 0.0658f
C20431 a_21038_6146# a_21342_6186# 0.0931f
C20432 vcm a_18938_11166# 0.1f
C20433 col[21] rowoff_n[10] 0.0901f
C20434 a_33086_11166# a_34090_11166# 0.843f
C20435 row_n[14] a_2475_16210# 0.405f
C20436 VDD a_15014_1126# 0.035f
C20437 col[5] a_2275_14202# 0.0899f
C20438 a_2275_15206# a_19942_15182# 0.136f
C20439 col[10] a_2275_3158# 0.0899f
C20440 VDD a_4370_10524# 0.0779f
C20441 col_n[31] a_34394_10202# 0.084f
C20442 col[27] a_30074_8154# 0.367f
C20443 ctop a_19030_15182# 4.11f
C20444 row_n[4] a_12002_6146# 0.282f
C20445 a_2475_3158# a_33998_3134# 0.264f
C20446 a_17934_3134# a_18026_3134# 0.326f
C20447 rowon_n[8] a_11910_10162# 0.118f
C20448 a_2275_3158# a_31382_3174# 0.144f
C20449 rowoff_n[8] a_35094_10162# 0.0135f
C20450 m2_34864_12994# rowoff_n[11] 0.278f
C20451 m2_20232_5390# a_20034_5142# 0.165f
C20452 col[25] a_2475_13198# 0.136f
C20453 rowoff_n[10] a_4370_12532# 0.0133f
C20454 a_22346_1166# vcm 0.16f
C20455 col[30] a_2475_2154# 0.136f
C20456 vcm a_33998_15182# 0.1f
C20457 a_24050_13174# a_24050_12170# 0.843f
C20458 a_2475_12194# a_12002_12170# 0.316f
C20459 VDD a_30074_5142# 0.483f
C20460 m2_18224_18442# VDD 0.0456f
C20461 row_n[15] a_32386_17230# 0.0117f
C20462 col_n[22] a_25358_8194# 0.084f
C20463 a_2275_17214# a_35002_17190# 0.136f
C20464 a_17934_17190# a_18330_17230# 0.0313f
C20465 VDD a_19430_14540# 0.0779f
C20466 a_34090_2130# m2_34864_1950# 0.843f
C20467 col_n[17] col[18] 7.13f
C20468 row_n[15] col[2] 0.0342f
C20469 row_n[11] ctop 0.186f
C20470 col_n[2] rowoff_n[15] 0.0471f
C20471 rowon_n[15] col[3] 0.0323f
C20472 row_n[14] col[0] 0.0322f
C20473 rowon_n[14] col[1] 0.0323f
C20474 col_n[3] a_5886_9158# 0.0765f
C20475 col[5] rowoff_n[11] 0.0901f
C20476 a_2275_9182# a_2874_9158# 0.136f
C20477 a_2475_9182# a_3878_9158# 0.264f
C20478 rowoff_n[14] a_20434_16548# 0.0133f
C20479 vcm a_14922_18194# 0.101f
C20480 m2_3164_17438# rowon_n[15] 0.0322f
C20481 a_2475_14202# a_27062_14178# 0.316f
C20482 a_14010_14178# a_15014_14178# 0.843f
C20483 col[22] a_2275_16210# 0.0899f
C20484 m2_9188_13422# rowon_n[11] 0.0322f
C20485 VDD a_10998_8154# 0.483f
C20486 row_n[7] a_32994_9158# 0.0437f
C20487 m2_15212_9406# rowon_n[7] 0.0322f
C20488 m2_1732_5966# m3_1864_5094# 0.0341f
C20489 m2_21236_5390# rowon_n[3] 0.0322f
C20490 rowon_n[11] a_32082_13174# 0.248f
C20491 col[27] a_2275_5166# 0.0899f
C20492 VDD a_34490_18556# 0.0858f
C20493 m2_11196_3382# a_10998_3134# 0.165f
C20494 col[16] a_19030_6146# 0.367f
C20495 vcm a_17022_3134# 0.56f
C20496 a_32994_7150# a_33086_7150# 0.326f
C20497 col[23] a_25966_8154# 0.0682f
C20498 a_2275_11190# a_18026_11166# 0.399f
C20499 VDD a_2275_2154# 1.96f
C20500 col_n[31] a_34090_2130# 0.305f
C20501 m2_22816_18014# a_22954_18194# 0.225f
C20502 a_4974_16186# a_4974_15182# 0.843f
C20503 row_n[11] a_9994_13174# 0.282f
C20504 VDD a_26058_12170# 0.483f
C20505 m2_14784_18014# m3_13912_18146# 0.0341f
C20506 rowon_n[15] a_9902_17190# 0.118f
C20507 m2_35292_14426# rowon_n[12] 0.0322f
C20508 col_n[11] a_14314_6186# 0.084f
C20509 col_n[12] a_2475_12194# 0.0531f
C20510 a_27974_4138# a_28370_4178# 0.0313f
C20511 rowoff_n[1] a_5978_3134# 0.294f
C20512 col_n[21] a_24354_18234# 0.084f
C20513 row_n[1] a_20034_3134# 0.282f
C20514 col_n[17] a_2475_1150# 0.0486f
C20515 vcm a_32082_7150# 0.56f
C20516 rowon_n[5] a_19942_7150# 0.118f
C20517 a_2275_8178# a_8290_8194# 0.144f
C20518 rowoff_n[12] a_26970_14178# 0.202f
C20519 a_2475_8178# a_10906_8154# 0.264f
C20520 a_17934_13174# a_18426_13536# 0.0658f
C20521 a_2275_13198# a_33086_13174# 0.399f
C20522 a_17022_13174# a_17326_13214# 0.0931f
C20523 row_n[3] a_7286_5182# 0.0117f
C20524 col[2] a_2475_9182# 0.136f
C20525 VDD a_6982_15182# 0.483f
C20526 a_2475_5166# a_1957_5166# 0.0734f
C20527 m2_16792_946# m3_17928_1078# 0.0341f
C20528 col[5] a_7986_4138# 0.367f
C20529 vcm a_13006_10162# 0.56f
C20530 rowoff_n[15] a_8386_17552# 0.0133f
C20531 a_2475_10186# a_25966_10162# 0.264f
C20532 a_2275_10186# a_23350_10202# 0.144f
C20533 a_13918_10162# a_14010_10162# 0.326f
C20534 col[15] a_18026_16186# 0.367f
C20535 col_n[9] a_2275_15206# 0.113f
C20536 row_n[14] a_30986_16186# 0.0437f
C20537 col[12] a_14922_6146# 0.0682f
C20538 col_n[14] a_2275_4162# 0.113f
C20539 m2_6752_18014# ctop 0.0422f
C20540 col[22] a_24962_18194# 0.0682f
C20541 col_n[30] a_33086_12170# 0.251f
C20542 a_15014_3134# a_15014_2130# 0.843f
C20543 col_n[27] a_29982_2130# 0.0765f
C20544 col_n[29] a_2475_14202# 0.0531f
C20545 vcm a_3270_4178# 0.155f
C20546 a_2275_7174# a_16930_7150# 0.136f
C20547 a_8898_7150# a_9294_7190# 0.0313f
C20548 m2_1732_17010# vcm 0.316f
C20549 col_n[10] a_13310_16226# 0.084f
C20550 col[4] a_2275_1150# 0.0899f
C20551 vcm a_28066_14178# 0.56f
C20552 VDD a_24962_4138# 0.181f
C20553 col[25] a_2475_18218# 0.136f
C20554 a_32994_17190# a_33486_17552# 0.0658f
C20555 a_32082_17190# a_32386_17230# 0.0931f
C20556 col[19] a_2475_11190# 0.136f
C20557 col_n[21] a_24450_10524# 0.0283f
C20558 row_n[8] a_18026_10162# 0.282f
C20559 rowoff_n[7] a_7894_9158# 0.202f
C20560 rowon_n[12] a_17934_14178# 0.118f
C20561 a_2475_4162# a_8990_4138# 0.316f
C20562 a_4974_4138# a_5978_4138# 0.843f
C20563 m3_21944_18146# ctop 0.209f
C20564 m2_2160_16434# row_n[14] 0.0194f
C20565 vcm a_18330_8194# 0.155f
C20566 m2_8184_12418# row_n[10] 0.0128f
C20567 rowoff_n[13] a_14922_15182# 0.202f
C20568 m2_14208_8402# row_n[6] 0.0128f
C20569 a_2275_9182# a_31990_9158# 0.136f
C20570 m2_20232_4386# row_n[2] 0.0128f
C20571 sample a_2161_4162# 0.0858f
C20572 m2_1732_13998# a_2161_14202# 0.0454f
C20573 row_n[10] a_5278_12210# 0.0117f
C20574 rowon_n[2] a_27974_4138# 0.118f
C20575 ctop a_31078_3134# 4.11f
C20576 col_n[26] a_2275_17214# 0.113f
C20577 vcm a_8990_17190# 0.56f
C20578 a_28978_14178# a_29070_14178# 0.326f
C20579 VDD a_5886_7150# 0.181f
C20580 col[4] a_6982_14178# 0.367f
C20581 rowoff_n[5] a_16930_7150# 0.202f
C20582 col_n[31] a_2275_6170# 0.113f
C20583 m2_1732_2954# m3_1864_2082# 0.0341f
C20584 col_n[29] rowoff_n[14] 0.0471f
C20585 a_2275_18218# a_9994_18194# 0.0924f
C20586 row_n[0] a_15318_2170# 0.0117f
C20587 col[11] a_13918_16186# 0.0682f
C20588 vcm a_11910_2130# 0.1f
C20589 m2_34864_6970# m2_35292_7398# 0.165f
C20590 sample_n rowoff_n[10] 0.14f
C20591 col_n[19] a_22042_10162# 0.251f
C20592 a_30074_7150# a_30074_6146# 0.843f
C20593 a_2475_6170# a_24050_6146# 0.316f
C20594 col[16] a_2275_14202# 0.0899f
C20595 rowoff_n[3] a_25966_5142# 0.202f
C20596 row_n[2] a_5886_4138# 0.0437f
C20597 col_n[26] a_28978_12170# 0.0765f
C20598 vcm a_33390_12210# 0.155f
C20599 a_23958_11166# a_24354_11206# 0.0313f
C20600 col[21] a_2275_3158# 0.0899f
C20601 VDD a_31478_2492# 0.0779f
C20602 m2_29268_17438# row_n[15] 0.0128f
C20603 m2_34864_17010# a_2475_17214# 0.282f
C20604 m2_34864_12994# row_n[11] 0.267f
C20605 rowon_n[6] a_4974_8154# 0.248f
C20606 m2_18800_18014# a_19030_17190# 0.843f
C20607 ctop a_12002_6146# 4.11f
C20608 VDD a_20946_11166# 0.181f
C20609 a_2275_3158# a_15014_3134# 0.399f
C20610 a_7986_3134# a_8290_3174# 0.0931f
C20611 a_2475_18218# a_7986_18194# 0.0299f
C20612 a_8898_3134# a_9390_3496# 0.0658f
C20613 rowoff_n[8] a_17422_10524# 0.0133f
C20614 rowoff_n[1] a_35002_3134# 0.202f
C20615 m2_1732_13998# rowoff_n[12] 0.415f
C20616 a_28978_1126# a_2275_1150# 0.136f
C20617 col_n[10] a_13406_8516# 0.0283f
C20618 vcm a_26970_6146# 0.1f
C20619 a_20034_8154# a_21038_8154# 0.843f
C20620 vcm a_14314_15222# 0.155f
C20621 VDD a_12402_5504# 0.0779f
C20622 col_n[23] col[23] 0.489f
C20623 row_n[13] col[9] 0.0342f
C20624 rowon_n[12] col[8] 0.0323f
C20625 rowon_n[9] col[2] 0.0323f
C20626 row_n[9] col[1] 0.0342f
C20627 col_n[13] rowoff_n[15] 0.0471f
C20628 rowon_n[10] col[4] 0.0323f
C20629 row_n[10] col[3] 0.0342f
C20630 col_n[6] a_2475_10186# 0.0531f
C20631 rowon_n[14] col[12] 0.0323f
C20632 rowon_n[11] col[6] 0.0323f
C20633 rowon_n[15] col[14] 0.0323f
C20634 rowon_n[2] rowon_n[1] 0.0632f
C20635 rowon_n[5] ctop 0.203f
C20636 row_n[12] col[7] 0.0342f
C20637 a_24354_1166# VDD 0.0149f
C20638 rowon_n[13] col[10] 0.0323f
C20639 row_n[14] col[11] 0.0342f
C20640 rowon_n[8] col[0] 0.0318f
C20641 row_n[11] col[5] 0.0342f
C20642 row_n[15] col[13] 0.0342f
C20643 row_n[15] a_16018_17190# 0.282f
C20644 ctop a_27062_10162# 4.11f
C20645 a_2475_17214# a_17934_17190# 0.264f
C20646 a_2275_17214# a_15318_17230# 0.144f
C20647 a_9902_17190# a_9994_17190# 0.326f
C20648 rowoff_n[6] a_26458_8516# 0.0133f
C20649 col[16] rowoff_n[11] 0.0901f
C20650 row_n[5] a_26058_7150# 0.282f
C20651 a_2275_5166# a_30074_5142# 0.399f
C20652 rowon_n[9] a_25966_11166# 0.118f
C20653 a_29982_1126# a_30474_1488# 0.0658f
C20654 vcm a_7894_9158# 0.1f
C20655 a_10998_10162# a_10998_9158# 0.843f
C20656 rowoff_n[14] a_2161_16210# 0.0226f
C20657 col_n[8] a_10998_8154# 0.251f
C20658 m2_34288_16434# a_34090_16186# 0.165f
C20659 rowoff_n[4] a_35494_6508# 0.0133f
C20660 m2_28840_946# a_2475_1150# 0.286f
C20661 a_4882_14178# a_5278_14218# 0.0313f
C20662 a_2275_14202# a_8898_14178# 0.136f
C20663 col_n[15] a_17934_10162# 0.0765f
C20664 m3_12908_1078# a_13006_2130# 0.0302f
C20665 row_n[7] a_13310_9198# 0.0117f
C20666 VDD a_27462_9520# 0.0779f
C20667 ctop a_7986_13174# 4.11f
C20668 VDD a_16930_18194# 0.343f
C20669 a_2275_2154# a_20338_2170# 0.144f
C20670 a_2475_2154# a_22954_2130# 0.264f
C20671 col_n[3] a_2275_13198# 0.113f
C20672 m2_21812_946# VDD 1f
C20673 rowoff_n[9] a_27062_11166# 0.294f
C20674 col_n[8] a_2275_2154# 0.113f
C20675 a_23046_7150# a_23350_7190# 0.0931f
C20676 a_23958_7150# a_24450_7512# 0.0658f
C20677 rowon_n[13] a_2874_15182# 0.118f
C20678 vcm a_22954_13174# 0.1f
C20679 VDD a_19030_3134# 0.483f
C20680 col_n[9] a_12402_18556# 0.0283f
C20681 m2_26832_18014# a_2275_18218# 0.28f
C20682 col[28] a_31078_7150# 0.367f
C20683 a_2275_16210# a_23958_16186# 0.136f
C20684 rowon_n[3] a_13006_5142# 0.248f
C20685 m2_11772_946# col_n[9] 0.331f
C20686 VDD a_8386_12532# 0.0779f
C20687 col_n[23] a_2475_12194# 0.0531f
C20688 a_30074_1126# m2_29844_946# 0.0249f
C20689 col[0] rowoff_n[12] 0.0901f
C20690 ctop a_23046_17190# 4.06f
C20691 col_n[28] a_2475_1150# 0.0531f
C20692 a_19942_4138# a_20034_4138# 0.326f
C20693 a_2275_4162# a_2275_3158# 0.0715f
C20694 row_n[1] a_1957_3158# 0.187f
C20695 m2_3164_6394# a_2966_6146# 0.165f
C20696 m2_25252_14426# a_25054_14178# 0.165f
C20697 col[13] a_2475_9182# 0.136f
C20698 a_26058_14178# a_26058_13174# 0.843f
C20699 a_2475_13198# a_16018_13174# 0.316f
C20700 VDD a_34090_7150# 0.483f
C20701 col_n[23] a_26362_7190# 0.084f
C20702 a_19942_18194# a_20338_18234# 0.0313f
C20703 m2_22816_18014# a_2475_18218# 0.286f
C20704 VDD a_23446_16548# 0.0779f
C20705 col_n[4] a_6890_8154# 0.0765f
C20706 a_14922_1126# a_15318_1166# 0.0313f
C20707 row_n[12] a_24050_14178# 0.282f
C20708 a_30986_1126# col_n[28] 0.0772f
C20709 m2_4744_18014# col_n[2] 0.243f
C20710 vcm a_5978_1126# 0.165f
C20711 col_n[20] a_2275_15206# 0.113f
C20712 m2_4168_7398# rowon_n[5] 0.0322f
C20713 m2_10192_3382# rowon_n[1] 0.0322f
C20714 m2_29844_946# m2_30272_1374# 0.165f
C20715 col_n[25] a_2275_4162# 0.113f
C20716 row_n[2] a_34090_4138# 0.282f
C20717 a_4882_10162# a_5374_10524# 0.0658f
C20718 a_2275_10186# a_6982_10162# 0.399f
C20719 a_3970_10162# a_4274_10202# 0.0931f
C20720 row_n[14] a_11302_16226# 0.0117f
C20721 rowon_n[6] a_33998_8154# 0.118f
C20722 a_2475_15206# a_31078_15182# 0.316f
C20723 a_16018_15182# a_17022_15182# 0.843f
C20724 VDD a_15014_10162# 0.483f
C20725 row_n[4] a_21342_6186# 0.0117f
C20726 col[17] a_20034_5142# 0.367f
C20727 col[10] a_2275_12194# 0.0899f
C20728 col[15] a_2275_1150# 0.0899f
C20729 col[27] a_30074_17190# 0.367f
C20730 col[24] a_26970_7150# 0.0682f
C20731 vcm a_21038_5142# 0.56f
C20732 a_34090_8154# a_34394_8194# 0.0931f
C20733 a_35002_8154# a_35094_8154# 0.0991f
C20734 rowoff_n[10] a_15014_12170# 0.294f
C20735 a_33390_1166# vcm 0.16f
C20736 m2_16216_12418# a_16018_12170# 0.165f
C20737 m2_19228_16434# rowon_n[14] 0.0322f
C20738 m2_25252_12418# rowon_n[10] 0.0322f
C20739 row_n[6] a_11910_8154# 0.0437f
C20740 m2_31276_8402# rowon_n[6] 0.0322f
C20741 a_2275_12194# a_22042_12170# 0.399f
C20742 rowon_n[10] a_10998_12170# 0.248f
C20743 col[30] a_2475_11190# 0.136f
C20744 a_6982_17190# a_6982_16186# 0.843f
C20745 VDD a_30074_14178# 0.483f
C20746 col_n[12] a_15318_5182# 0.084f
C20747 rowon_n[0] a_21038_2130# 0.248f
C20748 rowoff_n[0] a_6982_2130# 0.294f
C20749 col_n[22] a_25358_17230# 0.084f
C20750 a_29982_5142# a_30378_5182# 0.0313f
C20751 m2_8760_946# ctop 0.0428f
C20752 col_n[3] a_5886_18194# 0.0762f
C20753 m2_34864_7974# a_35094_8154# 0.0249f
C20754 vcm a_2475_8178# 1.08f
C20755 a_2475_9182# a_14922_9158# 0.264f
C20756 rowoff_n[14] a_31078_16186# 0.294f
C20757 a_2275_9182# a_12306_9198# 0.144f
C20758 a_19030_14178# a_19334_14218# 0.0931f
C20759 a_19942_14178# a_20434_14540# 0.0658f
C20760 VDD a_10998_17190# 0.484f
C20761 a_26058_2130# a_27062_2130# 0.843f
C20762 col[27] a_2275_14202# 0.0899f
C20763 m3_20940_1078# VDD 0.0157f
C20764 col[6] a_8990_3134# 0.367f
C20765 vcm a_26362_3174# 0.155f
C20766 row_n[9] a_32082_11166# 0.282f
C20767 a_2275_6170# a_5886_6146# 0.136f
C20768 m2_7180_10410# a_6982_10162# 0.165f
C20769 rowon_n[13] a_31990_15182# 0.118f
C20770 col[16] a_19030_15182# 0.367f
C20771 vcm a_17022_12170# 0.56f
C20772 col[13] a_15926_5142# 0.0682f
C20773 a_2475_11190# a_29982_11166# 0.264f
C20774 a_2275_11190# a_27366_11206# 0.144f
C20775 a_15926_11166# a_16018_11166# 0.326f
C20776 VDD a_13918_2130# 0.181f
C20777 col[23] a_25966_17190# 0.0682f
C20778 row_n[11] a_19334_13214# 0.0117f
C20779 VDD a_2275_11190# 1.96f
C20780 col_n[31] a_34090_11166# 0.251f
C20781 m2_28840_18014# m3_28972_18146# 3.79f
C20782 a_17022_4138# a_17022_3134# 0.843f
C20783 col_n[1] a_4274_3174# 0.084f
C20784 row_n[1] a_29374_3174# 0.0117f
C20785 m2_26256_6394# a_26058_6146# 0.165f
C20786 row_n[13] a_9902_15182# 0.0437f
C20787 col_n[11] a_14314_15222# 0.084f
C20788 vcm a_7286_6186# 0.155f
C20789 rowoff_n[11] a_2874_13174# 0.202f
C20790 a_10906_8154# a_11302_8194# 0.0313f
C20791 a_2275_8178# a_20946_8154# 0.136f
C20792 rowon_n[9] col[13] 0.0323f
C20793 rowon_n[5] col[5] 0.0323f
C20794 rowon_n[7] col[9] 0.0323f
C20795 rowon_n[12] col[19] 0.0323f
C20796 row_n[9] col[12] 0.0342f
C20797 row_n[14] col[22] 0.0342f
C20798 rowon_n[6] col[7] 0.0323f
C20799 row_n[6] col[6] 0.0342f
C20800 row_n[12] col[18] 0.0342f
C20801 rowon_n[10] col[15] 0.0323f
C20802 rowon_n[13] col[21] 0.0323f
C20803 rowon_n[14] col[23] 0.0323f
C20804 row_n[10] col[14] 0.0342f
C20805 row_n[5] col[4] 0.0342f
C20806 row_n[13] col[20] 0.0342f
C20807 rowon_n[3] col[1] 0.0323f
C20808 row_n[8] col[10] 0.0342f
C20809 row_n[4] col[2] 0.0342f
C20810 col_n[28] col[29] 7.1f
C20811 row_n[15] col[24] 0.0342f
C20812 row_n[11] col[16] 0.0342f
C20813 row_n[3] col[0] 0.0322f
C20814 rowon_n[11] col[17] 0.0323f
C20815 rowon_n[15] col[25] 0.0323f
C20816 row_n[0] ctop 0.181f
C20817 col_n[24] rowoff_n[15] 0.0471f
C20818 rowon_n[8] col[11] 0.0323f
C20819 sw sw_n 0.23f
C20820 row_n[7] col[8] 0.0342f
C20821 rowon_n[4] col[3] 0.0323f
C20822 col_n[17] a_2475_10186# 0.0531f
C20823 ctop a_20034_1126# 0.561f
C20824 vcm a_32082_16186# 0.56f
C20825 VDD a_28978_6146# 0.181f
C20826 row_n[3] a_19942_5142# 0.0437f
C20827 col[27] rowoff_n[11] 0.0901f
C20828 rowon_n[7] a_19030_9158# 0.248f
C20829 col_n[22] a_25454_9520# 0.0283f
C20830 a_35002_18194# a_35494_18556# 0.0658f
C20831 rowoff_n[6] a_8898_8154# 0.202f
C20832 m2_3164_6394# row_n[4] 0.0128f
C20833 m2_8184_2378# row_n[0] 0.0128f
C20834 col[7] a_2475_7174# 0.136f
C20835 a_2475_5166# a_13006_5142# 0.316f
C20836 a_6982_5142# a_7986_5142# 0.843f
C20837 m2_32856_946# m3_31984_1078# 0.0341f
C20838 col_n[0] a_3366_3496# 0.0283f
C20839 vcm a_22346_10202# 0.155f
C20840 rowoff_n[15] a_19030_17190# 0.294f
C20841 a_2275_10186# a_34394_10202# 0.144f
C20842 rowoff_n[4] a_17934_6146# 0.202f
C20843 col[5] a_7986_13174# 0.367f
C20844 col[2] a_4882_3134# 0.0682f
C20845 a_30986_15182# a_31078_15182# 0.326f
C20846 VDD a_9902_9158# 0.181f
C20847 col[12] a_14922_15182# 0.0682f
C20848 col_n[14] a_2275_13198# 0.113f
C20849 col_n[19] a_2275_2154# 0.113f
C20850 col_n[20] a_23046_9158# 0.251f
C20851 m2_18224_15430# row_n[13] 0.0128f
C20852 a_2275_2154# a_3970_2130# 0.399f
C20853 m2_24248_11414# row_n[9] 0.0128f
C20854 m2_30272_7398# row_n[5] 0.0128f
C20855 m2_17220_4386# a_17022_4138# 0.165f
C20856 m2_35292_3382# row_n[1] 0.0128f
C20857 vcm a_15926_4138# 0.1f
C20858 a_2475_7174# a_28066_7150# 0.316f
C20859 col_n[27] a_29982_11166# 0.0765f
C20860 rowoff_n[9] a_9390_11528# 0.0133f
C20861 rowoff_n[2] a_26970_4138# 0.202f
C20862 rowon_n[1] a_6890_3134# 0.118f
C20863 a_32082_8154# a_32082_7150# 0.843f
C20864 vcm a_3270_13214# 0.155f
C20865 a_25966_12170# a_26362_12210# 0.0313f
C20866 VDD a_35494_4500# 0.106f
C20867 col[11] rowoff_n[12] 0.0901f
C20868 col[4] a_2275_10186# 0.0899f
C20869 ctop a_16018_8154# 4.11f
C20870 a_2275_16210# a_4274_16226# 0.144f
C20871 a_2475_16210# a_6890_16186# 0.264f
C20872 VDD a_24962_13174# 0.181f
C20873 row_n[8] a_27366_10202# 0.0117f
C20874 m2_2736_1950# m2_2736_946# 0.843f
C20875 rowoff_n[7] a_18426_9520# 0.0133f
C20876 col_n[11] a_14410_7512# 0.0283f
C20877 a_2275_4162# a_19030_4138# 0.399f
C20878 a_9994_4138# a_10298_4178# 0.0931f
C20879 a_10906_4138# a_11398_4500# 0.0658f
C20880 m3_34996_3086# ctop 0.209f
C20881 col[24] a_2475_9182# 0.136f
C20882 vcm a_30986_8154# 0.1f
C20883 a_22042_9158# a_23046_9158# 0.843f
C20884 rowoff_n[13] a_25454_15544# 0.0133f
C20885 row_n[10] a_17934_12170# 0.0437f
C20886 vcm a_18330_17230# 0.155f
C20887 rowon_n[14] a_17022_16186# 0.248f
C20888 VDD a_16418_7512# 0.0779f
C20889 rowoff_n[5] a_27462_7512# 0.0133f
C20890 sample a_2161_13198# 0.0858f
C20891 ctop a_31078_12170# 4.11f
C20892 a_2275_18218# a_19334_18234# 0.145f
C20893 a_11910_18194# a_12002_18194# 0.0991f
C20894 row_n[0] a_27974_2130# 0.0437f
C20895 VDD a_5886_16186# 0.181f
C20896 col_n[31] a_2275_15206# 0.113f
C20897 a_2475_1150# a_11910_1126# 0.264f
C20898 a_2275_1150# a_9294_1166# 0.145f
C20899 a_6890_1126# a_6982_1126# 0.0991f
C20900 rowon_n[4] a_27062_6146# 0.248f
C20901 a_2275_6170# a_34090_6146# 0.399f
C20902 col_n[9] a_12002_7150# 0.251f
C20903 vcm a_11910_11166# 0.1f
C20904 a_13006_11166# a_13006_10162# 0.843f
C20905 VDD a_7986_1126# 0.035f
C20906 col_n[16] a_18938_9158# 0.0765f
C20907 col[21] a_2275_12194# 0.0899f
C20908 a_6890_15182# a_7286_15222# 0.0313f
C20909 a_2275_15206# a_12914_15182# 0.136f
C20910 VDD a_31478_11528# 0.0779f
C20911 col[26] a_2275_1150# 0.0899f
C20912 ctop a_12002_15182# 4.11f
C20913 row_n[4] a_4974_6146# 0.282f
C20914 a_2475_3158# a_26970_3134# 0.264f
C20915 rowon_n[8] a_4882_10162# 0.118f
C20916 a_2275_3158# a_24354_3174# 0.144f
C20917 rowoff_n[8] a_28066_10162# 0.294f
C20918 vcm a_2966_5142# 0.56f
C20919 a_25054_8154# a_25358_8194# 0.0931f
C20920 rowoff_n[11] a_31990_13174# 0.202f
C20921 a_25966_8154# a_26458_8516# 0.0658f
C20922 col_n[10] a_13406_17552# 0.0283f
C20923 m2_1732_11990# a_2475_12194# 0.139f
C20924 vcm a_26970_15182# 0.1f
C20925 a_2475_12194# a_4974_12170# 0.316f
C20926 col[29] a_32082_6146# 0.367f
C20927 VDD a_23046_5142# 0.483f
C20928 m2_4168_18442# VDD 0.0456f
C20929 row_n[15] a_25358_17230# 0.0117f
C20930 a_2275_17214# a_27974_17190# 0.136f
C20931 VDD a_12402_14540# 0.0779f
C20932 rowon_n[0] a_2966_2130# 0.0141f
C20933 m3_32988_18146# a_33086_17190# 0.0303f
C20934 col_n[11] a_2475_8178# 0.0531f
C20935 a_21950_5142# a_22042_5142# 0.326f
C20936 rowoff_n[14] a_13406_16548# 0.0133f
C20937 col_n[24] a_27366_6186# 0.084f
C20938 vcm a_7894_18194# 0.101f
C20939 a_28066_15182# a_28066_14178# 0.843f
C20940 a_2475_14202# a_20034_14178# 0.316f
C20941 col_n[8] a_10998_17190# 0.251f
C20942 m2_16792_946# a_18026_1126# 0.843f
C20943 row_n[7] a_25966_9158# 0.0437f
C20944 VDD a_3970_8154# 0.483f
C20945 col_n[5] a_7894_7150# 0.0765f
C20946 col[1] a_2475_5166# 0.136f
C20947 rowon_n[11] a_25054_13174# 0.248f
C20948 VDD a_27462_18556# 0.0858f
C20949 a_16930_2130# a_17326_2170# 0.0313f
C20950 a_2275_2154# a_32994_2130# 0.136f
C20951 m3_16924_18146# VDD 0.0277f
C20952 vcm a_9994_3134# 0.56f
C20953 rowon_n[1] a_35094_3134# 0.0141f
C20954 a_2275_11190# a_10998_11166# 0.399f
C20955 a_6890_11166# a_7382_11528# 0.0658f
C20956 col_n[8] a_2275_11190# 0.113f
C20957 a_5978_11166# a_6282_11206# 0.0931f
C20958 m2_17796_18014# a_18026_18194# 0.0249f
C20959 row_n[11] a_2874_13174# 0.0436f
C20960 a_18026_16186# a_19030_16186# 0.843f
C20961 a_2475_16210# a_35094_16186# 0.0299f
C20962 VDD a_19030_12170# 0.483f
C20963 m2_4744_18014# m3_5880_18146# 0.0341f
C20964 col[18] a_21038_4138# 0.367f
C20965 rowon_n[15] a_2161_17214# 0.0177f
C20966 m2_8184_14426# rowon_n[12] 0.0322f
C20967 col[28] a_31078_16186# 0.367f
C20968 m2_14208_10410# rowon_n[8] 0.0322f
C20969 m2_20232_6394# rowon_n[4] 0.0322f
C20970 col[25] a_27974_6146# 0.0682f
C20971 rowon_n[11] col[28] 0.0323f
C20972 rowon_n[13] sample_n 0.0692f
C20973 rowon_n[5] col[16] 0.0323f
C20974 row_n[8] col[21] 0.0342f
C20975 row_n[11] col[27] 0.0342f
C20976 col_n[28] a_2475_10186# 0.0531f
C20977 rowon_n[9] col[24] 0.0323f
C20978 rowon_n[2] col[10] 0.0323f
C20979 row_n[0] col[5] 0.0342f
C20980 row_n[12] col[29] 0.0342f
C20981 row_n[2] col[9] 0.0342f
C20982 row_n[1] col[7] 0.0342f
C20983 rowon_n[0] col[6] 0.0323f
C20984 row_n[1] a_13006_3134# 0.282f
C20985 rowon_n[3] col[12] 0.0323f
C20986 row_n[5] col[15] 0.0342f
C20987 rowon_n[8] col[22] 0.0323f
C20988 row_n[4] col[13] 0.0342f
C20989 rowon_n[7] col[20] 0.0323f
C20990 rowon_n[12] col[30] 0.0323f
C20991 row_n[6] col[17] 0.0342f
C20992 rowon_n[10] col[26] 0.0323f
C20993 ctop col[2] 0.124f
C20994 row_n[7] col[19] 0.0342f
C20995 row_n[10] col[25] 0.0342f
C20996 row_n[13] col[31] 0.0342f
C20997 en_C0_n col[1] 0.142f
C20998 rowon_n[6] col[18] 0.0323f
C20999 row_n[9] col[23] 0.0342f
C21000 row_n[3] col[11] 0.0342f
C21001 rowon_n[1] col[8] 0.0323f
C21002 rowon_n[4] col[14] 0.0323f
C21003 vcm a_25054_7150# 0.56f
C21004 rowon_n[5] a_12914_7150# 0.118f
C21005 rowoff_n[12] a_19942_14178# 0.202f
C21006 a_2275_13198# a_26058_13174# 0.399f
C21007 col_n[13] a_16322_4178# 0.084f
C21008 VDD a_34090_16186# 0.483f
C21009 col_n[23] a_26362_16226# 0.084f
C21010 col[18] a_2475_7174# 0.136f
C21011 row_n[12] a_33390_14218# 0.0117f
C21012 col_n[4] a_6890_17190# 0.0765f
C21013 vcm a_15318_1166# 0.16f
C21014 m2_34864_15002# rowon_n[13] 0.231f
C21015 a_31990_6146# a_32386_6186# 0.0313f
C21016 m2_7756_946# m3_7888_1078# 3.79f
C21017 vcm a_5978_10162# 0.56f
C21018 a_2475_10186# a_18938_10162# 0.264f
C21019 a_2275_10186# a_16322_10202# 0.144f
C21020 row_n[14] a_23958_16186# 0.0437f
C21021 col_n[25] a_2275_13198# 0.113f
C21022 m2_21812_946# col_n[19] 0.331f
C21023 a_21038_15182# a_21342_15222# 0.0931f
C21024 a_21950_15182# a_22442_15544# 0.0658f
C21025 col_n[30] a_2275_2154# 0.113f
C21026 row_n[4] a_33998_6146# 0.0437f
C21027 rowon_n[8] a_33086_10162# 0.248f
C21028 a_28066_3134# a_29070_3134# 0.843f
C21029 col[7] a_9994_2130# 0.367f
C21030 m2_19804_18014# col[17] 0.347f
C21031 m2_1732_3958# a_2966_4138# 0.843f
C21032 col[17] a_20034_14178# 0.367f
C21033 vcm a_30378_5182# 0.155f
C21034 a_2275_7174# a_9902_7150# 0.136f
C21035 col[14] a_16930_4138# 0.0682f
C21036 col[15] a_2275_10186# 0.0899f
C21037 m2_21812_18014# vcm 0.353f
C21038 col[22] rowoff_n[12] 0.0901f
C21039 col[24] a_26970_16186# 0.0682f
C21040 vcm a_21038_14178# 0.56f
C21041 a_17934_12170# a_18026_12170# 0.326f
C21042 a_2275_12194# a_31382_12210# 0.144f
C21043 a_2475_12194# a_33998_12170# 0.264f
C21044 VDD a_17934_4138# 0.181f
C21045 row_n[8] a_10998_10162# 0.282f
C21046 col_n[2] a_5278_2170# 0.084f
C21047 col_n[12] a_15318_14218# 0.084f
C21048 rowon_n[12] a_10906_14178# 0.118f
C21049 a_19030_5142# a_19030_4138# 0.843f
C21050 m2_31852_946# ctop 0.0429f
C21051 m2_34864_6970# a_2275_7174# 0.278f
C21052 vcm a_11302_8194# 0.155f
C21053 m2_29844_18014# m2_30848_18014# 0.843f
C21054 rowoff_n[13] a_7894_15182# 0.202f
C21055 a_2275_9182# a_24962_9158# 0.136f
C21056 a_12914_9158# a_13310_9198# 0.0313f
C21057 m2_31276_15430# a_31078_15182# 0.165f
C21058 rowon_n[2] a_20946_4138# 0.118f
C21059 vcm a_2475_17214# 1.08f
C21060 ctop a_24050_3134# 4.11f
C21061 VDD a_32994_8154# 0.181f
C21062 col_n[23] a_26458_8516# 0.0283f
C21063 rowoff_n[5] a_9902_7150# 0.202f
C21064 col_n[5] a_2475_6170# 0.0531f
C21065 a_2275_18218# a_2874_18194# 0.136f
C21066 row_n[0] a_8290_2170# 0.0117f
C21067 a_31990_2130# a_32482_2492# 0.0658f
C21068 a_31078_2130# a_31382_2170# 0.0931f
C21069 vcm a_4882_2130# 0.1f
C21070 col[6] rowoff_n[13] 0.0901f
C21071 a_2475_6170# a_17022_6146# 0.316f
C21072 a_8990_6146# a_9994_6146# 0.843f
C21073 col[6] a_8990_12170# 0.367f
C21074 vcm a_26362_12210# 0.155f
C21075 rowoff_n[3] a_18938_5142# 0.202f
C21076 m2_1732_17010# row_n[15] 0.292f
C21077 col[3] a_5886_2130# 0.0682f
C21078 VDD a_24450_2492# 0.0779f
C21079 m2_7180_13422# row_n[11] 0.0128f
C21080 m2_13204_9406# row_n[7] 0.0128f
C21081 m2_19228_5390# row_n[3] 0.0128f
C21082 ctop a_4974_6146# 4.11f
C21083 m2_34864_6970# rowoff_n[5] 0.278f
C21084 col[13] a_15926_14178# 0.0682f
C21085 row_n[11] a_31990_13174# 0.0437f
C21086 a_32994_16186# a_33086_16186# 0.326f
C21087 VDD a_13918_11166# 0.181f
C21088 rowon_n[15] a_31078_17190# 0.248f
C21089 col_n[21] a_24050_8154# 0.251f
C21090 a_2275_3158# a_7986_3134# 0.399f
C21091 rowoff_n[8] a_10394_10524# 0.0133f
C21092 rowoff_n[1] a_27974_3134# 0.202f
C21093 col_n[2] a_2275_9182# 0.113f
C21094 col_n[28] a_30986_10162# 0.0765f
C21095 m2_34864_5966# a_35002_6146# 0.225f
C21096 vcm a_19942_6146# 0.1f
C21097 col_n[1] a_4274_12210# 0.084f
C21098 a_34090_9158# a_34090_8154# 0.843f
C21099 a_2475_8178# a_32082_8154# 0.316f
C21100 sample a_1957_2154# 0.345f
C21101 m2_22240_13422# a_22042_13174# 0.165f
C21102 m3_1864_1078# m2_1732_946# 3.79f
C21103 m3_2868_2082# m2_2736_946# 0.0341f
C21104 vcm a_7286_15222# 0.155f
C21105 a_27974_13174# a_28370_13214# 0.0313f
C21106 VDD a_5374_5504# 0.0779f
C21107 row_n[15] a_8990_17190# 0.282f
C21108 ctop a_20034_10162# 4.11f
C21109 col_n[22] a_2475_8178# 0.0531f
C21110 m2_34288_14426# row_n[12] 0.0128f
C21111 a_2275_17214# a_8290_17230# 0.144f
C21112 a_2475_17214# a_10906_17190# 0.264f
C21113 rowoff_n[6] a_19430_8516# 0.0133f
C21114 VDD a_28978_15182# 0.181f
C21115 col_n[12] a_15414_6508# 0.0283f
C21116 col_n[22] a_25454_18556# 0.0283f
C21117 a_2275_5166# a_23046_5142# 0.399f
C21118 a_12002_5142# a_12306_5182# 0.0931f
C21119 row_n[5] a_19030_7150# 0.282f
C21120 a_12914_5142# a_13406_5504# 0.0658f
C21121 rowon_n[9] a_18938_11166# 0.118f
C21122 vcm a_35002_10162# 0.101f
C21123 a_24050_10162# a_25054_10162# 0.843f
C21124 col[7] a_2475_16210# 0.136f
C21125 rowoff_n[4] a_28466_6508# 0.0133f
C21126 col[12] a_2475_5166# 0.136f
C21127 col_n[0] a_3366_12532# 0.0283f
C21128 m2_11772_946# a_2275_1150# 0.28f
C21129 m2_28840_946# a_29070_2130# 0.843f
C21130 a_2475_14202# a_1957_14202# 0.0734f
C21131 VDD a_20434_9520# 0.0779f
C21132 row_n[7] a_6282_9198# 0.0117f
C21133 col[2] a_4882_12170# 0.0682f
C21134 m3_1864_11118# a_2966_11166# 0.0302f
C21135 VDD a_9902_18194# 0.343f
C21136 a_2275_2154# a_13310_2170# 0.144f
C21137 a_2475_2154# a_15926_2130# 0.264f
C21138 a_8898_2130# a_8990_2130# 0.326f
C21139 col_n[10] a_13006_6146# 0.251f
C21140 m2_6176_1374# VDD 0.0194f
C21141 col_n[19] a_2275_11190# 0.113f
C21142 rowoff_n[9] a_20034_11166# 0.294f
C21143 m2_13204_11414# a_13006_11166# 0.165f
C21144 col_n[17] a_19942_8154# 0.0765f
C21145 vcm a_15926_13174# 0.1f
C21146 a_15014_12170# a_15014_11166# 0.843f
C21147 VDD a_12002_3134# 0.483f
C21148 m2_12776_18014# a_2275_18218# 0.28f
C21149 m2_4744_18014# a_5278_18234# 0.087f
C21150 a_8898_16186# a_9294_16226# 0.0313f
C21151 a_2275_16210# a_16930_16186# 0.136f
C21152 VDD a_35494_13536# 0.106f
C21153 rowon_n[3] a_5978_5142# 0.248f
C21154 row_n[8] sample_n 0.0596f
C21155 row_n[0] col[16] 0.0342f
C21156 rowon_n[4] col[25] 0.0323f
C21157 row_n[7] col[30] 0.0342f
C21158 col[3] col[4] 0.0355f
C21159 rowon_n[3] col[23] 0.0323f
C21160 rowon_n[5] col[27] 0.0323f
C21161 row_n[4] col[24] 0.0342f
C21162 row_n[3] col[22] 0.0342f
C21163 rowon_n[2] col[21] 0.0323f
C21164 rowon_n[0] col[17] 0.0323f
C21165 ctop col[13] 0.123f
C21166 rowon_n[1] col[19] 0.0323f
C21167 row_n[2] col[20] 0.0342f
C21168 row_n[1] col[18] 0.0342f
C21169 rowon_n[7] col[31] 0.0323f
C21170 rowon_n[6] col[29] 0.0323f
C21171 row_n[5] col[26] 0.0342f
C21172 row_n[6] col[28] 0.0342f
C21173 ctop a_16018_17190# 4.06f
C21174 col[9] a_2275_8178# 0.0899f
C21175 rowoff_n[7] a_29070_9158# 0.294f
C21176 a_2475_4162# a_30986_4138# 0.264f
C21177 col_n[1] a_4370_4500# 0.0283f
C21178 a_2275_4162# a_28370_4178# 0.144f
C21179 m2_32280_7398# a_32082_7150# 0.165f
C21180 col_n[11] a_14410_16548# 0.0283f
C21181 a_27062_9158# a_27366_9198# 0.0931f
C21182 a_27974_9158# a_28466_9520# 0.0658f
C21183 col[30] a_33086_5142# 0.367f
C21184 vcm a_30986_17190# 0.1f
C21185 a_4974_13174# a_5978_13174# 0.843f
C21186 a_2475_13198# a_8990_13174# 0.316f
C21187 col[29] a_2475_7174# 0.136f
C21188 VDD a_27062_7150# 0.483f
C21189 m2_8760_18014# a_2475_18218# 0.286f
C21190 a_2275_18218# a_31990_18194# 0.136f
C21191 VDD a_16418_16548# 0.0779f
C21192 a_2275_1150# a_21950_1126# 0.136f
C21193 row_n[12] a_17022_14178# 0.282f
C21194 vcm a_33086_2130# 0.56f
C21195 a_23958_6146# a_24050_6146# 0.326f
C21196 m2_22816_946# m2_23244_1374# 0.165f
C21197 m2_4168_9406# a_3970_9158# 0.165f
C21198 col_n[0] a_2475_4162# 0.0532f
C21199 col_n[25] a_28370_5182# 0.084f
C21200 row_n[2] a_27062_4138# 0.282f
C21201 VDD a_17326_1166# 0.0149f
C21202 row_n[14] a_4274_16226# 0.0117f
C21203 col_n[9] a_12002_16186# 0.251f
C21204 rowon_n[6] a_26970_8154# 0.118f
C21205 col_n[6] a_8898_6146# 0.0765f
C21206 a_2475_15206# a_24050_15182# 0.316f
C21207 a_30074_16186# a_30074_15182# 0.843f
C21208 col_n[16] a_18938_18194# 0.0762f
C21209 VDD a_7986_10162# 0.483f
C21210 m2_1732_3958# col[0] 0.0137f
C21211 row_n[4] a_14314_6186# 0.0117f
C21212 a_2475_18218# a_29982_18194# 0.264f
C21213 col[26] a_2275_10186# 0.0899f
C21214 a_18938_3134# a_19334_3174# 0.0313f
C21215 m2_23244_5390# a_23046_5142# 0.165f
C21216 vcm a_14010_5142# 0.56f
C21217 rowoff_n[10] a_7986_12170# 0.294f
C21218 a_27974_1126# vcm 0.0989f
C21219 row_n[6] a_4882_8154# 0.0437f
C21220 m2_3164_8402# rowon_n[6] 0.0322f
C21221 vcm a_2966_14178# 0.56f
C21222 m2_9188_4386# rowon_n[2] 0.0322f
C21223 a_7986_12170# a_8290_12210# 0.0931f
C21224 a_2275_12194# a_15014_12170# 0.399f
C21225 a_8898_12170# a_9390_12532# 0.0658f
C21226 rowon_n[10] a_3970_12170# 0.248f
C21227 m2_25828_18014# VDD 1f
C21228 col[19] a_22042_3134# 0.367f
C21229 a_20034_17190# a_21038_17190# 0.843f
C21230 VDD a_23046_14178# 0.483f
C21231 col[29] a_32082_15182# 0.367f
C21232 a_2275_1150# m2_2736_946# 0.281f
C21233 col[26] a_28978_5142# 0.0682f
C21234 rowon_n[0] a_14010_2130# 0.248f
C21235 col_n[11] a_2475_17214# 0.0531f
C21236 vcm a_29070_9158# 0.56f
C21237 a_2475_9182# a_7894_9158# 0.264f
C21238 a_2275_9182# a_5278_9198# 0.144f
C21239 a_4882_9158# a_4974_9158# 0.326f
C21240 a_3878_9158# a_4274_9198# 0.0313f
C21241 rowoff_n[14] a_24050_16186# 0.294f
C21242 col_n[16] a_2475_6170# 0.0531f
C21243 rowon_n[2] a_2275_4162# 1.79f
C21244 col_n[14] a_17326_3174# 0.084f
C21245 a_2275_14202# a_30074_14178# 0.399f
C21246 m2_18224_17438# rowon_n[15] 0.0322f
C21247 m2_34864_13998# ctop 0.0422f
C21248 m2_24248_13422# rowon_n[11] 0.0322f
C21249 m2_30272_9406# rowon_n[7] 0.0322f
C21250 col_n[24] a_27366_15222# 0.084f
C21251 m2_35292_5390# rowon_n[3] 0.0322f
C21252 col[17] rowoff_n[13] 0.0901f
C21253 VDD a_3970_17190# 0.484f
C21254 col_n[5] a_7894_16186# 0.0765f
C21255 col[1] a_2475_14202# 0.136f
C21256 m2_14208_3382# a_14010_3134# 0.165f
C21257 vcm a_19334_3174# 0.155f
C21258 VDD rowoff_n[6] 1.51f
C21259 col_n[0] rowoff_n[8] 0.0471f
C21260 col[6] a_2475_3158# 0.136f
C21261 vcm rowoff_n[9] 0.533f
C21262 sample rowoff_n[7] 0.0775f
C21263 row_n[9] a_25054_11166# 0.282f
C21264 rowon_n[13] a_24962_15182# 0.118f
C21265 vcm a_9994_12170# 0.56f
C21266 a_2275_11190# a_20338_11206# 0.144f
C21267 a_2475_11190# a_22954_11166# 0.264f
C21268 VDD a_6890_2130# 0.181f
C21269 m2_23820_18014# a_24354_18234# 0.087f
C21270 row_n[11] a_12306_13214# 0.0117f
C21271 a_23046_16186# a_23350_16226# 0.0931f
C21272 a_23958_16186# a_24450_16548# 0.0658f
C21273 rowon_n[3] a_35002_5142# 0.118f
C21274 m2_19804_18014# m3_18932_18146# 0.0341f
C21275 col_n[13] a_2275_9182# 0.113f
C21276 col[18] a_21038_13174# 0.367f
C21277 a_30074_4138# a_31078_4138# 0.843f
C21278 col[15] a_17934_3134# 0.0682f
C21279 row_n[1] a_22346_3174# 0.0117f
C21280 row_n[13] a_2161_15206# 0.0221f
C21281 vcm a_35398_7190# 0.161f
C21282 col[25] a_27974_15182# 0.0682f
C21283 a_2275_8178# a_13918_8154# 0.136f
C21284 rowoff_n[12] a_30474_14540# 0.0133f
C21285 col_n[0] a_3270_9198# 0.084f
C21286 vcm a_25054_16186# 0.56f
C21287 a_2275_13198# a_2275_12194# 0.0715f
C21288 a_19942_13174# a_20034_13174# 0.326f
C21289 VDD a_21950_6146# 0.181f
C21290 col[3] a_2275_6170# 0.0899f
C21291 row_n[3] a_12914_5142# 0.0437f
C21292 col[1] rowoff_n[14] 0.0901f
C21293 col_n[3] a_6282_1166# 0.0839f
C21294 rowon_n[7] a_12002_9158# 0.248f
C21295 col_n[13] a_16322_13214# 0.084f
C21296 col[18] a_2475_16210# 0.136f
C21297 a_3878_5142# a_4370_5504# 0.0658f
C21298 a_2966_5142# a_3270_5182# 0.0931f
C21299 a_21038_6146# a_21038_5142# 0.843f
C21300 a_2475_5166# a_5978_5142# 0.316f
C21301 m2_22816_946# m3_23952_1078# 0.0341f
C21302 m3_32988_18146# m3_33992_18146# 0.202f
C21303 m2_34864_946# m3_34996_2082# 0.0341f
C21304 col[23] a_2475_5166# 0.136f
C21305 vcm a_15318_10202# 0.155f
C21306 a_14922_10162# a_15318_10202# 0.0313f
C21307 rowoff_n[15] a_12002_17190# 0.294f
C21308 a_2275_10186# a_28978_10162# 0.136f
C21309 col_n[24] a_27462_7512# 0.0283f
C21310 rowoff_n[4] a_10906_6146# 0.202f
C21311 ctop a_28066_5142# 4.11f
C21312 VDD a_2161_9182# 0.187f
C21313 col_n[30] a_2275_11190# 0.113f
C21314 a_33998_3134# a_34490_3496# 0.0658f
C21315 a_33086_3134# a_33390_3174# 0.0931f
C21316 m2_2160_7398# row_n[5] 0.0194f
C21317 m2_8184_3382# row_n[1] 0.0128f
C21318 m2_1732_9982# m2_2160_10410# 0.165f
C21319 vcm a_8898_4138# 0.1f
C21320 rowoff_n[2] a_19942_4138# 0.202f
C21321 a_2475_7174# a_21038_7150# 0.316f
C21322 col[7] a_9994_11166# 0.367f
C21323 a_10998_7150# a_12002_7150# 0.843f
C21324 rowoff_n[9] a_1957_11190# 0.0219f
C21325 col[4] a_6890_1126# 0.0682f
C21326 row_n[6] a_33086_8154# 0.282f
C21327 vcm a_30378_14218# 0.155f
C21328 col[14] a_16930_13174# 0.0682f
C21329 VDD col_n[1] 4.83f
C21330 VDD a_28466_4500# 0.0779f
C21331 sample vcm 16.6f
C21332 rowon_n[10] a_32994_12170# 0.118f
C21333 row_n[2] col[31] 0.0342f
C21334 rowon_n[1] col[30] 0.0323f
C21335 rowon_n[2] sample_n 0.0692f
C21336 ctop col[24] 0.123f
C21337 row_n[0] col[27] 0.0342f
C21338 row_n[1] col[29] 0.0342f
C21339 rowon_n[0] col[28] 0.0323f
C21340 ctop a_8990_8154# 4.11f
C21341 col[20] a_2275_8178# 0.0899f
C21342 col_n[22] a_25054_7150# 0.251f
C21343 a_34090_17190# a_34394_17230# 0.0931f
C21344 a_35002_17190# a_35094_17190# 0.0991f
C21345 VDD a_17934_13174# 0.181f
C21346 row_n[8] a_20338_10202# 0.0117f
C21347 rowoff_n[0] a_28978_2130# 0.202f
C21348 rowoff_n[7] a_11398_9520# 0.0133f
C21349 col_n[29] a_31990_9158# 0.0765f
C21350 a_2275_4162# a_12002_4138# 0.399f
C21351 col_n[2] a_5278_11206# 0.084f
C21352 m3_34996_17142# ctop 0.209f
C21353 m2_17220_16434# row_n[14] 0.0128f
C21354 m2_23244_12418# row_n[10] 0.0128f
C21355 vcm a_23958_8154# 0.1f
C21356 a_2475_9182# a_2475_8178# 0.0666f
C21357 m2_29268_8402# row_n[6] 0.0128f
C21358 rowoff_n[13] a_18426_15544# 0.0133f
C21359 m2_34864_3958# row_n[2] 0.267f
C21360 row_n[10] a_10906_12170# 0.0437f
C21361 vcm a_11302_17230# 0.155f
C21362 a_29982_14178# a_30378_14218# 0.0313f
C21363 rowon_n[14] a_9994_16186# 0.248f
C21364 VDD a_9390_7512# 0.0779f
C21365 rowoff_n[5] a_20434_7512# 0.0133f
C21366 col_n[13] a_16418_5504# 0.0283f
C21367 ctop a_24050_12170# 4.11f
C21368 a_2275_18218# a_12306_18234# 0.145f
C21369 col_n[23] a_26458_17552# 0.0283f
C21370 VDD a_32994_17190# 0.181f
C21371 row_n[0] a_20946_2130# 0.0437f
C21372 col_n[5] a_2475_15206# 0.0531f
C21373 a_2475_1150# a_4882_1126# 0.264f
C21374 a_2874_1126# a_3366_1488# 0.0658f
C21375 a_2275_1150# a_3878_1126# 0.106f
C21376 rowon_n[4] a_20034_6146# 0.248f
C21377 col_n[10] a_2475_4162# 0.0531f
C21378 m2_1732_1950# a_2275_2154# 0.191f
C21379 a_2275_6170# a_27062_6146# 0.399f
C21380 a_14922_6146# a_15414_6508# 0.0658f
C21381 a_14010_6146# a_14314_6186# 0.0931f
C21382 rowoff_n[3] a_29470_5504# 0.0133f
C21383 vcm a_4882_11166# 0.1f
C21384 a_26058_11166# a_27062_11166# 0.843f
C21385 a_2275_15206# a_5886_15182# 0.136f
C21386 VDD a_24450_11528# 0.0779f
C21387 col[3] a_5886_11166# 0.0682f
C21388 col[0] a_2475_1150# 0.148f
C21389 ctop a_4974_15182# 4.11f
C21390 col_n[11] a_14010_5142# 0.251f
C21391 a_2475_3158# a_19942_3134# 0.264f
C21392 a_10906_3134# a_10998_3134# 0.326f
C21393 a_2275_3158# a_17326_3174# 0.144f
C21394 rowoff_n[8] a_21038_10162# 0.294f
C21395 col_n[21] a_24050_17190# 0.251f
C21396 a_33086_1126# a_2475_1150# 0.0299f
C21397 row_n[13] a_31078_15182# 0.282f
C21398 col_n[18] a_20946_7150# 0.0765f
C21399 m2_34864_13998# m2_34864_12994# 0.843f
C21400 rowoff_n[11] a_24962_13174# 0.202f
C21401 col_n[2] a_2275_18218# 0.113f
C21402 col_n[7] a_2275_7174# 0.113f
C21403 vcm a_19942_15182# 0.1f
C21404 a_17022_13174# a_17022_12170# 0.843f
C21405 VDD a_16018_5142# 0.483f
C21406 sample a_1957_11190# 0.345f
C21407 a_29982_1126# VDD 0.405f
C21408 row_n[15] a_18330_17230# 0.0117f
C21409 a_2275_17214# a_20946_17190# 0.136f
C21410 a_10906_17190# a_11302_17230# 0.0313f
C21411 VDD a_5374_14540# 0.0779f
C21412 rowoff_n[6] a_30074_8154# 0.294f
C21413 a_23046_2130# m2_23244_2378# 0.165f
C21414 col_n[2] a_5374_3496# 0.0283f
C21415 col_n[22] a_2475_17214# 0.0531f
C21416 col_n[12] a_15414_15544# 0.0283f
C21417 a_2275_5166# a_32386_5182# 0.144f
C21418 row_n[5] a_28370_7190# 0.0117f
C21419 a_2475_5166# a_35002_5142# 0.264f
C21420 col_n[27] a_2475_6170# 0.0531f
C21421 m3_22948_1078# m3_23952_1078# 0.202f
C21422 col[31] a_34090_4138# 0.367f
C21423 a_31990_1126# a_32082_1126# 0.0991f
C21424 a_29070_10162# a_29374_10202# 0.0931f
C21425 rowoff_n[14] a_6378_16548# 0.0133f
C21426 a_29982_10162# a_30474_10524# 0.0658f
C21427 m2_12776_946# a_13006_1126# 0.0249f
C21428 col[28] rowoff_n[13] 0.0901f
C21429 m3_15920_1078# a_16018_2130# 0.0302f
C21430 a_2475_14202# a_13006_14178# 0.316f
C21431 a_6982_14178# a_7986_14178# 0.843f
C21432 VDD a_31078_9158# 0.483f
C21433 row_n[7] a_18938_9158# 0.0437f
C21434 col[12] a_2475_14202# 0.136f
C21435 rowon_n[11] a_18026_13174# 0.248f
C21436 VDD a_20434_18556# 0.0858f
C21437 col_n[4] rowoff_n[2] 0.0471f
C21438 col_n[3] rowoff_n[1] 0.0471f
C21439 col_n[2] rowoff_n[0] 0.0471f
C21440 col_n[10] rowoff_n[8] 0.0471f
C21441 col_n[9] rowoff_n[7] 0.0471f
C21442 col_n[8] rowoff_n[6] 0.0471f
C21443 col_n[11] rowoff_n[9] 0.0471f
C21444 col_n[6] rowoff_n[4] 0.0471f
C21445 col_n[5] rowoff_n[3] 0.0471f
C21446 col_n[7] rowoff_n[5] 0.0471f
C21447 col[17] a_2475_3158# 0.136f
C21448 a_2275_2154# a_25966_2130# 0.136f
C21449 m2_34864_3958# a_34090_4138# 0.843f
C21450 m2_29268_1374# VDD 0.0194f
C21451 vcm a_2874_3134# 0.1f
C21452 col_n[26] a_29374_4178# 0.084f
C21453 a_25966_7150# a_26058_7150# 0.326f
C21454 rowon_n[1] a_28066_3134# 0.248f
C21455 col_n[10] a_13006_15182# 0.251f
C21456 col_n[7] a_9902_5142# 0.0765f
C21457 a_2275_11190# a_3970_11166# 0.399f
C21458 col_n[24] a_2275_9182# 0.113f
C21459 col_n[17] a_19942_17190# 0.0765f
C21460 a_2475_16210# a_28066_16186# 0.316f
C21461 a_32082_17190# a_32082_16186# 0.843f
C21462 VDD a_12002_12170# 0.483f
C21463 a_20946_4138# a_21342_4178# 0.0313f
C21464 row_n[1] a_5978_3134# 0.282f
C21465 col[9] a_2275_17214# 0.0899f
C21466 rowon_n[5] a_5886_7150# 0.118f
C21467 vcm a_18026_7150# 0.56f
C21468 col[14] a_2275_6170# 0.0899f
C21469 rowoff_n[12] a_12914_14178# 0.202f
C21470 col_n[1] a_4370_13536# 0.0283f
C21471 m2_28264_14426# a_28066_14178# 0.165f
C21472 col[12] rowoff_n[14] 0.0901f
C21473 col[20] a_23046_2130# 0.367f
C21474 a_2275_13198# a_19030_13174# 0.399f
C21475 a_9994_13174# a_10298_13214# 0.0931f
C21476 a_10906_13174# a_11398_13536# 0.0658f
C21477 VDD a_3878_6146# 0.181f
C21478 col[30] a_33086_14178# 0.367f
C21479 col[27] a_29982_4138# 0.0682f
C21480 col[29] a_2475_16210# 0.136f
C21481 VDD a_27062_16186# 0.483f
C21482 row_n[12] a_26362_14218# 0.0117f
C21483 vcm a_8290_1166# 0.16f
C21484 m2_7180_15430# rowon_n[13] 0.0322f
C21485 m2_13204_11414# rowon_n[9] 0.0322f
C21486 m2_19228_7398# rowon_n[5] 0.0322f
C21487 m2_25252_3382# rowon_n[1] 0.0322f
C21488 vcm a_33086_11166# 0.56f
C21489 col_n[15] a_18330_2170# 0.0839f
C21490 a_2275_10186# a_9294_10202# 0.144f
C21491 a_2475_10186# a_11910_10162# 0.264f
C21492 a_6890_10162# a_6982_10162# 0.326f
C21493 row_n[14] a_16930_16186# 0.0437f
C21494 col_n[25] a_28370_14218# 0.084f
C21495 col_n[0] a_2475_13198# 0.0532f
C21496 a_2275_15206# a_34090_15182# 0.399f
C21497 col_n[4] a_2475_2154# 0.0531f
C21498 col_n[6] a_8898_15182# 0.0765f
C21499 row_n[4] a_26970_6146# 0.0437f
C21500 rowon_n[8] a_26058_10162# 0.248f
C21501 a_7986_3134# a_7986_2130# 0.843f
C21502 vcm a_23350_5182# 0.155f
C21503 VDD col_n[12] 5.17f
C21504 vcm col_n[9] 1.94f
C21505 col_n[4] col_n[5] 0.0101f
C21506 a_2475_7174# a_2966_7150# 0.317f
C21507 a_2161_7174# a_2275_7174# 0.183f
C21508 col[14] col[15] 0.0355f
C21509 m2_7756_18014# vcm 0.353f
C21510 m2_19228_12418# a_19030_12170# 0.165f
C21511 m2_34288_16434# rowon_n[14] 0.0322f
C21512 col[31] a_2275_8178# 0.0899f
C21513 vcm a_14010_14178# 0.56f
C21514 a_2475_12194# a_26970_12170# 0.264f
C21515 a_2275_12194# a_24354_12210# 0.144f
C21516 VDD a_10906_4138# 0.181f
C21517 a_25966_17190# a_26458_17552# 0.0658f
C21518 a_25054_17190# a_25358_17230# 0.0931f
C21519 col[19] a_22042_12170# 0.367f
C21520 row_n[8] a_3970_10162# 0.282f
C21521 col[16] a_18938_2130# 0.0682f
C21522 a_32082_5142# a_33086_5142# 0.843f
C21523 col[26] a_28978_14178# 0.0682f
C21524 col_n[1] a_2275_5166# 0.113f
C21525 m2_22816_18014# m2_23820_18014# 0.843f
C21526 vcm a_4274_8194# 0.155f
C21527 a_2275_9182# a_17934_9158# 0.136f
C21528 m2_5748_946# col_n[3] 0.331f
C21529 rowon_n[2] a_13918_4138# 0.118f
C21530 ctop a_17022_3134# 4.11f
C21531 vcm a_29070_18194# 0.165f
C21532 a_21950_14178# a_22042_14178# 0.326f
C21533 col_n[16] a_2475_15206# 0.0531f
C21534 VDD a_25966_8154# 0.181f
C21535 rowoff_n[5] a_2161_7174# 0.0226f
C21536 col_n[21] a_2475_4162# 0.0531f
C21537 col_n[14] a_17326_12210# 0.084f
C21538 row_n[0] a_2275_2154# 19.2f
C21539 rowon_n[4] a_1957_6170# 0.0172f
C21540 m3_34996_1078# VDD 0.0192f
C21541 row_n[9] a_35398_11206# 0.0117f
C21542 vcm a_31990_3134# 0.1f
C21543 a_23046_7150# a_23046_6146# 0.843f
C21544 a_2475_6170# a_9994_6146# 0.316f
C21545 m2_10192_10410# a_9994_10162# 0.165f
C21546 col_n[25] a_28466_6508# 0.0283f
C21547 rowoff_n[3] a_11910_5142# 0.202f
C21548 vcm a_19334_12210# 0.155f
C21549 col[6] a_2475_12194# 0.136f
C21550 a_2275_11190# a_32994_11166# 0.136f
C21551 a_16930_11166# a_17326_11206# 0.0313f
C21552 VDD a_17422_2492# 0.0779f
C21553 col[11] a_2475_1150# 0.136f
C21554 m2_34864_8978# VDD 0.772f
C21555 ctop a_32082_7150# 4.11f
C21556 row_n[11] a_24962_13174# 0.0437f
C21557 VDD a_6890_11166# 0.181f
C21558 m2_33860_18014# m3_33992_18146# 3.79f
C21559 rowon_n[15] a_24050_17190# 0.248f
C21560 col_n[13] a_2275_18218# 0.113f
C21561 rowoff_n[1] a_20946_3134# 0.202f
C21562 col[8] a_10998_10162# 0.367f
C21563 rowoff_n[8] a_2966_10162# 0.294f
C21564 row_n[1] a_35002_3134# 0.0437f
C21565 m2_29268_6394# a_29070_6146# 0.165f
C21566 col_n[18] a_2275_7174# 0.113f
C21567 vcm a_12914_6146# 0.1f
C21568 rowon_n[5] a_34090_7150# 0.248f
C21569 a_2475_8178# a_25054_8154# 0.316f
C21570 a_13006_8154# a_14010_8154# 0.843f
C21571 col[15] a_17934_12170# 0.0682f
C21572 vcm a_35398_16226# 0.161f
C21573 col_n[23] a_26058_6146# 0.251f
C21574 VDD a_32482_6508# 0.0779f
C21575 col_n[0] a_3270_18234# 0.084f
C21576 ctop a_13006_10162# 4.11f
C21577 row_n[15] a_2475_17214# 0.405f
C21578 m2_6176_14426# row_n[12] 0.0128f
C21579 rowoff_n[6] a_12402_8516# 0.0133f
C21580 VDD a_21950_15182# 0.181f
C21581 col_n[30] a_32994_8154# 0.0765f
C21582 m2_12200_10410# row_n[8] 0.0128f
C21583 col[3] a_2275_15206# 0.0899f
C21584 m2_18224_6394# row_n[4] 0.0128f
C21585 col[8] a_2275_4162# 0.0899f
C21586 col_n[3] a_6282_10202# 0.084f
C21587 a_2275_5166# a_16018_5142# 0.399f
C21588 row_n[5] a_12002_7150# 0.282f
C21589 m2_2736_1950# vcm 0.353f
C21590 m3_1864_8106# m3_1864_7102# 0.202f
C21591 rowon_n[9] a_11910_11166# 0.118f
C21592 vcm a_27974_10162# 0.1f
C21593 a_3970_10162# a_3970_9158# 0.843f
C21594 col[23] a_2475_14202# 0.136f
C21595 rowoff_n[4] a_21438_6508# 0.0133f
C21596 col_n[14] a_17422_4500# 0.0283f
C21597 col_n[20] rowoff_n[7] 0.0471f
C21598 col_n[16] rowoff_n[3] 0.0471f
C21599 a_31990_15182# a_32386_15222# 0.0313f
C21600 col_n[13] rowoff_n[0] 0.0471f
C21601 col_n[21] rowoff_n[8] 0.0471f
C21602 col[28] a_2475_3158# 0.136f
C21603 col_n[15] rowoff_n[2] 0.0471f
C21604 col_n[22] rowoff_n[9] 0.0471f
C21605 col_n[17] rowoff_n[4] 0.0471f
C21606 col_n[18] rowoff_n[5] 0.0471f
C21607 col_n[19] rowoff_n[6] 0.0471f
C21608 col_n[14] rowoff_n[1] 0.0471f
C21609 m2_1732_17010# ctop 0.0424f
C21610 VDD a_13406_9520# 0.0779f
C21611 col_n[24] a_27462_16548# 0.0283f
C21612 ctop a_28066_14178# 4.11f
C21613 col_n[0] a_2475_18218# 0.053f
C21614 VDD a_2161_18218# 0.227f
C21615 a_2275_2154# a_6282_2170# 0.144f
C21616 a_2475_2154# a_8898_2130# 0.264f
C21617 m2_33284_15430# row_n[13] 0.0128f
C21618 m2_20232_4386# a_20034_4138# 0.165f
C21619 rowoff_n[9] a_13006_11166# 0.294f
C21620 a_16018_7150# a_16322_7190# 0.0931f
C21621 rowoff_n[2] a_30474_4500# 0.0133f
C21622 a_2275_7174# a_31078_7150# 0.399f
C21623 a_16930_7150# a_17422_7512# 0.0658f
C21624 vcm a_8898_13174# 0.1f
C21625 a_28066_12170# a_29070_12170# 0.843f
C21626 VDD a_4974_3134# 0.483f
C21627 col[4] a_6890_10162# 0.0682f
C21628 a_2275_16210# a_9902_16186# 0.136f
C21629 VDD a_28466_13536# 0.0779f
C21630 col_n[12] a_15014_4138# 0.251f
C21631 ctop a_8990_17190# 4.06f
C21632 col[20] a_2275_17214# 0.0899f
C21633 row_n[8] a_32994_10162# 0.0437f
C21634 rowoff_n[7] a_22042_9158# 0.294f
C21635 col_n[22] a_25054_16186# 0.251f
C21636 col[25] a_2275_6170# 0.0899f
C21637 col_n[19] a_21950_6146# 0.0765f
C21638 rowon_n[12] a_32082_14178# 0.248f
C21639 a_2475_4162# a_23958_4138# 0.264f
C21640 a_12914_4138# a_13006_4138# 0.326f
C21641 a_2275_4162# a_21342_4178# 0.144f
C21642 m3_12908_1078# ctop 0.21f
C21643 col[23] rowoff_n[14] 0.0901f
C21644 col_n[29] a_31990_18194# 0.0762f
C21645 rowoff_n[13] a_29070_15182# 0.294f
C21646 col_n[6] rowoff_n[10] 0.0471f
C21647 col_n[0] a_2966_10162# 0.251f
C21648 vcm a_23958_17190# 0.1f
C21649 a_19030_14178# a_19030_13174# 0.843f
C21650 VDD a_20034_7150# 0.483f
C21651 rowoff_n[5] a_31078_7150# 0.294f
C21652 a_12914_18194# a_13310_18234# 0.0313f
C21653 col_n[3] a_6378_2492# 0.0283f
C21654 a_2275_18218# a_24962_18194# 0.136f
C21655 VDD a_9390_16548# 0.0779f
C21656 col_n[13] a_16418_14540# 0.0283f
C21657 a_7894_1126# a_8290_1166# 0.0313f
C21658 a_2275_1150# a_14922_1126# 0.136f
C21659 row_n[12] a_9994_14178# 0.282f
C21660 vcm a_26058_2130# 0.56f
C21661 a_2966_6146# a_2966_5142# 0.843f
C21662 col_n[10] a_2475_13198# 0.0531f
C21663 row_n[2] a_20034_4138# 0.282f
C21664 col_n[15] a_2475_2154# 0.0531f
C21665 a_31990_11166# a_32482_11528# 0.0658f
C21666 a_31078_11166# a_31382_11206# 0.0931f
C21667 VDD a_10298_1166# 0.0149f
C21668 rowon_n[6] a_19942_8154# 0.118f
C21669 a_8990_15182# a_9994_15182# 0.843f
C21670 a_2475_15206# a_17022_15182# 0.316f
C21671 rowon_n[0] m2_30272_2378# 0.0322f
C21672 row_n[4] a_7286_6186# 0.0117f
C21673 vcm col_n[20] 1.94f
C21674 VDD col_n[23] 5.17f
C21675 col_n[27] a_30378_3174# 0.084f
C21676 col[7] rowoff_n[15] 0.0901f
C21677 a_2275_3158# a_29982_3134# 0.136f
C21678 col_n[1] a_3970_2130# 0.25f
C21679 col[0] a_2475_10186# 0.148f
C21680 a_2475_18218# a_22954_18194# 0.264f
C21681 col_n[11] a_14010_14178# 0.251f
C21682 vcm a_6982_5142# 0.56f
C21683 col_n[8] a_10906_4138# 0.0765f
C21684 rowoff_n[11] a_35494_13536# 0.0133f
C21685 a_27974_8154# a_28066_8154# 0.326f
C21686 col_n[18] a_20946_16186# 0.0765f
C21687 a_2275_12194# a_7986_12170# 0.399f
C21688 m2_11772_18014# VDD 1.07f
C21689 row_n[15] a_30986_17190# 0.0437f
C21690 col_n[7] a_2275_16210# 0.113f
C21691 a_2475_17214# a_32082_17190# 0.316f
C21692 VDD a_16018_14178# 0.483f
C21693 col_n[12] a_2275_5166# 0.113f
C21694 rowon_n[0] a_6982_2130# 0.248f
C21695 a_22954_5142# a_23350_5182# 0.0313f
C21696 col_n[2] a_5374_12532# 0.0283f
C21697 vcm a_22042_9158# 0.56f
C21698 col_n[27] a_2475_15206# 0.0531f
C21699 rowoff_n[14] a_17022_16186# 0.294f
C21700 col[31] a_34090_13174# 0.367f
C21701 col[2] a_2275_2154# 0.0899f
C21702 col[28] a_30986_3134# 0.0682f
C21703 m2_20808_946# a_20946_1126# 0.225f
C21704 a_12002_14178# a_12306_14218# 0.0931f
C21705 a_12914_14178# a_13406_14540# 0.0658f
C21706 a_2275_14202# a_23046_14178# 0.399f
C21707 m2_2160_9406# rowon_n[7] 0.0219f
C21708 m2_8184_5390# rowon_n[3] 0.0322f
C21709 m2_9764_946# vcm 0.353f
C21710 VDD a_31078_18194# 0.0356f
C21711 a_19030_2130# a_20034_2130# 0.843f
C21712 m3_31984_18146# VDD 0.0636f
C21713 col[17] a_2475_12194# 0.136f
C21714 row_n[9] a_18026_11166# 0.282f
C21715 vcm a_12306_3174# 0.155f
C21716 col[22] a_2475_1150# 0.136f
C21717 m2_1732_15002# sample_n 0.0522f
C21718 col_n[16] a_19334_1166# 0.0572f
C21719 rowon_n[13] a_17934_15182# 0.118f
C21720 col_n[26] a_29374_13214# 0.084f
C21721 vcm a_2874_12170# 0.1f
C21722 a_2275_11190# a_13310_11206# 0.144f
C21723 a_2475_11190# a_15926_11166# 0.264f
C21724 a_8898_11166# a_8990_11166# 0.326f
C21725 VDD a_33998_3134# 0.181f
C21726 col_n[7] a_9902_14178# 0.0765f
C21727 row_n[11] a_5278_13214# 0.0117f
C21728 rowon_n[3] a_27974_5142# 0.118f
C21729 col_n[24] a_2275_18218# 0.113f
C21730 m2_9764_18014# m3_10900_18146# 0.0341f
C21731 m2_23244_14426# rowon_n[12] 0.0322f
C21732 col_n[29] a_2275_7174# 0.113f
C21733 m2_29268_10410# rowon_n[8] 0.0322f
C21734 m2_34864_5966# rowon_n[4] 0.231f
C21735 a_9994_4138# a_9994_3134# 0.843f
C21736 rowoff_n[1] a_2275_3158# 0.151f
C21737 row_n[1] a_15318_3174# 0.0117f
C21738 vcm a_27366_7190# 0.155f
C21739 rowoff_n[12] a_23446_14540# 0.0133f
C21740 a_2275_8178# a_6890_8154# 0.136f
C21741 m2_1732_12994# a_2161_13198# 0.0454f
C21742 vcm a_18026_16186# 0.56f
C21743 a_2475_13198# a_30986_13174# 0.264f
C21744 a_2275_13198# a_28370_13214# 0.144f
C21745 col[14] a_2275_15206# 0.0899f
C21746 VDD a_14922_6146# 0.181f
C21747 row_n[3] a_5886_5142# 0.0437f
C21748 col[19] a_2275_4162# 0.0899f
C21749 col[20] a_23046_11166# 0.367f
C21750 rowon_n[7] a_4974_9158# 0.248f
C21751 a_27974_18194# a_28466_18556# 0.0658f
C21752 col[17] a_19942_1126# 0.0703f
C21753 VDD a_3878_15182# 0.181f
C21754 a_22954_1126# a_23446_1488# 0.0658f
C21755 col[27] a_29982_13174# 0.0682f
C21756 vcm a_20946_1126# 0.0989f
C21757 a_33998_6146# a_34394_6186# 0.0313f
C21758 m2_12776_946# m3_12908_1078# 3.79f
C21759 m3_18932_18146# m3_19936_18146# 0.202f
C21760 col_n[29] rowoff_n[5] 0.0471f
C21761 col_n[28] rowoff_n[4] 0.0471f
C21762 vcm a_8290_10202# 0.155f
C21763 col_n[31] rowoff_n[7] 0.0471f
C21764 col_n[27] rowoff_n[3] 0.0471f
C21765 col_n[30] rowoff_n[6] 0.0471f
C21766 col_n[26] rowoff_n[2] 0.0471f
C21767 col_n[25] rowoff_n[1] 0.0471f
C21768 col_n[24] rowoff_n[0] 0.0471f
C21769 rowoff_n[15] a_4974_17190# 0.294f
C21770 a_2275_10186# a_21950_10162# 0.136f
C21771 m2_34864_16006# a_2475_16210# 0.282f
C21772 rowoff_n[4] a_3366_6508# 0.0133f
C21773 ctop a_21038_5142# 4.11f
C21774 m2_11772_946# a_12002_2130# 0.843f
C21775 col_n[15] a_18330_11206# 0.084f
C21776 col_n[10] a_2475_18218# 0.0529f
C21777 a_23958_15182# a_24050_15182# 0.326f
C21778 VDD a_29982_10162# 0.181f
C21779 col_n[4] a_2475_11190# 0.0531f
C21780 vcm a_34394_5182# 0.155f
C21781 col_n[26] a_29470_5504# 0.0283f
C21782 a_25054_8154# a_25054_7150# 0.843f
C21783 a_2475_7174# a_14010_7150# 0.316f
C21784 rowoff_n[2] a_12914_4138# 0.202f
C21785 rowoff_n[10] a_29982_12170# 0.202f
C21786 row_n[6] a_26058_8154# 0.282f
C21787 vcm a_23350_14218# 0.155f
C21788 a_18938_12170# a_19334_12210# 0.0313f
C21789 VDD a_21438_4500# 0.0779f
C21790 rowon_n[10] a_25966_12170# 0.118f
C21791 col[31] a_2275_17214# 0.0899f
C21792 ctop a_2475_8178# 0.0488f
C21793 VDD a_10906_13174# 0.181f
C21794 row_n[8] a_13310_10202# 0.0117f
C21795 col[9] a_12002_9158# 0.367f
C21796 rowoff_n[0] a_21950_2130# 0.202f
C21797 rowoff_n[7] a_4370_9520# 0.0133f
C21798 vcm m2_34864_1950# 0.408f
C21799 a_2275_4162# a_4974_4138# 0.399f
C21800 a_2874_4138# a_3270_4178# 0.0313f
C21801 a_3878_4138# a_3970_4138# 0.326f
C21802 m3_8892_18146# ctop 0.209f
C21803 col_n[17] rowoff_n[10] 0.0471f
C21804 col[16] a_18938_11166# 0.0682f
C21805 vcm a_16930_8154# 0.1f
C21806 m2_33860_18014# m2_34288_18442# 0.165f
C21807 m2_1732_7974# row_n[6] 0.292f
C21808 a_15014_9158# a_16018_9158# 0.843f
C21809 a_2475_9182# a_29070_9158# 0.316f
C21810 rowoff_n[13] a_11398_15544# 0.0133f
C21811 col_n[1] a_2275_14202# 0.113f
C21812 m2_7180_4386# row_n[2] 0.0128f
C21813 col_n[24] a_27062_5142# 0.251f
C21814 m2_34288_15430# a_34090_15182# 0.165f
C21815 col_n[6] a_2275_3158# 0.113f
C21816 vcm a_4274_17230# 0.155f
C21817 rowon_n[14] a_2874_16186# 0.118f
C21818 m3_20940_1078# a_20034_1126# 0.0341f
C21819 VDD a_1957_7174# 0.196f
C21820 col_n[31] a_33998_7150# 0.0765f
C21821 rowoff_n[5] a_13406_7512# 0.0133f
C21822 ctop a_17022_12170# 4.11f
C21823 a_4882_18194# a_4974_18194# 0.0991f
C21824 a_3878_18194# a_4274_18234# 0.0313f
C21825 a_2275_18218# a_5278_18234# 0.145f
C21826 row_n[0] a_13918_2130# 0.0437f
C21827 VDD a_25966_17190# 0.181f
C21828 col_n[4] a_7286_9198# 0.084f
C21829 col[0] a_2966_7150# 0.367f
C21830 a_33998_2130# a_34090_2130# 0.326f
C21831 rowon_n[4] a_13006_6146# 0.248f
C21832 col_n[21] a_2475_13198# 0.0531f
C21833 col_n[26] a_2475_2154# 0.0531f
C21834 a_2275_6170# a_20034_6146# 0.399f
C21835 m2_34864_9982# vcm 0.408f
C21836 row_n[2] a_1957_4162# 0.187f
C21837 rowoff_n[3] a_22442_5504# 0.0133f
C21838 vcm a_31990_12170# 0.1f
C21839 col_n[15] a_18426_3496# 0.0283f
C21840 a_5978_11166# a_5978_10162# 0.843f
C21841 VDD a_28066_2130# 0.483f
C21842 m2_16216_17438# row_n[15] 0.0128f
C21843 m2_6176_17438# a_5978_17190# 0.165f
C21844 m2_22240_13422# row_n[11] 0.0128f
C21845 m2_28264_9406# row_n[7] 0.0128f
C21846 col_n[25] a_28466_15544# 0.0283f
C21847 m2_34288_5390# row_n[3] 0.0128f
C21848 col_n[0] rowon_n[15] 0.111f
C21849 sample row_n[15] 0.423f
C21850 vcm col_n[31] 1.95f
C21851 VDD rowon_n[14] 3.04f
C21852 VDD a_17422_11528# 0.0779f
C21853 col[11] a_2475_10186# 0.136f
C21854 col[18] rowoff_n[15] 0.0901f
C21855 m2_34864_17010# m3_34996_16138# 0.0341f
C21856 col[25] col[26] 0.0414f
C21857 ctop a_32082_16186# 4.11f
C21858 col_n[1] rowoff_n[11] 0.0471f
C21859 a_2475_3158# a_12914_3134# 0.264f
C21860 a_2275_3158# a_10298_3174# 0.144f
C21861 rowoff_n[8] a_14010_10162# 0.294f
C21862 rowoff_n[1] a_31478_3496# 0.0133f
C21863 a_26058_1126# a_2475_1150# 0.0299f
C21864 m2_3164_5390# a_2966_5142# 0.165f
C21865 row_n[13] a_24050_15182# 0.282f
C21866 rowoff_n[11] a_17934_13174# 0.202f
C21867 a_2275_8178# a_35094_8154# 0.0924f
C21868 a_18938_8154# a_19430_8516# 0.0658f
C21869 a_18026_8154# a_18330_8194# 0.0931f
C21870 m2_25252_13422# a_25054_13174# 0.165f
C21871 col_n[18] a_2275_16210# 0.113f
C21872 col[5] a_7894_9158# 0.0682f
C21873 vcm a_12914_15182# 0.1f
C21874 a_30074_13174# a_31078_13174# 0.843f
C21875 VDD a_8990_5142# 0.483f
C21876 col_n[23] a_2275_5166# 0.113f
C21877 row_n[3] a_34090_5142# 0.282f
C21878 col_n[13] a_16018_3134# 0.251f
C21879 row_n[15] a_11302_17230# 0.0117f
C21880 m2_13780_18014# col[11] 0.347f
C21881 rowon_n[7] a_33998_9158# 0.118f
C21882 a_2275_17214# a_13918_17190# 0.136f
C21883 col_n[23] a_26058_15182# 0.251f
C21884 rowoff_n[6] a_23046_8154# 0.294f
C21885 VDD a_32482_15544# 0.0779f
C21886 col_n[20] a_22954_5142# 0.0765f
C21887 col_n[30] a_32994_17190# 0.0765f
C21888 a_2275_5166# a_25358_5182# 0.144f
C21889 a_14922_5142# a_15014_5142# 0.326f
C21890 row_n[5] a_21342_7190# 0.0117f
C21891 a_2475_5166# a_27974_5142# 0.264f
C21892 col[8] a_2275_13198# 0.0899f
C21893 m3_8892_1078# m3_9896_1078# 0.202f
C21894 col[13] a_2275_2154# 0.0899f
C21895 rowoff_n[15] a_33998_17190# 0.202f
C21896 rowoff_n[4] a_32082_6146# 0.294f
C21897 a_2475_14202# a_5978_14178# 0.316f
C21898 m2_20808_946# a_2275_1150# 0.28f
C21899 a_21038_15182# a_21038_14178# 0.843f
C21900 a_2966_14178# a_3270_14218# 0.0931f
C21901 a_3878_14178# a_4370_14540# 0.0658f
C21902 col_n[4] a_7382_1488# 0.0283f
C21903 VDD a_24050_9158# 0.483f
C21904 row_n[7] a_11910_9158# 0.0437f
C21905 rowon_n[11] a_10998_13174# 0.248f
C21906 col_n[14] a_17422_13536# 0.0283f
C21907 col[28] a_2475_12194# 0.136f
C21908 VDD a_13406_18556# 0.0858f
C21909 a_2275_2154# a_18938_2130# 0.136f
C21910 a_9902_2130# a_10298_2170# 0.0313f
C21911 m2_13780_946# VDD 1f
C21912 vcm a_30074_4138# 0.56f
C21913 rowon_n[1] a_21038_3134# 0.248f
C21914 m2_16216_11414# a_16018_11166# 0.165f
C21915 a_33998_12170# a_34490_12532# 0.0658f
C21916 a_33086_12170# a_33390_12210# 0.0931f
C21917 m2_8760_18014# a_8898_18194# 0.225f
C21918 m2_1732_11990# VDD 0.856f
C21919 a_10998_16186# a_12002_16186# 0.843f
C21920 a_2475_16210# a_21038_16186# 0.316f
C21921 VDD a_4974_12170# 0.483f
C21922 col_n[28] a_31382_2170# 0.084f
C21923 col_n[12] a_15014_13174# 0.251f
C21924 a_2275_4162# a_33998_4138# 0.136f
C21925 col_n[9] a_11910_3134# 0.0765f
C21926 m2_29844_18014# col_n[27] 0.243f
C21927 m2_34864_6970# a_35094_7150# 0.0249f
C21928 vcm a_10998_7150# 0.56f
C21929 col[25] a_2275_15206# 0.0899f
C21930 col_n[19] a_21950_15182# 0.0765f
C21931 a_29982_9158# a_30074_9158# 0.326f
C21932 rowoff_n[12] a_5886_14178# 0.202f
C21933 col[30] a_2275_4162# 0.0899f
C21934 row_n[10] a_32082_12170# 0.282f
C21935 a_2275_13198# a_12002_13174# 0.399f
C21936 rowon_n[14] a_31990_16186# 0.118f
C21937 VDD a_20034_16186# 0.483f
C21938 row_n[12] a_19334_14218# 0.0117f
C21939 col_n[3] a_6378_11528# 0.0283f
C21940 rowon_n[9] rowoff_n[9] 20.2f
C21941 vcm a_2275_1150# 7.17f
C21942 a_24962_6146# a_25358_6186# 0.0313f
C21943 m2_7180_9406# a_6982_9158# 0.165f
C21944 col_n[21] a_2475_18218# 0.0529f
C21945 vcm a_26058_11166# 0.56f
C21946 row_n[2] a_29374_4178# 0.0117f
C21947 a_2874_10162# a_3366_10524# 0.0658f
C21948 a_2275_10186# a_3878_10162# 0.136f
C21949 a_2475_10186# a_4882_10162# 0.264f
C21950 col[29] a_31990_2130# 0.0682f
C21951 VDD a_22954_1126# 0.405f
C21952 row_n[14] a_9902_16186# 0.0437f
C21953 ctop a_2966_5142# 4.06f
C21954 col_n[15] a_2475_11190# 0.0531f
C21955 a_14922_15182# a_15414_15544# 0.0658f
C21956 a_14010_15182# a_14314_15222# 0.0931f
C21957 a_2275_15206# a_27062_15182# 0.399f
C21958 m2_34864_13998# m3_34996_13126# 0.0341f
C21959 row_n[4] a_19942_6146# 0.0437f
C21960 a_21038_3134# a_22042_3134# 0.843f
C21961 rowon_n[8] a_19030_10162# 0.248f
C21962 m2_26256_5390# a_26058_5142# 0.165f
C21963 vcm a_16322_5182# 0.155f
C21964 col_n[27] a_30378_12210# 0.084f
C21965 col_n[1] a_3970_11166# 0.251f
C21966 m2_6176_16434# rowon_n[14] 0.0322f
C21967 col[5] a_2475_8178# 0.136f
C21968 m2_12200_12418# rowon_n[10] 0.0322f
C21969 m2_18224_8402# rowon_n[6] 0.0322f
C21970 vcm a_6982_14178# 0.56f
C21971 m2_24248_4386# rowon_n[2] 0.0322f
C21972 a_2475_12194# a_19942_12170# 0.264f
C21973 a_10906_12170# a_10998_12170# 0.326f
C21974 col_n[8] a_10906_13174# 0.0765f
C21975 a_2275_12194# a_17326_12210# 0.144f
C21976 VDD a_3366_4500# 0.0779f
C21977 m2_33284_18442# VDD 0.0456f
C21978 col_n[28] rowoff_n[10] 0.0471f
C21979 rowoff_n[0] a_3878_2130# 0.202f
C21980 col_n[12] a_2275_14202# 0.113f
C21981 a_12002_5142# a_12002_4138# 0.843f
C21982 col_n[17] a_2275_3158# 0.113f
C21983 vcm a_31382_9198# 0.155f
C21984 m2_15788_18014# m2_16792_18014# 0.843f
C21985 a_5886_9158# a_6282_9198# 0.0313f
C21986 a_2275_9182# a_10906_9158# 0.136f
C21987 rowon_n[2] a_6890_4138# 0.118f
C21988 vcm a_22042_18194# 0.165f
C21989 ctop a_9994_3134# 4.11f
C21990 col[21] a_24050_10162# 0.367f
C21991 m2_33284_17438# rowon_n[15] 0.0322f
C21992 a_2275_14202# a_32386_14218# 0.144f
C21993 a_2475_14202# a_35002_14178# 0.264f
C21994 VDD a_18938_8154# 0.181f
C21995 m2_32856_946# vcm 0.352f
C21996 col[2] a_2275_11190# 0.0899f
C21997 col[28] a_30986_12170# 0.0682f
C21998 a_24962_2130# a_25454_2492# 0.0658f
C21999 a_24050_2130# a_24354_2170# 0.0931f
C22000 m2_17220_3382# a_17022_3134# 0.165f
C22001 m3_7888_1078# VDD 0.0157f
C22002 row_n[9] a_27366_11206# 0.0117f
C22003 vcm a_24962_3134# 0.1f
C22004 a_2475_6170# a_2874_6146# 0.264f
C22005 a_1957_6170# a_2275_6170# 0.158f
C22006 vcm a_12306_12210# 0.155f
C22007 rowoff_n[3] a_4882_5142# 0.202f
C22008 col_n[0] row_n[10] 0.298f
C22009 col_n[7] row_n[14] 0.298f
C22010 col_n[6] rowon_n[13] 0.111f
C22011 col_n[2] rowon_n[11] 0.111f
C22012 col_n[4] rowon_n[12] 0.111f
C22013 VDD row_n[9] 3.29f
C22014 col_n[10] rowon_n[15] 0.111f
C22015 vcm rowon_n[10] 0.65f
C22016 col_n[5] row_n[13] 0.298f
C22017 sample rowon_n[9] 0.0935f
C22018 col_n[9] row_n[15] 0.298f
C22019 col_n[1] row_n[11] 0.298f
C22020 col_n[3] row_n[12] 0.298f
C22021 col_n[8] rowon_n[14] 0.111f
C22022 a_2275_11190# a_25966_11166# 0.136f
C22023 col[22] a_2475_10186# 0.136f
C22024 VDD a_10394_2492# 0.0779f
C22025 col[29] rowoff_n[15] 0.0901f
C22026 col_n[16] a_19334_10202# 0.084f
C22027 m2_4744_18014# a_4974_17190# 0.843f
C22028 m2_27836_18014# a_27974_18194# 0.225f
C22029 ctop a_25054_7150# 4.11f
C22030 row_n[11] a_17934_13174# 0.0437f
C22031 a_25966_16186# a_26058_16186# 0.326f
C22032 VDD a_33998_12170# 0.181f
C22033 m2_1732_17010# m3_1864_18146# 0.0341f
C22034 m2_24824_18014# m3_23952_18146# 0.0341f
C22035 col_n[12] rowoff_n[11] 0.0471f
C22036 rowon_n[15] a_17022_17190# 0.248f
C22037 col_n[27] a_30474_4500# 0.0283f
C22038 rowoff_n[1] a_13918_3134# 0.202f
C22039 row_n[1] a_27974_3134# 0.0437f
C22040 col_n[29] a_2275_16210# 0.113f
C22041 vcm a_5886_6146# 0.1f
C22042 rowon_n[5] a_27062_7150# 0.248f
C22043 a_27062_9158# a_27062_8154# 0.843f
C22044 a_2475_8178# a_18026_8154# 0.316f
C22045 rowoff_n[12] a_34090_14178# 0.294f
C22046 vcm a_27366_16226# 0.155f
C22047 a_20946_13174# a_21342_13214# 0.0313f
C22048 VDD a_25454_6508# 0.0779f
C22049 ctop a_5978_10162# 4.11f
C22050 VDD a_14922_15182# 0.181f
C22051 col[10] a_13006_8154# 0.367f
C22052 rowoff_n[6] a_5374_8516# 0.0133f
C22053 col[19] a_2275_13198# 0.0899f
C22054 col[24] a_2275_2154# 0.0899f
C22055 col[17] a_19942_10162# 0.0682f
C22056 a_2275_5166# a_8990_5142# 0.399f
C22057 row_n[5] a_4974_7150# 0.282f
C22058 a_5886_5142# a_6378_5504# 0.0658f
C22059 a_4974_5142# a_5278_5182# 0.0931f
C22060 m2_27836_946# m3_28972_1078# 0.0341f
C22061 m3_1864_15134# m3_1864_14130# 0.202f
C22062 col_n[25] a_28066_4138# 0.251f
C22063 rowon_n[9] a_4882_11166# 0.118f
C22064 vcm a_20946_10162# 0.1f
C22065 a_17022_10162# a_18026_10162# 0.843f
C22066 a_2475_10186# a_33086_10162# 0.316f
C22067 rowoff_n[4] a_14410_6508# 0.0133f
C22068 m2_21812_18014# ctop 0.0422f
C22069 VDD a_6378_9520# 0.0779f
C22070 col_n[5] a_8290_8194# 0.084f
C22071 m2_34864_10986# m3_34996_10114# 0.0341f
C22072 ctop a_21038_14178# 4.11f
C22073 a_32386_1166# col_n[29] 0.084f
C22074 m2_5172_15430# row_n[13] 0.0128f
C22075 m2_11196_11414# row_n[9] 0.0128f
C22076 m2_17220_7398# row_n[5] 0.0128f
C22077 m2_23244_3382# row_n[1] 0.0128f
C22078 a_2275_7174# a_24050_7150# 0.399f
C22079 rowoff_n[2] a_23446_4500# 0.0133f
C22080 rowon_n[1] a_2966_3134# 0.248f
C22081 rowoff_n[9] a_5978_11166# 0.294f
C22082 col_n[16] a_19430_2492# 0.0283f
C22083 col_n[9] a_2475_9182# 0.0531f
C22084 m2_1732_10986# a_2475_11190# 0.139f
C22085 vcm a_34394_14218# 0.155f
C22086 col_n[26] a_29470_14540# 0.0283f
C22087 a_7986_12170# a_7986_11166# 0.843f
C22088 VDD a_32082_4138# 0.483f
C22089 a_2475_16210# a_2966_16186# 0.317f
C22090 a_2161_16210# a_2275_16210# 0.183f
C22091 VDD a_21438_13536# 0.0779f
C22092 ctop a_2475_17214# 0.0463f
C22093 row_n[8] a_25966_10162# 0.0437f
C22094 rowoff_n[0] a_32482_2492# 0.0133f
C22095 rowoff_n[7] a_15014_9158# 0.294f
C22096 rowon_n[12] a_25054_14178# 0.248f
C22097 a_2475_4162# a_16930_4138# 0.264f
C22098 a_2275_4162# a_14314_4178# 0.144f
C22099 m3_1864_9110# ctop 0.21f
C22100 m2_32280_16434# row_n[14] 0.0128f
C22101 m2_1732_17010# m2_1732_16006# 0.843f
C22102 col[6] a_8898_8154# 0.0682f
C22103 a_20034_9158# a_20338_9198# 0.0931f
C22104 a_20946_9158# a_21438_9520# 0.0658f
C22105 rowoff_n[13] a_22042_15182# 0.294f
C22106 rowon_n[2] a_35094_4138# 0.0141f
C22107 col_n[14] a_17022_2130# 0.251f
C22108 a_32994_1126# col[30] 0.0682f
C22109 vcm a_16930_17190# 0.1f
C22110 a_32082_14178# a_33086_14178# 0.843f
C22111 VDD a_13006_7150# 0.483f
C22112 rowoff_n[5] a_24050_7150# 0.294f
C22113 col_n[24] a_27062_14178# 0.251f
C22114 col_n[6] a_2275_12194# 0.113f
C22115 col_n[21] a_23958_4138# 0.0765f
C22116 row_n[6] rowoff_n[5] 0.085f
C22117 a_2275_18218# a_17934_18194# 0.136f
C22118 col_n[11] a_2275_1150# 0.113f
C22119 VDD a_1957_16210# 0.196f
C22120 col_n[31] a_33998_16186# 0.0765f
C22121 a_2275_1150# a_7894_1126# 0.136f
C22122 row_n[12] a_2874_14178# 0.0436f
C22123 col_n[4] a_7286_18234# 0.084f
C22124 vcm a_19030_2130# 0.56f
C22125 a_2475_6170# a_31990_6146# 0.264f
C22126 a_2275_6170# a_29374_6186# 0.144f
C22127 a_16930_6146# a_17022_6146# 0.326f
C22128 col[0] a_2966_16186# 0.367f
C22129 row_n[2] a_13006_4138# 0.282f
C22130 rowoff_n[3] a_33086_5142# 0.294f
C22131 col_n[26] a_2475_11190# 0.0531f
C22132 VDD a_3270_1166# 0.0149f
C22133 m2_23820_18014# a_24050_17190# 0.843f
C22134 rowon_n[6] a_12914_8154# 0.118f
C22135 col_n[15] a_18426_12532# 0.0283f
C22136 a_2475_15206# a_9994_15182# 0.316f
C22137 a_23046_16186# a_23046_15182# 0.843f
C22138 VDD a_28066_11166# 0.483f
C22139 a_11910_3134# a_12306_3174# 0.0313f
C22140 a_2275_3158# a_22954_3134# 0.136f
C22141 a_2475_18218# a_15926_18194# 0.264f
C22142 col[16] a_2475_8178# 0.136f
C22143 row_n[13] a_33390_15222# 0.0117f
C22144 vcm a_34090_6146# 0.56f
C22145 rowoff_n[11] a_28466_13536# 0.0133f
C22146 col_n[0] a_2874_8154# 0.0765f
C22147 a_33486_1488# VDD 0.0985f
C22148 col[5] a_7894_18194# 0.0682f
C22149 row_n[15] a_23958_17190# 0.0437f
C22150 a_13006_17190# a_14010_17190# 0.843f
C22151 a_2475_17214# a_25054_17190# 0.316f
C22152 col_n[23] a_2275_14202# 0.113f
C22153 VDD a_8990_14178# 0.483f
C22154 a_26058_2130# m2_26256_2378# 0.165f
C22155 col_n[13] a_16018_12170# 0.251f
C22156 col_n[28] a_2275_3158# 0.113f
C22157 col_n[10] a_12914_2130# 0.0765f
C22158 row_n[5] a_33998_7150# 0.0437f
C22159 col_n[20] a_22954_14178# 0.0765f
C22160 m2_30848_946# col[28] 0.425f
C22161 rowon_n[9] a_33086_11166# 0.248f
C22162 vcm a_15014_9158# 0.56f
C22163 rowoff_n[14] a_9994_16186# 0.294f
C22164 a_31990_10162# a_32082_10162# 0.326f
C22165 col[13] a_2275_11190# 0.0899f
C22166 a_2275_14202# a_16018_14178# 0.399f
C22167 m2_34864_7974# m3_34996_7102# 0.0341f
C22168 VDD a_24050_18194# 0.0356f
C22169 col_n[4] a_7382_10524# 0.0283f
C22170 a_2475_2154# a_30074_2130# 0.316f
C22171 a_33086_3134# a_33086_2130# 0.843f
C22172 m2_1732_2954# a_2966_3134# 0.843f
C22173 m3_3872_18146# VDD 0.0678f
C22174 col_n[17] rowon_n[13] 0.111f
C22175 sample row_n[4] 0.423f
C22176 col_n[10] row_n[10] 0.298f
C22177 col_n[1] rowon_n[5] 0.111f
C22178 col_n[18] row_n[14] 0.298f
C22179 row_n[9] a_10998_11166# 0.282f
C22180 col_n[9] rowon_n[9] 0.111f
C22181 col_n[6] row_n[8] 0.298f
C22182 col_n[3] rowon_n[6] 0.111f
C22183 col_n[19] rowon_n[14] 0.111f
C22184 col_n[16] row_n[13] 0.298f
C22185 col_n[7] rowon_n[8] 0.111f
C22186 col_n[21] rowon_n[15] 0.111f
C22187 col_n[14] row_n[12] 0.298f
C22188 col_n[8] row_n[9] 0.298f
C22189 vcm row_n[5] 0.616f
C22190 vcm a_5278_3174# 0.155f
C22191 col_n[12] row_n[11] 0.298f
C22192 col_n[26] col_n[27] 0.0102f
C22193 col_n[0] rowon_n[4] 0.111f
C22194 col_n[15] rowon_n[12] 0.111f
C22195 VDD rowon_n[3] 3.04f
C22196 col_n[20] row_n[15] 0.298f
C22197 col_n[5] rowon_n[7] 0.111f
C22198 col_n[2] row_n[6] 0.298f
C22199 col_n[11] rowon_n[10] 0.111f
C22200 col_n[4] row_n[7] 0.298f
C22201 col_n[13] rowon_n[11] 0.111f
C22202 rowoff_n[9] a_35002_11166# 0.202f
C22203 a_26970_7150# a_27366_7190# 0.0313f
C22204 m2_1732_12994# vcm 0.316f
C22205 rowon_n[13] a_10906_15182# 0.118f
C22206 vcm a_30074_13174# 0.56f
C22207 a_2475_11190# a_8898_11166# 0.264f
C22208 a_2275_11190# a_6282_11206# 0.144f
C22209 col_n[23] rowoff_n[11] 0.0471f
C22210 VDD a_26970_3134# 0.181f
C22211 a_16018_16186# a_16322_16226# 0.0931f
C22212 a_2275_16210# a_31078_16186# 0.399f
C22213 a_16930_16186# a_17422_16548# 0.0658f
C22214 rowon_n[3] a_20946_5142# 0.118f
C22215 m2_1732_9982# rowon_n[8] 0.236f
C22216 col_n[3] a_2475_7174# 0.0531f
C22217 m2_7180_6394# rowon_n[4] 0.0322f
C22218 m2_12200_2378# rowon_n[0] 0.0322f
C22219 a_23046_4138# a_24050_4138# 0.843f
C22220 col_n[2] a_4974_10162# 0.251f
C22221 row_n[1] a_8290_3174# 0.0117f
C22222 col_n[28] a_31382_11206# 0.084f
C22223 m2_34864_5966# a_2275_6170# 0.278f
C22224 vcm a_20338_7190# 0.155f
C22225 a_35002_9158# a_35398_9198# 0.0313f
C22226 rowoff_n[12] a_16418_14540# 0.0133f
C22227 col_n[9] a_11910_12170# 0.0765f
C22228 m2_31276_14426# a_31078_14178# 0.165f
C22229 vcm a_10998_16186# 0.56f
C22230 ctop a_33086_2130# 4.06f
C22231 a_2475_13198# a_23958_13174# 0.264f
C22232 a_2275_13198# a_21342_13214# 0.144f
C22233 a_12914_13174# a_13006_13174# 0.326f
C22234 VDD a_7894_6146# 0.181f
C22235 col[30] a_2275_13198# 0.0899f
C22236 row_n[12] a_31990_14178# 0.0437f
C22237 vcm a_13918_1126# 0.0989f
C22238 m2_34864_4962# m2_35292_5390# 0.165f
C22239 m2_22240_15430# rowon_n[13] 0.0322f
C22240 a_14010_6146# a_14010_5142# 0.843f
C22241 m2_28264_11414# rowon_n[9] 0.0322f
C22242 m2_34288_7398# rowon_n[5] 0.0322f
C22243 m3_4876_18146# m3_5880_18146# 0.202f
C22244 vcm a_2275_10186# 6.49f
C22245 col_n[7] rowoff_n[12] 0.0471f
C22246 a_7894_10162# a_8290_10202# 0.0313f
C22247 a_2275_10186# a_14922_10162# 0.136f
C22248 col[22] a_25054_9158# 0.367f
C22249 ctop a_14010_5142# 4.11f
C22250 a_2966_15182# a_2966_14178# 0.843f
C22251 VDD a_22954_10162# 0.181f
C22252 col[29] a_31990_11166# 0.0682f
C22253 ctop a_2966_14178# 4.06f
C22254 a_26058_3134# a_26362_3174# 0.0931f
C22255 a_26970_3134# a_27462_3496# 0.0658f
C22256 col_n[20] a_2475_9182# 0.0531f
C22257 m2_34864_4962# a_35002_5142# 0.225f
C22258 vcm a_28978_5142# 0.1f
C22259 a_3970_7150# a_4974_7150# 0.843f
C22260 rowoff_n[2] a_5886_4138# 0.202f
C22261 a_2475_7174# a_6982_7150# 0.316f
C22262 rowoff_n[10] a_22954_12170# 0.202f
C22263 col_n[17] a_20338_9198# 0.084f
C22264 m2_22240_12418# a_22042_12170# 0.165f
C22265 row_n[6] a_19030_8154# 0.282f
C22266 vcm a_16322_14218# 0.155f
C22267 a_2275_12194# a_29982_12170# 0.136f
C22268 VDD a_14410_4500# 0.0779f
C22269 rowon_n[10] a_18938_12170# 0.118f
C22270 col[5] a_2475_17214# 0.136f
C22271 ctop a_29070_9158# 4.11f
C22272 row_n[0] m2_28264_2378# 0.0128f
C22273 a_27974_17190# a_28066_17190# 0.326f
C22274 VDD a_3366_13536# 0.0779f
C22275 col[10] a_2475_6170# 0.136f
C22276 row_n[8] a_6282_10202# 0.0117f
C22277 col_n[28] a_31478_3496# 0.0283f
C22278 rowoff_n[0] a_14922_2130# 0.202f
C22279 rowon_n[0] a_28978_2130# 0.118f
C22280 m2_26832_18014# m2_27260_18442# 0.165f
C22281 vcm a_9902_8154# 0.1f
C22282 a_2475_9182# a_22042_9158# 0.316f
C22283 a_29070_10162# a_29070_9158# 0.843f
C22284 rowoff_n[13] a_4370_15544# 0.0133f
C22285 col_n[17] a_2275_12194# 0.113f
C22286 row_n[2] rowoff_n[2] 0.209f
C22287 ctop rowoff_n[9] 0.177f
C22288 vcm a_31382_18234# 0.16f
C22289 col_n[22] a_2275_1150# 0.113f
C22290 a_22954_14178# a_23350_14218# 0.0313f
C22291 VDD a_29470_8516# 0.0779f
C22292 rowoff_n[5] a_6378_7512# 0.0133f
C22293 m2_34864_4962# m3_34996_4090# 0.0341f
C22294 col[11] a_14010_7150# 0.367f
C22295 ctop a_9994_12170# 4.11f
C22296 VDD a_18938_17190# 0.181f
C22297 row_n[0] a_6890_2130# 0.0437f
C22298 col[18] a_20946_9158# 0.0682f
C22299 rowon_n[4] a_5978_6146# 0.248f
C22300 col_n[26] a_29070_3134# 0.251f
C22301 a_7894_6146# a_8386_6508# 0.0658f
C22302 col[7] a_2275_9182# 0.0899f
C22303 a_6982_6146# a_7286_6186# 0.0931f
C22304 a_2275_6170# a_13006_6146# 0.399f
C22305 m2_13204_10410# a_13006_10162# 0.165f
C22306 rowoff_n[3] a_15414_5504# 0.0133f
C22307 vcm a_24962_12170# 0.1f
C22308 a_19030_11166# a_20034_11166# 0.843f
C22309 VDD a_21038_2130# 0.483f
C22310 col_n[6] a_9294_7190# 0.084f
C22311 m2_6176_5390# row_n[3] 0.0128f
C22312 VDD a_10394_11528# 0.0779f
C22313 col[27] a_2475_8178# 0.136f
C22314 ctop a_25054_16186# 4.11f
C22315 a_2275_3158# a_3270_3174# 0.144f
C22316 a_2475_3158# a_5886_3134# 0.264f
C22317 rowoff_n[8] a_6982_10162# 0.294f
C22318 rowoff_n[1] a_24450_3496# 0.0133f
C22319 m2_32280_6394# a_32082_6146# 0.165f
C22320 row_n[13] a_17022_15182# 0.282f
C22321 rowoff_n[11] a_10906_13174# 0.202f
C22322 col_n[27] a_30474_13536# 0.0283f
C22323 a_2275_8178# a_28066_8154# 0.399f
C22324 vcm a_5886_15182# 0.1f
C22325 a_9994_13174# a_9994_12170# 0.843f
C22326 VDD a_2475_5166# 26.1f
C22327 row_n[3] a_27062_5142# 0.282f
C22328 row_n[15] a_4274_17230# 0.0117f
C22329 rowon_n[7] a_26970_9158# 0.118f
C22330 m2_21236_14426# row_n[12] 0.0128f
C22331 a_2275_17214# a_6890_17190# 0.136f
C22332 rowoff_n[6] a_16018_8154# 0.294f
C22333 VDD a_25454_15544# 0.0779f
C22334 m2_27260_10410# row_n[8] 0.0128f
C22335 m2_33284_6394# row_n[4] 0.0128f
C22336 col[0] a_2874_5142# 0.0682f
C22337 col[10] a_13006_17190# 0.367f
C22338 a_2275_5166# a_18330_5182# 0.144f
C22339 row_n[5] a_14314_7190# 0.0117f
C22340 col[7] a_9902_7150# 0.0682f
C22341 a_2475_5166# a_20946_5142# 0.264f
C22342 m2_4168_8402# a_3970_8154# 0.165f
C22343 col[24] a_2275_11190# 0.0899f
C22344 a_24962_1126# a_25054_1126# 0.0991f
C22345 a_22954_10162# a_23446_10524# 0.0658f
C22346 col_n[15] a_18026_1126# 0.303f
C22347 a_22042_10162# a_22346_10202# 0.0931f
C22348 rowoff_n[15] a_26970_17190# 0.202f
C22349 rowoff_n[4] a_25054_6146# 0.294f
C22350 col_n[25] a_28066_13174# 0.251f
C22351 m2_6752_946# a_2475_1150# 0.286f
C22352 col_n[22] a_24962_3134# 0.0765f
C22353 a_33998_15182# a_34394_15222# 0.0313f
C22354 VDD a_17022_9158# 0.483f
C22355 row_n[7] a_4882_9158# 0.0437f
C22356 rowon_n[11] a_3970_13174# 0.248f
C22357 col_n[11] row_n[5] 0.298f
C22358 col_n[26] rowon_n[12] 0.111f
C22359 col_n[31] row_n[15] 0.298f
C22360 col_n[17] row_n[8] 0.298f
C22361 col_n[21] row_n[10] 0.298f
C22362 vcm sw 0.0365f
C22363 col_n[3] row_n[1] 0.298f
C22364 col_n[1] row_n[0] 0.297f
C22365 col_n[25] row_n[12] 0.298f
C22366 col_n[7] row_n[3] 0.298f
C22367 col_n[15] row_n[7] 0.298f
C22368 col_n[18] rowon_n[8] 0.111f
C22369 col_n[22] rowon_n[10] 0.111f
C22370 col_n[6] rowon_n[2] 0.111f
C22371 col_n[16] rowon_n[7] 0.111f
C22372 col_n[30] rowon_n[14] 0.111f
C22373 col_n[9] row_n[4] 0.298f
C22374 col_n[24] rowon_n[11] 0.111f
C22375 col_n[29] row_n[14] 0.298f
C22376 VDD a_6378_18556# 0.0858f
C22377 col_n[10] rowon_n[4] 0.111f
C22378 col_n[28] rowon_n[13] 0.111f
C22379 col_n[13] row_n[6] 0.298f
C22380 col_n[2] rowon_n[0] 0.111f
C22381 col_n[8] rowon_n[3] 0.111f
C22382 VDD en_C0_n 0.206f
C22383 col_n[12] rowon_n[5] 0.111f
C22384 col_n[27] row_n[13] 0.298f
C22385 col_n[19] row_n[9] 0.298f
C22386 col_n[4] rowon_n[1] 0.111f
C22387 col_n[23] row_n[11] 0.298f
C22388 col_n[14] rowon_n[6] 0.111f
C22389 col_n[20] rowon_n[9] 0.111f
C22390 col_n[5] row_n[2] 0.298f
C22391 col_n[5] a_8290_17230# 0.084f
C22392 a_2275_2154# a_11910_2130# 0.136f
C22393 m2_23244_4386# a_23046_4138# 0.165f
C22394 vcm a_23046_4138# 0.56f
C22395 rowoff_n[2] a_34090_4138# 0.294f
C22396 rowon_n[1] a_14010_3134# 0.248f
C22397 a_18938_7150# a_19030_7150# 0.326f
C22398 a_2275_7174# a_33390_7190# 0.144f
C22399 col_n[16] a_19430_11528# 0.0283f
C22400 m2_3740_18014# a_3970_18194# 0.0249f
C22401 col_n[14] a_2475_7174# 0.0531f
C22402 a_2475_16210# a_14010_16186# 0.316f
C22403 a_25054_17190# a_25054_16186# 0.843f
C22404 VDD a_32082_13174# 0.483f
C22405 rowon_n[3] a_2275_5166# 1.79f
C22406 a_22346_1166# m2_21812_946# 0.087f
C22407 a_2275_4162# a_26970_4138# 0.136f
C22408 a_13918_4138# a_14314_4178# 0.0313f
C22409 m3_27968_1078# ctop 0.21f
C22410 vcm a_3970_7150# 0.56f
C22411 col[4] a_2475_4162# 0.136f
C22412 row_n[10] a_25054_12170# 0.282f
C22413 col[6] a_8898_17190# 0.0682f
C22414 rowon_n[14] a_24962_16186# 0.118f
C22415 a_3878_13174# a_3970_13174# 0.326f
C22416 a_2275_13198# a_4974_13174# 0.399f
C22417 a_2874_13174# a_3270_13214# 0.0313f
C22418 col_n[14] a_17022_11166# 0.251f
C22419 col_n[11] a_13918_1126# 0.0765f
C22420 row_n[0] a_35094_2130# 0.0123f
C22421 VDD a_13006_16186# 0.483f
C22422 a_2475_1150# a_19030_1126# 0.31f
C22423 row_n[12] a_12306_14218# 0.0117f
C22424 col_n[21] a_23958_13174# 0.0765f
C22425 rowon_n[4] a_35002_6146# 0.118f
C22426 col_n[11] a_2275_10186# 0.113f
C22427 col_n[18] rowoff_n[12] 0.0471f
C22428 vcm a_28370_2170# 0.155f
C22429 vcm a_19030_11166# 0.56f
C22430 row_n[2] a_22346_4178# 0.0117f
C22431 a_33998_11166# a_34090_11166# 0.326f
C22432 VDD a_15926_1126# 0.405f
C22433 row_n[14] a_2161_16210# 0.0221f
C22434 a_2275_15206# a_20034_15182# 0.399f
C22435 col_n[5] a_8386_9520# 0.0283f
C22436 col_n[31] a_2475_9182# 0.0531f
C22437 col[1] a_2275_7174# 0.0899f
C22438 row_n[4] a_12914_6146# 0.0437f
C22439 a_2475_3158# a_34090_3134# 0.316f
C22440 rowon_n[8] a_12002_10162# 0.248f
C22441 vcm a_9294_5182# 0.155f
C22442 a_28978_8154# a_29374_8194# 0.0313f
C22443 m2_33860_946# sw_n 0.535f
C22444 col[16] a_2475_17214# 0.136f
C22445 vcm a_34090_15182# 0.56f
C22446 col[21] a_2475_6170# 0.136f
C22447 a_2275_12194# a_10298_12210# 0.144f
C22448 a_2475_12194# a_12914_12170# 0.264f
C22449 VDD a_30986_5142# 0.181f
C22450 col_n[0] a_2874_17190# 0.0765f
C22451 m2_19228_18442# VDD 0.0456f
C22452 a_18938_17190# a_19430_17552# 0.0658f
C22453 a_2275_17214# a_35094_17190# 0.0924f
C22454 a_18026_17190# a_18330_17230# 0.0931f
C22455 a_35002_2130# m2_34864_1950# 0.225f
C22456 col_n[2] rowoff_n[13] 0.0471f
C22457 col_n[3] a_5978_9158# 0.251f
C22458 col_n[29] a_32386_10202# 0.084f
C22459 a_25054_5142# a_26058_5142# 0.843f
C22460 col_n[28] a_2275_12194# 0.113f
C22461 col_n[10] a_12914_11166# 0.0765f
C22462 col[5] rowoff_n[9] 0.0901f
C22463 col[3] rowoff_n[7] 0.0901f
C22464 col[1] rowoff_n[5] 0.0901f
C22465 col[2] rowoff_n[6] 0.0901f
C22466 col[4] rowoff_n[8] 0.0901f
C22467 col[0] rowoff_n[4] 0.0901f
C22468 m2_8760_18014# m2_9764_18014# 0.843f
C22469 vcm a_24354_9198# 0.155f
C22470 a_2874_9158# a_2966_9158# 0.326f
C22471 vcm a_15014_18194# 0.165f
C22472 m2_5172_17438# rowon_n[15] 0.0322f
C22473 a_2475_14202# a_27974_14178# 0.264f
C22474 a_2275_14202# a_25358_14218# 0.144f
C22475 a_14922_14178# a_15014_14178# 0.326f
C22476 m2_11196_13422# rowon_n[11] 0.0322f
C22477 row_n[7] a_33086_9158# 0.282f
C22478 VDD a_11910_8154# 0.181f
C22479 m2_17220_9406# rowon_n[7] 0.0322f
C22480 m2_23244_5390# rowon_n[3] 0.0322f
C22481 rowon_n[11] a_32994_13174# 0.118f
C22482 VDD a_33390_18234# 0.019f
C22483 col[18] a_2275_9182# 0.0899f
C22484 vcm a_17934_3134# 0.1f
C22485 row_n[9] a_20338_11206# 0.0117f
C22486 a_16018_7150# a_16018_6146# 0.843f
C22487 col_n[1] a_3878_9158# 0.0765f
C22488 col[23] a_26058_8154# 0.367f
C22489 vcm a_5278_12210# 0.155f
C22490 a_2275_11190# a_18938_11166# 0.136f
C22491 a_9902_11166# a_10298_11206# 0.0313f
C22492 m2_22816_18014# a_23046_18194# 0.0249f
C22493 col[30] a_32994_10162# 0.0682f
C22494 ctop a_18026_7150# 4.11f
C22495 row_n[11] a_10906_13174# 0.0437f
C22496 VDD a_26970_12170# 0.181f
C22497 m2_14784_18014# m3_15920_18146# 0.0341f
C22498 rowon_n[15] a_9994_17190# 0.248f
C22499 a_28978_4138# a_29470_4500# 0.0658f
C22500 a_28066_4138# a_28370_4178# 0.0931f
C22501 rowoff_n[1] a_6890_3134# 0.202f
C22502 row_n[1] a_20946_3134# 0.0437f
C22503 col_n[3] a_2475_16210# 0.0531f
C22504 col_n[18] a_21342_8194# 0.084f
C22505 vcm a_32994_7150# 0.1f
C22506 rowon_n[5] a_20034_7150# 0.248f
C22507 col_n[8] a_2475_5166# 0.0531f
C22508 a_2475_8178# a_10998_8154# 0.316f
C22509 rowoff_n[12] a_27062_14178# 0.294f
C22510 a_5978_8154# a_6982_8154# 0.843f
C22511 vcm a_20338_16226# 0.155f
C22512 a_2275_13198# a_33998_13174# 0.136f
C22513 VDD a_18426_6508# 0.0779f
C22514 ctop a_33086_11166# 4.11f
C22515 a_29982_18194# a_30074_18194# 0.0991f
C22516 m3_34996_9110# a_34090_9158# 0.0303f
C22517 col_n[29] a_32482_2492# 0.0283f
C22518 VDD a_7894_15182# 0.181f
C22519 a_1957_5166# a_2161_5166# 0.115f
C22520 a_2475_5166# a_2275_5166# 2.76f
C22521 vcm a_13918_10162# 0.1f
C22522 a_2475_10186# a_26058_10162# 0.316f
C22523 a_31078_11166# a_31078_10162# 0.843f
C22524 row_n[14] a_31078_16186# 0.282f
C22525 rowoff_n[4] a_7382_6508# 0.0133f
C22526 col[12] a_15014_6146# 0.367f
C22527 col_n[1] col[2] 7.13f
C22528 col_n[12] row_n[0] 0.298f
C22529 col_n[27] rowon_n[7] 0.111f
C22530 col_n[31] rowon_n[9] 0.111f
C22531 col_n[19] rowon_n[3] 0.111f
C22532 col_n[23] rowon_n[5] 0.111f
C22533 col_n[15] rowon_n[1] 0.111f
C22534 col_n[18] row_n[3] 0.298f
C22535 vcm col[3] 5.46f
C22536 col_n[20] row_n[4] 0.298f
C22537 col_n[24] row_n[6] 0.298f
C22538 col_n[9] ctop 0.0594f
C22539 col_n[22] row_n[5] 0.298f
C22540 col_n[17] rowon_n[2] 0.111f
C22541 col_n[16] row_n[2] 0.298f
C22542 a_24962_15182# a_25358_15222# 0.0313f
C22543 col_n[21] rowon_n[4] 0.111f
C22544 col_n[28] row_n[8] 0.298f
C22545 col_n[13] rowon_n[0] 0.111f
C22546 col_n[26] row_n[7] 0.298f
C22547 col_n[29] rowon_n[8] 0.111f
C22548 col_n[25] rowon_n[6] 0.111f
C22549 col_n[14] row_n[1] 0.298f
C22550 VDD col[6] 3.83f
C22551 col_n[30] row_n[9] 0.298f
C22552 VDD a_33486_10524# 0.0779f
C22553 m2_7756_18014# ctop 0.0422f
C22554 col_n[5] a_2275_8178# 0.113f
C22555 col[19] a_21950_8154# 0.0682f
C22556 ctop a_14010_14178# 4.11f
C22557 col_n[27] a_30074_2130# 0.251f
C22558 a_2275_7174# a_17022_7150# 0.399f
C22559 rowoff_n[2] a_16418_4500# 0.0133f
C22560 rowoff_n[10] a_33486_12532# 0.0133f
C22561 a_9902_7150# a_10394_7512# 0.0658f
C22562 a_8990_7150# a_9294_7190# 0.0931f
C22563 col_n[25] a_2475_7174# 0.0531f
C22564 row_n[6] a_28370_8194# 0.0117f
C22565 vcm a_28978_14178# 0.1f
C22566 col_n[7] a_10298_6186# 0.084f
C22567 a_21038_12170# a_22042_12170# 0.843f
C22568 VDD a_25054_4138# 0.483f
C22569 col_n[17] a_20338_18234# 0.084f
C22570 VDD a_14410_13536# 0.0779f
C22571 row_n[8] a_18938_10162# 0.0437f
C22572 rowoff_n[0] a_25454_2492# 0.0133f
C22573 rowoff_n[7] a_7986_9158# 0.294f
C22574 col[10] a_2475_15206# 0.136f
C22575 rowon_n[12] a_18026_14178# 0.248f
C22576 a_2475_4162# a_9902_4138# 0.264f
C22577 a_2275_4162# a_7286_4178# 0.144f
C22578 a_5886_4138# a_5978_4138# 0.326f
C22579 m3_23952_18146# ctop 0.209f
C22580 col_n[28] a_31478_12532# 0.0283f
C22581 col[15] a_2475_4162# 0.136f
C22582 m2_4168_16434# row_n[14] 0.0128f
C22583 m2_10192_12418# row_n[10] 0.0128f
C22584 rowoff_n[13] a_15014_15182# 0.294f
C22585 a_2275_9182# a_32082_9158# 0.399f
C22586 m2_16216_8402# row_n[6] 0.0128f
C22587 m2_22240_4386# row_n[2] 0.0128f
C22588 rowon_n[2] a_28066_4138# 0.248f
C22589 vcm a_9902_17190# 0.1f
C22590 a_12002_14178# a_12002_13174# 0.843f
C22591 VDD a_5978_7150# 0.483f
C22592 rowoff_n[5] a_17022_7150# 0.294f
C22593 col[1] a_3970_4138# 0.367f
C22594 a_5886_18194# a_6282_18234# 0.0313f
C22595 col_n[29] rowoff_n[12] 0.0471f
C22596 col_n[22] a_2275_10186# 0.113f
C22597 a_2275_18218# a_10906_18194# 0.136f
C22598 VDD a_29470_17552# 0.0779f
C22599 col[11] a_14010_16186# 0.367f
C22600 col[8] a_10906_6146# 0.0682f
C22601 m2_34864_2954# a_34090_3134# 0.843f
C22602 vcm a_12002_2130# 0.56f
C22603 col[18] a_20946_18194# 0.0682f
C22604 a_2475_6170# a_24962_6146# 0.264f
C22605 a_2275_6170# a_22346_6186# 0.144f
C22606 rowoff_n[3] a_26058_5142# 0.294f
C22607 col_n[26] a_29070_12170# 0.251f
C22608 row_n[2] a_5978_4138# 0.282f
C22609 a_24962_11166# a_25454_11528# 0.0658f
C22610 col[7] a_2275_18218# 0.0899f
C22611 a_24050_11166# a_24354_11206# 0.0931f
C22612 m2_31276_17438# row_n[15] 0.0128f
C22613 col_n[23] a_25966_2130# 0.0765f
C22614 rowon_n[6] a_5886_8154# 0.118f
C22615 m2_9188_17438# a_8990_17190# 0.165f
C22616 col[12] a_2275_7174# 0.0899f
C22617 a_2475_15206# a_2874_15182# 0.264f
C22618 a_1957_15206# a_2275_15206# 0.158f
C22619 VDD a_21038_11166# 0.483f
C22620 col_n[6] a_9294_16226# 0.084f
C22621 a_2275_3158# a_15926_3134# 0.136f
C22622 a_2475_18218# a_8898_18194# 0.264f
C22623 col[27] a_2475_17214# 0.136f
C22624 rowoff_n[1] a_35094_3134# 0.0135f
C22625 en_bit_n[2] a_18938_1126# 0.0724f
C22626 a_29070_1126# a_2275_1150# 0.0924f
C22627 row_n[13] a_26362_15222# 0.0117f
C22628 vcm a_27062_6146# 0.56f
C22629 rowoff_n[11] a_21438_13536# 0.0133f
C22630 a_20946_8154# a_21038_8154# 0.326f
C22631 m2_28264_13422# a_28066_13174# 0.165f
C22632 col_n[17] a_20434_10524# 0.0283f
C22633 m2_2736_1950# ctop 0.0845f
C22634 col_n[13] rowoff_n[13] 0.0471f
C22635 a_26458_1488# VDD 0.0977f
C22636 row_n[15] a_16930_17190# 0.0437f
C22637 a_2475_17214# a_18026_17190# 0.316f
C22638 VDD a_2475_14202# 26.1f
C22639 col_n[2] a_2475_3158# 0.0531f
C22640 col[11] rowoff_n[4] 0.0901f
C22641 col[12] rowoff_n[5] 0.0901f
C22642 col[10] rowoff_n[3] 0.0901f
C22643 col[7] rowoff_n[0] 0.0901f
C22644 col[14] rowoff_n[7] 0.0901f
C22645 col[16] rowoff_n[9] 0.0901f
C22646 col[8] rowoff_n[1] 0.0901f
C22647 col[13] rowoff_n[6] 0.0901f
C22648 col[15] rowoff_n[8] 0.0901f
C22649 col[9] rowoff_n[2] 0.0901f
C22650 col[0] a_2874_14178# 0.0682f
C22651 a_15926_5142# a_16322_5182# 0.0313f
C22652 row_n[5] a_26970_7150# 0.0437f
C22653 a_2275_5166# a_30986_5142# 0.136f
C22654 rowon_n[9] a_26058_11166# 0.248f
C22655 vcm a_7986_9158# 0.56f
C22656 rowoff_n[14] a_2874_16186# 0.202f
C22657 col[7] a_9902_16186# 0.0682f
C22658 col_n[15] a_18026_10162# 0.251f
C22659 m2_33860_946# a_34090_2130# 0.752f
C22660 m2_29844_946# a_2475_1150# 0.286f
C22661 a_5886_14178# a_6378_14540# 0.0658f
C22662 a_2275_14202# a_8990_14178# 0.399f
C22663 a_4974_14178# a_5278_14218# 0.0931f
C22664 col[29] a_2275_9182# 0.0899f
C22665 col_n[22] a_24962_12170# 0.0765f
C22666 VDD a_17022_18194# 0.0356f
C22667 a_2475_2154# a_23046_2130# 0.316f
C22668 a_12002_2130# a_13006_2130# 0.843f
C22669 m2_22816_946# VDD 1f
C22670 vcm a_32386_4178# 0.155f
C22671 row_n[9] a_3970_11166# 0.282f
C22672 rowoff_n[9] a_27974_11166# 0.202f
C22673 m2_19228_11414# a_19030_11166# 0.165f
C22674 col_n[0] a_2275_6170# 0.113f
C22675 vcm a_23046_13174# 0.56f
C22676 VDD a_19942_3134# 0.181f
C22677 VDD rowoff_n[14] 1.51f
C22678 m2_9764_18014# a_10298_18234# 0.087f
C22679 m2_27836_18014# a_2275_18218# 0.28f
C22680 col_n[6] a_9390_8516# 0.0283f
C22681 a_2275_16210# a_24050_16186# 0.399f
C22682 rowon_n[3] a_13918_5142# 0.118f
C22683 col[0] rowoff_n[10] 0.0901f
C22684 a_33486_1488# col_n[30] 0.0283f
C22685 col_n[14] a_2475_16210# 0.0531f
C22686 col_n[19] a_2475_5166# 0.0531f
C22687 m2_14784_946# col[12] 0.425f
C22688 row_n[1] a_2275_3158# 19.2f
C22689 vcm a_13310_7190# 0.155f
C22690 rowon_n[5] a_1957_7174# 0.0172f
C22691 rowoff_n[12] a_9390_14540# 0.0133f
C22692 a_30986_9158# a_31382_9198# 0.0313f
C22693 row_n[10] a_35398_12210# 0.0117f
C22694 ctop a_26058_2130# 4.06f
C22695 vcm a_3970_16186# 0.56f
C22696 a_2475_13198# a_16930_13174# 0.264f
C22697 a_2275_13198# a_14314_13214# 0.144f
C22698 VDD a_35002_7150# 0.258f
C22699 col[4] a_2475_13198# 0.136f
C22700 col[9] a_2475_2154# 0.136f
C22701 m2_23820_18014# a_2475_18218# 0.286f
C22702 a_20946_18194# a_21438_18556# 0.0658f
C22703 col_n[4] a_6982_8154# 0.251f
C22704 col_n[30] a_33390_9198# 0.084f
C22705 a_15926_1126# a_16418_1488# 0.0658f
C22706 row_n[12] a_24962_14178# 0.0437f
C22707 col_n[11] a_13918_10162# 0.0765f
C22708 vcm a_6890_1126# 0.0989f
C22709 a_27062_6146# a_28066_6146# 0.843f
C22710 m2_6176_7398# rowon_n[5] 0.0322f
C22711 m2_12200_3382# rowon_n[1] 0.0322f
C22712 m2_10192_9406# a_9994_9158# 0.165f
C22713 col_n[28] rowon_n[2] 0.111f
C22714 col_n[24] rowon_n[0] 0.111f
C22715 VDD col[17] 3.83f
C22716 vcm col[14] 5.46f
C22717 col_n[27] row_n[2] 0.298f
C22718 col_n[30] rowon_n[3] 0.111f
C22719 col_n[20] ctop 0.0594f
C22720 col_n[7] col[7] 0.489f
C22721 col_n[23] row_n[0] 0.298f
C22722 vcm a_28370_11206# 0.155f
C22723 col_n[26] rowon_n[1] 0.111f
C22724 col_n[31] row_n[4] 0.298f
C22725 col_n[25] row_n[1] 0.298f
C22726 col_n[29] row_n[3] 0.298f
C22727 row_n[2] a_35002_4138# 0.0437f
C22728 rowon_n[10] rowon_n[9] 0.0632f
C22729 m2_7756_18014# col[5] 0.347f
C22730 a_2275_10186# a_7894_10162# 0.136f
C22731 col_n[16] a_2275_8178# 0.113f
C22732 rowon_n[6] a_34090_8154# 0.248f
C22733 ctop a_6982_5142# 4.11f
C22734 a_2475_15206# a_31990_15182# 0.264f
C22735 a_16930_15182# a_17022_15182# 0.326f
C22736 a_2275_15206# a_29374_15222# 0.144f
C22737 VDD a_15926_10162# 0.181f
C22738 col_n[5] a_8386_18556# 0.0283f
C22739 col[1] a_2275_16210# 0.0899f
C22740 m2_29268_5390# a_29070_5142# 0.165f
C22741 col[24] a_27062_7150# 0.367f
C22742 col[6] a_2275_5166# 0.0899f
C22743 vcm a_21950_5142# 0.1f
C22744 rowoff_n[10] a_15926_12170# 0.202f
C22745 a_18026_8154# a_18026_7150# 0.843f
C22746 m2_21236_16434# rowon_n[14] 0.0322f
C22747 m2_27260_12418# rowon_n[10] 0.0322f
C22748 col[31] a_33998_9158# 0.0682f
C22749 row_n[6] a_12002_8154# 0.282f
C22750 m2_33284_8402# rowon_n[6] 0.0322f
C22751 vcm a_9294_14218# 0.155f
C22752 a_11910_12170# a_12306_12210# 0.0313f
C22753 a_2275_12194# a_22954_12170# 0.136f
C22754 rowon_n[10] a_11910_12170# 0.118f
C22755 VDD a_7382_4500# 0.0779f
C22756 ctop a_22042_9158# 4.11f
C22757 col[21] a_2475_15206# 0.136f
C22758 VDD a_30986_14178# 0.181f
C22759 col[26] a_2475_4162# 0.136f
C22760 rowoff_n[0] a_7894_2130# 0.202f
C22761 rowon_n[0] a_21950_2130# 0.118f
C22762 col_n[19] a_22346_7190# 0.084f
C22763 a_30074_5142# a_30378_5182# 0.0931f
C22764 a_30986_5142# a_31478_5504# 0.0658f
C22765 m2_9764_946# ctop 0.0428f
C22766 m2_19804_18014# m2_20232_18442# 0.165f
C22767 vcm a_2161_8178# 0.0169f
C22768 rowoff_n[14] a_31990_16186# 0.202f
C22769 a_2475_9182# a_15014_9158# 0.316f
C22770 a_7986_9158# a_8990_9158# 0.843f
C22771 a_26970_1126# col_n[24] 0.0765f
C22772 vcm a_24354_18234# 0.16f
C22773 VDD a_22442_8516# 0.0779f
C22774 m2_23820_18014# col_n[21] 0.243f
C22775 VDD a_11910_17190# 0.181f
C22776 a_26970_2130# a_27062_2130# 0.326f
C22777 m2_20232_3382# a_20034_3134# 0.165f
C22778 m3_22948_1078# VDD 0.0157f
C22779 row_n[9] a_32994_11166# 0.0437f
C22780 col[18] a_2275_18218# 0.0899f
C22781 a_2275_6170# a_5978_6146# 0.399f
C22782 rowon_n[13] a_32082_15182# 0.248f
C22783 col[23] a_2275_7174# 0.0899f
C22784 rowoff_n[3] a_8386_5504# 0.0133f
C22785 vcm a_17934_12170# 0.1f
C22786 col[13] a_16018_5142# 0.367f
C22787 a_33086_12170# a_33086_11166# 0.843f
C22788 col_n[1] a_3878_18194# 0.0762f
C22789 a_2475_11190# a_30074_11166# 0.316f
C22790 VDD a_14010_2130# 0.483f
C22791 col[23] a_26058_17190# 0.367f
C22792 m2_28840_18014# a_29374_18234# 0.087f
C22793 col[20] a_22954_7150# 0.0682f
C22794 a_26970_16186# a_27366_16226# 0.0313f
C22795 VDD a_2966_11166# 0.485f
C22796 m2_29844_18014# m3_28972_18146# 0.0341f
C22797 ctop a_18026_16186# 4.11f
C22798 rowoff_n[1] a_17422_3496# 0.0133f
C22799 row_n[13] a_9994_15182# 0.282f
C22800 rowoff_n[11] a_3366_13536# 0.0133f
C22801 a_2275_8178# a_21038_8154# 0.399f
C22802 col_n[8] a_11302_5182# 0.084f
C22803 a_10998_8154# a_11302_8194# 0.0931f
C22804 a_11910_8154# a_12402_8516# 0.0658f
C22805 col_n[24] rowoff_n[13] 0.0471f
C22806 col_n[18] a_21342_17230# 0.084f
C22807 vcm a_32994_16186# 0.1f
C22808 col_n[8] a_2475_14202# 0.0531f
C22809 a_23046_13174# a_24050_13174# 0.843f
C22810 VDD a_29070_6146# 0.483f
C22811 row_n[3] a_20034_5142# 0.282f
C22812 col_n[13] a_2475_3158# 0.0531f
C22813 col[23] rowoff_n[5] 0.0901f
C22814 col[26] rowoff_n[8] 0.0901f
C22815 col[20] rowoff_n[2] 0.0901f
C22816 col[19] rowoff_n[1] 0.0901f
C22817 col[25] rowoff_n[7] 0.0901f
C22818 col[27] rowoff_n[9] 0.0901f
C22819 col[24] rowoff_n[6] 0.0901f
C22820 col[22] rowoff_n[4] 0.0901f
C22821 col[21] rowoff_n[3] 0.0901f
C22822 col[18] rowoff_n[0] 0.0901f
C22823 rowon_n[7] a_19942_9158# 0.118f
C22824 a_35002_18194# a_35398_18234# 0.0313f
C22825 rowoff_n[6] a_8990_8154# 0.294f
C22826 VDD a_18426_15544# 0.0779f
C22827 m2_5172_6394# row_n[4] 0.0128f
C22828 m2_10192_2378# row_n[0] 0.0128f
C22829 col[4] a_2475_18218# 0.136f
C22830 col_n[29] a_32482_11528# 0.0283f
C22831 row_n[5] a_7286_7190# 0.0117f
C22832 a_2275_5166# a_11302_5182# 0.144f
C22833 a_2475_5166# a_13918_5142# 0.264f
C22834 a_7894_5142# a_7986_5142# 0.326f
C22835 m2_32856_946# m3_33992_1078# 0.0341f
C22836 rowoff_n[15] a_19942_17190# 0.202f
C22837 rowoff_n[4] a_18026_6146# 0.294f
C22838 a_14010_15182# a_14010_14178# 0.843f
C22839 col[2] a_4974_3134# 0.367f
C22840 VDD a_9994_9158# 0.483f
C22841 col[12] a_15014_15182# 0.367f
C22842 col[9] a_11910_5142# 0.0682f
C22843 col_n[5] a_2275_17214# 0.113f
C22844 a_2275_2154# a_4882_2130# 0.136f
C22845 col[19] a_21950_17190# 0.0682f
C22846 m2_20232_15430# row_n[13] 0.0128f
C22847 m2_26256_11414# row_n[9] 0.0128f
C22848 col_n[10] a_2275_6170# 0.113f
C22849 m2_32280_7398# row_n[5] 0.0128f
C22850 vcm a_16018_4138# 0.56f
C22851 rowon_n[1] a_6982_3134# 0.248f
C22852 a_2475_7174# a_28978_7150# 0.264f
C22853 a_2275_7174# a_26362_7190# 0.144f
C22854 col_n[8] rowoff_n[14] 0.0471f
C22855 rowoff_n[2] a_27062_4138# 0.294f
C22856 col_n[27] a_30074_11166# 0.251f
C22857 ctop m2_34864_1950# 0.0422f
C22858 a_26970_12170# a_27462_12532# 0.0658f
C22859 a_26058_12170# a_26362_12210# 0.0931f
C22860 VDD a_35398_4178# 0.0882f
C22861 col[11] rowoff_n[10] 0.0901f
C22862 col_n[25] a_2475_16210# 0.0531f
C22863 col_n[7] a_10298_15222# 0.084f
C22864 a_3970_16186# a_4974_16186# 0.843f
C22865 a_2475_16210# a_6982_16186# 0.316f
C22866 VDD a_25054_13174# 0.483f
C22867 col_n[30] a_2475_5166# 0.0531f
C22868 col[0] a_2275_3158# 0.099f
C22869 a_2275_4162# a_19942_4138# 0.136f
C22870 m3_2868_2082# ctop 0.418f
C22871 col_n[18] a_21438_9520# 0.0283f
C22872 vcm a_31078_8154# 0.56f
C22873 a_22954_9158# a_23046_9158# 0.326f
C22874 col[15] a_2475_13198# 0.136f
C22875 row_n[10] a_18026_12170# 0.282f
C22876 m2_1732_16006# sample 0.2f
C22877 col[20] a_2475_2154# 0.136f
C22878 rowon_n[14] a_17934_16186# 0.118f
C22879 m2_34864_9982# ctop 0.0422f
C22880 VDD a_5978_16186# 0.483f
C22881 row_n[0] a_28066_2130# 0.282f
C22882 a_2475_1150# a_12002_1126# 0.0299f
C22883 row_n[12] a_5278_14218# 0.0117f
C22884 rowon_n[4] a_27974_6146# 0.118f
C22885 col[1] a_3970_13174# 0.367f
C22886 rowon_n[7] row_n[7] 18.9f
C22887 vcm col[25] 5.46f
C22888 VDD col[28] 3.83f
C22889 col_n[12] col[13] 7.13f
C22890 col_n[31] ctop 0.264f
C22891 vcm a_21342_2170# 0.155f
C22892 col_n[27] a_2275_8178# 0.113f
C22893 a_17934_6146# a_18330_6186# 0.0313f
C22894 a_2275_6170# a_35002_6146# 0.136f
C22895 col[8] a_10906_15182# 0.0682f
C22896 m2_10768_946# m2_11772_946# 0.843f
C22897 row_n[2] a_15318_4178# 0.0117f
C22898 vcm a_12002_11166# 0.56f
C22899 col_n[16] a_19030_9158# 0.251f
C22900 VDD a_8898_1126# 0.405f
C22901 a_2275_15206# a_13006_15182# 0.399f
C22902 a_6982_15182# a_7286_15222# 0.0931f
C22903 a_7894_15182# a_8386_15544# 0.0658f
C22904 col_n[23] a_25966_11166# 0.0765f
C22905 col[12] a_2275_16210# 0.0899f
C22906 row_n[4] a_5886_6146# 0.0437f
C22907 col[17] a_2275_5166# 0.0899f
C22908 rowon_n[8] a_4974_10162# 0.248f
C22909 a_14010_3134# a_15014_3134# 0.843f
C22910 a_2475_3158# a_27062_3134# 0.316f
C22911 rowoff_n[8] a_28978_10162# 0.202f
C22912 vcm a_3878_5142# 0.1f
C22913 rowoff_n[11] a_32082_13174# 0.294f
C22914 m2_1732_11990# a_2161_12194# 0.0454f
C22915 vcm a_27062_15182# 0.56f
C22916 col_n[7] a_10394_7512# 0.0283f
C22917 a_2275_12194# a_3270_12210# 0.144f
C22918 a_2475_12194# a_5886_12170# 0.264f
C22919 VDD a_23958_5142# 0.181f
C22920 m2_5172_18442# VDD 0.0456f
C22921 a_2275_17214# a_28066_17190# 0.399f
C22922 a_29070_2130# m2_29268_2378# 0.165f
C22923 rowon_n[0] a_3878_2130# 0.118f
C22924 a_4974_5142# a_4974_4138# 0.843f
C22925 col_n[2] a_2475_12194# 0.0531f
C22926 col_n[7] a_2475_1150# 0.0531f
C22927 m2_1732_18014# m2_2736_18014# 0.843f
C22928 vcm a_17326_9198# 0.155f
C22929 a_32994_10162# a_33390_10202# 0.0313f
C22930 m2_34864_15002# a_2475_15206# 0.282f
C22931 ctop a_30074_4138# 4.11f
C22932 vcm a_7986_18194# 0.165f
C22933 m2_18224_1374# a_18026_1126# 0.165f
C22934 m3_21944_1078# a_22042_2130# 0.0302f
C22935 a_2475_14202# a_20946_14178# 0.264f
C22936 a_2275_14202# a_18330_14218# 0.144f
C22937 VDD a_4882_8154# 0.181f
C22938 row_n[7] a_26058_9158# 0.282f
C22939 col_n[5] a_7986_7150# 0.251f
C22940 rowon_n[11] a_25966_13174# 0.118f
C22941 col[29] a_2275_18218# 0.0899f
C22942 VDD a_26362_18234# 0.019f
C22943 col_n[12] a_14922_9158# 0.0765f
C22944 a_2275_2154# a_33086_2130# 0.399f
C22945 a_17022_2130# a_17326_2170# 0.0931f
C22946 a_17934_2130# a_18426_2492# 0.0658f
C22947 m3_18932_18146# VDD 0.0878f
C22948 vcm a_10906_3134# 0.1f
C22949 m2_1732_7974# m2_2160_8402# 0.165f
C22950 row_n[9] a_13310_11206# 0.0117f
C22951 a_29070_7150# a_30074_7150# 0.843f
C22952 vcm a_32386_13214# 0.155f
C22953 a_2275_11190# a_11910_11166# 0.136f
C22954 VDD a_30474_3496# 0.0779f
C22955 col_n[0] a_2275_15206# 0.113f
C22956 ctop a_10998_7150# 4.11f
C22957 a_18938_16186# a_19030_16186# 0.326f
C22958 a_2275_16210# a_33390_16226# 0.144f
C22959 VDD a_19942_12170# 0.181f
C22960 col_n[4] a_2275_4162# 0.113f
C22961 m2_5748_18014# m3_5880_18146# 3.79f
C22962 col_n[6] a_9390_17552# 0.0283f
C22963 rowon_n[15] a_2874_17190# 0.118f
C22964 m2_10192_14426# rowon_n[12] 0.0322f
C22965 m2_16216_10410# rowon_n[8] 0.0322f
C22966 m2_22240_6394# rowon_n[4] 0.0322f
C22967 col[25] a_28066_6146# 0.367f
C22968 row_n[14] rowoff_n[13] 0.085f
C22969 row_n[1] a_13918_3134# 0.0437f
C22970 vcm a_25966_7150# 0.1f
C22971 rowon_n[5] a_13006_7150# 0.248f
C22972 col_n[19] a_2475_14202# 0.0531f
C22973 rowoff_n[12] a_20034_14178# 0.294f
C22974 a_20034_9158# a_20034_8154# 0.843f
C22975 a_2275_8178# a_2966_8154# 0.399f
C22976 a_2475_8178# a_3970_8154# 0.316f
C22977 col_n[24] a_2475_3158# 0.0531f
C22978 m2_34288_14426# a_34090_14178# 0.165f
C22979 col[31] rowoff_n[2] 0.0901f
C22980 sample_n rowoff_n[3] 0.14f
C22981 col[30] rowoff_n[1] 0.0901f
C22982 col[29] rowoff_n[0] 0.0901f
C22983 ctop a_2275_1150# 0.125f
C22984 vcm a_13310_16226# 0.155f
C22985 a_13918_13174# a_14314_13214# 0.0313f
C22986 a_2275_13198# a_26970_13174# 0.136f
C22987 VDD a_11398_6508# 0.0779f
C22988 row_n[3] a_1957_5166# 0.187f
C22989 ctop a_26058_11166# 4.11f
C22990 col[15] a_2475_18218# 0.136f
C22991 VDD a_35002_16186# 0.257f
C22992 col_n[20] a_23350_6186# 0.084f
C22993 col[9] a_2475_11190# 0.136f
C22994 col_n[4] a_6982_17190# 0.251f
C22995 col_n[30] a_33390_18234# 0.084f
C22996 a_32082_6146# a_32386_6186# 0.0931f
C22997 a_32994_6146# a_33486_6508# 0.0658f
C22998 m2_34864_3958# rowoff_n[2] 0.278f
C22999 m2_8760_946# m3_7888_1078# 0.0341f
C23000 vcm a_6890_10162# 0.1f
C23001 a_9994_10162# a_10998_10162# 0.843f
C23002 a_2475_10186# a_19030_10162# 0.316f
C23003 row_n[14] a_24050_16186# 0.282f
C23004 m2_6176_16434# a_5978_16186# 0.165f
C23005 col_n[16] a_2275_17214# 0.113f
C23006 VDD a_26458_10524# 0.0779f
C23007 ctop a_6982_14178# 4.11f
C23008 col_n[21] a_2275_6170# 0.113f
C23009 row_n[4] a_34090_6146# 0.282f
C23010 m2_24824_946# col[22] 0.425f
C23011 col_n[19] rowoff_n[14] 0.0471f
C23012 a_28978_3134# a_29070_3134# 0.326f
C23013 rowon_n[8] a_33998_10162# 0.118f
C23014 m2_3164_4386# a_2966_4138# 0.165f
C23015 m2_34864_11990# m2_34864_10986# 0.843f
C23016 rowoff_n[2] a_9390_4500# 0.0133f
C23017 col[14] a_17022_4138# 0.367f
C23018 rowoff_n[10] a_26458_12532# 0.0133f
C23019 a_2275_7174# a_9994_7150# 0.399f
C23020 m2_22816_18014# vcm 0.353f
C23021 col[22] rowoff_n[10] 0.0901f
C23022 m2_25252_12418# a_25054_12170# 0.165f
C23023 col[24] a_27062_16186# 0.367f
C23024 row_n[6] a_21342_8194# 0.0117f
C23025 col[6] a_2275_14202# 0.0899f
C23026 vcm a_21950_14178# 0.1f
C23027 col[21] a_23958_6146# 0.0682f
C23028 a_2475_12194# a_34090_12170# 0.316f
C23029 VDD a_18026_4138# 0.483f
C23030 col[11] a_2275_3158# 0.0899f
C23031 col[31] a_33998_18194# 0.0682f
C23032 a_28978_17190# a_29374_17230# 0.0313f
C23033 VDD a_7382_13536# 0.0779f
C23034 row_n[8] a_11910_10162# 0.0437f
C23035 rowoff_n[0] a_18426_2492# 0.0133f
C23036 rowon_n[12] a_10998_14178# 0.248f
C23037 col[26] a_2475_13198# 0.136f
C23038 col_n[9] a_12306_4178# 0.084f
C23039 m2_32856_946# ctop 0.0456f
C23040 col[31] a_2475_2154# 0.136f
C23041 col_n[19] a_22346_16226# 0.084f
C23042 a_13918_9158# a_14410_9520# 0.0658f
C23043 a_13006_9158# a_13310_9198# 0.0931f
C23044 a_2275_9182# a_25054_9158# 0.399f
C23045 rowoff_n[13] a_7986_15182# 0.294f
C23046 rowon_n[2] a_21038_4138# 0.248f
C23047 vcm a_2161_17214# 0.0169f
C23048 a_25054_14178# a_26058_14178# 0.843f
C23049 VDD a_33086_8154# 0.483f
C23050 rowoff_n[5] a_9994_7150# 0.294f
C23051 col_n[3] rowoff_n[15] 0.0471f
C23052 rowon_n[10] ctop 0.203f
C23053 rowon_n[14] col[2] 0.0323f
C23054 rowon_n[13] col[0] 0.0318f
C23055 row_n[15] col[3] 0.0342f
C23056 rowon_n[15] col[4] 0.0323f
C23057 row_n[14] col[1] 0.0342f
C23058 col_n[18] col[18] 0.489f
C23059 a_2874_18194# a_2966_18194# 0.0991f
C23060 VDD a_22442_17552# 0.0779f
C23061 col_n[30] a_33486_10524# 0.0283f
C23062 vcm a_4974_2130# 0.56f
C23063 col[6] rowoff_n[11] 0.0901f
C23064 a_2275_6170# a_15318_6186# 0.144f
C23065 a_9902_6146# a_9994_6146# 0.326f
C23066 a_2475_6170# a_17934_6146# 0.264f
C23067 m2_16216_10410# a_16018_10162# 0.165f
C23068 rowoff_n[3] a_19030_5142# 0.294f
C23069 col[3] a_5978_2130# 0.367f
C23070 m2_3164_17438# row_n[15] 0.0128f
C23071 m2_9188_13422# row_n[11] 0.0128f
C23072 col[23] a_2275_16210# 0.0899f
C23073 m2_15212_9406# row_n[7] 0.0128f
C23074 m2_21236_5390# row_n[3] 0.0128f
C23075 col[13] a_16018_14178# 0.367f
C23076 col[28] a_2275_5166# 0.0899f
C23077 row_n[11] a_32082_13174# 0.282f
C23078 a_16018_16186# a_16018_15182# 0.843f
C23079 VDD a_14010_11166# 0.483f
C23080 m2_1732_946# m2_2736_946# 0.843f
C23081 col[10] a_12914_4138# 0.0682f
C23082 rowon_n[15] a_31990_17190# 0.118f
C23083 col[20] a_22954_16186# 0.0682f
C23084 a_2275_3158# a_8898_3134# 0.136f
C23085 a_4882_3134# a_5278_3174# 0.0313f
C23086 rowoff_n[1] a_28066_3134# 0.294f
C23087 col_n[28] a_31078_10162# 0.251f
C23088 m2_34864_5966# a_35094_6146# 0.0249f
C23089 row_n[13] a_19334_15222# 0.0117f
C23090 vcm a_20034_6146# 0.56f
C23091 a_2475_8178# a_32994_8154# 0.264f
C23092 a_2275_8178# a_30378_8194# 0.144f
C23093 rowoff_n[11] a_14410_13536# 0.0133f
C23094 m3_1864_1078# m2_2736_946# 0.0341f
C23095 a_28066_13174# a_28370_13214# 0.0931f
C23096 col_n[8] a_11302_14218# 0.084f
C23097 a_28978_13174# a_29470_13536# 0.0658f
C23098 row_n[3] a_29374_5182# 0.0117f
C23099 row_n[15] a_9902_17190# 0.0437f
C23100 col[1] a_3878_2130# 0.0682f
C23101 a_5978_17190# a_6982_17190# 0.843f
C23102 m2_35292_14426# row_n[12] 0.0128f
C23103 a_2475_17214# a_10998_17190# 0.316f
C23104 VDD a_29070_15182# 0.483f
C23105 col_n[13] a_2475_12194# 0.0531f
C23106 col_n[18] a_2475_1150# 0.0531f
C23107 col_n[19] a_22442_8516# 0.0283f
C23108 a_2275_5166# a_23958_5142# 0.136f
C23109 row_n[5] a_19942_7150# 0.0437f
C23110 m2_7180_8402# a_6982_8154# 0.165f
C23111 rowon_n[9] a_19030_11166# 0.248f
C23112 vcm a_35094_10162# 0.165f
C23113 a_25966_1126# a_26362_1166# 0.0313f
C23114 a_24962_10162# a_25054_10162# 0.326f
C23115 rowoff_n[15] a_30474_17552# 0.0133f
C23116 a_2475_14202# a_2275_14202# 2.76f
C23117 a_1957_14202# a_2161_14202# 0.115f
C23118 m2_4744_946# a_5278_1166# 0.087f
C23119 m2_12776_946# a_2275_1150# 0.28f
C23120 col[3] a_2475_9182# 0.136f
C23121 col[2] a_4974_12170# 0.367f
C23122 VDD a_9994_18194# 0.0356f
C23123 a_2475_2154# a_16018_2130# 0.316f
C23124 a_26058_3134# a_26058_2130# 0.843f
C23125 m2_26256_4386# a_26058_4138# 0.165f
C23126 col[9] a_11910_14178# 0.0682f
C23127 m2_7180_1374# VDD 0.0194f
C23128 vcm a_25358_4178# 0.155f
C23129 a_19942_7150# a_20338_7190# 0.0313f
C23130 rowoff_n[9] a_20946_11166# 0.202f
C23131 col_n[17] a_20034_8154# 0.251f
C23132 col_n[10] a_2275_15206# 0.113f
C23133 vcm a_16018_13174# 0.56f
C23134 col_n[15] a_2275_4162# 0.113f
C23135 VDD a_12914_3134# 0.181f
C23136 m2_13780_18014# a_2275_18218# 0.28f
C23137 col_n[24] a_26970_10162# 0.0765f
C23138 a_8990_16186# a_9294_16226# 0.0931f
C23139 a_2275_16210# a_17022_16186# 0.399f
C23140 a_9902_16186# a_10394_16548# 0.0658f
C23141 VDD a_35398_13214# 0.0882f
C23142 rowon_n[3] a_6890_5142# 0.118f
C23143 a_25966_1126# m2_25828_946# 0.225f
C23144 rowoff_n[7] a_29982_9158# 0.202f
C23145 col_n[30] a_2475_14202# 0.0531f
C23146 a_2475_4162# a_31078_4138# 0.316f
C23147 a_16018_4138# a_17022_4138# 0.843f
C23148 col[0] a_2275_12194# 0.099f
C23149 col[5] a_2275_1150# 0.0899f
C23150 vcm a_6282_7190# 0.155f
C23151 rowoff_n[12] a_1957_14202# 0.0219f
C23152 col_n[8] a_11398_6508# 0.0283f
C23153 row_n[10] a_27366_12210# 0.0117f
C23154 col[26] a_2475_18218# 0.136f
C23155 col_n[18] a_21438_18556# 0.0283f
C23156 vcm a_31078_17190# 0.56f
C23157 ctop a_19030_2130# 4.11f
C23158 a_2475_13198# a_9902_13174# 0.264f
C23159 a_5886_13174# a_5978_13174# 0.326f
C23160 a_2275_13198# a_7286_13214# 0.144f
C23161 VDD a_27974_7150# 0.181f
C23162 col[20] a_2475_11190# 0.136f
C23163 a_2275_18218# a_32082_18194# 0.0924f
C23164 m2_9764_18014# a_2475_18218# 0.286f
C23165 a_2275_1150# a_22042_1126# 0.0924f
C23166 row_n[12] a_17934_14178# 0.0437f
C23167 vcm a_33998_2130# 0.098f
C23168 a_6982_6146# a_6982_5142# 0.843f
C23169 m3_33992_1078# sw 0.0243f
C23170 vcm a_21342_11206# 0.155f
C23171 row_n[2] a_27974_4138# 0.0437f
C23172 col_n[27] a_2275_17214# 0.113f
C23173 VDD a_19430_1488# 0.0914f
C23174 rowon_n[6] a_27062_8154# 0.248f
C23175 col_n[6] a_8990_6146# 0.251f
C23176 m2_34864_4962# VDD 0.772f
C23177 ctop a_34090_6146# 4.06f
C23178 a_2475_15206# a_24962_15182# 0.264f
C23179 a_2275_15206# a_22346_15222# 0.144f
C23180 col_n[30] rowoff_n[14] 0.0471f
C23181 VDD a_8898_10162# 0.181f
C23182 col_n[13] a_15926_8154# 0.0765f
C23183 a_19942_3134# a_20434_3496# 0.0658f
C23184 a_19030_3134# a_19334_3174# 0.0931f
C23185 a_2475_18218# a_30074_18194# 0.0299f
C23186 col_n[0] m2_2736_946# 0.331f
C23187 col[17] a_2275_14202# 0.0899f
C23188 vcm a_14922_5142# 0.1f
C23189 a_31078_8154# a_32082_8154# 0.843f
C23190 rowoff_n[10] a_8898_12170# 0.202f
C23191 a_28066_1126# vcm 0.165f
C23192 col[22] a_2275_3158# 0.0899f
C23193 row_n[6] a_4974_8154# 0.282f
C23194 m2_5172_8402# rowon_n[6] 0.0322f
C23195 vcm a_3878_14178# 0.1f
C23196 a_2275_12194# a_15926_12170# 0.136f
C23197 m2_11196_4386# rowon_n[2] 0.0322f
C23198 VDD a_34490_5504# 0.0779f
C23199 rowon_n[10] a_4882_12170# 0.118f
C23200 m2_26832_18014# VDD 1.1f
C23201 ctop a_15014_9158# 4.11f
C23202 col_n[7] a_10394_16548# 0.0283f
C23203 a_20946_17190# a_21038_17190# 0.326f
C23204 VDD a_23958_14178# 0.181f
C23205 a_2966_1126# m2_2736_946# 0.0249f
C23206 col[26] a_29070_5142# 0.367f
C23207 rowon_n[0] a_14922_2130# 0.118f
C23208 m2_12776_18014# m2_13204_18442# 0.165f
C23209 vcm a_29982_9158# 0.1f
C23210 a_22042_10162# a_22042_9158# 0.843f
C23211 rowoff_n[14] a_24962_16186# 0.202f
C23212 a_2475_9182# a_7986_9158# 0.316f
C23213 rowon_n[2] a_2966_4138# 0.248f
C23214 rowon_n[12] col[9] 0.0323f
C23215 col_n[23] col[24] 7.13f
C23216 rowon_n[8] col[1] 0.0323f
C23217 row_n[9] col[2] 0.0342f
C23218 rowon_n[9] col[3] 0.0323f
C23219 col_n[7] a_2475_10186# 0.0531f
C23220 rowon_n[14] col[13] 0.0323f
C23221 row_n[11] col[6] 0.0342f
C23222 row_n[13] col[10] 0.0342f
C23223 row_n[8] col[0] 0.0322f
C23224 rowon_n[13] col[11] 0.0323f
C23225 row_n[5] ctop 0.186f
C23226 vcm a_17326_18234# 0.16f
C23227 row_n[14] col[12] 0.0342f
C23228 row_n[10] col[4] 0.0342f
C23229 row_n[15] col[14] 0.0342f
C23230 col_n[14] rowoff_n[15] 0.0471f
C23231 rowon_n[15] col[15] 0.0323f
C23232 rowon_n[11] col[7] 0.0323f
C23233 rowon_n[10] col[5] 0.0323f
C23234 row_n[12] col[8] 0.0342f
C23235 m2_20232_17438# rowon_n[15] 0.0322f
C23236 a_15926_14178# a_16322_14218# 0.0313f
C23237 a_2275_14202# a_30986_14178# 0.136f
C23238 m2_1732_12994# ctop 0.0428f
C23239 VDD a_15414_8516# 0.0779f
C23240 m2_26256_13422# rowon_n[11] 0.0322f
C23241 m2_32280_9406# rowon_n[7] 0.0322f
C23242 col_n[21] a_24354_5182# 0.084f
C23243 ctop a_30074_13174# 4.11f
C23244 VDD a_4882_17190# 0.181f
C23245 col[17] rowoff_n[11] 0.0901f
C23246 col_n[5] a_7986_16186# 0.251f
C23247 col_n[2] a_4882_6146# 0.0765f
C23248 col_n[12] a_14922_18194# 0.0762f
C23249 row_n[9] a_25966_11166# 0.0437f
C23250 a_35002_7150# a_35494_7512# 0.0658f
C23251 m2_1732_9982# a_2475_10186# 0.139f
C23252 rowon_n[13] a_25054_15182# 0.248f
C23253 vcm a_10906_12170# 0.1f
C23254 a_2475_11190# a_23046_11166# 0.316f
C23255 a_12002_11166# a_13006_11166# 0.843f
C23256 VDD a_6982_2130# 0.483f
C23257 rowon_n[3] a_35094_5142# 0.0141f
C23258 VDD a_30474_12532# 0.0779f
C23259 m2_19804_18014# m3_20940_18146# 0.0341f
C23260 ctop a_10998_16186# 4.11f
C23261 col_n[4] a_2275_13198# 0.113f
C23262 a_30986_4138# a_31078_4138# 0.326f
C23263 col_n[9] a_2275_2154# 0.113f
C23264 rowoff_n[1] a_10394_3496# 0.0133f
C23265 col[15] a_18026_3134# 0.367f
C23266 row_n[13] a_2874_15182# 0.0436f
C23267 vcm a_1957_6170# 0.139f
C23268 col[25] a_28066_15182# 0.367f
C23269 a_2275_8178# a_14010_8154# 0.399f
C23270 col[22] a_24962_5142# 0.0682f
C23271 vcm a_25966_16186# 0.1f
C23272 VDD a_22042_6146# 0.483f
C23273 col_n[24] a_2475_12194# 0.0531f
C23274 row_n[3] a_13006_5142# 0.282f
C23275 col[1] rowoff_n[12] 0.0901f
C23276 ctop a_2275_10186# 0.0683f
C23277 rowon_n[7] a_12914_9158# 0.118f
C23278 col_n[29] a_2475_1150# 0.0531f
C23279 a_30986_18194# a_31382_18234# 0.0313f
C23280 rowoff_n[6] a_2475_8178# 3.9f
C23281 VDD a_11398_15544# 0.0779f
C23282 col_n[10] a_13310_3174# 0.084f
C23283 m3_4876_18146# a_4974_17190# 0.0303f
C23284 a_2475_5166# a_6890_5142# 0.264f
C23285 col_n[20] a_23350_15222# 0.084f
C23286 a_2275_5166# a_4274_5182# 0.144f
C23287 m2_23820_946# m3_23952_1078# 3.79f
C23288 m3_33992_18146# m3_34996_18146# 0.202f
C23289 a_15926_10162# a_16418_10524# 0.0658f
C23290 a_2275_10186# a_29070_10162# 0.399f
C23291 col[14] a_2475_9182# 0.136f
C23292 rowoff_n[15] a_12914_17190# 0.202f
C23293 a_15014_10162# a_15318_10202# 0.0931f
C23294 row_n[14] a_33390_16226# 0.0117f
C23295 rowoff_n[4] a_10998_6146# 0.294f
C23296 m2_16792_946# a_17022_2130# 0.843f
C23297 a_27062_15182# a_28066_15182# 0.843f
C23298 VDD a_2874_9158# 0.182f
C23299 col_n[31] a_34490_9520# 0.0283f
C23300 col_n[21] a_2275_15206# 0.113f
C23301 m2_4168_7398# row_n[5] 0.0128f
C23302 m2_10192_3382# row_n[1] 0.0128f
C23303 vcm a_8990_4138# 0.56f
C23304 col_n[26] a_2275_4162# 0.113f
C23305 a_2275_7174# a_19334_7190# 0.144f
C23306 rowoff_n[2] a_20034_4138# 0.294f
C23307 rowoff_n[9] a_2275_11190# 0.151f
C23308 a_11910_7150# a_12002_7150# 0.326f
C23309 a_2475_7174# a_21950_7150# 0.264f
C23310 row_n[6] a_33998_8154# 0.0437f
C23311 col[14] a_17022_13174# 0.367f
C23312 rowon_n[10] a_33086_12170# 0.248f
C23313 col[11] a_13918_3134# 0.0682f
C23314 a_18026_17190# a_18026_16186# 0.843f
C23315 col[21] a_23958_15182# 0.0682f
C23316 VDD a_18026_13174# 0.483f
C23317 col[11] a_2275_12194# 0.0899f
C23318 rowoff_n[0] a_29070_2130# 0.294f
C23319 col[16] a_2275_1150# 0.0896f
C23320 col_n[29] a_32082_9158# 0.251f
C23321 a_6890_4138# a_7286_4178# 0.0313f
C23322 a_2275_4162# a_12914_4138# 0.136f
C23323 m3_34996_16138# ctop 0.209f
C23324 m2_19228_16434# row_n[14] 0.0128f
C23325 m2_25252_12418# row_n[10] 0.0128f
C23326 vcm a_24050_8154# 0.56f
C23327 a_2275_9182# a_35398_9198# 0.145f
C23328 m2_31276_8402# row_n[6] 0.0128f
C23329 col_n[9] a_12306_13214# 0.084f
C23330 row_n[10] a_10998_12170# 0.282f
C23331 col[31] a_2475_11190# 0.136f
C23332 a_30074_14178# a_30378_14218# 0.0931f
C23333 rowon_n[14] a_10906_16186# 0.118f
C23334 a_30986_14178# a_31478_14540# 0.0658f
C23335 row_n[0] a_21038_2130# 0.282f
C23336 VDD a_33086_17190# 0.484f
C23337 a_2475_1150# a_4974_1126# 0.0299f
C23338 col_n[20] a_23446_7512# 0.0283f
C23339 rowon_n[4] a_20946_6146# 0.118f
C23340 m2_2736_1950# a_2275_2154# 0.281f
C23341 vcm a_14314_2170# 0.155f
C23342 a_2275_6170# a_27974_6146# 0.136f
C23343 col_n[1] a_2475_8178# 0.0531f
C23344 m2_1732_10986# sample_n 0.0522f
C23345 row_n[2] a_8290_4178# 0.0117f
C23346 vcm a_4974_11166# 0.56f
C23347 a_26970_11166# a_27062_11166# 0.326f
C23348 m2_12200_17438# a_12002_17190# 0.165f
C23349 a_2275_15206# a_5978_15182# 0.399f
C23350 col[3] a_5978_11166# 0.367f
C23351 col[28] a_2275_14202# 0.0899f
C23352 col[10] a_12914_13174# 0.0682f
C23353 a_2475_3158# a_20034_3134# 0.316f
C23354 a_28066_4138# a_28066_3134# 0.843f
C23355 rowoff_n[8] a_21950_10162# 0.202f
C23356 m2_34864_4962# a_2275_5166# 0.278f
C23357 a_35002_1126# a_2475_1150# 0.264f
C23358 a_31382_1166# a_2275_1150# 0.145f
C23359 col_n[18] a_21038_7150# 0.251f
C23360 row_n[13] a_31990_15182# 0.0437f
C23361 vcm a_29374_6186# 0.155f
C23362 rowoff_n[11] a_25054_13174# 0.294f
C23363 a_21950_8154# a_22346_8194# 0.0313f
C23364 m2_31276_13422# a_31078_13174# 0.165f
C23365 col_n[25] a_27974_9158# 0.0765f
C23366 vcm a_20034_15182# 0.56f
C23367 VDD a_16930_5142# 0.181f
C23368 a_30074_1126# VDD 0.035f
C23369 a_2275_17214# a_21038_17190# 0.399f
C23370 a_11910_17190# a_12402_17552# 0.0658f
C23371 a_10998_17190# a_11302_17230# 0.0931f
C23372 rowoff_n[6] a_30986_8154# 0.202f
C23373 col[1] a_3878_11166# 0.0682f
C23374 a_18026_5142# a_19030_5142# 0.843f
C23375 a_2475_5166# a_35094_5142# 0.0299f
C23376 col_n[9] a_12402_5504# 0.0283f
C23377 m3_23952_1078# m3_24956_1078# 0.202f
C23378 row_n[3] col[1] 0.0342f
C23379 row_n[15] col[25] 0.0342f
C23380 rowon_n[9] col[14] 0.0323f
C23381 col_n[18] a_2475_10186# 0.0531f
C23382 rowon_n[15] col[26] 0.0323f
C23383 rowon_n[4] col[4] 0.0323f
C23384 rowon_n[13] col[22] 0.0323f
C23385 row_n[5] col[5] 0.0342f
C23386 rowon_n[14] col[24] 0.0323f
C23387 rowon_n[11] col[18] 0.0323f
C23388 row_n[4] col[3] 0.0342f
C23389 rowon_n[3] col[2] 0.0323f
C23390 row_n[14] col[23] 0.0342f
C23391 rowon_n[6] col[8] 0.0323f
C23392 rowon_n[7] col[10] 0.0323f
C23393 sw ctop 0.435f
C23394 row_n[8] col[11] 0.0342f
C23395 rowon_n[5] col[6] 0.0323f
C23396 rowon_n[12] col[20] 0.0323f
C23397 col_n[29] col[29] 0.539f
C23398 row_n[11] col[17] 0.0342f
C23399 row_n[6] col[7] 0.0342f
C23400 row_n[12] col[19] 0.0342f
C23401 col_n[25] rowoff_n[15] 0.0471f
C23402 row_n[10] col[15] 0.0342f
C23403 row_n[7] col[9] 0.0342f
C23404 rowon_n[2] col[0] 0.0318f
C23405 rowon_n[8] col[12] 0.0323f
C23406 rowon_n[10] col[16] 0.0323f
C23407 row_n[13] col[21] 0.0342f
C23408 row_n[9] col[13] 0.0342f
C23409 col_n[19] a_22442_17552# 0.0283f
C23410 vcm a_10298_9198# 0.155f
C23411 ctop a_23046_4138# 4.11f
C23412 col[28] rowoff_n[11] 0.0901f
C23413 a_2475_14202# a_13918_14178# 0.264f
C23414 a_7894_14178# a_7986_14178# 0.326f
C23415 a_2275_14202# a_11302_14218# 0.144f
C23416 VDD a_31990_9158# 0.181f
C23417 row_n[7] a_19030_9158# 0.282f
C23418 rowon_n[11] a_18938_13174# 0.118f
C23419 VDD a_19334_18234# 0.019f
C23420 a_2275_2154# a_26058_2130# 0.399f
C23421 col[8] a_2475_7174# 0.136f
C23422 m2_34864_3958# a_35002_4138# 0.225f
C23423 m2_30272_1374# VDD 0.0194f
C23424 row_n[9] a_6282_11206# 0.0117f
C23425 rowoff_n[9] a_31478_11528# 0.0133f
C23426 rowon_n[1] a_28978_3134# 0.118f
C23427 a_8990_7150# a_8990_6146# 0.843f
C23428 m2_22240_11414# a_22042_11166# 0.165f
C23429 col_n[7] a_9994_5142# 0.251f
C23430 vcm a_25358_13214# 0.155f
C23431 a_2966_11166# a_3970_11166# 0.843f
C23432 a_2275_11190# a_4882_11166# 0.136f
C23433 VDD a_23446_3496# 0.0779f
C23434 col_n[17] a_20034_17190# 0.251f
C23435 m2_13780_18014# a_13918_18194# 0.225f
C23436 col_n[14] a_16930_7150# 0.0765f
C23437 ctop a_3970_7150# 4.11f
C23438 col_n[15] a_2275_13198# 0.113f
C23439 m3_1864_5094# a_2966_5142# 0.0302f
C23440 a_2275_16210# a_26362_16226# 0.144f
C23441 a_2475_16210# a_28978_16186# 0.264f
C23442 VDD a_12914_12170# 0.181f
C23443 col_n[20] a_2275_2154# 0.113f
C23444 a_21038_4138# a_21342_4178# 0.0931f
C23445 a_21950_4138# a_22442_4500# 0.0658f
C23446 row_n[1] a_6890_3134# 0.0437f
C23447 vcm a_18938_7150# 0.1f
C23448 rowon_n[5] a_5978_7150# 0.248f
C23449 a_33086_9158# a_34090_9158# 0.843f
C23450 rowoff_n[12] a_13006_14178# 0.294f
C23451 col[12] rowoff_n[12] 0.0901f
C23452 col[5] a_2275_10186# 0.0899f
C23453 vcm a_6282_16226# 0.155f
C23454 a_2275_13198# a_19942_13174# 0.136f
C23455 col_n[8] a_11398_15544# 0.0283f
C23456 VDD a_4370_6508# 0.0779f
C23457 col_n[31] a_34394_6186# 0.084f
C23458 col[27] a_30074_4138# 0.367f
C23459 ctop a_19030_11166# 4.11f
C23460 a_22954_18194# a_23046_18194# 0.0991f
C23461 VDD a_27974_16186# 0.181f
C23462 a_17934_1126# a_18026_1126# 0.361f
C23463 m2_9188_15430# rowon_n[13] 0.0322f
C23464 col[25] a_2475_9182# 0.136f
C23465 m2_15212_11414# rowon_n[9] 0.0322f
C23466 m2_21236_7398# rowon_n[5] 0.0322f
C23467 m2_34864_5966# vcm 0.408f
C23468 m2_27260_3382# rowon_n[1] 0.0322f
C23469 m2_13204_9406# a_13006_9158# 0.165f
C23470 vcm a_33998_11166# 0.1f
C23471 a_24050_11166# a_24050_10162# 0.843f
C23472 a_2475_10186# a_12002_10162# 0.316f
C23473 row_n[14] a_17022_16186# 0.282f
C23474 a_2275_15206# a_35002_15182# 0.136f
C23475 a_17934_15182# a_18330_15222# 0.0313f
C23476 col_n[22] a_25358_4178# 0.084f
C23477 VDD a_19430_10524# 0.0779f
C23478 col_n[6] a_8990_15182# 0.251f
C23479 ctop a_34090_15182# 4.06f
C23480 col_n[3] a_5886_5142# 0.0765f
C23481 row_n[4] a_27062_6146# 0.282f
C23482 rowon_n[8] a_26970_10162# 0.118f
C23483 col_n[13] a_15926_17190# 0.0765f
C23484 m2_32280_5390# a_32082_5142# 0.165f
C23485 a_2475_7174# a_3878_7150# 0.264f
C23486 a_2275_7174# a_2874_7150# 0.136f
C23487 rowoff_n[10] a_19430_12532# 0.0133f
C23488 rowoff_n[2] a_1957_4162# 0.0219f
C23489 m2_8760_18014# vcm 0.353f
C23490 m2_35292_16434# rowon_n[14] 0.0322f
C23491 row_n[6] a_14314_8194# 0.0117f
C23492 vcm a_14922_14178# 0.1f
C23493 a_14010_12170# a_15014_12170# 0.843f
C23494 a_2475_12194# a_27062_12170# 0.316f
C23495 VDD a_10998_4138# 0.483f
C23496 col[22] a_2275_12194# 0.0899f
C23497 col[27] a_2275_1150# 0.0899f
C23498 VDD a_34490_14540# 0.0779f
C23499 row_n[8] a_4882_10162# 0.0437f
C23500 col[16] a_19030_2130# 0.367f
C23501 rowoff_n[0] a_11398_2492# 0.0133f
C23502 rowon_n[12] a_3970_14178# 0.248f
C23503 a_32994_5142# a_33086_5142# 0.326f
C23504 col[26] a_29070_14178# 0.367f
C23505 col[23] a_25966_4138# 0.0682f
C23506 m2_4168_7398# a_3970_7150# 0.165f
C23507 a_2275_9182# a_18026_9158# 0.399f
C23508 rowoff_n[14] a_35494_16548# 0.0133f
C23509 rowon_n[2] a_14010_4138# 0.248f
C23510 vcm a_29982_18194# 0.101f
C23511 a_4974_14178# a_4974_13174# 0.843f
C23512 VDD a_26058_8154# 0.483f
C23513 rowoff_n[5] a_2874_7150# 0.202f
C23514 m2_8760_946# col[6] 0.425f
C23515 row_n[0] a_2966_2130# 0.0122f
C23516 col_n[11] a_14314_2170# 0.084f
C23517 VDD a_15414_17552# 0.0779f
C23518 col_n[12] a_2475_8178# 0.0531f
C23519 a_27974_2130# a_28370_2170# 0.0313f
C23520 rowon_n[4] a_2275_6170# 1.79f
C23521 col_n[21] a_24354_14218# 0.084f
C23522 m2_23244_3382# a_23046_3134# 0.165f
C23523 vcm a_32082_3134# 0.56f
C23524 a_2275_6170# a_8290_6186# 0.144f
C23525 a_2475_6170# a_10906_6146# 0.264f
C23526 col_n[2] a_4882_15182# 0.0765f
C23527 rowoff_n[3] a_12002_5142# 0.294f
C23528 a_2275_11190# a_33086_11166# 0.399f
C23529 a_17022_11166# a_17326_11206# 0.0931f
C23530 a_17934_11166# a_18426_11528# 0.0658f
C23531 m2_9764_18014# a_9994_17190# 0.843f
C23532 m2_32856_18014# a_32994_18194# 0.225f
C23533 m2_1732_7974# VDD 0.856f
C23534 a_29070_16186# a_30074_16186# 0.843f
C23535 row_n[11] a_25054_13174# 0.282f
C23536 col[2] a_2475_5166# 0.136f
C23537 VDD a_6982_11166# 0.483f
C23538 m2_34864_18014# m3_33992_18146# 0.0341f
C23539 rowon_n[15] a_24962_17190# 0.118f
C23540 a_2475_3158# a_1957_3158# 0.0734f
C23541 row_n[1] a_35094_3134# 0.0123f
C23542 rowoff_n[1] a_21038_3134# 0.294f
C23543 rowoff_n[8] a_3878_10162# 0.202f
C23544 row_n[13] a_12306_15222# 0.0117f
C23545 rowon_n[5] a_35002_7150# 0.118f
C23546 vcm a_13006_6146# 0.56f
C23547 a_2475_8178# a_25966_8154# 0.264f
C23548 a_2275_8178# a_23350_8194# 0.144f
C23549 a_13918_8154# a_14010_8154# 0.326f
C23550 rowoff_n[11] a_7382_13536# 0.0133f
C23551 col_n[9] a_2275_11190# 0.113f
C23552 col[15] a_18026_12170# 0.367f
C23553 col[12] a_14922_2130# 0.0682f
C23554 vcm a_1957_15206# 0.139f
C23555 col[22] a_24962_14178# 0.0682f
C23556 row_n[3] a_22346_5182# 0.0117f
C23557 row_n[15] a_2161_17214# 0.0221f
C23558 m2_8184_14426# row_n[12] 0.0128f
C23559 a_2275_17214# a_2966_17190# 0.399f
C23560 a_2475_17214# a_3970_17190# 0.316f
C23561 VDD a_22042_15182# 0.483f
C23562 m2_14208_10410# row_n[8] 0.0128f
C23563 col_n[30] a_33086_8154# 0.251f
C23564 a_2275_2154# m2_34864_1950# 0.278f
C23565 m2_20232_6394# row_n[4] 0.0128f
C23566 row_n[8] col[22] 0.0342f
C23567 row_n[5] col[16] 0.0342f
C23568 row_n[11] col[28] 0.0342f
C23569 rowon_n[7] col[21] 0.0323f
C23570 rowon_n[3] col[13] 0.0323f
C23571 rowon_n[9] col[25] 0.0323f
C23572 rowon_n[4] col[15] 0.0323f
C23573 rowon_n[6] col[19] 0.0323f
C23574 rowon_n[10] col[27] 0.0323f
C23575 row_n[12] col[30] 0.0342f
C23576 row_n[10] col[26] 0.0342f
C23577 row_n[6] col[18] 0.0342f
C23578 row_n[7] col[20] 0.0342f
C23579 row_n[4] col[14] 0.0342f
C23580 ctop col[3] 0.123f
C23581 row_n[1] col[8] 0.0342f
C23582 rowon_n[11] col[29] 0.0323f
C23583 rowon_n[0] col[7] 0.0323f
C23584 rowon_n[8] col[23] 0.0323f
C23585 row_n[2] col[10] 0.0342f
C23586 rowon_n[1] col[9] 0.0323f
C23587 row_n[9] col[24] 0.0342f
C23588 row_n[0] col[6] 0.0342f
C23589 row_n[13] sample_n 0.0596f
C23590 rowon_n[12] col[31] 0.0323f
C23591 row_n[3] col[12] 0.0342f
C23592 rowon_n[2] col[11] 0.0323f
C23593 rowon_n[5] col[17] 0.0323f
C23594 col_n[29] a_2475_10186# 0.0531f
C23595 a_2275_5166# a_16930_5142# 0.136f
C23596 row_n[5] a_12914_7150# 0.0437f
C23597 a_8898_5142# a_9294_5182# 0.0313f
C23598 m3_34996_8106# m3_34996_7102# 0.202f
C23599 col_n[10] a_13310_12210# 0.084f
C23600 rowon_n[9] a_12002_11166# 0.248f
C23601 vcm a_28066_10162# 0.56f
C23602 rowoff_n[15] a_23446_17552# 0.0133f
C23603 a_32994_15182# a_33486_15544# 0.0658f
C23604 a_32082_15182# a_32386_15222# 0.0931f
C23605 col[19] a_2475_7174# 0.136f
C23606 col_n[21] a_24450_6508# 0.0283f
C23607 VDD a_2874_18194# 0.343f
C23608 col_n[31] a_34490_18556# 0.0283f
C23609 a_4974_2130# a_5978_2130# 0.843f
C23610 a_2475_2154# a_8990_2130# 0.316f
C23611 m2_34864_15002# row_n[13] 0.267f
C23612 vcm a_18330_4178# 0.155f
C23613 rowoff_n[9] a_13918_11166# 0.202f
C23614 a_2275_7174# a_31990_7150# 0.136f
C23615 col_n[26] a_2275_13198# 0.113f
C23616 vcm a_8990_13174# 0.56f
C23617 a_28978_12170# a_29070_12170# 0.326f
C23618 VDD a_5886_3134# 0.181f
C23619 col_n[31] a_2275_2154# 0.113f
C23620 col[4] a_6982_10162# 0.367f
C23621 m2_17796_18014# col_n[15] 0.243f
C23622 a_2275_16210# a_9994_16186# 0.399f
C23623 col[11] a_13918_12170# 0.0682f
C23624 row_n[8] a_33086_10162# 0.282f
C23625 rowoff_n[7] a_22954_9158# 0.202f
C23626 rowon_n[12] a_32994_14178# 0.118f
C23627 col_n[19] a_22042_6146# 0.251f
C23628 a_2475_4162# a_24050_4138# 0.316f
C23629 a_30074_5142# a_30074_4138# 0.843f
C23630 m3_14916_1078# ctop 0.21f
C23631 col[23] rowoff_n[12] 0.0901f
C23632 col[16] a_2275_10186# 0.0899f
C23633 col_n[26] a_28978_8154# 0.0765f
C23634 vcm a_33390_8194# 0.155f
C23635 a_23958_9158# a_24354_9198# 0.0313f
C23636 rowoff_n[13] a_29982_15182# 0.202f
C23637 row_n[10] a_20338_12210# 0.0117f
C23638 ctop a_12002_2130# 4.06f
C23639 vcm a_24050_17190# 0.56f
C23640 VDD a_20946_7150# 0.181f
C23641 rowoff_n[5] a_31990_7150# 0.202f
C23642 a_13918_18194# a_14410_18556# 0.0658f
C23643 a_2275_18218# a_25054_18194# 0.0924f
C23644 row_n[0] a_30378_2170# 0.0117f
C23645 a_2275_1150# a_15014_1126# 0.0924f
C23646 a_8898_1126# a_9390_1488# 0.0658f
C23647 row_n[12] a_10906_14178# 0.0437f
C23648 col_n[10] a_13406_4500# 0.0283f
C23649 vcm a_26970_2130# 0.1f
C23650 col_n[20] a_23446_16548# 0.0283f
C23651 a_20034_6146# a_21038_6146# 0.843f
C23652 m2_14784_946# m2_15212_1374# 0.165f
C23653 row_n[2] a_20946_4138# 0.0437f
C23654 vcm a_14314_11206# 0.155f
C23655 col_n[1] a_2475_17214# 0.0531f
C23656 VDD a_12402_1488# 0.0977f
C23657 m2_28840_18014# a_29070_17190# 0.843f
C23658 rowon_n[6] a_20034_8154# 0.248f
C23659 col_n[6] a_2475_6170# 0.0531f
C23660 ctop a_27062_6146# 4.11f
C23661 a_9902_15182# a_9994_15182# 0.326f
C23662 a_2475_15206# a_17934_15182# 0.264f
C23663 a_2275_15206# a_15318_15222# 0.144f
C23664 rowon_n[0] m2_32280_2378# 0.0322f
C23665 a_2475_18218# a_23046_18194# 0.0299f
C23666 a_2275_3158# a_30074_3134# 0.399f
C23667 col[7] rowoff_n[13] 0.0901f
C23668 rowoff_n[8] a_32482_10524# 0.0133f
C23669 vcm a_7894_5142# 0.1f
C23670 col_n[8] a_10998_4138# 0.251f
C23671 a_10998_8154# a_10998_7150# 0.843f
C23672 col_n[18] a_21038_16186# 0.251f
C23673 vcm a_29374_15222# 0.155f
C23674 col_n[15] a_17934_6146# 0.0765f
C23675 a_4882_12170# a_5278_12210# 0.0313f
C23676 a_2275_12194# a_8898_12170# 0.136f
C23677 VDD a_27462_5504# 0.0779f
C23678 col_n[25] a_27974_18194# 0.0762f
C23679 m2_12776_18014# VDD 0.993f
C23680 row_n[15] a_31078_17190# 0.282f
C23681 ctop a_7986_9158# 4.11f
C23682 a_2475_17214# a_32994_17190# 0.264f
C23683 a_2275_17214# a_30378_17230# 0.144f
C23684 VDD a_16930_14178# 0.181f
C23685 a_32082_2130# m2_32280_2378# 0.165f
C23686 rowon_n[0] a_7894_2130# 0.118f
C23687 col_n[3] a_2275_9182# 0.113f
C23688 a_23046_5142# a_23350_5182# 0.0931f
C23689 a_23958_5142# a_24450_5504# 0.0658f
C23690 vcm a_22954_9158# 0.1f
C23691 m2_5748_18014# m2_6176_18442# 0.165f
C23692 rowoff_n[14] a_17934_16186# 0.202f
C23693 col_n[9] a_12402_14540# 0.0283f
C23694 vcm a_10298_18234# 0.16f
C23695 m3_24956_1078# a_25054_2130# 0.0302f
C23696 a_2275_14202# a_23958_14178# 0.136f
C23697 col[28] a_31078_3134# 0.367f
C23698 m2_20808_946# a_21038_1126# 0.0249f
C23699 col_n[23] a_2475_8178# 0.0531f
C23700 VDD a_8386_8516# 0.0779f
C23701 row_n[7] a_28370_9198# 0.0117f
C23702 m2_4168_9406# rowon_n[7] 0.0322f
C23703 m2_10192_5390# rowon_n[3] 0.0322f
C23704 ctop a_23046_13174# 4.11f
C23705 m2_10768_946# vcm 0.353f
C23706 VDD a_31990_18194# 0.343f
C23707 a_2275_2154# a_2275_1150# 0.0693f
C23708 a_19942_2130# a_20034_2130# 0.326f
C23709 m3_33992_18146# VDD 0.0317f
C23710 row_n[9] a_18938_11166# 0.0437f
C23711 col[8] a_2475_16210# 0.136f
C23712 rowon_n[13] a_18026_15182# 0.248f
C23713 col[13] a_2475_5166# 0.136f
C23714 a_26058_12170# a_26058_11166# 0.843f
C23715 a_2475_11190# a_16018_11166# 0.316f
C23716 col_n[23] a_26362_3174# 0.084f
C23717 VDD a_34090_3134# 0.483f
C23718 col_n[7] a_9994_14178# 0.251f
C23719 a_19942_16186# a_20338_16226# 0.0313f
C23720 rowon_n[3] a_28066_5142# 0.248f
C23721 col_n[4] a_6890_4138# 0.0765f
C23722 VDD a_23446_12532# 0.0779f
C23723 m2_10768_18014# m3_10900_18146# 3.79f
C23724 ctop a_3970_16186# 4.11f
C23725 col_n[14] a_16930_16186# 0.0765f
C23726 m2_25252_14426# rowon_n[12] 0.0322f
C23727 m2_31276_10410# rowon_n[8] 0.0322f
C23728 col_n[20] a_2275_11190# 0.113f
C23729 rowoff_n[1] a_2966_3134# 0.294f
C23730 m2_1732_15002# m2_1732_13998# 0.843f
C23731 a_3970_8154# a_4274_8194# 0.0931f
C23732 a_2275_8178# a_6982_8154# 0.399f
C23733 a_4882_8154# a_5374_8516# 0.0658f
C23734 vcm a_18938_16186# 0.1f
C23735 a_2475_13198# a_31078_13174# 0.316f
C23736 a_16018_13174# a_17022_13174# 0.843f
C23737 VDD a_15014_6146# 0.483f
C23738 row_n[3] a_5978_5142# 0.282f
C23739 rowon_n[0] col[18] 0.0323f
C23740 rowon_n[5] col[28] 0.0323f
C23741 row_n[6] col[29] 0.0342f
C23742 row_n[2] col[21] 0.0342f
C23743 row_n[0] col[17] 0.0342f
C23744 row_n[1] col[19] 0.0342f
C23745 rowon_n[3] col[24] 0.0323f
C23746 rowon_n[1] col[20] 0.0323f
C23747 row_n[5] col[27] 0.0342f
C23748 ctop col[14] 0.123f
C23749 row_n[7] col[31] 0.0342f
C23750 rowon_n[2] col[22] 0.0323f
C23751 row_n[3] col[23] 0.0342f
C23752 row_n[4] col[25] 0.0342f
C23753 rowon_n[4] col[26] 0.0323f
C23754 rowon_n[6] col[30] 0.0323f
C23755 rowon_n[7] sample_n 0.0692f
C23756 rowon_n[7] a_5886_9158# 0.118f
C23757 VDD a_4370_15544# 0.0779f
C23758 col[17] a_20034_1126# 0.428f
C23759 col[10] a_2275_8178# 0.0899f
C23760 col_n[31] a_34394_15222# 0.084f
C23761 m2_1732_8978# rowoff_n[7] 0.415f
C23762 col[27] a_30074_13174# 0.367f
C23763 col[24] a_26970_3134# 0.0682f
C23764 vcm a_21038_1126# 0.165f
C23765 a_34090_6146# a_34394_6186# 0.0931f
C23766 a_35002_6146# a_35094_6146# 0.0991f
C23767 m2_13780_946# m3_12908_1078# 0.0341f
C23768 m3_19936_18146# m3_20940_18146# 0.202f
C23769 rowoff_n[15] a_5886_17190# 0.202f
C23770 a_2275_10186# a_22042_10162# 0.399f
C23771 row_n[14] a_26362_16226# 0.0117f
C23772 col[30] a_2475_7174# 0.136f
C23773 m2_9188_16434# a_8990_16186# 0.165f
C23774 rowoff_n[4] a_3970_6146# 0.294f
C23775 a_6982_15182# a_6982_14178# 0.843f
C23776 VDD a_30074_10162# 0.483f
C23777 col_n[12] a_15318_1166# 0.0839f
C23778 col_n[22] a_25358_13214# 0.084f
C23779 a_29982_3134# a_30378_3174# 0.0313f
C23780 col_n[3] a_5886_14178# 0.0765f
C23781 vcm a_2475_4162# 1.08f
C23782 a_2475_7174# a_14922_7150# 0.264f
C23783 a_2275_7174# a_12306_7190# 0.144f
C23784 rowoff_n[2] a_13006_4138# 0.294f
C23785 rowoff_n[10] a_30074_12170# 0.294f
C23786 m2_28264_12418# a_28066_12170# 0.165f
C23787 row_n[6] a_26970_8154# 0.0437f
C23788 a_19030_12170# a_19334_12210# 0.0931f
C23789 a_19942_12170# a_20434_12532# 0.0658f
C23790 rowon_n[10] a_26058_12170# 0.248f
C23791 a_31078_17190# a_32082_17190# 0.843f
C23792 VDD a_10998_13174# 0.483f
C23793 col[27] a_2275_10186# 0.0899f
C23794 rowoff_n[0] a_22042_2130# 0.294f
C23795 m2_1732_15002# col[0] 0.0137f
C23796 vcm m2_1732_946# 0.321f
C23797 a_2275_4162# a_5886_4138# 0.136f
C23798 m3_10900_18146# ctop 0.209f
C23799 col[16] a_19030_11166# 0.367f
C23800 col[13] a_15926_1126# 0.0682f
C23801 vcm a_17022_8154# 0.56f
C23802 a_2275_9182# a_27366_9198# 0.144f
C23803 a_2475_9182# a_29982_9158# 0.264f
C23804 m2_3164_8402# row_n[6] 0.0128f
C23805 a_15926_9158# a_16018_9158# 0.326f
C23806 m2_9188_4386# row_n[2] 0.0128f
C23807 row_n[10] a_3970_12170# 0.282f
C23808 col[23] a_25966_13174# 0.0682f
C23809 VDD a_2275_7174# 1.96f
C23810 col_n[31] a_34090_7150# 0.251f
C23811 VDD a_26058_17190# 0.484f
C23812 row_n[0] a_14010_2130# 0.282f
C23813 rowon_n[4] a_13918_6146# 0.118f
C23814 col_n[11] a_14314_11206# 0.084f
C23815 col_n[12] a_2475_17214# 0.0531f
C23816 vcm a_7286_2170# 0.155f
C23817 a_2275_6170# a_20946_6146# 0.136f
C23818 a_10906_6146# a_11302_6186# 0.0313f
C23819 m2_1732_8978# vcm 0.316f
C23820 col_n[17] a_2475_6170# 0.0531f
C23821 m2_19228_10410# a_19030_10162# 0.165f
C23822 row_n[2] a_2275_4162# 19.2f
C23823 vcm a_32082_12170# 0.56f
C23824 m2_18224_17438# row_n[15] 0.0128f
C23825 VDD a_28978_2130# 0.181f
C23826 rowon_n[6] a_1957_8178# 0.0172f
C23827 m2_24248_13422# row_n[11] 0.0128f
C23828 m2_30272_9406# row_n[7] 0.0128f
C23829 m2_35292_5390# row_n[3] 0.0128f
C23830 a_35002_16186# a_35494_16548# 0.0658f
C23831 col_n[22] a_25454_5504# 0.0283f
C23832 row_n[11] a_35398_13214# 0.0117f
C23833 col[18] rowoff_n[13] 0.0901f
C23834 col[2] a_2475_14202# 0.136f
C23835 a_2475_3158# a_13006_3134# 0.316f
C23836 sample rowoff_n[6] 0.0775f
C23837 col_n[1] rowoff_n[9] 0.0471f
C23838 VDD rowoff_n[5] 1.51f
C23839 a_6982_3134# a_7986_3134# 0.843f
C23840 col_n[0] rowoff_n[7] 0.0471f
C23841 vcm rowoff_n[8] 0.533f
C23842 col[7] a_2475_3158# 0.136f
C23843 rowoff_n[8] a_14922_10162# 0.202f
C23844 a_26970_1126# a_2475_1150# 0.264f
C23845 a_24354_1166# a_2275_1150# 0.145f
C23846 row_n[13] a_24962_15182# 0.0437f
C23847 vcm a_22346_6186# 0.155f
C23848 a_2275_8178# a_34394_8194# 0.144f
C23849 rowoff_n[11] a_18026_13174# 0.294f
C23850 col[5] a_7986_9158# 0.367f
C23851 vcm a_13006_15182# 0.56f
C23852 a_30986_13174# a_31078_13174# 0.326f
C23853 VDD a_9902_5142# 0.181f
C23854 row_n[3] a_35002_5142# 0.0437f
C23855 col[12] a_14922_11166# 0.0682f
C23856 col_n[14] a_2275_9182# 0.113f
C23857 rowon_n[7] a_34090_9158# 0.248f
C23858 a_2275_17214# a_14010_17190# 0.399f
C23859 rowoff_n[6] a_23958_8154# 0.202f
C23860 col_n[20] a_23046_5142# 0.251f
C23861 col_n[30] a_33086_17190# 0.251f
C23862 m2_34864_2954# m2_35292_3382# 0.165f
C23863 col_n[27] a_29982_7150# 0.0765f
C23864 a_2475_5166# a_28066_5142# 0.316f
C23865 a_32082_6146# a_32082_5142# 0.843f
C23866 m3_9896_1078# m3_10900_1078# 0.202f
C23867 m2_10192_8402# a_9994_8154# 0.165f
C23868 vcm a_3270_9198# 0.155f
C23869 rowoff_n[15] a_34090_17190# 0.294f
C23870 a_25966_10162# a_26362_10202# 0.0313f
C23871 col[4] a_2275_6170# 0.0899f
C23872 rowoff_n[4] a_32994_6146# 0.202f
C23873 ctop a_16018_4138# 4.11f
C23874 col[2] rowoff_n[14] 0.0901f
C23875 m2_21812_946# a_2275_1150# 0.28f
C23876 m2_8760_946# a_8898_1126# 0.225f
C23877 a_2475_14202# a_6890_14178# 0.264f
C23878 a_2275_14202# a_4274_14218# 0.144f
C23879 row_n[7] a_12002_9158# 0.282f
C23880 VDD a_24962_9158# 0.181f
C23881 rowon_n[11] a_11910_13174# 0.118f
C23882 VDD a_12306_18234# 0.019f
C23883 col_n[11] a_14410_3496# 0.0283f
C23884 a_9994_2130# a_10298_2170# 0.0931f
C23885 a_2275_2154# a_19030_2130# 0.399f
C23886 a_10906_2130# a_11398_2492# 0.0658f
C23887 col[19] a_2475_16210# 0.136f
C23888 col_n[21] a_24450_15544# 0.0283f
C23889 m2_29268_4386# a_29070_4138# 0.165f
C23890 m2_14784_946# VDD 1f
C23891 col[24] a_2475_5166# 0.136f
C23892 vcm a_30986_4138# 0.1f
C23893 rowon_n[1] a_21950_3134# 0.118f
C23894 rowoff_n[9] a_24450_11528# 0.0133f
C23895 a_22042_7150# a_23046_7150# 0.843f
C23896 vcm a_18330_13214# 0.155f
C23897 VDD a_16418_3496# 0.0779f
C23898 sample a_2161_9182# 0.0858f
C23899 m2_8760_18014# a_8990_18194# 0.0249f
C23900 ctop a_31078_8154# 4.11f
C23901 a_11910_16186# a_12002_16186# 0.326f
C23902 a_2275_16210# a_19334_16226# 0.144f
C23903 a_2475_16210# a_21950_16186# 0.264f
C23904 VDD a_5886_12170# 0.181f
C23905 col_n[31] a_2275_11190# 0.113f
C23906 a_27366_1166# m2_26832_946# 0.087f
C23907 rowoff_n[7] a_33486_9520# 0.0133f
C23908 a_2275_4162# a_34090_4138# 0.399f
C23909 col_n[9] a_12002_3134# 0.251f
C23910 vcm a_11910_7150# 0.1f
C23911 col_n[19] a_22042_15182# 0.251f
C23912 a_13006_9158# a_13006_8154# 0.843f
C23913 rowoff_n[12] a_5978_14178# 0.294f
C23914 col_n[16] a_18938_5142# 0.0765f
C23915 row_n[10] a_32994_12170# 0.0437f
C23916 VDD col_n[2] 5.17f
C23917 col_n[0] vcm 1.94f
C23918 row_n[2] sample_n 0.0596f
C23919 rowon_n[0] col[29] 0.0323f
C23920 col[9] col[10] 0.0355f
C23921 rowon_n[1] col[31] 0.0323f
C23922 row_n[0] col[28] 0.0342f
C23923 row_n[1] col[30] 0.0342f
C23924 ctop col[25] 0.123f
C23925 vcm a_33390_17230# 0.155f
C23926 col_n[26] a_28978_17190# 0.0765f
C23927 m2_32856_18014# col[30] 0.347f
C23928 col[21] a_2275_8178# 0.0899f
C23929 a_2275_13198# a_12914_13174# 0.136f
C23930 rowon_n[14] a_32082_16186# 0.248f
C23931 a_6890_13174# a_7286_13214# 0.0313f
C23932 VDD a_31478_7512# 0.0779f
C23933 ctop a_12002_11166# 4.11f
C23934 a_2275_18218# a_35398_18234# 0.145f
C23935 VDD a_20946_16186# 0.181f
C23936 vcm a_2966_1126# 0.165f
C23937 a_25966_6146# a_26458_6508# 0.0658f
C23938 a_25054_6146# a_25358_6186# 0.0931f
C23939 m2_26832_946# m2_27836_946# 0.843f
C23940 col_n[10] a_13406_13536# 0.0283f
C23941 vcm a_26970_11166# 0.1f
C23942 a_2475_10186# a_4974_10162# 0.316f
C23943 VDD a_23046_1126# 0.035f
C23944 col[29] a_32082_2130# 0.367f
C23945 row_n[14] a_9994_16186# 0.282f
C23946 a_2275_15206# a_27974_15182# 0.136f
C23947 VDD a_12402_10524# 0.0779f
C23948 col_n[6] a_2475_15206# 0.0531f
C23949 ctop a_27062_15182# 4.11f
C23950 row_n[4] a_20034_6146# 0.282f
C23951 col_n[11] a_2475_4162# 0.0531f
C23952 a_21950_3134# a_22042_3134# 0.326f
C23953 rowon_n[8] a_19942_10162# 0.118f
C23954 rowoff_n[10] a_12402_12532# 0.0133f
C23955 a_30378_1166# vcm 0.16f
C23956 col_n[24] a_27366_2170# 0.084f
C23957 m2_8184_16434# rowon_n[14] 0.0322f
C23958 row_n[6] a_7286_8194# 0.0117f
C23959 m2_14208_12418# rowon_n[10] 0.0322f
C23960 m2_20232_8402# rowon_n[6] 0.0322f
C23961 vcm a_7894_14178# 0.1f
C23962 m2_26256_4386# rowon_n[2] 0.0322f
C23963 col_n[8] a_10998_13174# 0.251f
C23964 a_2475_12194# a_20034_12170# 0.316f
C23965 a_28066_13174# a_28066_12170# 0.843f
C23966 VDD a_3970_4138# 0.483f
C23967 col_n[5] a_7894_3134# 0.0765f
C23968 m2_34288_18442# VDD 0.0456f
C23969 col[1] a_2475_1150# 0.136f
C23970 col_n[15] a_17934_15182# 0.0765f
C23971 a_21950_17190# a_22346_17230# 0.0313f
C23972 VDD a_27462_14540# 0.0779f
C23973 rowoff_n[0] a_4370_2492# 0.0133f
C23974 en_bit_n[0] a_20338_1166# 0.0266f
C23975 col_n[3] a_2275_18218# 0.113f
C23976 a_6890_9158# a_7382_9520# 0.0658f
C23977 col_n[8] a_2275_7174# 0.113f
C23978 rowoff_n[14] a_28466_16548# 0.0133f
C23979 a_2275_9182# a_10998_9158# 0.399f
C23980 a_5978_9158# a_6282_9198# 0.0931f
C23981 rowon_n[2] a_6982_4138# 0.248f
C23982 vcm a_22954_18194# 0.101f
C23983 a_18026_14178# a_19030_14178# 0.843f
C23984 a_2475_14202# a_35094_14178# 0.0299f
C23985 m2_34864_17010# rowon_n[15] 0.231f
C23986 VDD a_19030_8154# 0.483f
C23987 m2_33860_946# vcm 0.158f
C23988 col[28] a_31078_12170# 0.367f
C23989 VDD a_8386_17552# 0.0779f
C23990 col_n[23] a_2475_17214# 0.0531f
C23991 col[25] a_27974_2130# 0.0682f
C23992 col_n[28] a_2475_6170# 0.0531f
C23993 m3_9896_1078# VDD 0.0157f
C23994 vcm a_25054_3134# 0.56f
C23995 rowoff_n[3] a_4974_5142# 0.294f
C23996 a_2275_11190# a_26058_11166# 0.399f
C23997 col[29] rowoff_n[13] 0.0901f
C23998 m2_27836_18014# a_28066_18194# 0.0249f
C23999 col[13] a_2475_14202# 0.136f
C24000 row_n[11] a_18026_13174# 0.282f
C24001 a_8990_16186# a_8990_15182# 0.843f
C24002 col_n[23] a_26362_12210# 0.084f
C24003 VDD a_34090_12170# 0.483f
C24004 col_n[3] rowoff_n[0] 0.0471f
C24005 col_n[7] rowoff_n[4] 0.0471f
C24006 col[18] a_2475_3158# 0.136f
C24007 col_n[4] rowoff_n[1] 0.0471f
C24008 col_n[5] rowoff_n[2] 0.0471f
C24009 col_n[6] rowoff_n[3] 0.0471f
C24010 col_n[9] rowoff_n[6] 0.0471f
C24011 col_n[8] rowoff_n[5] 0.0471f
C24012 col_n[11] rowoff_n[8] 0.0471f
C24013 m2_24824_18014# m3_25960_18146# 0.0341f
C24014 col_n[10] rowoff_n[7] 0.0471f
C24015 col_n[12] rowoff_n[9] 0.0471f
C24016 rowon_n[15] a_17934_17190# 0.118f
C24017 col_n[4] a_6890_13174# 0.0765f
C24018 a_31990_4138# a_32386_4178# 0.0313f
C24019 row_n[1] a_28066_3134# 0.282f
C24020 rowoff_n[1] a_14010_3134# 0.294f
C24021 row_n[13] a_5278_15222# 0.0117f
C24022 rowon_n[5] a_27974_7150# 0.118f
C24023 vcm a_5978_6146# 0.56f
C24024 a_2475_8178# a_18938_8154# 0.264f
C24025 a_2275_8178# a_16322_8194# 0.144f
C24026 rowoff_n[12] a_35002_14178# 0.202f
C24027 col_n[25] a_2275_9182# 0.113f
C24028 a_21038_13174# a_21342_13214# 0.0931f
C24029 a_21950_13174# a_22442_13536# 0.0658f
C24030 row_n[3] a_15318_5182# 0.0117f
C24031 VDD a_15014_15182# 0.483f
C24032 m3_7888_18146# a_7986_17190# 0.0303f
C24033 col[17] a_20034_10162# 0.367f
C24034 col[10] a_2275_17214# 0.0899f
C24035 row_n[5] a_5886_7150# 0.0437f
C24036 a_2275_5166# a_9902_5142# 0.136f
C24037 col[15] a_2275_6170# 0.0899f
C24038 m2_28840_946# m3_28972_1078# 3.79f
C24039 m3_34996_15134# m3_34996_14130# 0.202f
C24040 col[24] a_26970_12170# 0.0682f
C24041 rowon_n[9] a_4974_11166# 0.248f
C24042 col[13] rowoff_n[14] 0.0901f
C24043 vcm a_21038_10162# 0.56f
C24044 rowoff_n[15] a_16418_17552# 0.0133f
C24045 a_2275_10186# a_31382_10202# 0.144f
C24046 a_2475_10186# a_33998_10162# 0.264f
C24047 a_17934_10162# a_18026_10162# 0.326f
C24048 m2_22816_18014# ctop 0.0422f
C24049 col[30] a_2475_16210# 0.136f
C24050 col_n[12] a_15318_10202# 0.084f
C24051 a_19030_3134# a_19030_2130# 0.843f
C24052 m2_7180_15430# row_n[13] 0.0128f
C24053 m2_13204_11414# row_n[9] 0.0128f
C24054 m2_19228_7398# row_n[5] 0.0128f
C24055 m2_25252_3382# row_n[1] 0.0128f
C24056 vcm a_11302_4178# 0.155f
C24057 a_12914_7150# a_13310_7190# 0.0313f
C24058 a_2275_7174# a_24962_7150# 0.136f
C24059 rowon_n[1] a_3878_3134# 0.118f
C24060 rowoff_n[9] a_6890_11166# 0.202f
C24061 m2_1732_18014# sample_n 0.0513f
C24062 m2_1732_10986# a_2161_11190# 0.0454f
C24063 vcm a_2475_13198# 1.08f
C24064 VDD a_32994_4138# 0.181f
C24065 col_n[23] a_26458_4500# 0.0283f
C24066 col_n[5] a_2475_2154# 0.0531f
C24067 a_2475_16210# a_3878_16186# 0.264f
C24068 a_2275_16210# a_2874_16186# 0.136f
C24069 row_n[8] a_26058_10162# 0.282f
C24070 rowoff_n[7] a_15926_9158# 0.202f
C24071 rowon_n[12] a_25966_14178# 0.118f
C24072 a_8990_4138# a_9994_4138# 0.843f
C24073 a_2475_4162# a_17022_4138# 0.316f
C24074 m3_1864_8106# ctop 0.21f
C24075 VDD col_n[13] 5.17f
C24076 vcm col_n[10] 1.94f
C24077 analog_in col[31] 0.176f
C24078 m2_34288_16434# row_n[14] 0.0128f
C24079 vcm a_26362_8194# 0.155f
C24080 col[6] a_8990_8154# 0.367f
C24081 rowoff_n[13] a_22954_15182# 0.202f
C24082 row_n[10] a_13310_12210# 0.0117f
C24083 m2_34864_13998# a_2475_14202# 0.282f
C24084 col[13] a_15926_10162# 0.0682f
C24085 vcm a_17022_17190# 0.56f
C24086 ctop a_4974_2130# 4.06f
C24087 a_32994_14178# a_33086_14178# 0.326f
C24088 VDD a_13918_7150# 0.181f
C24089 rowoff_n[5] a_24962_7150# 0.202f
C24090 col_n[21] a_24050_4138# 0.251f
C24091 a_2275_18218# a_18026_18194# 0.0924f
C24092 VDD a_2275_16210# 1.96f
C24093 row_n[0] a_23350_2170# 0.0117f
C24094 col_n[31] a_34090_16186# 0.251f
C24095 a_2275_1150# a_7986_1126# 0.0924f
C24096 col_n[28] a_30986_6146# 0.0765f
C24097 col_n[2] a_2275_5166# 0.113f
C24098 vcm a_19942_2130# 0.1f
C24099 a_2475_6170# a_32082_6146# 0.316f
C24100 a_34090_7150# a_34090_6146# 0.843f
C24101 col_n[1] a_4274_8194# 0.084f
C24102 m2_7756_946# m2_8184_1374# 0.165f
C24103 vcm a_7286_11206# 0.155f
C24104 row_n[2] a_13918_4138# 0.0437f
C24105 rowoff_n[3] a_33998_5142# 0.202f
C24106 a_28370_1166# col_n[25] 0.084f
C24107 a_27974_11166# a_28370_11206# 0.0313f
C24108 VDD a_5374_1488# 0.0977f
C24109 rowon_n[6] a_13006_8154# 0.248f
C24110 col_n[17] a_2475_15206# 0.0531f
C24111 m2_15212_17438# a_15014_17190# 0.165f
C24112 ctop a_20034_6146# 4.11f
C24113 a_2475_15206# a_10906_15182# 0.264f
C24114 a_2275_15206# a_8290_15222# 0.144f
C24115 col_n[22] a_2475_4162# 0.0531f
C24116 VDD a_28978_11166# 0.181f
C24117 col_n[12] a_15414_2492# 0.0283f
C24118 col_n[22] a_25454_14540# 0.0283f
C24119 row_n[4] a_1957_6170# 0.187f
C24120 a_2275_3158# a_23046_3134# 0.399f
C24121 a_12002_3134# a_12306_3174# 0.0931f
C24122 a_12914_3134# a_13406_3496# 0.0658f
C24123 a_2475_18218# a_16018_18194# 0.0299f
C24124 rowoff_n[8] a_25454_10524# 0.0133f
C24125 vcm a_35002_6146# 0.101f
C24126 a_24050_8154# a_25054_8154# 0.843f
C24127 col[7] a_2475_12194# 0.136f
C24128 m2_34288_13422# a_34090_13174# 0.165f
C24129 col_n[0] a_3366_8516# 0.0283f
C24130 col[12] a_2475_1150# 0.136f
C24131 vcm a_22346_15222# 0.155f
C24132 a_2475_12194# a_1957_12194# 0.0734f
C24133 VDD a_20434_5504# 0.0779f
C24134 a_32386_1166# VDD 0.0149f
C24135 row_n[15] a_24050_17190# 0.282f
C24136 col[2] a_4882_8154# 0.0682f
C24137 a_2275_17214# a_23350_17230# 0.144f
C24138 a_13918_17190# a_14010_17190# 0.326f
C24139 a_2475_17214# a_25966_17190# 0.264f
C24140 VDD a_9902_14178# 0.181f
C24141 rowoff_n[6] a_34490_8516# 0.0133f
C24142 col_n[14] a_2275_18218# 0.113f
C24143 col_n[10] a_13006_2130# 0.251f
C24144 a_28978_1126# col[26] 0.0682f
C24145 col_n[19] a_2275_7174# 0.113f
C24146 row_n[5] a_34090_7150# 0.282f
C24147 col_n[20] a_23046_14178# 0.251f
C24148 col_n[17] a_19942_4138# 0.0765f
C24149 rowon_n[9] a_33998_11166# 0.118f
C24150 a_35002_1126# a_35494_1488# 0.0658f
C24151 vcm a_15926_9158# 0.1f
C24152 a_15014_10162# a_15014_9158# 0.843f
C24153 rowoff_n[14] a_10906_16186# 0.202f
C24154 col_n[27] a_29982_16186# 0.0765f
C24155 m2_6176_15430# a_5978_15182# 0.165f
C24156 vcm a_3270_18234# 0.16f
C24157 a_8898_14178# a_9294_14218# 0.0313f
C24158 a_2275_14202# a_16930_14178# 0.136f
C24159 row_n[7] a_21342_9198# 0.0117f
C24160 VDD a_35494_9520# 0.106f
C24161 col[4] a_2275_15206# 0.0899f
C24162 ctop a_16018_13174# 4.11f
C24163 col[9] a_2275_4162# 0.0899f
C24164 VDD a_24962_18194# 0.343f
C24165 a_2475_2154# a_30986_2130# 0.264f
C24166 a_2275_2154# a_28370_2170# 0.144f
C24167 m2_3164_3382# a_2966_3134# 0.165f
C24168 col_n[11] a_14410_12532# 0.0283f
C24169 m3_5880_18146# VDD 0.0308f
C24170 row_n[9] a_11910_11166# 0.0437f
C24171 rowoff_n[9] a_35094_11166# 0.0135f
C24172 a_27062_7150# a_27366_7190# 0.0931f
C24173 a_27974_7150# a_28466_7512# 0.0658f
C24174 m2_25252_11414# a_25054_11166# 0.165f
C24175 rowon_n[13] a_10998_15182# 0.248f
C24176 col[24] a_2475_14202# 0.136f
C24177 vcm a_30986_13174# 0.1f
C24178 a_4974_11166# a_5978_11166# 0.843f
C24179 a_2475_11190# a_8990_11166# 0.316f
C24180 col_n[16] rowoff_n[2] 0.0471f
C24181 col_n[19] rowoff_n[5] 0.0471f
C24182 VDD a_27062_3134# 0.483f
C24183 col_n[23] rowoff_n[9] 0.0471f
C24184 col_n[18] rowoff_n[4] 0.0471f
C24185 col_n[20] rowoff_n[6] 0.0471f
C24186 col[29] a_2475_3158# 0.136f
C24187 col_n[17] rowoff_n[3] 0.0471f
C24188 col_n[21] rowoff_n[7] 0.0471f
C24189 col_n[15] rowoff_n[1] 0.0471f
C24190 col_n[14] rowoff_n[0] 0.0471f
C24191 col_n[22] rowoff_n[8] 0.0471f
C24192 m2_14784_18014# a_15318_18234# 0.087f
C24193 a_2275_16210# a_31990_16186# 0.136f
C24194 rowon_n[3] a_21038_5142# 0.248f
C24195 VDD a_16418_12532# 0.0779f
C24196 vcm a_2475_18218# 1.08f
C24197 sample a_2161_18218# 0.0858f
C24198 ctop a_31078_17190# 4.06f
C24199 m2_3164_10410# rowon_n[8] 0.0322f
C24200 m2_9188_6394# rowon_n[4] 0.0322f
C24201 m2_14208_2378# rowon_n[0] 0.0322f
C24202 a_23958_4138# a_24050_4138# 0.326f
C24203 col_n[9] a_12002_12170# 0.251f
C24204 col_n[6] a_8898_2130# 0.0765f
C24205 ctop a_33998_2130# 0.0293f
C24206 vcm a_11910_16186# 0.1f
C24207 a_30074_14178# a_30074_13174# 0.843f
C24208 a_2475_13198# a_24050_13174# 0.316f
C24209 VDD a_7986_6146# 0.483f
C24210 col_n[16] a_18938_14178# 0.0765f
C24211 col[21] a_2275_17214# 0.0899f
C24212 a_23958_18194# a_24354_18234# 0.0313f
C24213 VDD a_31478_16548# 0.0779f
C24214 a_18938_1126# a_19334_1166# 0.0346f
C24215 col[26] a_2275_6170# 0.0899f
C24216 row_n[12] a_32082_14178# 0.282f
C24217 col[24] rowoff_n[14] 0.0901f
C24218 vcm a_14010_1126# 0.165f
C24219 m2_24248_15430# rowon_n[13] 0.0322f
C24220 m2_30272_11414# rowon_n[9] 0.0322f
C24221 m2_35292_7398# rowon_n[5] 0.0322f
C24222 m2_16216_9406# a_16018_9158# 0.165f
C24223 m3_5880_18146# m3_6884_18146# 0.202f
C24224 vcm a_2966_10162# 0.56f
C24225 col_n[7] rowoff_n[10] 0.0471f
C24226 a_7986_10162# a_8290_10202# 0.0931f
C24227 a_2275_10186# a_15014_10162# 0.399f
C24228 a_8898_10162# a_9390_10524# 0.0658f
C24229 row_n[14] a_19334_16226# 0.0117f
C24230 a_20034_15182# a_21038_15182# 0.843f
C24231 VDD a_23046_10162# 0.483f
C24232 col[29] a_32082_11166# 0.367f
C24233 row_n[4] a_29374_6186# 0.0117f
C24234 m2_34864_4962# a_35094_5142# 0.0249f
C24235 col_n[11] a_2475_13198# 0.0531f
C24236 vcm a_29070_5142# 0.56f
C24237 a_3878_7150# a_4274_7190# 0.0313f
C24238 rowoff_n[2] a_5978_4138# 0.294f
C24239 rowoff_n[10] a_23046_12170# 0.294f
C24240 a_4882_7150# a_4974_7150# 0.326f
C24241 a_2275_7174# a_5278_7190# 0.144f
C24242 a_2475_7174# a_7894_7150# 0.264f
C24243 col_n[16] a_2475_2154# 0.0531f
C24244 row_n[6] a_19942_8154# 0.0437f
C24245 a_2275_12194# a_30074_12170# 0.399f
C24246 rowon_n[10] a_19030_12170# 0.248f
C24247 col_n[24] a_27366_11206# 0.084f
C24248 row_n[0] m2_30272_2378# 0.0128f
C24249 a_10998_17190# a_10998_16186# 0.843f
C24250 VDD a_3970_13174# 0.483f
C24251 col_n[5] a_7894_12170# 0.0765f
C24252 VDD col_n[24] 5.17f
C24253 col_n[10] col_n[11] 0.0101f
C24254 vcm col_n[21] 1.94f
C24255 col[20] col[21] 0.0355f
C24256 col[8] rowoff_n[15] 0.0901f
C24257 col[1] a_2475_10186# 0.136f
C24258 rowoff_n[0] a_15014_2130# 0.294f
C24259 rowon_n[0] a_29070_2130# 0.248f
C24260 m2_7180_7398# a_6982_7150# 0.165f
C24261 vcm a_9994_8154# 0.56f
C24262 a_2275_9182# a_20338_9198# 0.144f
C24263 a_2475_9182# a_22954_9158# 0.264f
C24264 col_n[8] a_2275_16210# 0.113f
C24265 a_23958_14178# a_24450_14540# 0.0658f
C24266 a_23046_14178# a_23350_14218# 0.0931f
C24267 col_n[13] a_2275_5166# 0.113f
C24268 row_n[0] a_6982_2130# 0.282f
C24269 VDD a_19030_17190# 0.484f
C24270 col[18] a_21038_9158# 0.367f
C24271 a_30074_2130# a_31078_2130# 0.843f
C24272 rowon_n[4] a_6890_6146# 0.118f
C24273 m2_26256_3382# a_26058_3134# 0.165f
C24274 col[25] a_27974_11166# 0.0682f
C24275 vcm a_35398_3174# 0.161f
C24276 a_2275_6170# a_13918_6146# 0.136f
C24277 col_n[28] a_2475_15206# 0.0531f
C24278 col_n[0] a_3270_5182# 0.084f
C24279 vcm a_25054_12170# 0.56f
C24280 a_2275_11190# a_2275_10186# 0.0715f
C24281 a_19942_11166# a_20034_11166# 0.326f
C24282 col[3] a_2275_2154# 0.0899f
C24283 VDD a_21950_2130# 0.181f
C24284 m2_2160_9406# row_n[7] 0.0194f
C24285 m2_8184_5390# row_n[3] 0.0128f
C24286 row_n[11] a_27366_13214# 0.0117f
C24287 col_n[13] a_16322_9198# 0.084f
C24288 col[18] a_2475_12194# 0.136f
C24289 a_2966_3134# a_3270_3174# 0.0931f
C24290 a_3878_3134# a_4370_3496# 0.0658f
C24291 a_2475_3158# a_5978_3134# 0.316f
C24292 a_21038_4138# a_21038_3134# 0.843f
C24293 rowoff_n[8] a_7894_10162# 0.202f
C24294 col[23] a_2475_1150# 0.136f
C24295 row_n[13] a_17934_15182# 0.0437f
C24296 vcm a_15318_6186# 0.155f
C24297 a_2275_8178# a_28978_8154# 0.136f
C24298 a_14922_8154# a_15318_8194# 0.0313f
C24299 rowoff_n[11] a_10998_13174# 0.294f
C24300 col_n[24] a_27462_3496# 0.0283f
C24301 vcm a_5978_15182# 0.56f
C24302 VDD a_2161_5166# 0.187f
C24303 row_n[3] a_27974_5142# 0.0437f
C24304 col_n[25] a_2275_18218# 0.113f
C24305 a_3970_17190# a_4274_17230# 0.0931f
C24306 rowon_n[7] a_27062_9158# 0.248f
C24307 a_4882_17190# a_5374_17552# 0.0658f
C24308 a_2275_17214# a_6982_17190# 0.399f
C24309 m2_23244_14426# row_n[12] 0.0128f
C24310 col_n[30] a_2275_7174# 0.113f
C24311 rowoff_n[6] a_16930_8154# 0.202f
C24312 m2_29268_10410# row_n[8] 0.0128f
C24313 m2_34864_5966# row_n[4] 0.267f
C24314 a_10998_5142# a_12002_5142# 0.843f
C24315 col[7] a_9994_7150# 0.367f
C24316 a_2475_5166# a_21038_5142# 0.316f
C24317 vcm a_30378_10202# 0.155f
C24318 col[14] a_16930_9158# 0.0682f
C24319 rowoff_n[15] a_27062_17190# 0.294f
C24320 col[15] a_2275_15206# 0.0899f
C24321 rowoff_n[4] a_25966_6146# 0.202f
C24322 ctop a_8990_4138# 4.11f
C24323 col[20] a_2275_4162# 0.0899f
C24324 a_35002_15182# a_35094_15182# 0.0991f
C24325 a_34090_15182# a_34394_15222# 0.0931f
C24326 m2_7756_946# a_2475_1150# 0.286f
C24327 col_n[22] a_25054_3134# 0.251f
C24328 VDD a_17934_9158# 0.181f
C24329 row_n[7] a_4974_9158# 0.282f
C24330 col[18] a_19942_1126# 0.011f
C24331 rowon_n[11] a_4882_13174# 0.118f
C24332 col_n[29] a_31990_5142# 0.0765f
C24333 VDD a_5278_18234# 0.019f
C24334 a_2275_2154# a_12002_2130# 0.399f
C24335 col_n[2] a_5278_7190# 0.084f
C24336 vcm a_23958_4138# 0.1f
C24337 rowon_n[1] a_14922_3134# 0.118f
C24338 col_n[26] rowoff_n[1] 0.0471f
C24339 col_n[28] rowoff_n[3] 0.0471f
C24340 col_n[30] rowoff_n[5] 0.0471f
C24341 rowoff_n[2] a_35002_4138# 0.202f
C24342 a_2475_7174# a_2475_6170# 0.0666f
C24343 rowoff_n[9] a_17422_11528# 0.0133f
C24344 col_n[25] rowoff_n[0] 0.0471f
C24345 col_n[27] rowoff_n[2] 0.0471f
C24346 col_n[31] rowoff_n[6] 0.0471f
C24347 col_n[29] rowoff_n[4] 0.0471f
C24348 vcm a_11302_13214# 0.155f
C24349 a_29982_12170# a_30378_12210# 0.0313f
C24350 VDD a_9390_3496# 0.0779f
C24351 col_n[11] a_2475_18218# 0.0529f
C24352 col_n[13] a_16418_1488# 0.0283f
C24353 ctop a_24050_8154# 4.11f
C24354 a_2275_16210# a_12306_16226# 0.144f
C24355 a_2475_16210# a_14922_16186# 0.264f
C24356 rowon_n[3] a_2966_5142# 0.248f
C24357 col_n[23] a_26458_13536# 0.0283f
C24358 VDD a_32994_13174# 0.181f
C24359 col_n[5] a_2475_11190# 0.0531f
C24360 rowoff_n[7] a_26458_9520# 0.0133f
C24361 a_14010_4138# a_14314_4178# 0.0931f
C24362 a_14922_4138# a_15414_4500# 0.0658f
C24363 a_2275_4162# a_27062_4138# 0.399f
C24364 m3_29976_1078# ctop 0.21f
C24365 vcm a_4882_7150# 0.1f
C24366 a_26058_9158# a_27062_9158# 0.843f
C24367 rowoff_n[13] a_33486_15544# 0.0133f
C24368 row_n[10] a_25966_12170# 0.0437f
C24369 col[6] a_8990_17190# 0.367f
C24370 vcm a_26362_17230# 0.155f
C24371 rowon_n[14] a_25054_16186# 0.248f
C24372 a_2275_13198# a_5886_13174# 0.136f
C24373 col[3] a_5886_7150# 0.0682f
C24374 VDD a_24450_7512# 0.0779f
C24375 rowoff_n[5] a_35494_7512# 0.0133f
C24376 ctop a_4974_11166# 4.11f
C24377 a_2275_18218# a_27366_18234# 0.145f
C24378 a_15926_18194# a_16018_18194# 0.0991f
C24379 VDD a_13918_16186# 0.181f
C24380 row_n[0] a_34394_2170# 0.0117f
C24381 a_2475_1150# a_19942_1126# 0.285f
C24382 a_2275_1150# a_17326_1166# 0.145f
C24383 a_10906_1126# a_10998_1126# 0.0991f
C24384 rowon_n[4] a_35094_6146# 0.0141f
C24385 col_n[21] a_24050_13174# 0.251f
C24386 col_n[18] a_20946_3134# 0.0765f
C24387 col_n[18] rowoff_n[10] 0.0471f
C24388 col_n[28] a_30986_15182# 0.0765f
C24389 col_n[2] a_2275_14202# 0.113f
C24390 m2_1732_8978# a_2475_9182# 0.139f
C24391 vcm a_19942_11166# 0.1f
C24392 col_n[7] a_2275_3158# 0.113f
C24393 col_n[1] a_4274_17230# 0.084f
C24394 a_17022_11166# a_17022_10162# 0.843f
C24395 row_n[14] a_2874_16186# 0.0436f
C24396 VDD a_16018_1126# 0.035f
C24397 sample a_1957_7174# 0.345f
C24398 a_2275_15206# a_20946_15182# 0.136f
C24399 a_10906_15182# a_11302_15222# 0.0313f
C24400 VDD a_5374_10524# 0.0779f
C24401 ctop a_20034_15182# 4.11f
C24402 row_n[4] a_13006_6146# 0.282f
C24403 col_n[22] a_2475_13198# 0.0531f
C24404 col_n[12] a_15414_11528# 0.0283f
C24405 col_n[27] a_2475_2154# 0.0531f
C24406 a_2275_3158# a_32386_3174# 0.144f
C24407 a_2475_3158# a_35002_3134# 0.264f
C24408 rowon_n[8] a_12914_10162# 0.118f
C24409 rowoff_n[10] a_5374_12532# 0.0133f
C24410 a_29982_8154# a_30474_8516# 0.0658f
C24411 a_29070_8154# a_29374_8194# 0.0931f
C24412 a_23350_1166# vcm 0.16f
C24413 vcm a_35002_15182# 0.101f
C24414 a_6982_12170# a_7986_12170# 0.843f
C24415 a_2475_12194# a_13006_12170# 0.316f
C24416 VDD a_31078_5142# 0.483f
C24417 col_n[0] row_n[15] 0.298f
C24418 vcm rowon_n[15] 0.65f
C24419 sample rowon_n[14] 0.0935f
C24420 VDD row_n[14] 3.29f
C24421 m2_20232_18442# VDD 0.0456f
C24422 col[19] rowoff_n[15] 0.0901f
C24423 col[12] a_2475_10186# 0.136f
C24424 col_n[0] a_3366_17552# 0.0283f
C24425 row_n[15] a_33390_17230# 0.0117f
C24426 a_2275_17214# a_34394_17230# 0.144f
C24427 VDD a_20434_14540# 0.0779f
C24428 a_35094_2130# m2_34864_1950# 0.0249f
C24429 col_n[2] rowoff_n[11] 0.0471f
C24430 col[2] a_4882_17190# 0.0682f
C24431 a_25966_5142# a_26058_5142# 0.326f
C24432 col_n[10] a_13006_11166# 0.251f
C24433 m2_11772_18014# col_n[9] 0.243f
C24434 col_n[7] a_9902_1126# 0.0765f
C24435 col_n[19] a_2275_16210# 0.113f
C24436 a_2275_9182# a_3970_9158# 0.399f
C24437 rowoff_n[14] a_21438_16548# 0.0133f
C24438 col_n[24] a_2275_5166# 0.113f
C24439 col_n[17] a_19942_13174# 0.0765f
C24440 vcm a_15926_18194# 0.101f
C24441 m3_27968_1078# a_28066_2130# 0.0302f
C24442 m2_7180_17438# rowon_n[15] 0.0322f
C24443 a_32082_15182# a_32082_14178# 0.843f
C24444 a_2475_14202# a_28066_14178# 0.316f
C24445 m2_13204_13422# rowon_n[11] 0.0322f
C24446 VDD a_12002_8154# 0.483f
C24447 row_n[7] a_33998_9158# 0.0437f
C24448 m2_19228_9406# rowon_n[7] 0.0322f
C24449 m2_25252_5390# rowon_n[3] 0.0322f
C24450 rowon_n[11] a_33086_13174# 0.248f
C24451 VDD a_35494_18556# 0.114f
C24452 a_20946_2130# a_21342_2170# 0.0313f
C24453 col[9] a_2275_13198# 0.0899f
C24454 vcm a_18026_3134# 0.56f
C24455 col[14] a_2275_2154# 0.0899f
C24456 col_n[1] a_4370_9520# 0.0283f
C24457 a_10906_11166# a_11398_11528# 0.0658f
C24458 a_2275_11190# a_19030_11166# 0.399f
C24459 a_9994_11166# a_10298_11206# 0.0931f
C24460 VDD a_3878_2130# 0.181f
C24461 col[30] a_33086_10162# 0.367f
C24462 row_n[11] a_10998_13174# 0.282f
C24463 a_22042_16186# a_23046_16186# 0.843f
C24464 col[29] a_2475_12194# 0.136f
C24465 VDD a_27062_12170# 0.483f
C24466 m2_15788_18014# m3_15920_18146# 3.79f
C24467 rowon_n[15] a_10906_17190# 0.118f
C24468 row_n[1] a_21038_3134# 0.282f
C24469 rowoff_n[1] a_6982_3134# 0.294f
C24470 vcm a_33086_7150# 0.56f
C24471 rowon_n[5] a_20946_7150# 0.118f
C24472 rowoff_n[12] a_27974_14178# 0.202f
C24473 a_6890_8154# a_6982_8154# 0.326f
C24474 a_2475_8178# a_11910_8154# 0.264f
C24475 a_2275_8178# a_9294_8194# 0.144f
C24476 col_n[0] a_2475_9182# 0.0532f
C24477 col_n[25] a_28370_10202# 0.084f
C24478 m2_1732_11990# sample 0.2f
C24479 a_2275_13198# a_34090_13174# 0.399f
C24480 m2_34864_5966# ctop 0.0422f
C24481 row_n[3] a_8290_5182# 0.0117f
C24482 col_n[6] a_8898_11166# 0.0765f
C24483 VDD a_7986_15182# 0.483f
C24484 col[26] a_2275_15206# 0.0899f
C24485 a_2475_5166# a_2966_5142# 0.317f
C24486 a_2161_5166# a_2275_5166# 0.183f
C24487 col[31] a_2275_4162# 0.0899f
C24488 vcm a_14010_10162# 0.56f
C24489 a_2475_10186# a_26970_10162# 0.264f
C24490 a_2275_10186# a_24354_10202# 0.144f
C24491 rowoff_n[15] a_9390_17552# 0.0133f
C24492 row_n[14] a_31990_16186# 0.0437f
C24493 m2_12200_16434# a_12002_16186# 0.165f
C24494 a_25966_15182# a_26458_15544# 0.0658f
C24495 a_25054_15182# a_25358_15222# 0.0931f
C24496 m2_8760_18014# ctop 0.0422f
C24497 col[19] a_22042_8154# 0.367f
C24498 row_n[9] rowoff_n[9] 0.209f
C24499 col[26] a_28978_10162# 0.0682f
C24500 a_32082_3134# a_33086_3134# 0.843f
C24501 col_n[1] a_2275_1150# 0.0947f
C24502 m2_34864_3958# a_2275_4162# 0.278f
C24503 vcm a_4274_4178# 0.155f
C24504 a_2275_7174# a_17934_7150# 0.136f
C24505 col_n[22] a_2475_18218# 0.0529f
C24506 m2_31276_12418# a_31078_12170# 0.165f
C24507 vcm a_29070_14178# 0.56f
C24508 a_21950_12170# a_22042_12170# 0.326f
C24509 VDD a_25966_4138# 0.181f
C24510 col_n[16] a_2475_11190# 0.0531f
C24511 col_n[14] a_17326_8194# 0.084f
C24512 row_n[8] a_19030_10162# 0.282f
C24513 rowoff_n[7] a_8898_9158# 0.202f
C24514 m3_34996_16138# a_34090_16186# 0.0303f
C24515 rowon_n[12] a_18938_14178# 0.118f
C24516 a_2475_4162# a_9994_4138# 0.316f
C24517 a_23046_5142# a_23046_4138# 0.843f
C24518 m3_25960_18146# ctop 0.209f
C24519 col_n[25] a_28466_2492# 0.0283f
C24520 m2_6176_16434# row_n[14] 0.0128f
C24521 m2_12200_12418# row_n[10] 0.0128f
C24522 col[6] a_2475_8178# 0.136f
C24523 vcm a_19334_8194# 0.155f
C24524 rowoff_n[13] a_15926_15182# 0.202f
C24525 a_2275_9182# a_32994_9158# 0.136f
C24526 m2_18224_8402# row_n[6] 0.0128f
C24527 a_16930_9158# a_17326_9198# 0.0313f
C24528 m2_24248_4386# row_n[2] 0.0128f
C24529 row_n[10] a_6282_12210# 0.0117f
C24530 rowon_n[2] a_28978_4138# 0.118f
C24531 ctop a_32082_3134# 4.11f
C24532 vcm a_9994_17190# 0.56f
C24533 VDD a_6890_7150# 0.181f
C24534 rowoff_n[5] a_17934_7150# 0.202f
C24535 col_n[29] rowoff_n[10] 0.0471f
C24536 a_6890_18194# a_7382_18556# 0.0658f
C24537 a_2275_18218# a_10998_18194# 0.0924f
C24538 row_n[0] a_16322_2170# 0.0117f
C24539 col_n[13] a_2275_14202# 0.113f
C24540 col[8] a_10998_6146# 0.367f
C24541 m2_34864_2954# a_35002_3134# 0.225f
C24542 col_n[18] a_2275_3158# 0.113f
C24543 vcm a_12914_2130# 0.1f
C24544 m2_1732_5966# m2_2160_6394# 0.165f
C24545 a_13006_6146# a_14010_6146# 0.843f
C24546 a_2475_6170# a_25054_6146# 0.316f
C24547 col[15] a_17934_8154# 0.0682f
C24548 m2_22240_10410# a_22042_10162# 0.165f
C24549 row_n[2] a_6890_4138# 0.0437f
C24550 vcm a_35398_12210# 0.161f
C24551 rowoff_n[3] a_26970_5142# 0.202f
C24552 VDD a_32482_2492# 0.0779f
C24553 col_n[23] a_26058_2130# 0.251f
C24554 m2_33284_17438# row_n[15] 0.0128f
C24555 rowon_n[6] a_5978_8154# 0.248f
C24556 col_n[0] a_3270_14218# 0.084f
C24557 ctop a_13006_6146# 4.11f
C24558 VDD a_21950_11166# 0.181f
C24559 col_n[30] a_32994_4138# 0.0765f
C24560 col[3] a_2275_11190# 0.0899f
C24561 col_n[3] a_6282_6186# 0.084f
C24562 a_2275_3158# a_16018_3134# 0.399f
C24563 col_n[13] a_16322_18234# 0.084f
C24564 a_2475_18218# a_8990_18194# 0.0299f
C24565 rowoff_n[8] a_18426_10524# 0.0133f
C24566 en_bit_n[2] a_19030_1126# 0.208f
C24567 a_29982_1126# a_2275_1150# 0.136f
C24568 vcm a_27974_6146# 0.1f
C24569 a_3970_8154# a_3970_7150# 0.843f
C24570 VDD rowon_n[8] 3.04f
C24571 col_n[8] row_n[14] 0.298f
C24572 col_n[7] rowon_n[13] 0.111f
C24573 col_n[9] rowon_n[14] 0.111f
C24574 col_n[10] row_n[15] 0.298f
C24575 sample row_n[9] 0.423f
C24576 col_n[11] rowon_n[15] 0.111f
C24577 col_n[0] rowon_n[9] 0.111f
C24578 vcm row_n[10] 0.616f
C24579 col_n[6] row_n[13] 0.298f
C24580 col_n[5] rowon_n[12] 0.111f
C24581 col_n[21] col_n[22] 0.0101f
C24582 col_n[1] rowon_n[10] 0.111f
C24583 col_n[2] row_n[11] 0.298f
C24584 col_n[4] row_n[12] 0.298f
C24585 col_n[3] rowon_n[11] 0.111f
C24586 col[30] rowoff_n[15] 0.0901f
C24587 col[23] a_2475_10186# 0.136f
C24588 m3_34996_1078# m2_34864_1950# 0.0341f
C24589 vcm a_15318_15222# 0.155f
C24590 a_31990_13174# a_32386_13214# 0.0313f
C24591 VDD a_13406_5504# 0.0779f
C24592 col_n[24] a_27462_12532# 0.0283f
C24593 col_n[13] rowoff_n[11] 0.0471f
C24594 a_25358_1166# VDD 0.0149f
C24595 ctop a_28066_10162# 4.11f
C24596 row_n[15] a_17022_17190# 0.282f
C24597 a_2275_17214# a_16322_17230# 0.144f
C24598 a_2475_17214# a_18938_17190# 0.264f
C24599 rowoff_n[6] a_27462_8516# 0.0133f
C24600 VDD a_2161_14202# 0.187f
C24601 col_n[30] a_2275_16210# 0.113f
C24602 a_16930_5142# a_17422_5504# 0.0658f
C24603 a_16018_5142# a_16322_5182# 0.0931f
C24604 row_n[5] a_27062_7150# 0.282f
C24605 a_2275_5166# a_31078_5142# 0.399f
C24606 m2_13204_8402# a_13006_8154# 0.165f
C24607 rowon_n[9] a_26970_11166# 0.118f
C24608 vcm a_8898_9158# 0.1f
C24609 rowoff_n[14] a_3366_16548# 0.0133f
C24610 col[7] a_9994_16186# 0.367f
C24611 a_28066_10162# a_29070_10162# 0.843f
C24612 col[4] a_6890_6146# 0.0682f
C24613 col[14] a_16930_18194# 0.0682f
C24614 a_2275_14202# a_9902_14178# 0.136f
C24615 m2_9764_946# a_10298_1166# 0.087f
C24616 m2_30848_946# a_2475_1150# 0.286f
C24617 row_n[7] a_14314_9198# 0.0117f
C24618 VDD a_28466_9520# 0.0779f
C24619 col[20] a_2275_13198# 0.0899f
C24620 ctop a_8990_13174# 4.11f
C24621 col_n[22] a_25054_12170# 0.251f
C24622 VDD a_17934_18194# 0.343f
C24623 col_n[19] a_21950_2130# 0.0765f
C24624 col[25] a_2275_2154# 0.0899f
C24625 a_12914_2130# a_13006_2130# 0.326f
C24626 a_2475_2154# a_23958_2130# 0.264f
C24627 a_2275_2154# a_21342_2170# 0.144f
C24628 m2_32280_4386# a_32082_4138# 0.165f
C24629 col_n[29] a_31990_14178# 0.0765f
C24630 m2_23820_946# VDD 1f
C24631 row_n[9] a_4882_11166# 0.0437f
C24632 m2_34864_9982# m2_34864_8978# 0.843f
C24633 rowoff_n[9] a_28066_11166# 0.294f
C24634 col_n[2] a_5278_16226# 0.084f
C24635 rowon_n[13] a_3970_15182# 0.248f
C24636 col_n[0] a_2966_6146# 0.251f
C24637 vcm a_23958_13174# 0.1f
C24638 a_19030_12170# a_19030_11166# 0.843f
C24639 VDD rowoff_n[12] 1.51f
C24640 VDD a_20034_3134# 0.483f
C24641 m2_28840_18014# a_2275_18218# 0.28f
C24642 a_2275_16210# a_24962_16186# 0.136f
C24643 a_12914_16186# a_13310_16226# 0.0313f
C24644 VDD a_9390_12532# 0.0779f
C24645 rowon_n[3] a_14010_5142# 0.248f
C24646 a_30986_1126# m2_30848_946# 0.225f
C24647 col_n[13] a_16418_10524# 0.0283f
C24648 ctop a_24050_17190# 4.06f
C24649 a_2966_4138# a_2966_3134# 0.843f
C24650 row_n[1] a_2966_3134# 0.281f
C24651 col_n[10] a_2475_9182# 0.0531f
C24652 m2_4168_6394# a_3970_6146# 0.165f
C24653 rowon_n[5] a_2275_7174# 1.79f
C24654 a_31078_9158# a_31382_9198# 0.0931f
C24655 a_31990_9158# a_32482_9520# 0.0658f
C24656 vcm a_4882_16186# 0.1f
C24657 a_2475_13198# a_17022_13174# 0.316f
C24658 a_8990_13174# a_9994_13174# 0.843f
C24659 m2_24824_18014# a_2475_18218# 0.286f
C24660 VDD a_24450_16548# 0.0779f
C24661 col[3] a_5886_16186# 0.0682f
C24662 col[0] a_2475_6170# 0.148f
C24663 row_n[12] a_25054_14178# 0.282f
C24664 col_n[11] a_14010_10162# 0.251f
C24665 vcm a_6982_1126# 0.165f
C24666 a_27974_6146# a_28066_6146# 0.326f
C24667 m2_2160_11414# rowon_n[9] 0.0219f
C24668 m2_8184_7398# rowon_n[5] 0.0322f
C24669 m2_30848_946# m2_31276_1374# 0.165f
C24670 m2_14208_3382# rowon_n[1] 0.0322f
C24671 col_n[18] a_20946_12170# 0.0765f
C24672 row_n[2] a_35094_4138# 0.0123f
C24673 a_2275_10186# a_7986_10162# 0.399f
C24674 row_n[14] a_12306_16226# 0.0117f
C24675 rowon_n[6] a_35002_8154# 0.118f
C24676 col_n[7] a_2275_12194# 0.113f
C24677 a_2475_15206# a_32082_15182# 0.316f
C24678 a_34090_16186# a_34090_15182# 0.843f
C24679 rowon_n[5] rowoff_n[5] 20.2f
C24680 VDD a_16018_10162# 0.483f
C24681 col_n[12] a_2275_1150# 0.113f
C24682 sample a_1957_16210# 0.345f
C24683 row_n[4] a_22346_6186# 0.0117f
C24684 a_22954_3134# a_23350_3174# 0.0313f
C24685 col_n[2] a_5374_8516# 0.0283f
C24686 vcm a_22042_5142# 0.56f
C24687 col_n[27] a_2475_11190# 0.0531f
C24688 rowoff_n[10] a_16018_12170# 0.294f
C24689 a_29470_1488# col_n[26] 0.0283f
C24690 m2_23244_16434# rowon_n[14] 0.0322f
C24691 m2_29268_12418# rowon_n[10] 0.0322f
C24692 row_n[6] a_12914_8154# 0.0437f
C24693 col[31] a_34090_9158# 0.367f
C24694 m2_34864_7974# rowon_n[6] 0.231f
C24695 a_12914_12170# a_13406_12532# 0.0658f
C24696 a_2275_12194# a_23046_12170# 0.399f
C24697 a_12002_12170# a_12306_12210# 0.0931f
C24698 rowon_n[10] a_12002_12170# 0.248f
C24699 a_24050_17190# a_25054_17190# 0.843f
C24700 VDD a_31078_14178# 0.483f
C24701 rowoff_n[0] a_7986_2130# 0.294f
C24702 rowon_n[0] a_22042_2130# 0.248f
C24703 col[17] a_2475_8178# 0.136f
C24704 m2_10768_946# ctop 0.0428f
C24705 vcm a_2874_8154# 0.1f
C24706 col_n[26] a_29374_9198# 0.084f
C24707 a_2475_9182# a_15926_9158# 0.264f
C24708 a_2275_9182# a_13310_9198# 0.144f
C24709 rowoff_n[14] a_32082_16186# 0.294f
C24710 a_8898_9158# a_8990_9158# 0.326f
C24711 col_n[7] a_9902_10162# 0.0765f
C24712 col_n[24] a_2275_14202# 0.113f
C24713 m2_28840_946# col_n[26] 0.362f
C24714 col_n[29] a_2275_3158# 0.113f
C24715 VDD a_12002_17190# 0.484f
C24716 m3_24956_1078# VDD 0.0157f
C24717 vcm a_27366_3174# 0.155f
C24718 row_n[9] a_33086_11166# 0.282f
C24719 a_2275_6170# a_6890_6146# 0.136f
C24720 m2_26832_18014# col[24] 0.347f
C24721 rowon_n[13] a_32994_15182# 0.118f
C24722 vcm a_18026_12170# 0.56f
C24723 a_2475_11190# a_30986_11166# 0.264f
C24724 col_n[1] a_4370_18556# 0.0283f
C24725 col[14] a_2275_11190# 0.0899f
C24726 a_2275_11190# a_28370_11206# 0.144f
C24727 VDD a_14922_2130# 0.181f
C24728 col[20] a_23046_7150# 0.367f
C24729 a_27062_16186# a_27366_16226# 0.0931f
C24730 row_n[11] a_20338_13214# 0.0117f
C24731 a_27974_16186# a_28466_16548# 0.0658f
C24732 VDD a_3878_11166# 0.181f
C24733 m2_29844_18014# m3_30980_18146# 0.0341f
C24734 col[27] a_29982_9158# 0.0682f
C24735 VDD row_n[3] 3.29f
C24736 col_n[20] rowon_n[14] 0.111f
C24737 col_n[1] row_n[5] 0.298f
C24738 col_n[0] row_n[4] 0.298f
C24739 vcm rowon_n[4] 0.65f
C24740 col_n[15] row_n[12] 0.298f
C24741 col_n[8] rowon_n[8] 0.111f
C24742 col_n[2] rowon_n[5] 0.111f
C24743 col_n[21] row_n[15] 0.298f
C24744 col_n[16] rowon_n[12] 0.111f
C24745 col_n[11] row_n[10] 0.298f
C24746 col_n[5] row_n[7] 0.298f
C24747 col_n[4] rowon_n[6] 0.111f
C24748 col_n[14] rowon_n[11] 0.111f
C24749 col_n[19] row_n[14] 0.298f
C24750 col_n[12] rowon_n[10] 0.111f
C24751 col_n[10] rowon_n[9] 0.111f
C24752 col_n[3] row_n[6] 0.298f
C24753 col_n[13] row_n[11] 0.298f
C24754 col_n[9] row_n[9] 0.298f
C24755 col_n[22] rowon_n[15] 0.111f
C24756 sample rowon_n[3] 0.0935f
C24757 col_n[17] row_n[13] 0.298f
C24758 col_n[6] rowon_n[7] 0.111f
C24759 col_n[7] row_n[8] 0.298f
C24760 col_n[18] rowon_n[13] 0.111f
C24761 a_33998_4138# a_34394_4178# 0.0313f
C24762 row_n[1] a_30378_3174# 0.0117f
C24763 row_n[13] a_10906_15182# 0.0437f
C24764 vcm a_8290_6186# 0.155f
C24765 rowoff_n[11] a_3970_13174# 0.294f
C24766 a_2275_8178# a_21950_8154# 0.136f
C24767 col_n[24] rowoff_n[11] 0.0471f
C24768 vcm a_33086_16186# 0.56f
C24769 a_23958_13174# a_24050_13174# 0.326f
C24770 col_n[15] a_18330_7190# 0.084f
C24771 VDD a_29982_6146# 0.181f
C24772 row_n[3] a_20946_5142# 0.0437f
C24773 rowon_n[7] a_20034_9158# 0.248f
C24774 m2_1732_9982# row_n[8] 0.292f
C24775 rowoff_n[6] a_9902_8154# 0.202f
C24776 col_n[4] a_2475_7174# 0.0531f
C24777 m2_7180_6394# row_n[4] 0.0128f
C24778 m2_12200_2378# row_n[0] 0.0128f
C24779 m3_10900_18146# a_10998_17190# 0.0303f
C24780 a_2475_5166# a_14010_5142# 0.316f
C24781 a_25054_6146# a_25054_5142# 0.843f
C24782 m2_33860_946# m3_33992_1078# 1.11f
C24783 vcm a_23350_10202# 0.155f
C24784 a_18938_10162# a_19334_10202# 0.0313f
C24785 rowoff_n[15] a_20034_17190# 0.294f
C24786 rowoff_n[4] a_18938_6146# 0.202f
C24787 col[31] a_2275_13198# 0.0899f
C24788 ctop a_2475_4162# 0.0488f
C24789 m3_34996_3086# a_34090_3134# 0.0303f
C24790 VDD a_10906_9158# 0.181f
C24791 col[9] a_12002_5142# 0.367f
C24792 a_3878_2130# a_3970_2130# 0.326f
C24793 col[19] a_22042_17190# 0.367f
C24794 a_2275_2154# a_4974_2130# 0.399f
C24795 m2_22240_15430# row_n[13] 0.0128f
C24796 a_2874_2130# a_3270_2170# 0.0313f
C24797 m2_28264_11414# row_n[9] 0.0128f
C24798 m2_34288_7398# row_n[5] 0.0128f
C24799 col[16] a_18938_7150# 0.0682f
C24800 vcm a_16930_4138# 0.1f
C24801 rowoff_n[9] a_10394_11528# 0.0133f
C24802 a_2475_7174# a_29070_7150# 0.316f
C24803 col_n[1] a_2275_10186# 0.113f
C24804 rowon_n[1] a_7894_3134# 0.118f
C24805 rowoff_n[2] a_27974_4138# 0.202f
C24806 a_15014_7150# a_16018_7150# 0.843f
C24807 col_n[8] rowoff_n[12] 0.0471f
C24808 vcm a_4274_13214# 0.155f
C24809 VDD a_1957_3158# 0.196f
C24810 col_n[31] a_33998_3134# 0.0765f
C24811 ctop a_17022_8154# 4.11f
C24812 a_3878_16186# a_4274_16226# 0.0313f
C24813 a_4882_16186# a_4974_16186# 0.326f
C24814 a_2475_16210# a_7894_16186# 0.264f
C24815 a_2275_16210# a_5278_16226# 0.144f
C24816 VDD a_25966_13174# 0.181f
C24817 col_n[4] a_7286_5182# 0.084f
C24818 col[0] a_2966_3134# 0.367f
C24819 col_n[21] a_2475_9182# 0.0531f
C24820 row_n[8] a_28370_10202# 0.0117f
C24821 col_n[14] a_17326_17230# 0.084f
C24822 rowoff_n[7] a_19430_9520# 0.0133f
C24823 a_2275_4162# a_20034_4138# 0.399f
C24824 vcm a_31990_8154# 0.1f
C24825 a_5978_9158# a_5978_8154# 0.843f
C24826 rowoff_n[13] a_26458_15544# 0.0133f
C24827 row_n[10] a_18938_12170# 0.0437f
C24828 col_n[25] a_28466_11528# 0.0283f
C24829 col[6] a_2475_17214# 0.136f
C24830 vcm a_19334_17230# 0.155f
C24831 rowon_n[14] a_18026_16186# 0.248f
C24832 m2_1732_8978# ctop 0.0428f
C24833 VDD a_17422_7512# 0.0779f
C24834 rowoff_n[5] a_28466_7512# 0.0133f
C24835 col[11] a_2475_6170# 0.136f
C24836 ctop a_32082_12170# 4.11f
C24837 a_2275_18218# a_20338_18234# 0.145f
C24838 VDD a_6890_16186# 0.181f
C24839 row_n[0] a_28978_2130# 0.0437f
C24840 a_2475_1150# a_12914_1126# 0.264f
C24841 a_2275_1150# a_10298_1166# 0.145f
C24842 rowon_n[4] a_28066_6146# 0.248f
C24843 a_18938_6146# a_19430_6508# 0.0658f
C24844 a_2275_6170# a_35094_6146# 0.0924f
C24845 a_18026_6146# a_18330_6186# 0.0931f
C24846 col[8] a_10998_15182# 0.367f
C24847 col[5] a_7894_5142# 0.0682f
C24848 col_n[18] a_2275_12194# 0.113f
C24849 vcm a_12914_11166# 0.1f
C24850 ctop rowoff_n[8] 0.177f
C24851 a_30074_11166# a_31078_11166# 0.843f
C24852 row_n[2] rowoff_n[1] 0.085f
C24853 VDD a_8990_1126# 0.035f
C24854 col_n[23] a_2275_1150# 0.113f
C24855 col[15] a_17934_17190# 0.0682f
C24856 m2_18224_17438# a_18026_17190# 0.165f
C24857 a_2275_15206# a_13918_15182# 0.136f
C24858 col_n[23] a_26058_11166# 0.251f
C24859 VDD a_32482_11528# 0.0779f
C24860 col_n[20] a_22954_1126# 0.0765f
C24861 ctop a_13006_15182# 4.11f
C24862 row_n[4] a_5978_6146# 0.282f
C24863 col_n[30] a_32994_13174# 0.0765f
C24864 a_2275_3158# a_25358_3174# 0.144f
C24865 a_2475_3158# a_27974_3134# 0.264f
C24866 a_14922_3134# a_15014_3134# 0.326f
C24867 rowon_n[8] a_5886_10162# 0.118f
C24868 rowoff_n[8] a_29070_10162# 0.294f
C24869 col[8] a_2275_9182# 0.0899f
C24870 col_n[3] a_6282_15222# 0.084f
C24871 rowoff_n[11] a_32994_13174# 0.202f
C24872 vcm a_27974_15182# 0.1f
C24873 a_2966_12170# a_3270_12210# 0.0931f
C24874 a_21038_13174# a_21038_12170# 0.843f
C24875 a_3878_12170# a_4370_12532# 0.0658f
C24876 a_2475_12194# a_5978_12170# 0.316f
C24877 VDD a_24050_5142# 0.483f
C24878 m2_6176_18442# VDD 0.0456f
C24879 col_n[14] a_17422_9520# 0.0283f
C24880 row_n[15] a_26362_17230# 0.0117f
C24881 col[28] a_2475_8178# 0.136f
C24882 a_14922_17190# a_15318_17230# 0.0313f
C24883 a_2275_17214# a_28978_17190# 0.136f
C24884 VDD a_13406_14540# 0.0779f
C24885 rowoff_n[14] a_14410_16548# 0.0133f
C24886 a_33086_10162# a_33390_10202# 0.0931f
C24887 a_33998_10162# a_34490_10524# 0.0658f
C24888 m2_9188_15430# a_8990_15182# 0.165f
C24889 vcm a_8898_18194# 0.101f
C24890 a_10998_14178# a_12002_14178# 0.843f
C24891 a_2475_14202# a_21038_14178# 0.316f
C24892 row_n[7] a_26970_9158# 0.0437f
C24893 VDD a_4974_8154# 0.483f
C24894 col[4] a_6890_15182# 0.0682f
C24895 rowon_n[11] a_26058_13174# 0.248f
C24896 VDD a_28466_18556# 0.0858f
C24897 col_n[12] a_15014_9158# 0.251f
C24898 a_2275_2154# a_33998_2130# 0.136f
C24899 m3_20940_18146# VDD 0.0277f
C24900 vcm a_10998_3134# 0.56f
C24901 col[25] a_2275_11190# 0.0899f
C24902 col_n[19] a_21950_11166# 0.0765f
C24903 a_29982_7150# a_30074_7150# 0.326f
C24904 m2_28264_11414# a_28066_11166# 0.165f
C24905 a_2275_11190# a_12002_11166# 0.399f
C24906 m2_18800_18014# a_18938_18194# 0.225f
C24907 col_n[0] a_2966_15182# 0.251f
C24908 row_n[11] a_3970_13174# 0.282f
C24909 a_2475_16210# a_2475_15206# 0.0666f
C24910 VDD a_20034_12170# 0.483f
C24911 col_n[0] ctop 0.0568f
C24912 vcm sw_n 0.0315f
C24913 col_n[10] row_n[4] 0.298f
C24914 col_n[13] rowon_n[5] 0.111f
C24915 col_n[6] row_n[2] 0.298f
C24916 col_n[27] rowon_n[12] 0.111f
C24917 col_n[23] rowon_n[10] 0.111f
C24918 col_n[16] row_n[7] 0.298f
C24919 col_n[14] row_n[6] 0.298f
C24920 col_n[7] rowon_n[2] 0.111f
C24921 VDD en_bit_n[1] 0.206f
C24922 col_n[8] row_n[3] 0.298f
C24923 col_n[9] rowon_n[3] 0.111f
C24924 rowon_n[15] row_n[15] 18.9f
C24925 col_n[2] row_n[0] 0.298f
C24926 col_n[4] row_n[1] 0.298f
C24927 col_n[28] row_n[13] 0.298f
C24928 col_n[5] rowon_n[1] 0.111f
C24929 col_n[25] rowon_n[11] 0.111f
C24930 col_n[24] row_n[11] 0.298f
C24931 col_n[31] rowon_n[14] 0.111f
C24932 col_n[29] rowon_n[13] 0.111f
C24933 col_n[21] rowon_n[9] 0.111f
C24934 col_n[30] row_n[14] 0.298f
C24935 col_n[26] row_n[12] 0.298f
C24936 col_n[3] rowon_n[0] 0.111f
C24937 col_n[22] row_n[10] 0.298f
C24938 col_n[20] row_n[9] 0.298f
C24939 col_n[19] rowon_n[8] 0.111f
C24940 col_n[15] rowon_n[6] 0.111f
C24941 col_n[12] row_n[5] 0.298f
C24942 m2_6752_18014# m3_5880_18146# 0.0341f
C24943 col_n[18] row_n[8] 0.298f
C24944 col_n[11] rowon_n[4] 0.111f
C24945 col_n[17] rowon_n[7] 0.111f
C24946 m2_12200_14426# rowon_n[12] 0.0322f
C24947 col_n[3] a_6378_7512# 0.0283f
C24948 m2_18224_10410# rowon_n[8] 0.0322f
C24949 m2_24248_6394# rowon_n[4] 0.0322f
C24950 a_24962_4138# a_25358_4178# 0.0313f
C24951 row_n[1] a_14010_3134# 0.282f
C24952 vcm a_26058_7150# 0.56f
C24953 rowon_n[5] a_13918_7150# 0.118f
C24954 a_2874_8154# a_3366_8516# 0.0658f
C24955 rowoff_n[12] a_20946_14178# 0.202f
C24956 a_2275_8178# a_3878_8154# 0.136f
C24957 a_2475_8178# a_4882_8154# 0.264f
C24958 col_n[15] a_2475_7174# 0.0531f
C24959 a_14010_13174# a_14314_13214# 0.0931f
C24960 a_14922_13174# a_15414_13536# 0.0658f
C24961 a_2275_13198# a_27062_13174# 0.399f
C24962 row_n[3] a_2275_5166# 19.2f
C24963 rowon_n[7] a_1957_9182# 0.0172f
C24964 row_n[12] a_35398_14218# 0.0117f
C24965 vcm a_16322_1166# 0.16f
C24966 col_n[1] a_3970_7150# 0.251f
C24967 col_n[27] a_30378_8194# 0.084f
C24968 col[0] a_2475_15206# 0.148f
C24969 m2_1732_6970# sample_n 0.0522f
C24970 m2_8760_946# m3_9896_1078# 0.0341f
C24971 m2_19228_9406# a_19030_9158# 0.165f
C24972 col[5] a_2475_4162# 0.136f
C24973 vcm a_6982_10162# 0.56f
C24974 rowoff_n[15] a_1957_17214# 0.0219f
C24975 a_2275_10186# a_17326_10202# 0.144f
C24976 a_2475_10186# a_19942_10162# 0.264f
C24977 a_10906_10162# a_10998_10162# 0.326f
C24978 col_n[8] a_10906_9158# 0.0765f
C24979 row_n[14] a_24962_16186# 0.0437f
C24980 row_n[4] a_35002_6146# 0.0437f
C24981 col_n[19] rowoff_n[12] 0.0471f
C24982 col_n[12] a_2275_10186# 0.113f
C24983 a_12002_3134# a_12002_2130# 0.843f
C24984 rowon_n[8] a_34090_10162# 0.248f
C24985 vcm a_31382_5182# 0.155f
C24986 a_5886_7150# a_6282_7190# 0.0313f
C24987 a_2275_7174# a_10906_7150# 0.136f
C24988 m2_23820_18014# vcm 0.353f
C24989 col_n[2] a_5374_17552# 0.0283f
C24990 vcm a_22042_14178# 0.56f
C24991 col[21] a_24050_6146# 0.367f
C24992 a_2275_12194# a_32386_12210# 0.144f
C24993 a_2475_12194# a_35002_12170# 0.264f
C24994 VDD a_18938_4138# 0.181f
C24995 col[2] a_2275_7174# 0.0899f
C24996 col[28] a_30986_8154# 0.0682f
C24997 a_29982_17190# a_30474_17552# 0.0658f
C24998 a_29070_17190# a_29374_17230# 0.0931f
C24999 row_n[8] a_12002_10162# 0.282f
C25000 rowon_n[12] a_11910_14178# 0.118f
C25001 a_1957_4162# a_2275_4162# 0.158f
C25002 a_2475_4162# a_2874_4138# 0.264f
C25003 m2_33860_946# ctop 0.669f
C25004 m2_10192_7398# a_9994_7150# 0.165f
C25005 col[17] a_2475_17214# 0.136f
C25006 m2_30848_18014# m2_31852_18014# 0.843f
C25007 vcm a_12306_8194# 0.155f
C25008 rowoff_n[13] a_8898_15182# 0.202f
C25009 a_2275_9182# a_25966_9158# 0.136f
C25010 col[22] a_2475_6170# 0.136f
C25011 col_n[16] a_19334_6186# 0.084f
C25012 rowon_n[2] a_21950_4138# 0.118f
C25013 ctop a_25054_3134# 4.11f
C25014 col_n[26] a_29374_18234# 0.084f
C25015 vcm a_2874_17190# 0.1f
C25016 m3_17928_1078# a_18026_1126# 2.77f
C25017 a_25966_14178# a_26058_14178# 0.326f
C25018 VDD a_33998_8154# 0.181f
C25019 rowoff_n[5] a_10906_7150# 0.202f
C25020 col_n[3] rowoff_n[13] 0.0471f
C25021 a_2275_18218# a_3970_18194# 0.0924f
C25022 row_n[0] a_9294_2170# 0.0117f
C25023 m2_29268_3382# a_29070_3134# 0.165f
C25024 col_n[29] a_2275_12194# 0.113f
C25025 col[0] rowoff_n[3] 0.0901f
C25026 col[2] rowoff_n[5] 0.0901f
C25027 col[1] rowoff_n[4] 0.0901f
C25028 col[4] rowoff_n[7] 0.0901f
C25029 col[3] rowoff_n[6] 0.0901f
C25030 col[5] rowoff_n[8] 0.0901f
C25031 col[6] rowoff_n[9] 0.0901f
C25032 vcm a_5886_2130# 0.1f
C25033 a_27062_7150# a_27062_6146# 0.843f
C25034 a_2475_6170# a_18026_6146# 0.316f
C25035 vcm a_27366_12210# 0.155f
C25036 rowoff_n[3] a_19942_5142# 0.202f
C25037 a_20946_11166# a_21342_11206# 0.0313f
C25038 m2_5172_17438# row_n[15] 0.0128f
C25039 VDD a_25454_2492# 0.0779f
C25040 m2_14784_18014# a_15014_17190# 0.843f
C25041 m2_11196_13422# row_n[11] 0.0128f
C25042 m2_17220_9406# row_n[7] 0.0128f
C25043 m2_23244_5390# row_n[3] 0.0128f
C25044 ctop a_5978_6146# 4.11f
C25045 row_n[11] a_32994_13174# 0.0437f
C25046 VDD a_14922_11166# 0.181f
C25047 col[10] a_13006_4138# 0.367f
C25048 col[19] a_2275_9182# 0.0899f
C25049 rowon_n[15] a_32082_17190# 0.248f
C25050 col[20] a_23046_16186# 0.367f
C25051 col[17] a_19942_6146# 0.0682f
C25052 a_4974_3134# a_5278_3174# 0.0931f
C25053 a_2275_3158# a_8990_3134# 0.399f
C25054 a_5886_3134# a_6378_3496# 0.0658f
C25055 rowoff_n[8] a_11398_10524# 0.0133f
C25056 col[27] a_29982_18194# 0.0682f
C25057 rowoff_n[1] a_28978_3134# 0.202f
C25058 vcm a_20946_6146# 0.1f
C25059 a_17022_8154# a_18026_8154# 0.843f
C25060 a_2475_8178# a_33086_8154# 0.316f
C25061 m3_3872_1078# m2_2736_946# 0.0195f
C25062 vcm a_8290_15222# 0.155f
C25063 VDD a_6378_5504# 0.0779f
C25064 col_n[5] a_8290_4178# 0.084f
C25065 ctop a_21038_10162# 4.11f
C25066 row_n[15] a_9994_17190# 0.282f
C25067 col_n[15] a_18330_16226# 0.084f
C25068 a_6890_17190# a_6982_17190# 0.326f
C25069 a_2275_17214# a_9294_17230# 0.144f
C25070 a_2475_17214# a_11910_17190# 0.264f
C25071 rowoff_n[6] a_20434_8516# 0.0133f
C25072 VDD a_29982_15182# 0.181f
C25073 col_n[4] a_2475_16210# 0.0531f
C25074 row_n[5] a_20034_7150# 0.282f
C25075 a_2275_5166# a_24050_5142# 0.399f
C25076 col_n[9] a_2475_5166# 0.0531f
C25077 rowon_n[9] a_19942_11166# 0.118f
C25078 col_n[26] a_29470_10524# 0.0283f
C25079 a_26970_1126# a_27462_1488# 0.0658f
C25080 vcm a_34394_10202# 0.155f
C25081 a_7986_10162# a_7986_9158# 0.843f
C25082 rowoff_n[4] a_29470_6508# 0.0133f
C25083 m2_13780_946# a_2275_1150# 0.28f
C25084 a_2475_14202# a_2966_14178# 0.317f
C25085 a_2161_14202# a_2275_14202# 0.183f
C25086 VDD a_21438_9520# 0.0779f
C25087 row_n[7] a_7286_9198# 0.0117f
C25088 ctop a_2475_13198# 0.0488f
C25089 VDD a_10906_18194# 0.343f
C25090 a_2475_2154# a_16930_2130# 0.264f
C25091 a_2275_2154# a_14314_2170# 0.144f
C25092 col[9] a_12002_14178# 0.367f
C25093 m2_8184_1374# VDD 0.0194f
C25094 col[6] a_8898_4138# 0.0682f
C25095 a_20034_7150# a_20338_7190# 0.0931f
C25096 a_20946_7150# a_21438_7512# 0.0658f
C25097 rowoff_n[9] a_21038_11166# 0.294f
C25098 col[16] a_18938_16186# 0.0682f
C25099 vcm a_16930_13174# 0.1f
C25100 a_32082_12170# a_33086_12170# 0.843f
C25101 col_n[17] row_n[2] 0.298f
C25102 col_n[31] row_n[9] 0.298f
C25103 col_n[20] rowon_n[3] 0.111f
C25104 col_n[10] ctop 0.0594f
C25105 col_n[21] row_n[4] 0.298f
C25106 col_n[16] rowon_n[1] 0.111f
C25107 VDD col[7] 3.83f
C25108 col_n[13] row_n[0] 0.298f
C25109 col_n[14] rowon_n[0] 0.111f
C25110 col_n[18] rowon_n[2] 0.111f
C25111 col_n[23] row_n[5] 0.298f
C25112 col_n[22] rowon_n[4] 0.111f
C25113 col_n[25] row_n[6] 0.298f
C25114 col_n[26] rowon_n[6] 0.111f
C25115 col_n[2] col[2] 0.489f
C25116 col_n[29] row_n[8] 0.298f
C25117 vcm col[4] 5.46f
C25118 VDD a_13006_3134# 0.483f
C25119 col_n[28] rowon_n[7] 0.111f
C25120 col_n[27] row_n[7] 0.298f
C25121 col_n[19] row_n[3] 0.298f
C25122 col_n[15] row_n[1] 0.298f
C25123 col_n[24] rowon_n[5] 0.111f
C25124 col_n[30] rowon_n[8] 0.111f
C25125 col_n[24] a_27062_10162# 0.251f
C25126 m2_14784_18014# a_2275_18218# 0.28f
C25127 col_n[6] a_2275_8178# 0.113f
C25128 a_2275_16210# a_17934_16186# 0.136f
C25129 rowon_n[3] a_6982_5142# 0.248f
C25130 VDD a_1957_12194# 0.196f
C25131 col_n[31] a_33998_12170# 0.0765f
C25132 a_26058_1126# m2_25828_946# 0.0249f
C25133 ctop a_17022_17190# 4.06f
C25134 rowoff_n[7] a_30074_9158# 0.294f
C25135 col_n[4] a_7286_14218# 0.084f
C25136 a_2475_4162# a_31990_4138# 0.264f
C25137 a_16930_4138# a_17022_4138# 0.326f
C25138 a_2275_4162# a_29374_4178# 0.144f
C25139 col[0] a_2966_12170# 0.367f
C25140 col_n[26] a_2475_7174# 0.0531f
C25141 rowoff_n[12] a_2275_14202# 0.151f
C25142 vcm a_31990_17190# 0.1f
C25143 a_2475_13198# a_9994_13174# 0.316f
C25144 a_23046_14178# a_23046_13174# 0.843f
C25145 col_n[15] a_18426_8516# 0.0283f
C25146 VDD a_28066_7150# 0.483f
C25147 m2_10768_18014# a_2475_18218# 0.286f
C25148 a_2275_18218# a_32994_18194# 0.136f
C25149 a_16930_18194# a_17326_18234# 0.0313f
C25150 VDD a_17422_16548# 0.0779f
C25151 col[11] a_2475_15206# 0.136f
C25152 a_11910_1126# a_12306_1166# 0.0313f
C25153 a_2275_1150# a_22954_1126# 0.136f
C25154 row_n[12] a_18026_14178# 0.282f
C25155 col[16] a_2475_4162# 0.136f
C25156 vcm a_34090_2130# 0.56f
C25157 m2_23820_946# m2_24248_1374# 0.165f
C25158 col_n[0] a_2874_4138# 0.0765f
C25159 row_n[2] a_28066_4138# 0.282f
C25160 row_n[14] a_5278_16226# 0.0117f
C25161 rowon_n[6] a_27974_8154# 0.118f
C25162 m2_33860_18014# a_34090_17190# 0.843f
C25163 m2_1732_3958# VDD 0.856f
C25164 col[5] a_7894_14178# 0.0682f
C25165 a_2475_15206# a_25054_15182# 0.316f
C25166 a_13006_15182# a_14010_15182# 0.843f
C25167 col_n[30] rowoff_n[12] 0.0471f
C25168 col_n[23] a_2275_10186# 0.113f
C25169 VDD a_8990_10162# 0.483f
C25170 col_n[13] a_16018_8154# 0.251f
C25171 row_n[4] a_15318_6186# 0.0117f
C25172 col_n[20] a_22954_10162# 0.0765f
C25173 a_2475_18218# a_30986_18194# 0.264f
C25174 vcm a_15014_5142# 0.56f
C25175 a_31990_8154# a_32082_8154# 0.326f
C25176 rowoff_n[10] a_8990_12170# 0.294f
C25177 a_28978_1126# vcm 0.0989f
C25178 col[8] a_2275_18218# 0.0899f
C25179 m2_1732_11990# rowon_n[10] 0.236f
C25180 row_n[6] a_5886_8154# 0.0437f
C25181 col[13] a_2275_7174# 0.0899f
C25182 m2_7180_8402# rowon_n[6] 0.0322f
C25183 a_2275_12194# a_16018_12170# 0.399f
C25184 m2_13204_4386# rowon_n[2] 0.0322f
C25185 rowon_n[10] a_4974_12170# 0.248f
C25186 m2_27836_18014# VDD 1.06f
C25187 a_3970_17190# a_3970_16186# 0.843f
C25188 col_n[4] a_7382_6508# 0.0283f
C25189 VDD a_24050_14178# 0.483f
C25190 col_n[14] a_17422_18556# 0.0283f
C25191 rowon_n[0] a_15014_2130# 0.248f
C25192 col[28] a_2475_17214# 0.136f
C25193 a_26970_5142# a_27366_5182# 0.0313f
C25194 vcm a_30074_9158# 0.56f
C25195 a_2275_9182# a_6282_9198# 0.144f
C25196 a_2475_9182# a_8898_9158# 0.264f
C25197 rowoff_n[14] a_25054_16186# 0.294f
C25198 rowon_n[2] a_3878_4138# 0.118f
C25199 col_n[14] rowoff_n[13] 0.0471f
C25200 m3_2868_1078# a_3970_1126# 0.0379f
C25201 m2_22240_17438# rowon_n[15] 0.0322f
C25202 a_16018_14178# a_16322_14218# 0.0931f
C25203 a_2275_14202# a_31078_14178# 0.399f
C25204 m3_30980_1078# a_31078_2130# 0.0302f
C25205 a_16930_14178# a_17422_14540# 0.0658f
C25206 m2_28264_13422# rowon_n[11] 0.0322f
C25207 m2_34288_9406# rowon_n[7] 0.0322f
C25208 col_n[3] a_2475_3158# 0.0531f
C25209 col[11] rowoff_n[3] 0.0901f
C25210 col[13] rowoff_n[5] 0.0901f
C25211 col[17] rowoff_n[9] 0.0901f
C25212 col[12] rowoff_n[4] 0.0901f
C25213 col[10] rowoff_n[2] 0.0901f
C25214 col[9] rowoff_n[1] 0.0901f
C25215 col[8] rowoff_n[0] 0.0901f
C25216 col[15] rowoff_n[7] 0.0901f
C25217 col[16] rowoff_n[8] 0.0901f
C25218 col[14] rowoff_n[6] 0.0901f
C25219 VDD a_4974_17190# 0.484f
C25220 a_23046_2130# a_24050_2130# 0.843f
C25221 col_n[2] a_4974_6146# 0.251f
C25222 col_n[28] a_31382_7190# 0.084f
C25223 vcm a_20338_3174# 0.155f
C25224 row_n[9] a_26058_11166# 0.282f
C25225 a_35002_7150# a_35398_7190# 0.0313f
C25226 col_n[9] a_11910_8154# 0.0765f
C25227 m2_1732_9982# a_2161_10186# 0.0454f
C25228 rowon_n[13] a_25966_15182# 0.118f
C25229 vcm a_10998_12170# 0.56f
C25230 a_12914_11166# a_13006_11166# 0.326f
C25231 a_2275_11190# a_21342_11206# 0.144f
C25232 a_2475_11190# a_23958_11166# 0.264f
C25233 VDD a_7894_2130# 0.181f
C25234 m2_2736_18014# a_2966_17190# 0.843f
C25235 col[30] a_2275_9182# 0.0899f
C25236 row_n[11] a_13310_13214# 0.0117f
C25237 m2_20808_18014# m3_20940_18146# 3.79f
C25238 a_14010_4138# a_14010_3134# 0.843f
C25239 row_n[1] a_23350_3174# 0.0117f
C25240 col_n[3] a_6378_16548# 0.0283f
C25241 vcm a_2275_6170# 6.49f
C25242 a_7894_8154# a_8290_8194# 0.0313f
C25243 rowoff_n[12] a_31478_14540# 0.0133f
C25244 a_2275_8178# a_14922_8154# 0.136f
C25245 col[22] a_25054_5142# 0.367f
C25246 m2_34864_12994# a_2475_13198# 0.282f
C25247 sample rowoff_n[14] 0.0775f
C25248 vcm a_26058_16186# 0.56f
C25249 a_2966_13174# a_2966_12170# 0.843f
C25250 col[29] a_31990_7150# 0.0682f
C25251 VDD a_22954_6146# 0.181f
C25252 row_n[3] a_13918_5142# 0.0437f
C25253 m2_12776_946# col_n[10] 0.331f
C25254 col[1] rowoff_n[10] 0.0901f
C25255 ctop a_2966_10162# 4.06f
C25256 col_n[15] a_2475_16210# 0.0531f
C25257 a_31990_18194# a_32482_18556# 0.0658f
C25258 rowon_n[7] a_13006_9158# 0.248f
C25259 rowoff_n[6] a_2161_8178# 0.0226f
C25260 col_n[20] a_2475_5166# 0.0531f
C25261 a_3970_5142# a_4974_5142# 0.843f
C25262 a_2475_5166# a_6982_5142# 0.316f
C25263 row_n[5] a_1957_7174# 0.187f
C25264 m2_24824_946# m3_23952_1078# 0.0341f
C25265 col_n[17] a_20338_5182# 0.084f
C25266 vcm a_16322_10202# 0.155f
C25267 col_n[27] a_30378_17230# 0.084f
C25268 a_2275_10186# a_29982_10162# 0.136f
C25269 col_n[1] a_3970_16186# 0.251f
C25270 rowoff_n[15] a_13006_17190# 0.294f
C25271 m2_15212_16434# a_15014_16186# 0.165f
C25272 col[5] a_2475_13198# 0.136f
C25273 rowoff_n[4] a_11910_6146# 0.202f
C25274 ctop a_29070_5142# 4.11f
C25275 a_27974_15182# a_28066_15182# 0.326f
C25276 col_n[8] a_10906_18194# 0.0762f
C25277 VDD a_3366_9520# 0.0779f
C25278 col[10] a_2475_2154# 0.136f
C25279 m2_5748_18014# col_n[3] 0.243f
C25280 m2_6176_7398# row_n[5] 0.0128f
C25281 m2_12200_3382# row_n[1] 0.0128f
C25282 vcm a_9902_4138# 0.1f
C25283 rowoff_n[2] a_20946_4138# 0.202f
C25284 col_n[21] ctop 0.0594f
C25285 rowoff_n[9] a_2966_11166# 0.294f
C25286 col_n[17] en_bit_n[0] 0.186f
C25287 col_n[25] rowon_n[0] 0.111f
C25288 col_n[26] row_n[1] 0.298f
C25289 vcm col[15] 5.46f
C25290 col_n[31] rowon_n[3] 0.111f
C25291 col_n[27] rowon_n[1] 0.111f
C25292 col_n[7] col[8] 7.13f
C25293 col_n[28] row_n[2] 0.298f
C25294 a_29070_8154# a_29070_7150# 0.843f
C25295 col_n[30] row_n[3] 0.298f
C25296 VDD col[18] 3.83f
C25297 col_n[29] rowon_n[2] 0.111f
C25298 a_2475_7174# a_22042_7150# 0.316f
C25299 col_n[24] row_n[0] 0.298f
C25300 col_n[17] a_2275_8178# 0.113f
C25301 m2_34288_12418# a_34090_12170# 0.165f
C25302 row_n[6] a_34090_8154# 0.282f
C25303 vcm a_31382_14218# 0.155f
C25304 a_22954_12170# a_23350_12210# 0.0313f
C25305 VDD a_29470_4500# 0.0779f
C25306 rowon_n[10] a_33998_12170# 0.118f
C25307 col[11] a_14010_3134# 0.367f
C25308 ctop a_9994_8154# 4.11f
C25309 col[21] a_24050_15182# 0.367f
C25310 VDD a_18938_13174# 0.181f
C25311 col[18] a_20946_5142# 0.0682f
C25312 row_n[8] a_21342_10202# 0.0117f
C25313 rowoff_n[0] a_29982_2130# 0.202f
C25314 rowoff_n[7] a_12402_9520# 0.0133f
C25315 col[28] a_30986_17190# 0.0682f
C25316 col[2] a_2275_16210# 0.0899f
C25317 col[7] a_2275_5166# 0.0899f
C25318 a_2275_4162# a_13006_4138# 0.399f
C25319 a_6982_4138# a_7286_4178# 0.0931f
C25320 a_7894_4138# a_8386_4500# 0.0658f
C25321 m3_34996_15134# ctop 0.209f
C25322 m2_21236_16434# row_n[14] 0.0128f
C25323 vcm a_24962_8154# 0.1f
C25324 m2_27260_12418# row_n[10] 0.0128f
C25325 m2_33284_8402# row_n[6] 0.0128f
C25326 rowoff_n[13] a_19430_15544# 0.0133f
C25327 a_19030_9158# a_20034_9158# 0.843f
C25328 m2_6176_14426# a_5978_14178# 0.165f
C25329 row_n[10] a_11910_12170# 0.0437f
C25330 col_n[6] a_9294_3174# 0.084f
C25331 vcm a_12306_17230# 0.155f
C25332 rowon_n[14] a_10998_16186# 0.248f
C25333 VDD a_10394_7512# 0.0779f
C25334 col_n[16] a_19334_15222# 0.084f
C25335 col[22] a_2475_15206# 0.136f
C25336 rowoff_n[5] a_21438_7512# 0.0133f
C25337 col[27] a_2475_4162# 0.136f
C25338 ctop a_25054_12170# 4.11f
C25339 a_2275_18218# a_13310_18234# 0.145f
C25340 a_8898_18194# a_8990_18194# 0.0991f
C25341 VDD a_33998_17190# 0.181f
C25342 row_n[0] a_21950_2130# 0.0437f
C25343 a_2475_1150# a_5886_1126# 0.264f
C25344 a_2275_1150# a_3270_1166# 0.145f
C25345 rowon_n[4] a_21038_6146# 0.248f
C25346 m2_2736_1950# a_2966_2130# 0.0249f
C25347 a_2275_6170# a_28066_6146# 0.399f
C25348 col_n[27] a_30474_9520# 0.0283f
C25349 m2_25252_10410# a_25054_10162# 0.165f
C25350 rowoff_n[3] a_30474_5504# 0.0133f
C25351 vcm a_5886_11166# 0.1f
C25352 a_9994_11166# a_9994_10162# 0.843f
C25353 VDD a_2475_1150# 30.4f
C25354 a_2275_15206# a_6890_15182# 0.136f
C25355 VDD a_25454_11528# 0.0779f
C25356 col[0] a_2874_1126# 0.0682f
C25357 ctop a_5978_15182# 4.11f
C25358 col[10] a_13006_13174# 0.367f
C25359 col[7] a_9902_3134# 0.0682f
C25360 a_2475_3158# a_20946_3134# 0.264f
C25361 a_2275_3158# a_18330_3174# 0.144f
C25362 col[19] a_2275_18218# 0.0899f
C25363 rowoff_n[8] a_22042_10162# 0.294f
C25364 a_35094_1126# a_2475_1150# 0.0299f
C25365 col[17] a_19942_15182# 0.0682f
C25366 row_n[13] a_32082_15182# 0.282f
C25367 col[24] a_2275_7174# 0.0899f
C25368 m2_1732_12994# m2_1732_11990# 0.843f
C25369 a_22042_8154# a_22346_8194# 0.0931f
C25370 a_22954_8154# a_23446_8516# 0.0658f
C25371 rowoff_n[11] a_25966_13174# 0.202f
C25372 col_n[25] a_28066_9158# 0.251f
C25373 vcm a_20946_15182# 0.1f
C25374 a_33998_13174# a_34394_13214# 0.0313f
C25375 VDD a_17022_5142# 0.483f
C25376 a_30986_1126# VDD 0.405f
C25377 row_n[15] a_19334_17230# 0.0117f
C25378 a_2275_17214# a_21950_17190# 0.136f
C25379 rowoff_n[6] a_31078_8154# 0.294f
C25380 VDD a_6378_14540# 0.0779f
C25381 col_n[5] a_8290_13214# 0.084f
C25382 a_2275_5166# a_33390_5182# 0.144f
C25383 row_n[5] a_29374_7190# 0.0117f
C25384 a_18938_5142# a_19030_5142# 0.326f
C25385 m2_16216_8402# a_16018_8154# 0.165f
C25386 m3_24956_1078# m3_25960_1078# 0.202f
C25387 col_n[25] rowoff_n[13] 0.0471f
C25388 rowoff_n[14] a_7382_16548# 0.0133f
C25389 col_n[9] a_2475_14202# 0.0531f
C25390 col_n[16] a_19430_7512# 0.0283f
C25391 col_n[14] a_2475_3158# 0.0531f
C25392 col[19] rowoff_n[0] 0.0901f
C25393 col[24] rowoff_n[5] 0.0901f
C25394 col[28] rowoff_n[9] 0.0901f
C25395 m2_13780_946# a_13918_1126# 0.225f
C25396 col[22] rowoff_n[3] 0.0901f
C25397 col[20] rowoff_n[1] 0.0901f
C25398 col[21] rowoff_n[2] 0.0901f
C25399 col[23] rowoff_n[4] 0.0901f
C25400 col[25] rowoff_n[6] 0.0901f
C25401 col[27] rowoff_n[8] 0.0901f
C25402 col[26] rowoff_n[7] 0.0901f
C25403 a_2475_14202# a_14010_14178# 0.316f
C25404 a_25054_15182# a_25054_14178# 0.843f
C25405 VDD a_32082_9158# 0.483f
C25406 row_n[7] a_19942_9158# 0.0437f
C25407 rowon_n[11] a_19030_13174# 0.248f
C25408 col[5] a_2475_18218# 0.136f
C25409 VDD a_21438_18556# 0.0858f
C25410 a_2275_2154# a_26970_2130# 0.136f
C25411 a_13918_2130# a_14314_2170# 0.0313f
C25412 m2_34864_3958# a_35094_4138# 0.0249f
C25413 m2_31276_1374# VDD 0.0194f
C25414 vcm a_3970_3134# 0.56f
C25415 rowon_n[1] a_29070_3134# 0.248f
C25416 col[6] a_8898_13174# 0.0682f
C25417 a_2275_11190# a_4974_11166# 0.399f
C25418 a_3878_11166# a_3970_11166# 0.326f
C25419 a_2874_11166# a_3270_11206# 0.0313f
C25420 m2_13780_18014# a_14010_18194# 0.0249f
C25421 col_n[14] a_17022_7150# 0.251f
C25422 a_2475_16210# a_29070_16186# 0.316f
C25423 a_15014_16186# a_16018_16186# 0.843f
C25424 VDD a_13006_12170# 0.483f
C25425 a_32386_1166# m2_31852_946# 0.087f
C25426 col_n[6] a_2275_17214# 0.113f
C25427 col_n[21] a_23958_9158# 0.0765f
C25428 m2_1732_10986# col[0] 0.0137f
C25429 col_n[11] a_2275_6170# 0.113f
C25430 m2_2160_2378# rowon_n[0] 0.0219f
C25431 col_n[9] rowoff_n[14] 0.0471f
C25432 row_n[1] a_6982_3134# 0.282f
C25433 m2_7180_6394# a_6982_6146# 0.165f
C25434 vcm a_19030_7150# 0.56f
C25435 rowon_n[5] a_6890_7150# 0.118f
C25436 a_33998_9158# a_34090_9158# 0.326f
C25437 rowoff_n[12] a_13918_14178# 0.202f
C25438 col[12] rowoff_n[10] 0.0901f
C25439 col_n[26] a_2475_16210# 0.0531f
C25440 a_2275_13198# a_20034_13174# 0.399f
C25441 col_n[31] a_2475_5166# 0.0531f
C25442 col_n[5] a_8386_5504# 0.0283f
C25443 col[1] a_2275_3158# 0.0899f
C25444 col_n[15] a_18426_17552# 0.0283f
C25445 VDD a_28066_16186# 0.483f
C25446 row_n[12] a_27366_14218# 0.0117f
C25447 m2_11196_15430# rowon_n[13] 0.0322f
C25448 vcm a_9294_1166# 0.16f
C25449 a_28978_6146# a_29374_6186# 0.0313f
C25450 m2_17220_11414# rowon_n[9] 0.0322f
C25451 m2_1732_4962# vcm 0.316f
C25452 m2_23244_7398# rowon_n[5] 0.0322f
C25453 col[16] a_2475_13198# 0.136f
C25454 m2_29268_3382# rowon_n[1] 0.0322f
C25455 vcm a_34090_11166# 0.56f
C25456 col[21] a_2475_2154# 0.136f
C25457 a_2475_10186# a_12914_10162# 0.264f
C25458 a_2275_10186# a_10298_10202# 0.144f
C25459 row_n[14] a_17934_16186# 0.0437f
C25460 col_n[0] a_2874_13174# 0.0765f
C25461 a_2275_15206# a_35094_15182# 0.0924f
C25462 a_18026_15182# a_18330_15222# 0.0931f
C25463 a_18938_15182# a_19430_15544# 0.0658f
C25464 col_n[3] a_5978_5142# 0.251f
C25465 row_n[4] a_27974_6146# 0.0437f
C25466 m3_1864_12122# a_2966_12170# 0.0302f
C25467 col_n[29] a_32386_6186# 0.084f
C25468 rowon_n[15] ctop 0.203f
C25469 col_n[13] col[13] 0.489f
C25470 rowon_n[7] rowon_n[6] 0.0632f
C25471 VDD col[29] 3.83f
C25472 vcm col[26] 5.46f
C25473 col_n[13] a_16018_17190# 0.251f
C25474 a_25054_3134# a_26058_3134# 0.843f
C25475 rowon_n[8] a_27062_10162# 0.248f
C25476 col_n[28] a_2275_8178# 0.113f
C25477 col_n[10] a_12914_7150# 0.0765f
C25478 vcm a_24354_5182# 0.155f
C25479 a_2874_7150# a_2966_7150# 0.326f
C25480 rowoff_n[2] a_2275_4162# 0.151f
C25481 m2_9764_18014# vcm 0.353f
C25482 vcm a_15014_14178# 0.56f
C25483 a_2275_12194# a_25358_12210# 0.144f
C25484 a_2475_12194# a_27974_12170# 0.264f
C25485 a_14922_12170# a_15014_12170# 0.326f
C25486 VDD a_11910_4138# 0.181f
C25487 col[13] a_2275_16210# 0.0899f
C25488 col[18] a_2275_5166# 0.0899f
C25489 row_n[8] a_4974_10162# 0.282f
C25490 col_n[4] a_7382_15544# 0.0283f
C25491 rowon_n[12] a_4882_14178# 0.118f
C25492 col_n[1] a_3878_5142# 0.0765f
C25493 a_16018_5142# a_16018_4138# 0.843f
C25494 col[23] a_26058_4138# 0.367f
C25495 m2_23820_18014# m2_24824_18014# 0.843f
C25496 vcm a_5278_8194# 0.155f
C25497 a_9902_9158# a_10298_9198# 0.0313f
C25498 a_2275_9182# a_18938_9158# 0.136f
C25499 col[30] a_32994_6146# 0.0682f
C25500 rowon_n[2] a_14922_4138# 0.118f
C25501 ctop a_18026_3134# 4.11f
C25502 vcm a_30074_18194# 0.165f
C25503 VDD a_26970_8154# 0.181f
C25504 rowoff_n[5] a_3366_7512# 0.0133f
C25505 row_n[0] a_3878_2130# 0.0437f
C25506 a_28978_2130# a_29470_2492# 0.0658f
C25507 a_28066_2130# a_28370_2170# 0.0931f
C25508 rowon_n[4] a_2966_6146# 0.248f
C25509 col_n[3] a_2475_12194# 0.0531f
C25510 col_n[18] a_21342_4178# 0.084f
C25511 vcm a_32994_3134# 0.1f
C25512 col_n[8] a_2475_1150# 0.0531f
C25513 a_2475_6170# a_10998_6146# 0.316f
C25514 a_5978_6146# a_6982_6146# 0.843f
C25515 col_n[2] a_4974_15182# 0.251f
C25516 col_n[28] a_31382_16226# 0.084f
C25517 vcm a_20338_12210# 0.155f
C25518 rowoff_n[3] a_12914_5142# 0.202f
C25519 a_2275_11190# a_33998_11166# 0.136f
C25520 VDD a_18426_2492# 0.0779f
C25521 col_n[9] a_11910_17190# 0.0765f
C25522 m2_32856_18014# a_33086_18194# 0.0249f
C25523 ctop a_33086_7150# 4.11f
C25524 row_n[11] a_25966_13174# 0.0437f
C25525 a_29982_16186# a_30074_16186# 0.326f
C25526 VDD a_7894_11166# 0.181f
C25527 col[30] a_2275_18218# 0.0899f
C25528 rowon_n[15] a_25054_17190# 0.248f
C25529 a_1957_3158# a_2161_3158# 0.115f
C25530 a_2475_3158# a_2275_3158# 2.76f
C25531 rowoff_n[8] a_4370_10524# 0.0133f
C25532 row_n[1] a_34394_3174# 0.0117f
C25533 rowoff_n[1] a_21950_3134# 0.202f
C25534 rowon_n[5] a_35094_7150# 0.0141f
C25535 vcm a_13918_6146# 0.1f
C25536 a_31078_9158# a_31078_8154# 0.843f
C25537 a_2475_8178# a_26058_8154# 0.316f
C25538 col[12] a_15014_2130# 0.367f
C25539 vcm a_2275_15206# 6.49f
C25540 a_24962_13174# a_25358_13214# 0.0313f
C25541 VDD a_33486_6508# 0.0779f
C25542 col[22] a_25054_14178# 0.367f
C25543 col_n[5] a_2275_4162# 0.113f
C25544 col[19] a_21950_4138# 0.0682f
C25545 ctop a_14010_10162# 4.11f
C25546 row_n[15] a_2874_17190# 0.0436f
C25547 a_2874_17190# a_3366_17552# 0.0658f
C25548 m2_10192_14426# row_n[12] 0.0128f
C25549 a_2475_17214# a_4882_17190# 0.264f
C25550 a_2275_17214# a_3878_17190# 0.136f
C25551 col[29] a_31990_16186# 0.0682f
C25552 rowoff_n[6] a_13406_8516# 0.0133f
C25553 m2_16216_10410# row_n[8] 0.0128f
C25554 VDD a_22954_15182# 0.181f
C25555 m2_22240_6394# row_n[4] 0.0128f
C25556 rowon_n[13] rowoff_n[13] 20.2f
C25557 m3_13912_18146# a_14010_17190# 0.0303f
C25558 row_n[5] a_13006_7150# 0.282f
C25559 a_9902_5142# a_10394_5504# 0.0658f
C25560 a_8990_5142# a_9294_5182# 0.0931f
C25561 a_2275_5166# a_17022_5142# 0.399f
C25562 col_n[20] a_2475_14202# 0.0531f
C25563 m2_1732_7974# a_2475_8178# 0.139f
C25564 m3_1864_7102# m3_1864_6098# 0.202f
C25565 rowon_n[9] a_12914_11166# 0.118f
C25566 col_n[25] a_2475_3158# 0.0531f
C25567 col[31] rowoff_n[1] 0.0901f
C25568 col[30] rowoff_n[0] 0.0901f
C25569 sample_n rowoff_n[2] 0.14f
C25570 vcm a_28978_10162# 0.1f
C25571 col_n[7] a_10298_2170# 0.084f
C25572 en_C0_n a_2275_1150# 0.0363f
C25573 a_21038_10162# a_22042_10162# 0.843f
C25574 col_n[17] a_20338_14218# 0.084f
C25575 rowoff_n[4] a_22442_6508# 0.0133f
C25576 col[16] a_2475_18218# 0.136f
C25577 m2_24824_946# a_25054_2130# 0.843f
C25578 VDD a_14410_9520# 0.0779f
C25579 ctop a_29070_14178# 4.11f
C25580 col[10] a_2475_11190# 0.136f
C25581 VDD a_3366_18556# 0.0858f
C25582 a_5886_2130# a_5978_2130# 0.326f
C25583 a_2475_2154# a_9902_2130# 0.264f
C25584 a_2275_2154# a_7286_2170# 0.144f
C25585 col_n[28] a_31478_8516# 0.0283f
C25586 rowoff_n[2] a_31478_4500# 0.0133f
C25587 a_2275_7174# a_32082_7150# 0.399f
C25588 rowoff_n[9] a_14010_11166# 0.294f
C25589 vcm a_9902_13174# 0.1f
C25590 a_12002_12170# a_12002_11166# 0.843f
C25591 m2_22816_946# col_n[20] 0.331f
C25592 VDD a_5978_3134# 0.483f
C25593 col_n[17] a_2275_17214# 0.113f
C25594 m2_1732_18014# a_1957_18218# 0.245f
C25595 col_n[22] a_2275_6170# 0.113f
C25596 a_5886_16186# a_6282_16226# 0.0313f
C25597 a_2275_16210# a_10906_16186# 0.136f
C25598 VDD a_29470_13536# 0.0779f
C25599 col[11] a_14010_12170# 0.367f
C25600 col_n[20] rowoff_n[14] 0.0471f
C25601 row_n[8] a_33998_10162# 0.0437f
C25602 m2_20808_18014# col[18] 0.347f
C25603 col[8] a_10906_2130# 0.0682f
C25604 ctop a_9994_17190# 4.06f
C25605 rowoff_n[7] a_23046_9158# 0.294f
C25606 rowon_n[12] a_33086_14178# 0.248f
C25607 col[18] a_20946_14178# 0.0682f
C25608 a_2475_4162# a_24962_4138# 0.264f
C25609 a_2275_4162# a_22346_4178# 0.144f
C25610 m3_16924_1078# ctop 0.21f
C25611 col[23] rowoff_n[10] 0.0901f
C25612 col_n[26] a_29070_8154# 0.251f
C25613 a_24962_9158# a_25454_9520# 0.0658f
C25614 col[7] a_2275_14202# 0.0899f
C25615 rowoff_n[13] a_30074_15182# 0.294f
C25616 a_24050_9158# a_24354_9198# 0.0931f
C25617 col[12] a_2275_3158# 0.0899f
C25618 vcm a_24962_17190# 0.1f
C25619 a_1957_13198# a_2275_13198# 0.158f
C25620 a_2475_13198# a_2874_13174# 0.264f
C25621 VDD a_21038_7150# 0.483f
C25622 rowoff_n[5] a_32082_7150# 0.294f
C25623 col_n[6] a_9294_12210# 0.084f
C25624 a_2275_18218# a_25966_18194# 0.136f
C25625 VDD a_10394_16548# 0.0779f
C25626 row_n[12] a_10998_14178# 0.282f
C25627 a_2275_1150# a_15926_1126# 0.136f
C25628 col[27] a_2475_13198# 0.136f
C25629 vcm a_27062_2130# 0.56f
C25630 a_20946_6146# a_21038_6146# 0.326f
C25631 col_n[17] a_20434_6508# 0.0283f
C25632 row_n[2] a_21038_4138# 0.282f
C25633 col_n[27] a_30474_18556# 0.0283f
C25634 VDD a_11302_1166# 0.0149f
C25635 m2_21236_17438# a_21038_17190# 0.165f
C25636 rowon_n[6] a_20946_8154# 0.118f
C25637 a_27062_16186# a_27062_15182# 0.843f
C25638 a_2475_15206# a_18026_15182# 0.316f
C25639 row_n[15] col[4] 0.0342f
C25640 col_n[4] rowoff_n[15] 0.0471f
C25641 row_n[13] col[0] 0.0322f
C25642 VDD a_2475_10186# 26.1f
C25643 rowon_n[14] col[3] 0.0323f
C25644 col_n[18] col[19] 7.13f
C25645 rowon_n[4] row_n[4] 18.9f
C25646 rowon_n[15] col[5] 0.0323f
C25647 row_n[14] col[2] 0.0342f
C25648 rowon_n[13] col[1] 0.0323f
C25649 row_n[10] ctop 0.186f
C25650 m2_1732_13998# m3_1864_15134# 0.0341f
C25651 rowon_n[0] m2_34288_2378# 0.0322f
C25652 row_n[4] a_8290_6186# 0.0117f
C25653 a_2275_3158# a_30986_3134# 0.136f
C25654 col[7] rowoff_n[11] 0.0901f
C25655 a_15926_3134# a_16322_3174# 0.0313f
C25656 col[0] a_2874_10162# 0.0682f
C25657 a_2475_18218# a_23958_18194# 0.264f
C25658 vcm a_7986_5142# 0.56f
C25659 rowoff_n[10] a_2475_12194# 3.9f
C25660 col[7] a_9902_12170# 0.0682f
C25661 col[24] a_2275_16210# 0.0899f
C25662 a_2275_12194# a_8990_12170# 0.399f
C25663 a_5886_12170# a_6378_12532# 0.0658f
C25664 m2_1732_5966# rowoff_n[4] 0.415f
C25665 a_4974_12170# a_5278_12210# 0.0931f
C25666 col_n[15] a_18026_6146# 0.251f
C25667 col[29] a_2275_5166# 0.0899f
C25668 m2_13780_18014# VDD 1f
C25669 row_n[15] a_31990_17190# 0.0437f
C25670 col_n[22] a_24962_8154# 0.0765f
C25671 a_17022_17190# a_18026_17190# 0.843f
C25672 a_2475_17214# a_33086_17190# 0.316f
C25673 VDD a_17022_14178# 0.483f
C25674 rowon_n[0] a_7986_2130# 0.248f
C25675 col_n[0] a_2275_2154# 0.113f
C25676 vcm a_23046_9158# 0.56f
C25677 rowoff_n[14] a_18026_16186# 0.294f
C25678 m2_12200_15430# a_12002_15182# 0.165f
C25679 col_n[6] a_9390_4500# 0.0283f
C25680 a_2275_14202# a_24050_14178# 0.399f
C25681 col_n[16] a_19430_16548# 0.0283f
C25682 m2_6176_9406# rowon_n[7] 0.0322f
C25683 m2_12200_5390# rowon_n[3] 0.0322f
C25684 col_n[14] a_2475_12194# 0.0531f
C25685 m2_11772_946# vcm 0.353f
C25686 VDD a_32082_18194# 0.0356f
C25687 col_n[19] a_2475_1150# 0.0531f
C25688 m2_34864_2954# a_2275_3158# 0.278f
C25689 vcm a_13310_3174# 0.155f
C25690 row_n[9] a_19030_11166# 0.282f
C25691 a_30986_7150# a_31382_7190# 0.0313f
C25692 rowon_n[13] a_18938_15182# 0.118f
C25693 m2_31276_11414# a_31078_11166# 0.165f
C25694 vcm a_3970_12170# 0.56f
C25695 a_2275_11190# a_14314_11206# 0.144f
C25696 a_2475_11190# a_16930_11166# 0.264f
C25697 VDD a_35002_3134# 0.258f
C25698 m2_19804_18014# a_20338_18234# 0.087f
C25699 col[4] a_2475_9182# 0.136f
C25700 row_n[11] a_6282_13214# 0.0117f
C25701 a_20034_16186# a_20338_16226# 0.0931f
C25702 a_20946_16186# a_21438_16548# 0.0658f
C25703 col_n[30] a_33390_5182# 0.084f
C25704 rowon_n[3] a_28978_5142# 0.118f
C25705 col_n[4] a_6982_4138# 0.251f
C25706 m2_11772_18014# m3_10900_18146# 0.0341f
C25707 col_n[14] a_17022_16186# 0.251f
C25708 m2_27260_14426# rowon_n[12] 0.0322f
C25709 m2_33284_10410# rowon_n[8] 0.0322f
C25710 col_n[11] a_13918_6146# 0.0765f
C25711 a_27062_4138# a_28066_4138# 0.843f
C25712 col_n[21] a_23958_18194# 0.0762f
C25713 rowoff_n[1] a_3878_3134# 0.202f
C25714 row_n[1] a_16322_3174# 0.0117f
C25715 col_n[11] a_2275_15206# 0.113f
C25716 vcm a_28370_7190# 0.155f
C25717 rowoff_n[12] a_24450_14540# 0.0133f
C25718 a_2275_8178# a_7894_8154# 0.136f
C25719 col_n[16] a_2275_4162# 0.113f
C25720 vcm a_19030_16186# 0.56f
C25721 a_16930_13174# a_17022_13174# 0.326f
C25722 a_2475_13198# a_31990_13174# 0.264f
C25723 a_2275_13198# a_29374_13214# 0.144f
C25724 VDD a_15926_6146# 0.181f
C25725 row_n[3] a_6890_5142# 0.0437f
C25726 rowon_n[7] a_5978_9158# 0.248f
C25727 col_n[31] a_2475_14202# 0.0531f
C25728 col_n[5] a_8386_14540# 0.0283f
C25729 col[1] a_2275_12194# 0.0899f
C25730 col[24] a_27062_3134# 0.367f
C25731 col[6] a_2275_1150# 0.0899f
C25732 vcm a_21950_1126# 0.0989f
C25733 a_18026_6146# a_18026_5142# 0.843f
C25734 m3_20940_18146# m3_21944_18146# 0.202f
C25735 m2_13780_946# m3_14916_1078# 0.0341f
C25736 m2_22240_9406# a_22042_9158# 0.165f
C25737 col[31] a_33998_5142# 0.0682f
C25738 vcm a_9294_10202# 0.155f
C25739 col[27] a_2475_18218# 0.136f
C25740 a_11910_10162# a_12306_10202# 0.0313f
C25741 rowoff_n[15] a_5978_17190# 0.294f
C25742 a_2275_10186# a_22954_10162# 0.136f
C25743 rowoff_n[4] a_4882_6146# 0.202f
C25744 ctop a_22042_5142# 4.11f
C25745 col[21] a_2475_11190# 0.136f
C25746 VDD a_30986_10162# 0.181f
C25747 m2_1732_10986# m3_1864_12122# 0.0341f
C25748 col_n[19] a_22346_3174# 0.084f
C25749 a_30074_3134# a_30378_3174# 0.0931f
C25750 a_30986_3134# a_31478_3496# 0.0658f
C25751 col_n[29] a_32386_15222# 0.084f
C25752 col_n[3] a_5978_14178# 0.251f
C25753 vcm a_2161_4162# 0.0169f
C25754 a_2475_7174# a_15014_7150# 0.316f
C25755 a_7986_7150# a_8990_7150# 0.843f
C25756 rowoff_n[10] a_30986_12170# 0.202f
C25757 rowoff_n[2] a_13918_4138# 0.202f
C25758 col_n[28] a_2275_17214# 0.113f
C25759 col_n[10] a_12914_16186# 0.0765f
C25760 row_n[6] a_27062_8154# 0.282f
C25761 vcm a_24354_14218# 0.155f
C25762 rowon_n[10] a_26970_12170# 0.118f
C25763 VDD a_22442_4500# 0.0779f
C25764 col_n[31] rowoff_n[14] 0.0471f
C25765 m2_34864_16006# VDD 0.766f
C25766 a_31990_17190# a_32082_17190# 0.326f
C25767 VDD a_11910_13174# 0.181f
C25768 row_n[8] a_14314_10202# 0.0117f
C25769 rowoff_n[7] a_5374_9520# 0.0133f
C25770 rowoff_n[0] a_22954_2130# 0.202f
C25771 vcm m2_2736_946# 0.353f
C25772 col[18] a_2275_14202# 0.0899f
C25773 a_2275_4162# a_5978_4138# 0.399f
C25774 m3_12908_18146# ctop 0.209f
C25775 m2_13204_7398# a_13006_7150# 0.165f
C25776 col[23] a_2275_3158# 0.0899f
C25777 vcm a_17934_8154# 0.1f
C25778 m2_34864_18014# m2_35292_18442# 0.165f
C25779 a_2475_9182# a_30074_9158# 0.316f
C25780 a_33086_10162# a_33086_9158# 0.843f
C25781 m2_5172_8402# row_n[6] 0.0128f
C25782 rowoff_n[13] a_12402_15544# 0.0133f
C25783 col_n[1] a_3878_14178# 0.0765f
C25784 m2_11196_4386# row_n[2] 0.0128f
C25785 row_n[10] a_4882_12170# 0.0437f
C25786 col[23] a_26058_13174# 0.367f
C25787 col[20] a_22954_3134# 0.0682f
C25788 vcm a_5278_17230# 0.155f
C25789 a_26970_14178# a_27366_14218# 0.0313f
C25790 rowon_n[14] a_3970_16186# 0.248f
C25791 VDD a_2966_7150# 0.485f
C25792 col[30] a_32994_15182# 0.0682f
C25793 rowoff_n[5] a_14410_7512# 0.0133f
C25794 ctop a_18026_12170# 4.11f
C25795 a_2275_18218# a_6282_18234# 0.145f
C25796 row_n[0] a_14922_2130# 0.0437f
C25797 VDD a_26970_17190# 0.181f
C25798 rowon_n[4] a_14010_6146# 0.248f
C25799 m2_32280_3382# a_32082_3134# 0.165f
C25800 a_2275_6170# a_21038_6146# 0.399f
C25801 a_10998_6146# a_11302_6186# 0.0931f
C25802 col_n[8] a_11302_1166# 0.0839f
C25803 a_11910_6146# a_12402_6508# 0.0658f
C25804 col_n[18] a_21342_13214# 0.084f
C25805 rowoff_n[3] a_23446_5504# 0.0133f
C25806 row_n[2] a_2966_4138# 0.281f
C25807 vcm a_32994_12170# 0.1f
C25808 rowon_n[11] col[8] 0.0323f
C25809 row_n[15] col[15] 0.0342f
C25810 rowon_n[7] col[0] 0.0318f
C25811 row_n[13] col[11] 0.0342f
C25812 col_n[8] a_2475_10186# 0.0531f
C25813 rowon_n[9] col[4] 0.0323f
C25814 rowon_n[14] col[14] 0.0323f
C25815 rowon_n[10] col[6] 0.0323f
C25816 row_n[10] col[5] 0.0342f
C25817 rowon_n[4] ctop 0.203f
C25818 rowon_n[15] col[16] 0.0323f
C25819 rowon_n[12] col[10] 0.0323f
C25820 col_n[24] col[24] 0.489f
C25821 row_n[14] col[13] 0.0342f
C25822 rowon_n[13] col[12] 0.0323f
C25823 col_n[15] rowoff_n[15] 0.0471f
C25824 row_n[11] col[7] 0.0342f
C25825 row_n[12] col[9] 0.0342f
C25826 row_n[8] col[1] 0.0342f
C25827 row_n[9] col[3] 0.0342f
C25828 rowon_n[8] col[2] 0.0323f
C25829 a_23046_11166# a_24050_11166# 0.843f
C25830 VDD a_29070_2130# 0.483f
C25831 m2_20232_17438# row_n[15] 0.0128f
C25832 m2_26256_13422# row_n[11] 0.0128f
C25833 rowon_n[6] a_2275_8178# 1.79f
C25834 m2_32280_9406# row_n[7] 0.0128f
C25835 a_35002_16186# a_35398_16226# 0.0313f
C25836 VDD a_18426_11528# 0.0779f
C25837 col[18] rowoff_n[11] 0.0901f
C25838 ctop a_33086_16186# 4.11f
C25839 col_n[29] a_32482_7512# 0.0283f
C25840 a_2275_3158# a_11302_3174# 0.144f
C25841 a_2475_3158# a_13918_3134# 0.264f
C25842 a_7894_3134# a_7986_3134# 0.326f
C25843 rowoff_n[1] a_32482_3496# 0.0133f
C25844 rowoff_n[8] a_15014_10162# 0.294f
C25845 a_27062_1126# a_2475_1150# 0.0299f
C25846 m2_4168_5390# a_3970_5142# 0.165f
C25847 row_n[13] a_25054_15182# 0.282f
C25848 rowoff_n[11] a_18938_13174# 0.202f
C25849 vcm a_13918_15182# 0.1f
C25850 a_14010_13174# a_14010_12170# 0.843f
C25851 VDD a_9994_5142# 0.483f
C25852 row_n[3] a_35094_5142# 0.0123f
C25853 col[12] a_15014_11166# 0.367f
C25854 row_n[15] a_12306_17230# 0.0117f
C25855 rowon_n[7] a_35002_9158# 0.118f
C25856 a_7894_17190# a_8290_17230# 0.0313f
C25857 col[9] a_11910_1126# 0.0682f
C25858 a_2275_17214# a_14922_17190# 0.136f
C25859 rowoff_n[6] a_24050_8154# 0.294f
C25860 VDD a_33486_15544# 0.0779f
C25861 col_n[5] a_2275_13198# 0.113f
C25862 col[19] a_21950_13174# 0.0682f
C25863 col_n[10] a_2275_2154# 0.113f
C25864 row_n[5] a_22346_7190# 0.0117f
C25865 a_2275_5166# a_26362_5182# 0.144f
C25866 a_2475_5166# a_28978_5142# 0.264f
C25867 col_n[27] a_30074_7150# 0.251f
C25868 m3_10900_1078# m3_11904_1078# 0.202f
C25869 a_28978_1126# a_29070_1126# 0.0991f
C25870 rowoff_n[15] a_35002_17190# 0.202f
C25871 a_26970_10162# a_27462_10524# 0.0658f
C25872 a_26058_10162# a_26362_10202# 0.0931f
C25873 col_n[25] a_2475_12194# 0.0531f
C25874 rowoff_n[4] a_33086_6146# 0.294f
C25875 col_n[7] a_10298_11206# 0.084f
C25876 a_3970_14178# a_4974_14178# 0.843f
C25877 m2_22816_946# a_2275_1150# 0.28f
C25878 col[2] rowoff_n[12] 0.0901f
C25879 m2_8760_946# a_8990_1126# 0.0249f
C25880 a_2475_14202# a_6982_14178# 0.316f
C25881 col_n[30] a_2475_1150# 0.0481f
C25882 VDD a_25054_9158# 0.483f
C25883 row_n[7] a_12914_9158# 0.0437f
C25884 m2_1732_7974# m3_1864_9110# 0.0341f
C25885 rowon_n[11] a_12002_13174# 0.248f
C25886 VDD a_14410_18556# 0.0858f
C25887 a_2275_2154# a_19942_2130# 0.136f
C25888 col_n[18] a_21438_5504# 0.0283f
C25889 m2_15788_946# VDD 1f
C25890 vcm a_31078_4138# 0.56f
C25891 a_22954_7150# a_23046_7150# 0.326f
C25892 rowon_n[1] a_22042_3134# 0.248f
C25893 col_n[28] a_31478_17552# 0.0283f
C25894 col[15] a_2475_9182# 0.136f
C25895 a_2475_16210# a_22042_16186# 0.316f
C25896 a_29070_17190# a_29070_16186# 0.843f
C25897 VDD a_5978_12170# 0.483f
C25898 col[1] a_3970_9158# 0.367f
C25899 col_n[22] a_2275_15206# 0.113f
C25900 a_2275_4162# a_35002_4138# 0.136f
C25901 a_17934_4138# a_18330_4178# 0.0313f
C25902 col_n[27] a_2275_4162# 0.113f
C25903 col[8] a_10906_11166# 0.0682f
C25904 vcm a_12002_7150# 0.56f
C25905 rowoff_n[12] a_6890_14178# 0.202f
C25906 col_n[16] a_19030_5142# 0.251f
C25907 row_n[10] a_33086_12170# 0.282f
C25908 col_n[26] a_29070_17190# 0.251f
C25909 rowon_n[14] a_32994_16186# 0.118f
C25910 a_6982_13174# a_7286_13214# 0.0931f
C25911 a_7894_13174# a_8386_13536# 0.0658f
C25912 a_2275_13198# a_13006_13174# 0.399f
C25913 col_n[23] a_25966_7150# 0.0765f
C25914 col[12] a_2275_12194# 0.0899f
C25915 VDD a_21038_16186# 0.483f
C25916 col[17] a_2275_1150# 0.0896f
C25917 row_n[12] a_20338_14218# 0.0117f
C25918 vcm a_3878_1126# 0.0951f
C25919 m2_1732_2954# rowon_n[1] 0.236f
C25920 vcm a_27062_11166# 0.56f
C25921 col_n[7] a_10394_3496# 0.0283f
C25922 row_n[2] a_30378_4178# 0.0117f
C25923 a_2275_10186# a_3270_10202# 0.144f
C25924 a_2475_10186# a_5886_10162# 0.264f
C25925 row_n[14] a_10906_16186# 0.0437f
C25926 VDD a_23958_1126# 0.405f
C25927 col_n[17] a_20434_15544# 0.0283f
C25928 a_2275_15206# a_28066_15182# 0.399f
C25929 row_n[4] a_20946_6146# 0.0437f
C25930 a_4974_3134# a_4974_2130# 0.843f
C25931 rowon_n[8] a_20034_10162# 0.248f
C25932 col_n[2] a_2475_8178# 0.0531f
C25933 vcm a_17326_5182# 0.155f
C25934 a_32994_8154# a_33390_8194# 0.0313f
C25935 m2_10192_16434# rowon_n[14] 0.0322f
C25936 m2_16216_12418# rowon_n[10] 0.0322f
C25937 m2_22240_8402# rowon_n[6] 0.0322f
C25938 vcm a_7986_14178# 0.56f
C25939 a_2275_12194# a_18330_12210# 0.144f
C25940 m2_28264_4386# rowon_n[2] 0.0322f
C25941 a_2475_12194# a_20946_12170# 0.264f
C25942 VDD a_4882_4138# 0.181f
C25943 col_n[5] a_7986_3134# 0.251f
C25944 m2_35292_18442# VDD 0.0457f
C25945 col_n[15] a_18026_15182# 0.251f
C25946 a_22954_17190# a_23446_17552# 0.0658f
C25947 a_22042_17190# a_22346_17230# 0.0931f
C25948 col[29] a_2275_14202# 0.0899f
C25949 col_n[12] a_14922_5142# 0.0765f
C25950 col_n[22] a_24962_17190# 0.0765f
C25951 a_29070_5142# a_30074_5142# 0.843f
C25952 m2_16792_18014# m2_17796_18014# 0.843f
C25953 vcm a_32386_9198# 0.155f
C25954 a_2275_9182# a_11910_9158# 0.136f
C25955 rowon_n[2] a_7894_4138# 0.118f
C25956 col_n[0] a_2275_11190# 0.113f
C25957 vcm a_23046_18194# 0.165f
C25958 ctop a_10998_3134# 4.11f
C25959 m3_33992_1078# a_34090_2130# 0.0102f
C25960 a_2275_14202# a_33390_14218# 0.144f
C25961 a_18938_14178# a_19030_14178# 0.326f
C25962 VDD a_19942_8154# 0.181f
C25963 m2_1732_4962# m3_1864_6098# 0.0341f
C25964 col_n[6] a_9390_13536# 0.0283f
C25965 col[25] a_28066_2130# 0.367f
C25966 m3_11904_1078# VDD 0.0157f
C25967 row_n[9] a_28370_11206# 0.0117f
C25968 rowon_n[2] col[1] 0.0323f
C25969 col_n[26] rowoff_n[15] 0.0471f
C25970 rowon_n[12] col[21] 0.0323f
C25971 rowon_n[5] col[7] 0.0323f
C25972 vcm a_25966_3134# 0.1f
C25973 sw_n ctop 0.412f
C25974 rowon_n[6] col[9] 0.0323f
C25975 rowon_n[9] col[15] 0.0323f
C25976 row_n[11] col[18] 0.0342f
C25977 rowon_n[3] col[3] 0.0323f
C25978 row_n[7] col[10] 0.0342f
C25979 row_n[12] col[20] 0.0342f
C25980 row_n[10] col[16] 0.0342f
C25981 rowon_n[13] col[23] 0.0323f
C25982 row_n[14] col[24] 0.0342f
C25983 rowon_n[14] col[25] 0.0323f
C25984 col_n[29] col[30] 7.11f
C25985 rowon_n[7] col[11] 0.0323f
C25986 row_n[15] col[26] 0.0342f
C25987 row_n[2] col[0] 0.0322f
C25988 row_n[8] col[12] 0.0342f
C25989 row_n[5] col[6] 0.0342f
C25990 row_n[4] col[4] 0.0342f
C25991 rowon_n[10] col[17] 0.0323f
C25992 rowon_n[8] col[13] 0.0323f
C25993 row_n[9] col[14] 0.0342f
C25994 rowon_n[15] col[27] 0.0323f
C25995 rowon_n[11] col[19] 0.0323f
C25996 col_n[19] a_2475_10186# 0.0531f
C25997 row_n[3] col[2] 0.0342f
C25998 row_n[6] col[8] 0.0342f
C25999 row_n[13] col[22] 0.0342f
C26000 rowon_n[4] col[5] 0.0323f
C26001 a_20034_7150# a_20034_6146# 0.843f
C26002 a_2275_6170# a_2966_6146# 0.399f
C26003 a_2475_6170# a_3970_6146# 0.316f
C26004 rowoff_n[3] a_5886_5142# 0.202f
C26005 vcm a_13310_12210# 0.155f
C26006 a_13918_11166# a_14314_11206# 0.0313f
C26007 a_2275_11190# a_26970_11166# 0.136f
C26008 VDD a_11398_2492# 0.0779f
C26009 col[29] rowoff_n[11] 0.0901f
C26010 ctop a_26058_7150# 4.11f
C26011 row_n[11] a_18938_13174# 0.0437f
C26012 VDD a_35002_12170# 0.258f
C26013 m2_25828_18014# m3_25960_18146# 3.79f
C26014 col_n[20] a_23350_2170# 0.084f
C26015 rowon_n[15] a_18026_17190# 0.248f
C26016 col[9] a_2475_7174# 0.136f
C26017 col_n[4] a_6982_13174# 0.251f
C26018 col_n[30] a_33390_14218# 0.084f
C26019 a_32082_4138# a_32386_4178# 0.0931f
C26020 a_32994_4138# a_33486_4500# 0.0658f
C26021 row_n[1] a_28978_3134# 0.0437f
C26022 rowoff_n[1] a_14922_3134# 0.202f
C26023 col_n[11] a_13918_15182# 0.0765f
C26024 rowon_n[5] a_28066_7150# 0.248f
C26025 vcm a_6890_6146# 0.1f
C26026 rowoff_n[12] a_35094_14178# 0.0135f
C26027 a_9994_8154# a_10998_8154# 0.843f
C26028 a_2475_8178# a_19030_8154# 0.316f
C26029 vcm a_28370_16226# 0.155f
C26030 VDD a_26458_6508# 0.0779f
C26031 col_n[16] a_2275_13198# 0.113f
C26032 ctop a_6982_10162# 4.11f
C26033 col_n[21] a_2275_2154# 0.113f
C26034 a_33998_18194# a_34090_18194# 0.0991f
C26035 rowoff_n[6] a_6378_8516# 0.0133f
C26036 VDD a_15926_15182# 0.181f
C26037 a_2275_5166# a_9994_5142# 0.399f
C26038 row_n[5] a_5978_7150# 0.282f
C26039 m2_29844_946# m3_28972_1078# 0.0341f
C26040 m3_1864_14130# m3_1864_13126# 0.202f
C26041 col[24] a_27062_12170# 0.367f
C26042 rowon_n[9] a_5886_11166# 0.118f
C26043 col[13] rowoff_n[12] 0.0901f
C26044 col[6] a_2275_10186# 0.0899f
C26045 vcm a_21950_10162# 0.1f
C26046 col[21] a_23958_2130# 0.0682f
C26047 a_2475_10186# a_34090_10162# 0.316f
C26048 m2_18224_16434# a_18026_16186# 0.165f
C26049 rowoff_n[4] a_15414_6508# 0.0133f
C26050 col[31] a_33998_14178# 0.0682f
C26051 a_28978_15182# a_29374_15222# 0.0313f
C26052 VDD a_7382_9520# 0.0779f
C26053 m2_23820_18014# ctop 0.0422f
C26054 ctop a_22042_14178# 4.11f
C26055 m2_9188_15430# row_n[13] 0.0128f
C26056 col[26] a_2475_9182# 0.136f
C26057 m2_15212_11414# row_n[9] 0.0128f
C26058 m2_21236_7398# row_n[5] 0.0128f
C26059 m2_27260_3382# row_n[1] 0.0128f
C26060 col_n[19] a_22346_12210# 0.084f
C26061 a_13918_7150# a_14410_7512# 0.0658f
C26062 rowoff_n[9] a_6982_11166# 0.294f
C26063 a_13006_7150# a_13310_7190# 0.0931f
C26064 a_2275_7174# a_25054_7150# 0.399f
C26065 rowoff_n[2] a_24450_4500# 0.0133f
C26066 m2_34864_17010# vcm 0.408f
C26067 vcm a_2161_13198# 0.0169f
C26068 a_25054_12170# a_26058_12170# 0.843f
C26069 VDD a_33086_4138# 0.483f
C26070 a_2874_16186# a_2966_16186# 0.326f
C26071 VDD a_22442_13536# 0.0779f
C26072 col_n[30] a_33486_6508# 0.0283f
C26073 row_n[8] a_26970_10162# 0.0437f
C26074 rowoff_n[0] a_33486_2492# 0.0133f
C26075 rowoff_n[7] a_16018_9158# 0.294f
C26076 rowon_n[12] a_26058_14178# 0.248f
C26077 a_2275_4162# a_15318_4178# 0.144f
C26078 a_2475_4162# a_17934_4138# 0.264f
C26079 a_9902_4138# a_9994_4138# 0.326f
C26080 m3_1864_7102# ctop 0.21f
C26081 m2_35292_16434# row_n[14] 0.0128f
C26082 rowoff_n[13] a_23046_15182# 0.294f
C26083 m2_9188_14426# a_8990_14178# 0.165f
C26084 col[23] a_2275_12194# 0.0899f
C26085 col[13] a_16018_10162# 0.367f
C26086 vcm a_17934_17190# 0.1f
C26087 a_16018_14178# a_16018_13174# 0.843f
C26088 col[28] a_2275_1150# 0.0899f
C26089 VDD a_14010_7150# 0.483f
C26090 m2_1732_1950# m3_1864_3086# 0.0341f
C26091 rowoff_n[5] a_25054_7150# 0.294f
C26092 col[20] a_22954_12170# 0.0682f
C26093 a_2275_18218# a_18938_18194# 0.136f
C26094 a_9902_18194# a_10298_18234# 0.0313f
C26095 VDD a_2966_16186# 0.485f
C26096 a_2275_1150# a_8898_1126# 0.136f
C26097 a_4882_1126# a_5278_1166# 0.0313f
C26098 row_n[12] a_3970_14178# 0.282f
C26099 col_n[28] a_31078_6146# 0.251f
C26100 m2_6176_2378# a_5978_2130# 0.165f
C26101 vcm a_20034_2130# 0.56f
C26102 a_2275_6170# a_30378_6186# 0.144f
C26103 a_2475_6170# a_32994_6146# 0.264f
C26104 m2_28264_10410# a_28066_10162# 0.165f
C26105 m2_6752_946# col_n[4] 0.331f
C26106 row_n[2] a_14010_4138# 0.282f
C26107 rowoff_n[3] a_34090_5142# 0.294f
C26108 col_n[8] a_11302_10202# 0.084f
C26109 a_28978_11166# a_29470_11528# 0.0658f
C26110 a_28066_11166# a_28370_11206# 0.0931f
C26111 rowon_n[6] a_13918_8154# 0.118f
C26112 a_2475_15206# a_10998_15182# 0.316f
C26113 a_5978_15182# a_6982_15182# 0.843f
C26114 VDD a_29070_11166# 0.483f
C26115 col_n[13] a_2475_8178# 0.0531f
C26116 row_n[4] a_2275_6170# 19.2f
C26117 col_n[19] a_22442_4500# 0.0283f
C26118 a_2275_3158# a_23958_3134# 0.136f
C26119 rowon_n[8] a_1957_10186# 0.0172f
C26120 a_2475_18218# a_16930_18194# 0.264f
C26121 m2_34864_13998# rowoff_n[12] 0.278f
C26122 col_n[29] a_32482_16548# 0.0283f
C26123 row_n[13] a_35398_15222# 0.0117f
C26124 vcm a_35094_6146# 0.165f
C26125 rowoff_n[11] a_29470_13536# 0.0133f
C26126 a_24962_8154# a_25054_8154# 0.326f
C26127 m2_1732_7974# sample 0.2f
C26128 a_1957_12194# a_2161_12194# 0.115f
C26129 a_2475_12194# a_2275_12194# 2.76f
C26130 col[3] a_2475_5166# 0.136f
C26131 a_35494_1488# VDD 0.126f
C26132 row_n[15] a_24962_17190# 0.0437f
C26133 a_2475_17214# a_26058_17190# 0.316f
C26134 col[2] a_4974_8154# 0.367f
C26135 VDD a_9994_14178# 0.483f
C26136 col[9] a_11910_10162# 0.0682f
C26137 m2_1732_18014# col[0] 0.0137f
C26138 row_n[5] a_35002_7150# 0.0437f
C26139 a_19942_5142# a_20338_5182# 0.0313f
C26140 col_n[17] a_20034_4138# 0.251f
C26141 m2_19228_8402# a_19030_8154# 0.165f
C26142 col_n[10] a_2275_11190# 0.113f
C26143 rowon_n[9] a_34090_11166# 0.248f
C26144 vcm a_16018_9158# 0.56f
C26145 a_35002_1126# a_35398_1166# 0.0313f
C26146 rowoff_n[14] a_10998_16186# 0.294f
C26147 col_n[27] a_30074_16186# 0.251f
C26148 col_n[24] a_26970_6146# 0.0765f
C26149 a_2275_14202# a_17022_14178# 0.399f
C26150 a_8990_14178# a_9294_14218# 0.0931f
C26151 m2_14784_946# a_15318_1166# 0.087f
C26152 a_9902_14178# a_10394_14540# 0.0658f
C26153 VDD a_35398_9198# 0.0882f
C26154 rowon_n[10] col[28] 0.0323f
C26155 row_n[9] col[25] 0.0342f
C26156 rowon_n[7] col[22] 0.0323f
C26157 row_n[5] col[17] 0.0342f
C26158 rowon_n[11] col[30] 0.0323f
C26159 row_n[8] col[23] 0.0342f
C26160 row_n[11] col[29] 0.0342f
C26161 row_n[1] col[9] 0.0342f
C26162 row_n[0] col[7] 0.0342f
C26163 rowon_n[1] col[10] 0.0323f
C26164 rowon_n[3] col[14] 0.0323f
C26165 row_n[12] col[31] 0.0342f
C26166 rowon_n[5] col[18] 0.0323f
C26167 row_n[7] col[21] 0.0342f
C26168 rowon_n[8] col[24] 0.0323f
C26169 row_n[6] col[19] 0.0342f
C26170 row_n[2] col[11] 0.0342f
C26171 row_n[10] col[27] 0.0342f
C26172 row_n[4] col[15] 0.0342f
C26173 ctop col[4] 0.123f
C26174 rowon_n[6] col[20] 0.0323f
C26175 rowon_n[9] col[26] 0.0323f
C26176 row_n[3] col[13] 0.0342f
C26177 a_24354_1166# col_n[21] 0.0839f
C26178 rowon_n[0] col[8] 0.0323f
C26179 VDD a_25054_18194# 0.0356f
C26180 col_n[30] a_2475_10186# 0.0531f
C26181 rowon_n[2] col[12] 0.0323f
C26182 rowon_n[4] col[16] 0.0323f
C26183 rowon_n[12] sample_n 0.0692f
C26184 a_2475_2154# a_31078_2130# 0.316f
C26185 a_16018_2130# a_17022_2130# 0.843f
C26186 col[0] a_2275_8178# 0.099f
C26187 m3_7888_18146# VDD 0.0673f
C26188 vcm a_6282_3174# 0.155f
C26189 row_n[9] a_12002_11166# 0.282f
C26190 col_n[8] a_11398_2492# 0.0283f
C26191 rowon_n[13] a_11910_15182# 0.118f
C26192 col_n[18] a_21438_14540# 0.0283f
C26193 vcm a_31078_13174# 0.56f
C26194 a_2275_11190# a_7286_11206# 0.144f
C26195 a_2475_11190# a_9902_11166# 0.264f
C26196 a_5886_11166# a_5978_11166# 0.326f
C26197 VDD a_27974_3134# 0.181f
C26198 col[20] a_2475_7174# 0.136f
C26199 a_2275_16210# a_32082_16186# 0.399f
C26200 rowon_n[3] a_21950_5142# 0.118f
C26201 m2_1732_18014# m3_2868_18146# 0.0341f
C26202 m2_5172_10410# rowon_n[8] 0.0322f
C26203 m2_11196_6394# rowon_n[4] 0.0322f
C26204 m2_16216_2378# rowon_n[0] 0.0322f
C26205 a_6982_4138# a_6982_3134# 0.843f
C26206 row_n[1] a_9294_3174# 0.0117f
C26207 m2_10192_6394# a_9994_6146# 0.165f
C26208 vcm a_21342_7190# 0.155f
C26209 rowoff_n[12] a_17422_14540# 0.0133f
C26210 col_n[27] a_2275_13198# 0.113f
C26211 col_n[6] a_8990_2130# 0.251f
C26212 a_24962_1126# col[22] 0.0682f
C26213 ctop a_34090_2130# 4.05f
C26214 vcm a_12002_16186# 0.56f
C26215 a_2475_13198# a_24962_13174# 0.264f
C26216 a_2275_13198# a_22346_13214# 0.144f
C26217 col_n[16] a_19030_14178# 0.251f
C26218 VDD a_8898_6146# 0.181f
C26219 col_n[13] a_15926_4138# 0.0765f
C26220 a_24962_18194# a_25454_18556# 0.0658f
C26221 col_n[23] a_25966_16186# 0.0765f
C26222 a_19942_1126# a_20434_1488# 0.0667f
C26223 row_n[12] a_32994_14178# 0.0437f
C26224 a_19030_1126# a_19334_1166# 0.0997f
C26225 col[24] rowoff_n[12] 0.0901f
C26226 col[17] a_2275_10186# 0.0899f
C26227 vcm a_14922_1126# 0.0989f
C26228 m2_26256_15430# rowon_n[13] 0.0322f
C26229 m2_1732_3958# m2_2160_4386# 0.165f
C26230 a_31078_6146# a_32082_6146# 0.843f
C26231 m2_32280_11414# rowon_n[9] 0.0322f
C26232 m3_6884_18146# m3_7888_18146# 0.202f
C26233 m2_4744_946# m3_4876_1078# 3.79f
C26234 vcm a_3878_10162# 0.1f
C26235 a_2275_10186# a_15926_10162# 0.136f
C26236 ctop a_15014_5142# 4.11f
C26237 col_n[7] a_10394_12532# 0.0283f
C26238 m2_7756_946# a_7986_2130# 0.843f
C26239 a_20946_15182# a_21038_15182# 0.326f
C26240 VDD a_23958_10162# 0.181f
C26241 vcm a_29982_5142# 0.1f
C26242 rowoff_n[2] a_6890_4138# 0.202f
C26243 a_22042_8154# a_22042_7150# 0.843f
C26244 rowoff_n[10] a_23958_12170# 0.202f
C26245 a_2475_7174# a_7986_7150# 0.316f
C26246 col_n[2] a_2475_17214# 0.0531f
C26247 row_n[6] a_20034_8154# 0.282f
C26248 col_n[7] a_2475_6170# 0.0531f
C26249 vcm a_17326_14218# 0.155f
C26250 a_15926_12170# a_16322_12210# 0.0313f
C26251 a_2275_12194# a_30986_12170# 0.136f
C26252 VDD a_15414_4500# 0.0779f
C26253 rowon_n[10] a_19942_12170# 0.118f
C26254 ctop a_30074_9158# 4.11f
C26255 row_n[0] m2_32280_2378# 0.0128f
C26256 VDD a_4882_13174# 0.181f
C26257 col_n[5] a_7986_12170# 0.251f
C26258 col_n[2] a_4882_2130# 0.0765f
C26259 col[8] rowoff_n[13] 0.0901f
C26260 row_n[8] a_7286_10202# 0.0117f
C26261 rowon_n[0] a_29982_2130# 0.118f
C26262 rowoff_n[0] a_15926_2130# 0.202f
C26263 col_n[12] a_14922_14178# 0.0765f
C26264 a_35002_5142# a_35494_5504# 0.0658f
C26265 m2_27836_18014# m2_28264_18442# 0.165f
C26266 vcm a_10906_8154# 0.1f
C26267 a_12002_9158# a_13006_9158# 0.843f
C26268 a_2475_9182# a_23046_9158# 0.316f
C26269 rowoff_n[13] a_5374_15544# 0.0133f
C26270 vcm a_32386_18234# 0.16f
C26271 VDD a_30474_8516# 0.0779f
C26272 rowoff_n[5] a_7382_7512# 0.0133f
C26273 ctop a_10998_12170# 4.11f
C26274 VDD a_19942_17190# 0.181f
C26275 col_n[4] a_2275_9182# 0.113f
C26276 row_n[0] a_7894_2130# 0.0437f
C26277 a_30986_2130# a_31078_2130# 0.326f
C26278 rowon_n[4] a_6982_6146# 0.248f
C26279 vcm a_1957_2154# 0.139f
C26280 m2_34864_7974# m2_34864_6970# 0.843f
C26281 col[25] a_28066_11166# 0.367f
C26282 a_2275_6170# a_14010_6146# 0.399f
C26283 vcm a_25966_12170# 0.1f
C26284 rowoff_n[3] a_16418_5504# 0.0133f
C26285 VDD a_22042_2130# 0.483f
C26286 m2_34864_18014# a_35398_18234# 0.087f
C26287 col_n[24] a_2475_8178# 0.0531f
C26288 m2_4168_9406# row_n[7] 0.0128f
C26289 ctop a_2275_6170# 0.0683f
C26290 m2_10192_5390# row_n[3] 0.0128f
C26291 a_30986_16186# a_31382_16226# 0.0313f
C26292 VDD a_11398_11528# 0.0779f
C26293 ctop a_26058_16186# 4.11f
C26294 a_2275_3158# a_4274_3174# 0.144f
C26295 a_2475_3158# a_6890_3134# 0.264f
C26296 col_n[20] a_23350_11206# 0.084f
C26297 rowoff_n[1] a_25454_3496# 0.0133f
C26298 rowoff_n[8] a_7986_10162# 0.294f
C26299 m2_1732_15002# rowoff_n[13] 0.415f
C26300 col[9] a_2475_16210# 0.136f
C26301 row_n[13] a_18026_15182# 0.282f
C26302 a_15926_8154# a_16418_8516# 0.0658f
C26303 rowoff_n[11] a_11910_13174# 0.202f
C26304 a_15014_8154# a_15318_8194# 0.0931f
C26305 col[14] a_2475_5166# 0.136f
C26306 a_2275_8178# a_29070_8154# 0.399f
C26307 vcm a_6890_15182# 0.1f
C26308 a_27062_13174# a_28066_13174# 0.843f
C26309 VDD a_2874_5142# 0.182f
C26310 row_n[3] a_28066_5142# 0.282f
C26311 col_n[31] a_34490_5504# 0.0283f
C26312 row_n[15] a_5278_17230# 0.0117f
C26313 m2_25252_14426# row_n[12] 0.0128f
C26314 rowon_n[7] a_27974_9158# 0.118f
C26315 a_2275_17214# a_7894_17190# 0.136f
C26316 VDD a_26458_15544# 0.0779f
C26317 rowoff_n[6] a_17022_8154# 0.294f
C26318 m2_31276_10410# row_n[8] 0.0128f
C26319 col_n[21] a_2275_11190# 0.113f
C26320 m3_16924_18146# a_17022_17190# 0.0303f
C26321 a_11910_5142# a_12002_5142# 0.326f
C26322 a_2475_5166# a_21950_5142# 0.264f
C26323 a_2275_5166# a_19334_5182# 0.144f
C26324 row_n[5] a_15318_7190# 0.0117f
C26325 rowoff_n[15] a_27974_17190# 0.202f
C26326 col[14] a_17022_9158# 0.367f
C26327 rowoff_n[4] a_26058_6146# 0.294f
C26328 row_n[6] col[30] 0.0342f
C26329 rowon_n[6] col[31] 0.0323f
C26330 row_n[5] col[28] 0.0342f
C26331 rowon_n[4] col[27] 0.0323f
C26332 col[4] col[5] 0.0355f
C26333 row_n[2] col[22] 0.0342f
C26334 row_n[4] col[26] 0.0342f
C26335 m2_4744_946# a_3970_1126# 0.843f
C26336 rowon_n[3] col[25] 0.0323f
C26337 row_n[7] sample_n 0.0596f
C26338 rowon_n[0] col[19] 0.0323f
C26339 rowon_n[1] col[21] 0.0323f
C26340 rowon_n[5] col[29] 0.0323f
C26341 row_n[3] col[24] 0.0342f
C26342 ctop col[15] 0.124f
C26343 row_n[1] col[20] 0.0342f
C26344 rowon_n[2] col[23] 0.0323f
C26345 m2_8760_946# a_2475_1150# 0.286f
C26346 row_n[0] col[18] 0.0342f
C26347 col[21] a_23958_11166# 0.0682f
C26348 a_18026_15182# a_18026_14178# 0.843f
C26349 row_n[7] a_5886_9158# 0.0437f
C26350 VDD a_18026_9158# 0.483f
C26351 col[11] a_2275_8178# 0.0899f
C26352 rowon_n[11] a_4974_13174# 0.248f
C26353 col_n[29] a_32082_5142# 0.251f
C26354 VDD a_7382_18556# 0.0858f
C26355 a_6890_2130# a_7286_2170# 0.0313f
C26356 a_2275_2154# a_12914_2130# 0.136f
C26357 vcm a_24050_4138# 0.56f
C26358 rowon_n[1] a_15014_3134# 0.248f
C26359 rowoff_n[2] a_35094_4138# 0.0135f
C26360 a_2275_7174# a_35398_7190# 0.145f
C26361 col_n[9] a_12306_9198# 0.084f
C26362 col[31] a_2475_7174# 0.136f
C26363 a_30986_12170# a_31478_12532# 0.0658f
C26364 a_30074_12170# a_30378_12210# 0.0931f
C26365 m2_4744_18014# a_4882_18194# 0.225f
C26366 a_7986_16186# a_8990_16186# 0.843f
C26367 a_2475_16210# a_15014_16186# 0.316f
C26368 VDD a_33086_13174# 0.483f
C26369 rowon_n[3] a_3878_5142# 0.118f
C26370 col_n[20] a_23446_3496# 0.0283f
C26371 col_n[30] a_33486_15544# 0.0283f
C26372 a_2275_4162# a_27974_4138# 0.136f
C26373 col_n[1] a_2475_4162# 0.0531f
C26374 m3_31984_1078# ctop 0.21f
C26375 vcm a_4974_7150# 0.56f
C26376 a_26970_9158# a_27062_9158# 0.326f
C26377 row_n[10] a_26058_12170# 0.282f
C26378 rowon_n[14] a_25966_16186# 0.118f
C26379 a_2275_13198# a_5978_13174# 0.399f
C26380 col[3] a_5978_7150# 0.367f
C26381 col[28] a_2275_10186# 0.0899f
C26382 col[10] a_12914_9158# 0.0682f
C26383 VDD a_14010_16186# 0.483f
C26384 a_2475_1150# a_20034_1126# 0.31f
C26385 row_n[12] a_13310_14218# 0.0117f
C26386 col_n[18] a_21038_3134# 0.251f
C26387 vcm a_29374_2170# 0.155f
C26388 a_21950_6146# a_22346_6186# 0.0313f
C26389 col_n[28] a_31078_15182# 0.251f
C26390 m2_1732_8978# a_2161_9182# 0.0454f
C26391 col_n[25] a_27974_5142# 0.0765f
C26392 vcm a_20034_11166# 0.56f
C26393 row_n[2] a_23350_4178# 0.0117f
C26394 VDD a_16930_1126# 0.405f
C26395 m2_24248_17438# a_24050_17190# 0.165f
C26396 a_2275_15206# a_21038_15182# 0.399f
C26397 a_11910_15182# a_12402_15544# 0.0658f
C26398 a_10998_15182# a_11302_15222# 0.0931f
C26399 col[1] a_3878_7150# 0.0682f
C26400 row_n[4] a_13918_6146# 0.0437f
C26401 rowon_n[8] a_13006_10162# 0.248f
C26402 a_18026_3134# a_19030_3134# 0.843f
C26403 col_n[13] a_2475_17214# 0.0531f
C26404 a_2475_3158# a_35094_3134# 0.0299f
C26405 col_n[9] a_12402_1488# 0.0283f
C26406 col_n[18] a_2475_6170# 0.0531f
C26407 vcm a_10298_5182# 0.155f
C26408 col_n[19] a_22442_13536# 0.0283f
C26409 m2_34864_11990# a_2475_12194# 0.282f
C26410 row_n[6] a_1957_8178# 0.187f
C26411 vcm a_35094_15182# 0.165f
C26412 a_7894_12170# a_7986_12170# 0.326f
C26413 a_2275_12194# a_11302_12210# 0.144f
C26414 a_2475_12194# a_13918_12170# 0.264f
C26415 VDD a_31990_5142# 0.181f
C26416 col[19] rowoff_n[13] 0.0901f
C26417 m2_21236_18442# VDD 0.0456f
C26418 col[3] a_2475_14202# 0.136f
C26419 col[8] a_2475_3158# 0.136f
C26420 VDD rowoff_n[4] 1.51f
C26421 col_n[2] rowoff_n[9] 0.0471f
C26422 col_n[0] rowoff_n[6] 0.0471f
C26423 vcm rowoff_n[7] 0.533f
C26424 col_n[1] rowoff_n[8] 0.0471f
C26425 sample rowoff_n[5] 0.0775f
C26426 col[2] a_4974_17190# 0.367f
C26427 a_8990_5142# a_8990_4138# 0.843f
C26428 vcm a_25358_9198# 0.155f
C26429 m2_9764_18014# m2_10768_18014# 0.843f
C26430 a_2275_9182# a_4882_9158# 0.136f
C26431 a_2966_9158# a_3970_9158# 0.843f
C26432 col_n[17] a_20034_13174# 0.251f
C26433 m2_15212_15430# a_15014_15182# 0.165f
C26434 ctop a_3970_3134# 4.11f
C26435 col_n[14] a_16930_3134# 0.0765f
C26436 vcm a_16018_18194# 0.165f
C26437 col_n[15] a_2275_9182# 0.113f
C26438 a_2275_14202# a_26362_14218# 0.144f
C26439 a_2475_14202# a_28978_14178# 0.264f
C26440 m2_14784_18014# col[12] 0.347f
C26441 m2_9188_17438# rowon_n[15] 0.0322f
C26442 row_n[7] a_34090_9158# 0.282f
C26443 VDD a_12914_8154# 0.181f
C26444 m2_15212_13422# rowon_n[11] 0.0322f
C26445 m2_21236_9406# rowon_n[7] 0.0322f
C26446 col_n[24] a_26970_15182# 0.0765f
C26447 m2_27260_5390# rowon_n[3] 0.0322f
C26448 m2_20808_946# vcm 0.353f
C26449 rowon_n[11] a_33998_13174# 0.118f
C26450 VDD a_35398_18234# 0.103f
C26451 a_21038_2130# a_21342_2170# 0.0931f
C26452 a_21950_2130# a_22442_2492# 0.0658f
C26453 vcm a_18938_3134# 0.1f
C26454 row_n[9] a_21342_11206# 0.0117f
C26455 col[0] a_2275_17214# 0.099f
C26456 a_33086_7150# a_34090_7150# 0.843f
C26457 m2_34288_11414# a_34090_11166# 0.165f
C26458 col[5] a_2275_6170# 0.0899f
C26459 vcm a_6282_12210# 0.155f
C26460 a_2275_11190# a_19942_11166# 0.136f
C26461 col_n[8] a_11398_11528# 0.0283f
C26462 col[3] rowoff_n[14] 0.0901f
C26463 VDD a_4370_2492# 0.0779f
C26464 col_n[31] a_34394_2170# 0.0839f
C26465 m2_23820_18014# a_23958_18194# 0.225f
C26466 ctop a_19030_7150# 4.11f
C26467 row_n[11] a_11910_13174# 0.0437f
C26468 a_22954_16186# a_23046_16186# 0.326f
C26469 VDD a_27974_12170# 0.181f
C26470 m2_16792_18014# m3_15920_18146# 0.0341f
C26471 rowon_n[15] a_10998_17190# 0.248f
C26472 col[20] a_2475_16210# 0.136f
C26473 col[25] a_2475_5166# 0.136f
C26474 row_n[1] a_21950_3134# 0.0437f
C26475 rowoff_n[1] a_7894_3134# 0.202f
C26476 vcm a_33998_7150# 0.1f
C26477 rowon_n[5] a_21038_7150# 0.248f
C26478 a_2475_8178# a_12002_8154# 0.316f
C26479 a_24050_9158# a_24050_8154# 0.843f
C26480 rowoff_n[12] a_28066_14178# 0.294f
C26481 m2_6176_13422# a_5978_13174# 0.165f
C26482 vcm a_21342_16226# 0.155f
C26483 a_2275_13198# a_35002_13174# 0.136f
C26484 a_17934_13174# a_18330_13214# 0.0313f
C26485 VDD a_19430_6508# 0.0779f
C26486 m2_1732_4962# ctop 0.0428f
C26487 col_n[6] a_8990_11166# 0.251f
C26488 ctop a_34090_11166# 4.06f
C26489 col_n[3] a_5886_1126# 0.0765f
C26490 VDD a_8898_15182# 0.181f
C26491 col_n[13] a_15926_13174# 0.0765f
C26492 m2_30848_18014# col_n[28] 0.243f
C26493 a_2275_5166# a_2874_5142# 0.136f
C26494 a_2475_5166# a_3878_5142# 0.264f
C26495 m2_25252_9406# a_25054_9158# 0.165f
C26496 VDD col_n[3] 5.17f
C26497 rowon_n[0] col[30] 0.0323f
C26498 ctop col[26] 0.123f
C26499 rowon_n[1] sample_n 0.0692f
C26500 vcm a_14922_10162# 0.1f
C26501 row_n[0] col[29] 0.0342f
C26502 row_n[1] col[31] 0.0342f
C26503 a_2475_10186# a_27062_10162# 0.316f
C26504 a_14010_10162# a_15014_10162# 0.843f
C26505 col[22] a_2275_8178# 0.0899f
C26506 row_n[14] a_32082_16186# 0.282f
C26507 rowoff_n[4] a_8386_6508# 0.0133f
C26508 VDD a_34490_10524# 0.0779f
C26509 m2_9764_18014# ctop 0.0422f
C26510 ctop a_15014_14178# 4.11f
C26511 a_32994_3134# a_33086_3134# 0.326f
C26512 col[26] a_29070_10162# 0.367f
C26513 rowoff_n[2] a_17422_4500# 0.0133f
C26514 a_2275_7174# a_18026_7150# 0.399f
C26515 rowoff_n[10] a_34490_12532# 0.0133f
C26516 row_n[6] a_29374_8194# 0.0117f
C26517 vcm a_29982_14178# 0.1f
C26518 a_4974_12170# a_4974_11166# 0.843f
C26519 VDD a_26058_4138# 0.483f
C26520 col_n[7] a_2475_15206# 0.0531f
C26521 a_32994_17190# a_33390_17230# 0.0313f
C26522 VDD a_15414_13536# 0.0779f
C26523 col_n[12] a_2475_4162# 0.0531f
C26524 row_n[8] a_19942_10162# 0.0437f
C26525 col_n[21] a_24354_10202# 0.084f
C26526 rowoff_n[0] a_26458_2492# 0.0133f
C26527 rowoff_n[7] a_8990_9158# 0.294f
C26528 rowon_n[12] a_19030_14178# 0.248f
C26529 a_2475_4162# a_10906_4138# 0.264f
C26530 a_2275_4162# a_8290_4178# 0.144f
C26531 m3_27968_18146# ctop 0.209f
C26532 col_n[2] a_4882_11166# 0.0765f
C26533 m2_16216_7398# a_16018_7150# 0.165f
C26534 m2_8184_16434# row_n[14] 0.0128f
C26535 m2_14208_12418# row_n[10] 0.0128f
C26536 a_17022_9158# a_17326_9198# 0.0931f
C26537 a_2275_9182# a_33086_9158# 0.399f
C26538 m2_20232_8402# row_n[6] 0.0128f
C26539 rowoff_n[13] a_16018_15182# 0.294f
C26540 a_17934_9158# a_18426_9520# 0.0658f
C26541 m2_26256_4386# row_n[2] 0.0128f
C26542 rowon_n[2] a_29070_4138# 0.248f
C26543 vcm a_10906_17190# 0.1f
C26544 col[2] a_2475_1150# 0.136f
C26545 a_29070_14178# a_30074_14178# 0.843f
C26546 VDD a_6982_7150# 0.483f
C26547 rowoff_n[5] a_18026_7150# 0.294f
C26548 a_2275_18218# a_11910_18194# 0.136f
C26549 VDD a_30474_17552# 0.0779f
C26550 a_2475_1150# a_1957_1150# 0.0734f
C26551 m2_34864_2954# a_35094_3134# 0.0249f
C26552 col_n[4] a_2275_18218# 0.113f
C26553 vcm a_13006_2130# 0.56f
C26554 a_2475_6170# a_25966_6146# 0.264f
C26555 a_2275_6170# a_23350_6186# 0.144f
C26556 a_13918_6146# a_14010_6146# 0.326f
C26557 col[15] a_18026_8154# 0.367f
C26558 col_n[9] a_2275_7174# 0.113f
C26559 row_n[2] a_6982_4138# 0.282f
C26560 rowoff_n[3] a_27062_5142# 0.294f
C26561 vcm a_1957_11190# 0.139f
C26562 m2_34864_17010# row_n[15] 0.267f
C26563 col[22] a_24962_10162# 0.0682f
C26564 m2_19804_18014# a_20034_17190# 0.843f
C26565 rowon_n[6] a_6890_8154# 0.118f
C26566 a_2275_15206# a_2966_15182# 0.399f
C26567 a_20034_16186# a_20034_15182# 0.843f
C26568 a_2475_15206# a_3970_15182# 0.316f
C26569 col_n[30] a_33086_4138# 0.251f
C26570 VDD a_22042_11166# 0.483f
C26571 col_n[24] a_2475_17214# 0.0531f
C26572 ctop a_2275_15206# 0.0683f
C26573 col_n[29] a_2475_6170# 0.0531f
C26574 a_2275_3158# a_16930_3134# 0.136f
C26575 a_8898_3134# a_9294_3174# 0.0313f
C26576 a_2475_18218# a_9902_18194# 0.264f
C26577 col_n[10] a_13310_8194# 0.084f
C26578 a_30074_1126# a_2275_1150# 0.0924f
C26579 m2_7180_5390# a_6982_5142# 0.165f
C26580 row_n[13] a_27366_15222# 0.0117f
C26581 vcm a_28066_6146# 0.56f
C26582 rowoff_n[11] a_22442_13536# 0.0133f
C26583 col[30] rowoff_n[13] 0.0901f
C26584 a_32082_13174# a_32386_13214# 0.0931f
C26585 col[14] a_2475_14202# 0.136f
C26586 a_32994_13174# a_33486_13536# 0.0658f
C26587 col_n[12] rowoff_n[8] 0.0471f
C26588 col_n[10] rowoff_n[6] 0.0471f
C26589 col_n[13] rowoff_n[9] 0.0471f
C26590 col_n[11] rowoff_n[7] 0.0471f
C26591 col_n[4] rowoff_n[0] 0.0471f
C26592 col_n[8] rowoff_n[4] 0.0471f
C26593 col_n[7] rowoff_n[3] 0.0471f
C26594 a_27462_1488# VDD 0.0977f
C26595 col_n[6] rowoff_n[2] 0.0471f
C26596 col[19] a_2475_3158# 0.136f
C26597 col_n[5] rowoff_n[1] 0.0471f
C26598 col_n[9] rowoff_n[5] 0.0471f
C26599 row_n[15] a_17934_17190# 0.0437f
C26600 col_n[21] a_24450_2492# 0.0283f
C26601 a_9994_17190# a_10998_17190# 0.843f
C26602 a_2475_17214# a_19030_17190# 0.316f
C26603 VDD a_2874_14178# 0.182f
C26604 col_n[31] a_34490_14540# 0.0283f
C26605 row_n[5] a_27974_7150# 0.0437f
C26606 a_2275_5166# a_31990_5142# 0.136f
C26607 m2_1732_2954# sample_n 0.0522f
C26608 rowon_n[9] a_27062_11166# 0.248f
C26609 vcm a_8990_9158# 0.56f
C26610 col_n[26] a_2275_9182# 0.113f
C26611 a_29982_1126# a_30378_1166# 0.0313f
C26612 a_28978_10162# a_29070_10162# 0.326f
C26613 rowoff_n[14] a_3970_16186# 0.294f
C26614 col[4] a_6982_6146# 0.367f
C26615 m2_31852_946# a_2475_1150# 0.286f
C26616 a_2275_14202# a_9994_14178# 0.399f
C26617 col[11] a_13918_8154# 0.0682f
C26618 VDD a_18026_18194# 0.0356f
C26619 col_n[19] a_22042_2130# 0.251f
C26620 col[11] a_2275_17214# 0.0899f
C26621 a_30074_3134# a_30074_2130# 0.843f
C26622 a_2475_2154# a_24050_2130# 0.316f
C26623 col_n[29] a_32082_14178# 0.251f
C26624 col[16] a_2275_6170# 0.0899f
C26625 m2_24824_946# VDD 1f
C26626 col_n[26] a_28978_4138# 0.0765f
C26627 vcm a_33390_4178# 0.155f
C26628 row_n[9] a_4974_11166# 0.282f
C26629 rowoff_n[9] a_28978_11166# 0.202f
C26630 col[14] rowoff_n[14] 0.0901f
C26631 a_23958_7150# a_24354_7190# 0.0313f
C26632 rowon_n[13] a_4882_15182# 0.118f
C26633 vcm a_24050_13174# 0.56f
C26634 VDD a_20946_3134# 0.181f
C26635 col_n[9] a_12306_18234# 0.084f
C26636 VDD rowoff_n[10] 1.51f
C26637 m2_29844_18014# a_2275_18218# 0.28f
C26638 col[31] a_2475_16210# 0.136f
C26639 a_2275_16210# a_25054_16186# 0.399f
C26640 a_13918_16186# a_14410_16548# 0.0658f
C26641 a_13006_16186# a_13310_16226# 0.0931f
C26642 rowon_n[3] a_14922_5142# 0.118f
C26643 a_31078_1126# m2_30848_946# 0.0249f
C26644 a_20034_4138# a_21038_4138# 0.843f
C26645 col_n[20] a_23446_12532# 0.0283f
C26646 row_n[1] a_3878_3134# 0.0437f
C26647 rowon_n[5] a_2966_7150# 0.248f
C26648 vcm a_14314_7190# 0.155f
C26649 col_n[1] a_2475_13198# 0.0531f
C26650 rowoff_n[12] a_10394_14540# 0.0133f
C26651 col_n[6] a_2475_2154# 0.0531f
C26652 ctop a_27062_2130# 4.06f
C26653 vcm a_4974_16186# 0.56f
C26654 a_2475_13198# a_17934_13174# 0.264f
C26655 a_9902_13174# a_9994_13174# 0.326f
C26656 a_2275_13198# a_15318_13214# 0.144f
C26657 m2_25828_18014# a_2475_18218# 0.286f
C26658 col[3] a_5978_16186# 0.367f
C26659 row_n[12] a_25966_14178# 0.0437f
C26660 VDD col_n[14] 5.17f
C26661 vcm col_n[11] 1.94f
C26662 col_n[5] col_n[6] 0.0101f
C26663 col[15] col[16] 0.0337f
C26664 col[10] a_12914_18194# 0.0682f
C26665 vcm a_7894_1126# 0.0989f
C26666 m2_4168_11414# rowon_n[9] 0.0322f
C26667 a_10998_6146# a_10998_5142# 0.843f
C26668 m2_10192_7398# rowon_n[5] 0.0322f
C26669 m2_16216_3382# rowon_n[1] 0.0322f
C26670 col_n[18] a_21038_12170# 0.251f
C26671 vcm a_29374_11206# 0.155f
C26672 row_n[2] a_34394_4178# 0.0117f
C26673 col_n[15] a_17934_2130# 0.0765f
C26674 a_2275_10186# a_8898_10162# 0.136f
C26675 a_4882_10162# a_5278_10202# 0.0313f
C26676 rowon_n[6] a_35094_8154# 0.0141f
C26677 col_n[25] a_27974_14178# 0.0765f
C26678 ctop a_7986_5142# 4.11f
C26679 a_2275_15206# a_30378_15222# 0.144f
C26680 a_2475_15206# a_32994_15182# 0.264f
C26681 VDD a_16930_10162# 0.181f
C26682 col_n[3] a_2275_5166# 0.113f
C26683 a_23958_3134# a_24450_3496# 0.0658f
C26684 a_23046_3134# a_23350_3174# 0.0931f
C26685 col[1] a_3878_16186# 0.0682f
C26686 vcm a_22954_5142# 0.1f
C26687 rowoff_n[10] a_16930_12170# 0.202f
C26688 col_n[9] a_12402_10524# 0.0283f
C26689 m2_25252_16434# rowon_n[14] 0.0322f
C26690 row_n[6] a_13006_8154# 0.282f
C26691 col_n[18] a_2475_15206# 0.0531f
C26692 m2_31276_12418# rowon_n[10] 0.0322f
C26693 vcm a_10298_14218# 0.155f
C26694 a_2275_12194# a_23958_12170# 0.136f
C26695 VDD a_8386_4500# 0.0779f
C26696 col_n[23] a_2475_4162# 0.0531f
C26697 rowon_n[10] a_12914_12170# 0.118f
C26698 ctop a_23046_9158# 4.11f
C26699 a_24962_17190# a_25054_17190# 0.326f
C26700 VDD a_31990_14178# 0.181f
C26701 rowon_n[0] a_22954_2130# 0.118f
C26702 rowoff_n[0] a_8898_2130# 0.202f
C26703 col[8] a_2475_12194# 0.136f
C26704 m2_11772_946# ctop 0.0428f
C26705 m2_1732_6970# a_2475_7174# 0.139f
C26706 m2_20808_18014# m2_21236_18442# 0.165f
C26707 col[13] a_2475_1150# 0.136f
C26708 a_26058_10162# a_26058_9158# 0.843f
C26709 rowoff_n[14] a_32994_16186# 0.202f
C26710 a_2475_9182# a_16018_9158# 0.316f
C26711 vcm a_25358_18234# 0.16f
C26712 col_n[7] a_9994_10162# 0.251f
C26713 a_19942_14178# a_20338_14218# 0.0313f
C26714 VDD a_23446_8516# 0.0779f
C26715 col_n[14] a_16930_12170# 0.0765f
C26716 ctop a_3970_12170# 4.11f
C26717 col_n[15] a_2275_18218# 0.113f
C26718 VDD a_12914_17190# 0.181f
C26719 col_n[20] a_2275_7174# 0.113f
C26720 m2_31852_946# col[29] 0.425f
C26721 m3_26964_1078# VDD 0.0157f
C26722 row_n[9] a_33998_11166# 0.0437f
C26723 a_2275_6170# a_6982_6146# 0.399f
C26724 a_3970_6146# a_4274_6186# 0.0931f
C26725 a_4882_6146# a_5374_6508# 0.0658f
C26726 rowon_n[13] a_33086_15182# 0.248f
C26727 rowoff_n[3] a_9390_5504# 0.0133f
C26728 vcm a_18938_12170# 0.1f
C26729 a_16018_11166# a_17022_11166# 0.843f
C26730 a_2475_11190# a_31078_11166# 0.316f
C26731 VDD a_15014_2130# 0.483f
C26732 col[5] a_2275_15206# 0.0899f
C26733 col[10] a_2275_4162# 0.0899f
C26734 VDD a_4370_11528# 0.0779f
C26735 a_25454_1488# col_n[22] 0.0283f
C26736 m2_30848_18014# m3_30980_18146# 3.79f
C26737 col_n[31] a_34394_11206# 0.084f
C26738 ctop a_19030_16186# 4.11f
C26739 col[27] a_30074_9158# 0.367f
C26740 a_34090_4138# a_34394_4178# 0.0931f
C26741 a_35002_4138# a_35094_4138# 0.0991f
C26742 rowoff_n[1] a_18426_3496# 0.0133f
C26743 row_n[13] a_10998_15182# 0.282f
C26744 col[25] a_2475_14202# 0.136f
C26745 rowoff_n[11] a_4882_13174# 0.202f
C26746 a_2275_8178# a_22042_8154# 0.399f
C26747 col_n[21] rowoff_n[6] 0.0471f
C26748 col[30] a_2475_3158# 0.136f
C26749 col_n[22] rowoff_n[7] 0.0471f
C26750 col_n[18] rowoff_n[3] 0.0471f
C26751 col_n[16] rowoff_n[1] 0.0471f
C26752 col_n[15] rowoff_n[0] 0.0471f
C26753 col_n[23] rowoff_n[8] 0.0471f
C26754 col_n[17] rowoff_n[2] 0.0471f
C26755 col_n[24] rowoff_n[9] 0.0471f
C26756 col_n[19] rowoff_n[4] 0.0471f
C26757 col_n[20] rowoff_n[5] 0.0471f
C26758 vcm a_33998_16186# 0.1f
C26759 a_6982_13174# a_6982_12170# 0.843f
C26760 VDD a_30074_6146# 0.483f
C26761 row_n[3] a_21038_5142# 0.282f
C26762 col_n[1] a_2475_18218# 0.0529f
C26763 col_n[22] a_25358_9198# 0.084f
C26764 rowon_n[7] a_20946_9158# 0.118f
C26765 m2_3164_10410# row_n[8] 0.0128f
C26766 rowoff_n[6] a_9994_8154# 0.294f
C26767 VDD a_19430_15544# 0.0779f
C26768 m2_9188_6394# row_n[4] 0.0128f
C26769 m2_14208_2378# row_n[0] 0.0128f
C26770 col_n[3] a_5886_10162# 0.0765f
C26771 a_2275_5166# a_12306_5182# 0.144f
C26772 row_n[5] a_8290_7190# 0.0117f
C26773 a_2475_5166# a_14922_5142# 0.264f
C26774 m2_34864_946# m3_34568_1078# 0.0345f
C26775 m2_33860_946# m3_34996_1078# 0.027f
C26776 rowoff_n[15] a_20946_17190# 0.202f
C26777 a_19030_10162# a_19334_10202# 0.0931f
C26778 a_19942_10162# a_20434_10524# 0.0658f
C26779 m2_21236_16434# a_21038_16186# 0.165f
C26780 rowoff_n[4] a_19030_6146# 0.294f
C26781 a_31078_15182# a_32082_15182# 0.843f
C26782 VDD a_10998_9158# 0.483f
C26783 col[22] a_2275_17214# 0.0899f
C26784 col[27] a_2275_6170# 0.0899f
C26785 col[25] rowoff_n[14] 0.0901f
C26786 a_2275_2154# a_5886_2130# 0.136f
C26787 m2_24248_15430# row_n[13] 0.0128f
C26788 m2_30272_11414# row_n[9] 0.0128f
C26789 col[16] a_19030_7150# 0.367f
C26790 m2_35292_7398# row_n[5] 0.0128f
C26791 vcm a_17022_4138# 0.56f
C26792 a_2475_7174# a_29982_7150# 0.264f
C26793 col_n[8] rowoff_n[10] 0.0471f
C26794 a_15926_7150# a_16018_7150# 0.326f
C26795 a_2275_7174# a_27366_7190# 0.144f
C26796 rowoff_n[2] a_28066_4138# 0.294f
C26797 rowon_n[1] a_7986_3134# 0.248f
C26798 col[23] a_25966_9158# 0.0682f
C26799 ctop m2_2736_946# 0.0153f
C26800 VDD a_2275_3158# 1.96f
C26801 col_n[31] a_34090_3134# 0.251f
C26802 a_2475_16210# a_7986_16186# 0.316f
C26803 a_22042_17190# a_22042_16186# 0.843f
C26804 VDD a_26058_13174# 0.483f
C26805 col_n[11] a_14314_7190# 0.084f
C26806 col_n[12] a_2475_13198# 0.0531f
C26807 a_10906_4138# a_11302_4178# 0.0313f
C26808 a_2275_4162# a_20946_4138# 0.136f
C26809 m3_3872_1078# ctop 0.311f
C26810 col_n[17] a_2475_2154# 0.0531f
C26811 vcm a_32082_8154# 0.56f
C26812 row_n[10] a_19030_12170# 0.282f
C26813 m2_12200_14426# a_12002_14178# 0.165f
C26814 a_35002_14178# a_35494_14540# 0.0658f
C26815 rowon_n[14] a_18938_16186# 0.118f
C26816 vcm col_n[22] 1.94f
C26817 VDD col_n[25] 5.17f
C26818 col[9] rowoff_n[15] 0.0901f
C26819 m3_34996_10114# a_34090_10162# 0.0303f
C26820 col[2] a_2475_10186# 0.136f
C26821 row_n[0] a_29070_2130# 0.282f
C26822 VDD a_6982_16186# 0.483f
C26823 row_n[12] a_6282_14218# 0.0117f
C26824 a_2475_1150# a_13006_1126# 0.0299f
C26825 rowon_n[4] a_28978_6146# 0.118f
C26826 m2_9188_2378# a_8990_2130# 0.165f
C26827 vcm a_22346_2170# 0.155f
C26828 a_2275_6170# a_34394_6186# 0.144f
C26829 m2_11772_946# m2_12776_946# 0.843f
C26830 m2_31276_10410# a_31078_10162# 0.165f
C26831 col[5] a_7986_5142# 0.367f
C26832 row_n[2] a_16322_4178# 0.0117f
C26833 vcm a_13006_11166# 0.56f
C26834 a_30986_11166# a_31078_11166# 0.326f
C26835 col[15] a_18026_17190# 0.367f
C26836 VDD a_9902_1126# 0.405f
C26837 col_n[9] a_2275_16210# 0.113f
C26838 col[12] a_14922_7150# 0.0682f
C26839 col_n[14] a_2275_5166# 0.113f
C26840 a_2275_15206# a_14010_15182# 0.399f
C26841 rowon_n[0] m2_21236_2378# 0.0322f
C26842 row_n[4] a_6890_6146# 0.0437f
C26843 col_n[30] a_33086_13174# 0.251f
C26844 col_n[27] a_29982_3134# 0.0765f
C26845 a_2475_3158# a_28066_3134# 0.316f
C26846 a_32082_4138# a_32082_3134# 0.843f
C26847 rowon_n[8] a_5978_10162# 0.248f
C26848 rowoff_n[8] a_29982_10162# 0.202f
C26849 col_n[29] a_2475_15206# 0.0531f
C26850 vcm a_3270_5182# 0.155f
C26851 rowoff_n[11] a_33086_13174# 0.294f
C26852 a_25966_8154# a_26362_8194# 0.0313f
C26853 col_n[10] a_13310_17230# 0.084f
C26854 col[4] a_2275_2154# 0.0899f
C26855 vcm a_28066_15182# 0.56f
C26856 a_2275_12194# a_4274_12210# 0.144f
C26857 a_2475_12194# a_6890_12170# 0.264f
C26858 VDD a_24962_5142# 0.181f
C26859 m2_7180_18442# VDD 0.0456f
C26860 a_2275_17214# a_29070_17190# 0.399f
C26861 a_15014_17190# a_15318_17230# 0.0931f
C26862 a_15926_17190# a_16418_17552# 0.0658f
C26863 col[19] a_2475_12194# 0.136f
C26864 col_n[21] a_24450_11528# 0.0283f
C26865 col[24] a_2475_1150# 0.136f
C26866 a_22042_5142# a_23046_5142# 0.843f
C26867 m2_22240_8402# a_22042_8154# 0.165f
C26868 vcm a_18330_9198# 0.155f
C26869 m2_2736_18014# m2_3740_18014# 0.843f
C26870 sample a_2161_5166# 0.0858f
C26871 ctop a_31078_4138# 4.11f
C26872 col_n[26] a_2275_18218# 0.113f
C26873 vcm a_8990_18194# 0.165f
C26874 a_2475_14202# a_21950_14178# 0.264f
C26875 a_2275_14202# a_19334_14218# 0.144f
C26876 a_11910_14178# a_12002_14178# 0.326f
C26877 VDD a_5886_8154# 0.181f
C26878 row_n[7] a_27062_9158# 0.282f
C26879 col_n[31] a_2275_7174# 0.113f
C26880 col[4] a_6982_15182# 0.367f
C26881 rowon_n[11] a_26970_13174# 0.118f
C26882 VDD a_27366_18234# 0.019f
C26883 col[11] a_13918_17190# 0.0682f
C26884 a_2275_2154# a_34090_2130# 0.399f
C26885 m3_22948_18146# VDD 0.0885f
C26886 col_n[19] a_22042_11166# 0.251f
C26887 row_n[9] a_14314_11206# 0.0117f
C26888 vcm a_11910_3134# 0.1f
C26889 a_13006_7150# a_13006_6146# 0.843f
C26890 col_n[16] a_18938_1126# 0.0785f
C26891 col[16] a_2275_15206# 0.0899f
C26892 vcm a_33390_13214# 0.155f
C26893 col_n[26] a_28978_13174# 0.0765f
C26894 a_2275_11190# a_12914_11166# 0.136f
C26895 col[21] a_2275_4162# 0.0899f
C26896 a_6890_11166# a_7286_11206# 0.0313f
C26897 VDD a_31478_3496# 0.0779f
C26898 m2_18800_18014# a_19030_18194# 0.0249f
C26899 ctop a_12002_7150# 4.11f
C26900 row_n[11] a_4882_13174# 0.0437f
C26901 a_2275_16210# a_35398_16226# 0.145f
C26902 VDD a_20946_12170# 0.181f
C26903 m2_6752_18014# m3_7888_18146# 0.0341f
C26904 rowon_n[15] a_3970_17190# 0.248f
C26905 m2_14208_14426# rowon_n[12] 0.0322f
C26906 m2_20232_10410# rowon_n[8] 0.0322f
C26907 m2_26256_6394# rowon_n[4] 0.0322f
C26908 a_25966_4138# a_26458_4500# 0.0658f
C26909 a_25054_4138# a_25358_4178# 0.0931f
C26910 col_n[26] rowoff_n[0] 0.0471f
C26911 col_n[29] rowoff_n[3] 0.0471f
C26912 col_n[31] rowoff_n[5] 0.0471f
C26913 col_n[28] rowoff_n[2] 0.0471f
C26914 col_n[27] rowoff_n[1] 0.0471f
C26915 row_n[1] a_14922_3134# 0.0437f
C26916 col_n[30] rowoff_n[4] 0.0471f
C26917 col_n[10] a_13406_9520# 0.0283f
C26918 m2_13204_6394# a_13006_6146# 0.165f
C26919 rowon_n[5] a_14010_7150# 0.248f
C26920 vcm a_26970_7150# 0.1f
C26921 rowoff_n[12] a_21038_14178# 0.294f
C26922 a_2475_8178# a_4974_8154# 0.316f
C26923 col_n[12] a_2475_18218# 0.0529f
C26924 vcm a_14314_16226# 0.155f
C26925 a_2275_13198# a_27974_13174# 0.136f
C26926 VDD a_12402_6508# 0.0779f
C26927 row_n[3] a_2966_5142# 0.281f
C26928 col_n[6] a_2475_11190# 0.0531f
C26929 ctop a_27062_11166# 4.11f
C26930 rowon_n[7] a_2275_9182# 1.79f
C26931 a_26970_18194# a_27062_18194# 0.0991f
C26932 a_21950_1126# a_22042_1126# 0.0991f
C26933 m2_9764_946# m3_9896_1078# 3.79f
C26934 vcm a_7894_10162# 0.1f
C26935 a_28066_11166# a_28066_10162# 0.843f
C26936 col_n[8] a_10998_9158# 0.251f
C26937 rowoff_n[15] a_2275_17214# 0.151f
C26938 a_2475_10186# a_20034_10162# 0.316f
C26939 row_n[14] a_25054_16186# 0.282f
C26940 col_n[15] a_17934_11166# 0.0765f
C26941 a_21950_15182# a_22346_15222# 0.0313f
C26942 VDD a_27462_10524# 0.0779f
C26943 ctop a_7986_14178# 4.11f
C26944 row_n[4] a_35094_6146# 0.0123f
C26945 col_n[19] rowoff_n[10] 0.0471f
C26946 rowon_n[8] a_35002_10162# 0.118f
C26947 m2_4168_4386# a_3970_4138# 0.165f
C26948 col_n[3] a_2275_14202# 0.113f
C26949 m2_1732_10986# m2_1732_9982# 0.843f
C26950 rowoff_n[2] a_10394_4500# 0.0133f
C26951 a_6890_7150# a_7382_7512# 0.0658f
C26952 col_n[8] a_2275_3158# 0.113f
C26953 rowoff_n[10] a_27462_12532# 0.0133f
C26954 a_2275_7174# a_10998_7150# 0.399f
C26955 a_5978_7150# a_6282_7190# 0.0931f
C26956 m2_24824_18014# vcm 0.353f
C26957 row_n[6] a_22346_8194# 0.0117f
C26958 vcm a_22954_14178# 0.1f
C26959 a_2475_12194# a_35094_12170# 0.0299f
C26960 a_18026_12170# a_19030_12170# 0.843f
C26961 VDD a_19030_4138# 0.483f
C26962 col[28] a_31078_8154# 0.367f
C26963 VDD a_8386_13536# 0.0779f
C26964 col_n[23] a_2475_13198# 0.0531f
C26965 col_n[28] a_2475_2154# 0.0531f
C26966 row_n[8] a_12914_10162# 0.0437f
C26967 rowoff_n[0] a_19430_2492# 0.0133f
C26968 rowoff_n[7] a_2475_9182# 3.9f
C26969 rowon_n[12] a_12002_14178# 0.248f
C26970 rowoff_n[13] a_8990_15182# 0.294f
C26971 a_2275_9182# a_26058_9158# 0.399f
C26972 sample row_n[14] 0.423f
C26973 vcm row_n[15] 0.616f
C26974 col_n[1] rowon_n[15] 0.111f
C26975 rowon_n[2] a_22042_4138# 0.248f
C26976 col_n[0] rowon_n[14] 0.111f
C26977 VDD rowon_n[13] 3.04f
C26978 col[20] rowoff_n[15] 0.0901f
C26979 col[26] col[27] 0.0355f
C26980 col[13] a_2475_10186# 0.136f
C26981 a_8990_14178# a_8990_13174# 0.843f
C26982 VDD a_34090_8154# 0.483f
C26983 col_n[23] a_26362_8194# 0.084f
C26984 rowoff_n[5] a_10998_7150# 0.294f
C26985 col_n[3] rowoff_n[11] 0.0471f
C26986 a_2275_18218# a_4882_18194# 0.136f
C26987 col_n[4] a_6890_9158# 0.0765f
C26988 VDD a_23446_17552# 0.0779f
C26989 a_31990_2130# a_32386_2170# 0.0313f
C26990 vcm a_5978_2130# 0.56f
C26991 a_2475_6170# a_18938_6146# 0.264f
C26992 a_2275_6170# a_16322_6186# 0.144f
C26993 col_n[20] a_2275_16210# 0.113f
C26994 col_n[25] a_2275_5166# 0.113f
C26995 rowoff_n[3] a_20034_5142# 0.294f
C26996 a_21950_11166# a_22442_11528# 0.0658f
C26997 a_21038_11166# a_21342_11206# 0.0931f
C26998 m2_7180_17438# row_n[15] 0.0128f
C26999 m2_13204_13422# row_n[11] 0.0128f
C27000 m2_19228_9406# row_n[7] 0.0128f
C27001 m2_25252_5390# row_n[3] 0.0128f
C27002 row_n[11] a_33086_13174# 0.282f
C27003 a_33086_16186# a_34090_16186# 0.843f
C27004 VDD a_15014_11166# 0.483f
C27005 rowon_n[15] a_32994_17190# 0.118f
C27006 m2_1732_6970# col[0] 0.0137f
C27007 col[17] a_20034_6146# 0.367f
C27008 col[10] a_2275_13198# 0.0899f
C27009 a_2275_3158# a_9902_3134# 0.136f
C27010 col[15] a_2275_2154# 0.0899f
C27011 rowoff_n[1] a_29070_3134# 0.294f
C27012 col[24] a_26970_8154# 0.0682f
C27013 row_n[13] a_20338_15222# 0.0117f
C27014 vcm a_21038_6146# 0.56f
C27015 rowoff_n[11] a_15414_13536# 0.0133f
C27016 a_17934_8154# a_18026_8154# 0.326f
C27017 a_2475_8178# a_33998_8154# 0.264f
C27018 a_2275_8178# a_31382_8194# 0.144f
C27019 row_n[3] a_30378_5182# 0.0117f
C27020 col[30] a_2475_12194# 0.136f
C27021 row_n[15] a_10906_17190# 0.0437f
C27022 a_2475_17214# a_12002_17190# 0.316f
C27023 VDD a_30074_15182# 0.483f
C27024 col_n[12] a_15318_6186# 0.084f
C27025 col_n[22] a_25358_18234# 0.084f
C27026 m3_19936_18146# a_20034_17190# 0.0303f
C27027 row_n[5] a_20946_7150# 0.0437f
C27028 a_12914_5142# a_13310_5182# 0.0313f
C27029 a_2275_5166# a_24962_5142# 0.136f
C27030 rowon_n[9] a_20034_11166# 0.248f
C27031 vcm a_2475_9182# 1.08f
C27032 rowoff_n[15] a_31478_17552# 0.0133f
C27033 m2_29844_946# a_30074_2130# 0.843f
C27034 a_2275_14202# a_2874_14178# 0.136f
C27035 m2_14784_946# a_2275_1150# 0.28f
C27036 a_2475_14202# a_3878_14178# 0.264f
C27037 m2_34864_17010# ctop 0.0418f
C27038 VDD a_10998_18194# 0.0356f
C27039 a_8990_2130# a_9994_2130# 0.843f
C27040 a_2475_2154# a_17022_2130# 0.316f
C27041 col[27] a_2275_15206# 0.0899f
C27042 m2_9188_1374# VDD 0.0194f
C27043 vcm a_26362_4178# 0.155f
C27044 col[6] a_8990_4138# 0.367f
C27045 rowoff_n[9] a_21950_11166# 0.202f
C27046 col[16] a_19030_16186# 0.367f
C27047 vcm a_17022_13174# 0.56f
C27048 col[13] a_15926_6146# 0.0682f
C27049 a_32994_12170# a_33086_12170# 0.326f
C27050 VDD a_13918_3134# 0.181f
C27051 m2_5748_18014# a_6282_18234# 0.087f
C27052 m2_15788_18014# a_2275_18218# 0.28f
C27053 col[23] a_25966_18194# 0.0682f
C27054 a_2275_16210# a_18026_16186# 0.399f
C27055 VDD a_2275_12194# 1.95f
C27056 rowon_n[3] a_7894_5142# 0.118f
C27057 col_n[31] a_34090_12170# 0.251f
C27058 row_n[9] rowoff_n[8] 0.085f
C27059 col_n[28] a_30986_2130# 0.0765f
C27060 col_n[2] a_2275_1150# 0.113f
C27061 rowoff_n[7] a_30986_9158# 0.202f
C27062 a_34090_5142# a_34090_4138# 0.843f
C27063 a_2475_4162# a_32082_4138# 0.316f
C27064 col_n[1] a_4274_4178# 0.084f
C27065 col_n[23] a_2475_18218# 0.0529f
C27066 col_n[11] a_14314_16226# 0.084f
C27067 vcm a_7286_7190# 0.155f
C27068 a_27974_9158# a_28370_9198# 0.0313f
C27069 rowoff_n[12] a_2966_14178# 0.294f
C27070 m2_3164_1374# VDD 0.0194f
C27071 row_n[10] a_28370_12210# 0.0117f
C27072 col_n[17] a_2475_11190# 0.0531f
C27073 ctop a_20034_2130# 4.07f
C27074 vcm a_32082_17190# 0.56f
C27075 a_2475_13198# a_10906_13174# 0.264f
C27076 a_2275_13198# a_8290_13214# 0.144f
C27077 VDD a_28978_7150# 0.181f
C27078 a_2275_18218# a_33086_18194# 0.0924f
C27079 a_17934_18194# a_18426_18556# 0.0658f
C27080 m2_11772_18014# a_2475_18218# 0.286f
C27081 col_n[22] a_25454_10524# 0.0283f
C27082 a_2275_1150# a_23046_1126# 0.0924f
C27083 row_n[12] a_18938_14178# 0.0437f
C27084 a_12914_1126# a_13406_1488# 0.0658f
C27085 vcm a_35002_2130# 0.101f
C27086 a_24050_6146# a_25054_6146# 0.843f
C27087 col[7] a_2475_8178# 0.136f
C27088 col_n[0] a_3366_4500# 0.0283f
C27089 vcm a_22346_11206# 0.155f
C27090 row_n[2] a_28978_4138# 0.0437f
C27091 a_2475_10186# a_1957_10186# 0.0734f
C27092 VDD a_20434_1488# 0.0913f
C27093 rowon_n[6] a_28066_8154# 0.248f
C27094 m2_27260_17438# a_27062_17190# 0.165f
C27095 col[5] a_7986_14178# 0.367f
C27096 col[2] a_4882_4138# 0.0682f
C27097 a_2475_15206# a_25966_15182# 0.264f
C27098 a_13918_15182# a_14010_15182# 0.326f
C27099 a_2275_15206# a_23350_15222# 0.144f
C27100 col_n[30] rowoff_n[10] 0.0471f
C27101 VDD a_9902_10162# 0.181f
C27102 col[12] a_14922_16186# 0.0682f
C27103 col_n[14] a_2275_14202# 0.113f
C27104 col_n[19] a_2275_3158# 0.113f
C27105 col_n[20] a_23046_10162# 0.251f
C27106 a_2475_18218# a_31078_18194# 0.0299f
C27107 vcm a_15926_5142# 0.1f
C27108 rowoff_n[10] a_9902_12170# 0.202f
C27109 col_n[27] a_29982_12170# 0.0765f
C27110 a_15014_8154# a_15014_7150# 0.843f
C27111 a_29070_1126# vcm 0.165f
C27112 row_n[6] a_5978_8154# 0.282f
C27113 m2_3164_12418# rowon_n[10] 0.0322f
C27114 m2_9188_8402# rowon_n[6] 0.0322f
C27115 vcm a_3270_14218# 0.155f
C27116 a_8898_12170# a_9294_12210# 0.0313f
C27117 a_2275_12194# a_16930_12170# 0.136f
C27118 m2_15212_4386# rowon_n[2] 0.0322f
C27119 VDD a_35494_5504# 0.106f
C27120 rowon_n[10] a_5886_12170# 0.118f
C27121 col[4] a_2275_11190# 0.0899f
C27122 m2_28840_18014# VDD 0.993f
C27123 ctop a_16018_9158# 4.11f
C27124 VDD a_24962_14178# 0.181f
C27125 rowon_n[0] a_15926_2130# 0.118f
C27126 col_n[11] a_14410_8516# 0.0283f
C27127 a_27974_5142# a_28466_5504# 0.0658f
C27128 a_27062_5142# a_27366_5182# 0.0931f
C27129 col_n[4] rowon_n[11] 0.111f
C27130 vcm rowon_n[9] 0.65f
C27131 sample rowon_n[8] 0.0935f
C27132 col_n[12] rowon_n[15] 0.111f
C27133 col_n[1] row_n[10] 0.298f
C27134 col_n[5] row_n[12] 0.298f
C27135 col_n[9] row_n[14] 0.298f
C27136 col_n[0] row_n[9] 0.298f
C27137 col_n[7] row_n[13] 0.298f
C27138 col_n[11] row_n[15] 0.298f
C27139 col_n[3] row_n[11] 0.298f
C27140 VDD row_n[8] 3.29f
C27141 col_n[10] rowon_n[14] 0.111f
C27142 col_n[6] rowon_n[12] 0.111f
C27143 col_n[2] rowon_n[10] 0.111f
C27144 col_n[8] rowon_n[13] 0.111f
C27145 col[24] a_2475_10186# 0.136f
C27146 col[31] rowoff_n[15] 0.0901f
C27147 vcm a_30986_9158# 0.1f
C27148 m2_13780_18014# m2_14208_18442# 0.165f
C27149 a_4974_9158# a_5978_9158# 0.843f
C27150 rowoff_n[14] a_25966_16186# 0.202f
C27151 a_2475_9182# a_8990_9158# 0.316f
C27152 m2_18224_15430# a_18026_15182# 0.165f
C27153 vcm a_18330_18234# 0.16f
C27154 col_n[14] rowoff_n[11] 0.0471f
C27155 m3_4876_1078# a_3970_1126# 0.0341f
C27156 m2_24248_17438# rowon_n[15] 0.0322f
C27157 a_2275_14202# a_31990_14178# 0.136f
C27158 m2_30272_13422# rowon_n[11] 0.0322f
C27159 VDD a_16418_8516# 0.0779f
C27160 m2_35292_9406# rowon_n[7] 0.0322f
C27161 sample a_2161_14202# 0.0858f
C27162 ctop a_31078_13174# 4.11f
C27163 VDD a_5886_17190# 0.181f
C27164 col_n[31] a_2275_16210# 0.113f
C27165 a_23958_2130# a_24050_2130# 0.326f
C27166 row_n[9] a_26970_11166# 0.0437f
C27167 col_n[9] a_12002_8154# 0.251f
C27168 rowon_n[13] a_26058_15182# 0.248f
C27169 vcm a_11910_12170# 0.1f
C27170 rowoff_n[3] a_1957_5166# 0.0219f
C27171 a_30074_12170# a_30074_11166# 0.843f
C27172 a_2475_11190# a_24050_11166# 0.316f
C27173 VDD a_7986_2130# 0.483f
C27174 col_n[16] a_18938_10162# 0.0765f
C27175 m2_24824_18014# a_25358_18234# 0.087f
C27176 col[21] a_2275_13198# 0.0899f
C27177 a_23958_16186# a_24354_16226# 0.0313f
C27178 VDD a_31478_12532# 0.0779f
C27179 m2_21812_18014# m3_20940_18146# 0.0341f
C27180 col[26] a_2275_2154# 0.0899f
C27181 ctop a_12002_16186# 4.11f
C27182 rowoff_n[1] a_11398_3496# 0.0133f
C27183 row_n[13] a_3970_15182# 0.282f
C27184 vcm a_2966_6146# 0.56f
C27185 a_8898_8154# a_9390_8516# 0.0658f
C27186 a_2275_8178# a_15014_8154# 0.399f
C27187 a_7986_8154# a_8290_8194# 0.0931f
C27188 m2_9188_13422# a_8990_13174# 0.165f
C27189 col_n[10] a_13406_18556# 0.0283f
C27190 sample rowoff_n[12] 0.0775f
C27191 vcm a_26970_16186# 0.1f
C27192 a_20034_13174# a_21038_13174# 0.843f
C27193 VDD a_23046_6146# 0.483f
C27194 col[29] a_32082_7150# 0.367f
C27195 row_n[3] a_14010_5142# 0.282f
C27196 rowon_n[7] a_13918_9158# 0.118f
C27197 VDD a_12402_15544# 0.0779f
C27198 rowoff_n[6] a_2874_8154# 0.202f
C27199 m2_15788_946# col[13] 0.425f
C27200 col_n[11] a_2475_9182# 0.0531f
C27201 a_2275_5166# a_5278_5182# 0.144f
C27202 a_3878_5142# a_4274_5182# 0.0313f
C27203 row_n[5] a_2275_7174# 19.2f
C27204 a_2475_5166# a_7894_5142# 0.264f
C27205 a_4882_5142# a_4974_5142# 0.326f
C27206 m2_24824_946# m3_25960_1078# 0.0341f
C27207 m2_28264_9406# a_28066_9158# 0.165f
C27208 rowon_n[9] a_1957_11190# 0.0172f
C27209 a_2275_10186# a_30074_10162# 0.399f
C27210 rowoff_n[15] a_13918_17190# 0.202f
C27211 row_n[14] a_35398_16226# 0.0117f
C27212 col_n[24] a_27366_7190# 0.084f
C27213 rowoff_n[4] a_12002_6146# 0.294f
C27214 a_10998_15182# a_10998_14178# 0.843f
C27215 VDD a_3970_9158# 0.483f
C27216 col_n[5] a_7894_8154# 0.0765f
C27217 col[1] a_2475_6170# 0.136f
C27218 a_31990_1126# col_n[29] 0.0775f
C27219 m2_2160_11414# row_n[9] 0.0194f
C27220 m2_8184_7398# row_n[5] 0.0128f
C27221 m2_14208_3382# row_n[1] 0.0128f
C27222 vcm a_9994_4138# 0.56f
C27223 rowoff_n[2] a_21038_4138# 0.294f
C27224 a_2275_7174# a_20338_7190# 0.144f
C27225 a_2475_7174# a_22954_7150# 0.264f
C27226 rowoff_n[9] a_3878_11166# 0.202f
C27227 m2_8760_18014# col[6] 0.347f
C27228 row_n[6] a_35002_8154# 0.0437f
C27229 a_23046_12170# a_23350_12210# 0.0931f
C27230 col_n[8] a_2275_12194# 0.113f
C27231 a_23958_12170# a_24450_12532# 0.0658f
C27232 rowon_n[10] a_34090_12170# 0.248f
C27233 row_n[5] rowoff_n[5] 0.209f
C27234 col_n[13] a_2275_1150# 0.113f
C27235 VDD a_19030_13174# 0.483f
C27236 col[18] a_21038_5142# 0.367f
C27237 rowoff_n[0] a_30074_2130# 0.294f
C27238 col[28] a_31078_17190# 0.367f
C27239 col[25] a_27974_7150# 0.0682f
C27240 a_2275_4162# a_13918_4138# 0.136f
C27241 col_n[28] a_2475_11190# 0.0531f
C27242 m3_34996_14130# ctop 0.209f
C27243 m2_19228_7398# a_19030_7150# 0.165f
C27244 col_n[0] a_3270_1166# 0.0839f
C27245 m2_23244_16434# row_n[14] 0.0128f
C27246 vcm a_25054_8154# 0.56f
C27247 m2_29268_12418# row_n[10] 0.0128f
C27248 m2_34864_7974# row_n[6] 0.267f
C27249 a_19942_9158# a_20034_9158# 0.326f
C27250 a_2275_9182# a_2275_8178# 0.0715f
C27251 row_n[10] a_12002_12170# 0.282f
C27252 rowon_n[14] a_11910_16186# 0.118f
C27253 col_n[13] a_16322_5182# 0.084f
C27254 VDD a_34090_17190# 0.484f
C27255 col_n[23] a_26362_17230# 0.084f
C27256 row_n[0] a_22042_2130# 0.282f
C27257 col[18] a_2475_8178# 0.136f
C27258 a_2475_1150# a_5978_1126# 0.0299f
C27259 a_3878_1126# a_4370_1488# 0.0667f
C27260 rowon_n[4] a_21950_6146# 0.118f
C27261 col_n[4] a_6890_18194# 0.0762f
C27262 vcm a_15318_2170# 0.155f
C27263 a_14922_6146# a_15318_6186# 0.0313f
C27264 a_2275_6170# a_28978_6146# 0.136f
C27265 m2_4744_946# m2_5748_946# 0.843f
C27266 row_n[2] a_9294_4178# 0.0117f
C27267 vcm a_5978_11166# 0.56f
C27268 row_n[11] rowoff_n[10] 0.085f
C27269 VDD a_2161_1150# 0.23f
C27270 col_n[25] a_2275_14202# 0.113f
C27271 a_2275_15206# a_6982_15182# 0.399f
C27272 a_4882_15182# a_5374_15544# 0.0658f
C27273 a_3970_15182# a_4274_15222# 0.0931f
C27274 col_n[30] a_2275_3158# 0.113f
C27275 m2_24824_18014# col_n[22] 0.243f
C27276 m2_34864_16006# m3_34996_17142# 0.0341f
C27277 a_2475_3158# a_21038_3134# 0.316f
C27278 col[7] a_9994_3134# 0.367f
C27279 a_10998_3134# a_12002_3134# 0.843f
C27280 rowoff_n[8] a_22954_10162# 0.202f
C27281 m2_10192_5390# a_9994_5142# 0.165f
C27282 a_32386_1166# a_2275_1150# 0.145f
C27283 row_n[13] a_32994_15182# 0.0437f
C27284 col[17] a_20034_15182# 0.367f
C27285 vcm a_30378_6186# 0.155f
C27286 col[14] a_16930_5142# 0.0682f
C27287 rowoff_n[11] a_26058_13174# 0.294f
C27288 col[15] a_2275_11190# 0.0899f
C27289 col[24] a_26970_17190# 0.0682f
C27290 vcm a_21038_15182# 0.56f
C27291 a_34090_13174# a_34394_13214# 0.0931f
C27292 a_35002_13174# a_35094_13174# 0.0991f
C27293 VDD a_17934_5142# 0.181f
C27294 a_31078_1126# VDD 0.035f
C27295 a_2275_17214# a_22042_17190# 0.399f
C27296 rowoff_n[6] a_31990_8154# 0.202f
C27297 col_n[12] row_n[10] 0.298f
C27298 col_n[3] rowon_n[5] 0.111f
C27299 col_n[27] col_n[28] 0.0102f
C27300 col_n[22] row_n[15] 0.298f
C27301 col_n[17] rowon_n[12] 0.111f
C27302 col_n[11] rowon_n[9] 0.111f
C27303 col_n[16] row_n[12] 0.298f
C27304 sample row_n[3] 0.423f
C27305 col_n[2] a_5278_3174# 0.084f
C27306 col_n[2] row_n[5] 0.298f
C27307 VDD rowon_n[2] 3.04f
C27308 col_n[20] row_n[14] 0.298f
C27309 col_n[15] rowon_n[11] 0.111f
C27310 col_n[14] row_n[11] 0.298f
C27311 col_n[10] row_n[9] 0.298f
C27312 col_n[19] rowon_n[13] 0.111f
C27313 col_n[6] row_n[7] 0.298f
C27314 col_n[9] rowon_n[8] 0.111f
C27315 col_n[23] rowon_n[15] 0.111f
C27316 col_n[18] row_n[13] 0.298f
C27317 vcm row_n[4] 0.616f
C27318 col_n[21] rowon_n[14] 0.111f
C27319 col_n[7] rowon_n[7] 0.111f
C27320 col_n[0] rowon_n[3] 0.111f
C27321 col_n[13] rowon_n[10] 0.111f
C27322 col_n[4] row_n[6] 0.298f
C27323 col_n[8] row_n[8] 0.298f
C27324 col_n[1] rowon_n[4] 0.111f
C27325 col_n[5] rowon_n[6] 0.111f
C27326 col_n[12] a_15318_15222# 0.084f
C27327 a_2475_5166# a_2475_4162# 0.0666f
C27328 m3_25960_1078# m3_26964_1078# 0.202f
C27329 col_n[25] rowoff_n[11] 0.0471f
C27330 vcm a_11302_9198# 0.155f
C27331 a_29982_10162# a_30378_10202# 0.0313f
C27332 ctop a_24050_4138# 4.11f
C27333 m2_13780_946# a_14010_1126# 0.0249f
C27334 a_2475_14202# a_14922_14178# 0.264f
C27335 a_2275_14202# a_12306_14218# 0.144f
C27336 VDD a_32994_9158# 0.181f
C27337 row_n[7] a_20034_9158# 0.282f
C27338 col_n[23] a_26458_9520# 0.0283f
C27339 col_n[5] a_2475_7174# 0.0531f
C27340 rowon_n[11] a_19942_13174# 0.118f
C27341 VDD a_20338_18234# 0.019f
C27342 a_14922_2130# a_15414_2492# 0.0658f
C27343 a_2275_2154# a_27062_2130# 0.399f
C27344 a_14010_2130# a_14314_2170# 0.0931f
C27345 m2_32280_1374# VDD 0.0194f
C27346 vcm a_4882_3134# 0.1f
C27347 row_n[9] a_7286_11206# 0.0117f
C27348 rowoff_n[9] a_32482_11528# 0.0133f
C27349 rowon_n[1] a_29982_3134# 0.118f
C27350 a_26058_7150# a_27062_7150# 0.843f
C27351 col[6] a_8990_13174# 0.367f
C27352 vcm a_26362_13214# 0.155f
C27353 a_2275_11190# a_5886_11166# 0.136f
C27354 col[3] a_5886_3134# 0.0682f
C27355 VDD a_24450_3496# 0.0779f
C27356 m2_34864_11990# VDD 0.766f
C27357 col[13] a_15926_15182# 0.0682f
C27358 ctop a_4974_7150# 4.11f
C27359 a_2275_16210# a_27366_16226# 0.144f
C27360 a_15926_16186# a_16018_16186# 0.326f
C27361 a_2475_16210# a_29982_16186# 0.264f
C27362 VDD a_13918_12170# 0.181f
C27363 col_n[21] a_24050_9158# 0.251f
C27364 m2_3164_2378# rowon_n[0] 0.0322f
C27365 col_n[9] rowoff_n[12] 0.0471f
C27366 col_n[2] a_2275_10186# 0.113f
C27367 row_n[1] a_7894_3134# 0.0437f
C27368 col_n[28] a_30986_11166# 0.0765f
C27369 rowon_n[5] a_6982_7150# 0.248f
C27370 m2_34864_16006# m2_35292_16434# 0.165f
C27371 vcm a_19942_7150# 0.1f
C27372 col_n[1] a_4274_13214# 0.084f
C27373 a_17022_9158# a_17022_8154# 0.843f
C27374 rowoff_n[12] a_14010_14178# 0.294f
C27375 sample a_1957_3158# 0.345f
C27376 vcm a_7286_16226# 0.155f
C27377 a_2275_13198# a_20946_13174# 0.136f
C27378 a_10906_13174# a_11302_13214# 0.0313f
C27379 VDD a_5374_6508# 0.0779f
C27380 ctop a_20034_11166# 4.11f
C27381 col_n[22] a_2475_9182# 0.0531f
C27382 VDD a_28978_16186# 0.181f
C27383 col_n[12] a_15414_7512# 0.0283f
C27384 m2_13204_15430# rowon_n[13] 0.0322f
C27385 a_29982_6146# a_30474_6508# 0.0658f
C27386 a_29070_6146# a_29374_6186# 0.0931f
C27387 m2_19228_11414# rowon_n[9] 0.0322f
C27388 m2_25252_7398# rowon_n[5] 0.0322f
C27389 m2_31276_3382# rowon_n[1] 0.0322f
C27390 vcm a_35002_11166# 0.101f
C27391 a_2475_10186# a_13006_10162# 0.316f
C27392 col[7] a_2475_17214# 0.136f
C27393 a_6982_10162# a_7986_10162# 0.843f
C27394 row_n[14] a_18026_16186# 0.282f
C27395 m2_34864_17010# a_35398_17230# 0.087f
C27396 col_n[0] a_3366_13536# 0.0283f
C27397 col[12] a_2475_6170# 0.136f
C27398 a_2275_15206# a_34394_15222# 0.144f
C27399 VDD a_20434_10524# 0.0779f
C27400 m2_34864_12994# m3_34996_14130# 0.0341f
C27401 col[2] a_4882_13174# 0.0682f
C27402 row_n[4] a_28066_6146# 0.282f
C27403 a_25966_3134# a_26058_3134# 0.326f
C27404 rowon_n[8] a_27974_10162# 0.118f
C27405 col_n[10] a_13006_7150# 0.251f
C27406 col_n[19] a_2275_12194# 0.113f
C27407 rowoff_n[10] a_20434_12532# 0.0133f
C27408 rowoff_n[2] a_2966_4138# 0.294f
C27409 a_2275_7174# a_3970_7150# 0.399f
C27410 rowon_n[1] rowoff_n[1] 20.2f
C27411 ctop rowoff_n[7] 0.177f
C27412 m2_10768_18014# vcm 0.353f
C27413 col_n[24] a_2275_1150# 0.113f
C27414 col_n[17] a_19942_9158# 0.0765f
C27415 row_n[6] a_15318_8194# 0.0117f
C27416 vcm a_15926_14178# 0.1f
C27417 a_2475_12194# a_28066_12170# 0.316f
C27418 a_32082_13174# a_32082_12170# 0.843f
C27419 VDD a_12002_4138# 0.483f
C27420 a_25966_17190# a_26362_17230# 0.0313f
C27421 VDD a_35494_14540# 0.106f
C27422 row_n[8] a_5886_10162# 0.0437f
C27423 rowoff_n[0] a_12402_2492# 0.0133f
C27424 col[9] a_2275_9182# 0.0899f
C27425 rowon_n[12] a_4974_14178# 0.248f
C27426 col_n[1] a_4370_5504# 0.0283f
C27427 m2_20808_946# ctop 0.043f
C27428 col_n[11] a_14410_17552# 0.0283f
C27429 rowoff_n[13] a_2475_15206# 3.9f
C27430 a_9994_9158# a_10298_9198# 0.0931f
C27431 a_2275_9182# a_19030_9158# 0.399f
C27432 a_10906_9158# a_11398_9520# 0.0658f
C27433 col[30] a_33086_6146# 0.367f
C27434 rowon_n[2] a_15014_4138# 0.248f
C27435 vcm a_30986_18194# 0.101f
C27436 a_22042_14178# a_23046_14178# 0.843f
C27437 col[29] a_2475_8178# 0.136f
C27438 VDD a_27062_8154# 0.483f
C27439 rowoff_n[5] a_3970_7150# 0.294f
C27440 VDD a_16418_17552# 0.0779f
C27441 rowon_n[4] a_3878_6146# 0.118f
C27442 vcm a_33086_3134# 0.56f
C27443 a_2475_6170# a_11910_6146# 0.264f
C27444 a_2275_6170# a_9294_6186# 0.144f
C27445 a_6890_6146# a_6982_6146# 0.326f
C27446 col_n[25] a_28370_6186# 0.084f
C27447 col_n[0] a_2475_5166# 0.0532f
C27448 rowoff_n[3] a_13006_5142# 0.294f
C27449 a_2275_11190# a_34090_11166# 0.399f
C27450 col_n[9] a_12002_17190# 0.251f
C27451 col_n[6] a_8898_7150# 0.0765f
C27452 a_13006_16186# a_13006_15182# 0.843f
C27453 row_n[11] a_26058_13174# 0.282f
C27454 VDD a_7986_11166# 0.483f
C27455 m2_1732_17010# m3_1864_17142# 3.79f
C27456 rowon_n[15] a_25966_17190# 0.118f
C27457 a_2161_3158# a_2275_3158# 0.183f
C27458 a_2475_3158# a_2966_3134# 0.317f
C27459 col[26] a_2275_11190# 0.0899f
C27460 rowoff_n[1] a_22042_3134# 0.294f
C27461 row_n[13] a_13310_15222# 0.0117f
C27462 vcm a_14010_6146# 0.56f
C27463 a_2275_8178# a_24354_8194# 0.144f
C27464 a_2475_8178# a_26970_8154# 0.264f
C27465 rowoff_n[11] a_8386_13536# 0.0133f
C27466 vcm a_2966_15182# 0.56f
C27467 a_25966_13174# a_26458_13536# 0.0658f
C27468 a_25054_13174# a_25358_13214# 0.0931f
C27469 row_n[3] a_23350_5182# 0.0117f
C27470 col_n[13] row_n[5] 0.298f
C27471 col_n[7] row_n[2] 0.298f
C27472 col_n[3] row_n[0] 0.298f
C27473 col_n[22] rowon_n[9] 0.111f
C27474 col_n[8] rowon_n[2] 0.111f
C27475 col_n[25] row_n[11] 0.298f
C27476 col_n[29] row_n[13] 0.298f
C27477 col_n[15] row_n[6] 0.298f
C27478 col_n[21] row_n[9] 0.298f
C27479 col_n[11] row_n[4] 0.298f
C27480 col_n[19] row_n[8] 0.298f
C27481 col_n[6] rowon_n[1] 0.111f
C27482 col_n[23] row_n[10] 0.298f
C27483 col_n[24] rowon_n[10] 0.111f
C27484 col_n[16] rowon_n[6] 0.111f
C27485 col_n[20] rowon_n[8] 0.111f
C27486 col_n[28] rowon_n[12] 0.111f
C27487 col_n[30] rowon_n[13] 0.111f
C27488 col_n[17] row_n[7] 0.298f
C27489 col_n[27] row_n[12] 0.298f
C27490 col_n[9] row_n[3] 0.298f
C27491 col_n[12] rowon_n[4] 0.111f
C27492 col[19] a_22042_4138# 0.367f
C27493 col_n[14] rowon_n[5] 0.111f
C27494 VDD en_bit_n[2] 0.206f
C27495 vcm ctop 0.81f
C27496 col_n[31] row_n[14] 0.298f
C27497 rowon_n[15] rowon_n[14] 0.0632f
C27498 col_n[18] rowon_n[7] 0.111f
C27499 col_n[4] rowon_n[0] 0.111f
C27500 col_n[26] rowon_n[11] 0.111f
C27501 col_n[10] rowon_n[3] 0.111f
C27502 col_n[5] row_n[1] 0.298f
C27503 m2_12200_14426# row_n[12] 0.0128f
C27504 a_2475_17214# a_4974_17190# 0.316f
C27505 m2_18224_10410# row_n[8] 0.0128f
C27506 VDD a_23046_15182# 0.483f
C27507 col[29] a_32082_16186# 0.367f
C27508 m2_24248_6394# row_n[4] 0.0128f
C27509 col[26] a_28978_6146# 0.0682f
C27510 a_2275_5166# a_17934_5142# 0.136f
C27511 row_n[5] a_13918_7150# 0.0437f
C27512 m3_34996_7102# m3_34996_6098# 0.202f
C27513 m2_1732_7974# a_2161_8178# 0.0454f
C27514 rowon_n[9] a_13006_11166# 0.248f
C27515 vcm a_29070_10162# 0.56f
C27516 rowoff_n[15] a_24450_17552# 0.0133f
C27517 a_21950_10162# a_22042_10162# 0.326f
C27518 col_n[16] a_2475_7174# 0.0531f
C27519 m2_24248_16434# a_24050_16186# 0.165f
C27520 col_n[14] a_17326_4178# 0.084f
C27521 row_n[7] a_1957_9182# 0.187f
C27522 m2_34864_9982# m3_34996_11118# 0.0341f
C27523 col_n[24] a_27366_16226# 0.084f
C27524 VDD a_3970_18194# 0.0356f
C27525 col_n[5] a_7894_17190# 0.0765f
C27526 a_2475_2154# a_9994_2130# 0.316f
C27527 a_23046_3134# a_23046_2130# 0.843f
C27528 col[1] a_2475_15206# 0.136f
C27529 m2_1732_2954# rowoff_n[1] 0.415f
C27530 vcm a_19334_4178# 0.155f
C27531 col[6] a_2475_4162# 0.136f
C27532 a_16930_7150# a_17326_7190# 0.0313f
C27533 rowoff_n[9] a_14922_11166# 0.202f
C27534 a_2275_7174# a_32994_7150# 0.136f
C27535 m2_34864_10986# a_2475_11190# 0.282f
C27536 vcm a_9994_13174# 0.56f
C27537 VDD a_6890_3134# 0.181f
C27538 m2_1732_18014# a_2275_18218# 0.191f
C27539 a_2275_16210# a_10998_16186# 0.399f
C27540 a_5978_16186# a_6282_16226# 0.0931f
C27541 a_6890_16186# a_7382_16548# 0.0658f
C27542 m2_25828_946# col[23] 0.425f
C27543 col_n[20] rowoff_n[12] 0.0471f
C27544 col_n[13] a_2275_10186# 0.113f
C27545 col[8] a_10998_2130# 0.367f
C27546 row_n[8] a_34090_10162# 0.282f
C27547 rowoff_n[7] a_23958_9158# 0.202f
C27548 col[18] a_21038_14178# 0.367f
C27549 rowon_n[12] a_33998_14178# 0.118f
C27550 a_13006_4138# a_14010_4138# 0.843f
C27551 a_2475_4162# a_25054_4138# 0.316f
C27552 m3_18932_1078# ctop 0.266f
C27553 col[15] a_17934_4138# 0.0682f
C27554 vcm a_35398_8194# 0.161f
C27555 col[25] a_27974_16186# 0.0682f
C27556 rowoff_n[13] a_30986_15182# 0.202f
C27557 m2_15212_14426# a_15014_14178# 0.165f
C27558 row_n[10] a_21342_12210# 0.0117f
C27559 col_n[0] a_3270_10202# 0.084f
C27560 ctop a_13006_2130# 4.06f
C27561 vcm a_25054_17190# 0.56f
C27562 VDD a_21950_7150# 0.181f
C27563 col[3] a_2275_7174# 0.0899f
C27564 rowoff_n[5] a_32994_7150# 0.202f
C27565 col_n[3] a_6282_2170# 0.084f
C27566 a_2275_18218# a_26058_18194# 0.0924f
C27567 row_n[0] a_31382_2170# 0.0117f
C27568 a_2275_1150# a_16018_1126# 0.0924f
C27569 row_n[12] a_11910_14178# 0.0437f
C27570 col_n[13] a_16322_14218# 0.084f
C27571 m2_12200_2378# a_12002_2130# 0.165f
C27572 vcm a_27974_2130# 0.1f
C27573 col[18] a_2475_17214# 0.136f
C27574 a_3970_6146# a_3970_5142# 0.843f
C27575 m2_15788_946# m2_16216_1374# 0.165f
C27576 col[23] a_2475_6170# 0.136f
C27577 m2_34288_10410# a_34090_10162# 0.165f
C27578 vcm a_15318_11206# 0.155f
C27579 row_n[2] a_21950_4138# 0.0437f
C27580 a_31990_11166# a_32386_11206# 0.0313f
C27581 VDD a_13406_1488# 0.0977f
C27582 rowon_n[6] a_21038_8154# 0.248f
C27583 col_n[24] a_27462_8516# 0.0283f
C27584 ctop a_28066_6146# 4.11f
C27585 a_2475_15206# a_18938_15182# 0.264f
C27586 a_2275_15206# a_16322_15222# 0.144f
C27587 col_n[4] rowoff_n[13] 0.0471f
C27588 VDD a_2161_10186# 0.187f
C27589 m2_1732_13998# m3_1864_14130# 3.79f
C27590 rowon_n[0] m2_35292_2378# 0.0322f
C27591 col_n[30] a_2275_12194# 0.113f
C27592 col[0] rowoff_n[2] 0.0901f
C27593 col[7] rowoff_n[9] 0.0901f
C27594 col[6] rowoff_n[8] 0.0901f
C27595 col[2] rowoff_n[4] 0.0901f
C27596 a_2275_3158# a_31078_3134# 0.399f
C27597 col[1] rowoff_n[3] 0.0901f
C27598 col[5] rowoff_n[7] 0.0901f
C27599 a_16018_3134# a_16322_3174# 0.0931f
C27600 a_16930_3134# a_17422_3496# 0.0658f
C27601 col[4] rowoff_n[6] 0.0901f
C27602 col[3] rowoff_n[5] 0.0901f
C27603 a_2475_18218# a_24050_18194# 0.0299f
C27604 rowoff_n[8] a_33486_10524# 0.0133f
C27605 a_23350_1166# a_22954_1126# 0.0313f
C27606 vcm a_8898_5142# 0.1f
C27607 a_28066_8154# a_29070_8154# 0.843f
C27608 col[7] a_9994_12170# 0.367f
C27609 rowoff_n[10] a_2161_12194# 0.0226f
C27610 m2_6176_12418# a_5978_12170# 0.165f
C27611 col[4] a_6890_2130# 0.0682f
C27612 vcm a_30378_15222# 0.155f
C27613 a_2275_12194# a_9902_12170# 0.136f
C27614 col[14] a_16930_14178# 0.0682f
C27615 VDD a_28466_5504# 0.0779f
C27616 m2_14784_18014# VDD 1.1f
C27617 ctop a_8990_9158# 4.11f
C27618 col[20] a_2275_9182# 0.0899f
C27619 row_n[15] a_32082_17190# 0.282f
C27620 a_17934_17190# a_18026_17190# 0.326f
C27621 a_2475_17214# a_33998_17190# 0.264f
C27622 col_n[22] a_25054_8154# 0.251f
C27623 a_2275_17214# a_31382_17230# 0.144f
C27624 VDD a_17934_14178# 0.181f
C27625 col_n[29] a_31990_10162# 0.0765f
C27626 rowon_n[0] a_8898_2130# 0.118f
C27627 col_n[2] a_5278_12210# 0.084f
C27628 m2_25252_8402# a_25054_8154# 0.165f
C27629 vcm a_23958_9158# 0.1f
C27630 m2_6752_18014# m2_7180_18442# 0.165f
C27631 rowoff_n[14] a_18938_16186# 0.202f
C27632 a_19030_10162# a_19030_9158# 0.843f
C27633 vcm a_11302_18234# 0.16f
C27634 a_12914_14178# a_13310_14218# 0.0313f
C27635 m2_21812_946# a_21950_1126# 0.225f
C27636 a_2275_14202# a_24962_14178# 0.136f
C27637 row_n[7] a_29374_9198# 0.0117f
C27638 m2_2160_13422# rowon_n[11] 0.0219f
C27639 VDD a_9390_8516# 0.0779f
C27640 m2_34864_6970# m3_34996_8106# 0.0341f
C27641 m2_8184_9406# rowon_n[7] 0.0322f
C27642 col_n[13] a_16418_6508# 0.0283f
C27643 m2_14208_5390# rowon_n[3] 0.0322f
C27644 m2_12776_946# vcm 0.353f
C27645 ctop a_24050_13174# 4.11f
C27646 col_n[23] a_26458_18556# 0.0283f
C27647 VDD a_32994_18194# 0.343f
C27648 col_n[5] a_2475_16210# 0.0531f
C27649 col_n[10] a_2475_5166# 0.0531f
C27650 row_n[9] a_19942_11166# 0.0437f
C27651 a_31990_7150# a_32482_7512# 0.0658f
C27652 a_31078_7150# a_31382_7190# 0.0931f
C27653 m2_34864_12994# vcm 0.408f
C27654 rowon_n[13] a_19030_15182# 0.248f
C27655 vcm a_4882_12170# 0.1f
C27656 a_8990_11166# a_9994_11166# 0.843f
C27657 a_2475_11190# a_17022_11166# 0.316f
C27658 col[3] a_5886_12170# 0.0682f
C27659 rowon_n[3] a_29070_5142# 0.248f
C27660 VDD a_24450_12532# 0.0779f
C27661 m2_11772_18014# m3_12908_18146# 0.0341f
C27662 col[0] a_2475_2154# 0.148f
C27663 ctop a_4974_16186# 4.11f
C27664 m2_29268_14426# rowon_n[12] 0.0322f
C27665 m2_34864_9982# rowon_n[8] 0.231f
C27666 col_n[11] a_14010_6146# 0.251f
C27667 a_27974_4138# a_28066_4138# 0.326f
C27668 rowoff_n[1] a_4370_3496# 0.0133f
C27669 m2_16216_6394# a_16018_6146# 0.165f
C27670 col_n[18] a_20946_8154# 0.0765f
C27671 a_2275_8178# a_7986_8154# 0.399f
C27672 col_n[15] rowon_n[0] 0.111f
C27673 rowon_n[12] row_n[12] 18.9f
C27674 col_n[23] rowon_n[4] 0.111f
C27675 vcm col[5] 5.46f
C27676 col_n[28] row_n[7] 0.298f
C27677 col_n[27] rowon_n[6] 0.111f
C27678 col_n[29] rowon_n[7] 0.111f
C27679 col_n[11] ctop 0.0594f
C27680 col_n[16] row_n[1] 0.298f
C27681 col_n[30] row_n[8] 0.298f
C27682 VDD col[8] 3.83f
C27683 col_n[20] row_n[3] 0.298f
C27684 col_n[17] rowon_n[1] 0.111f
C27685 col_n[25] rowon_n[5] 0.111f
C27686 col_n[26] row_n[6] 0.298f
C27687 col_n[22] row_n[4] 0.298f
C27688 col_n[21] rowon_n[3] 0.111f
C27689 col_n[24] row_n[5] 0.298f
C27690 col_n[19] rowon_n[2] 0.111f
C27691 col_n[14] row_n[0] 0.298f
C27692 col_n[31] rowon_n[8] 0.111f
C27693 col_n[18] row_n[2] 0.298f
C27694 col_n[2] col[3] 7.13f
C27695 vcm a_19942_16186# 0.1f
C27696 col_n[7] a_2275_8178# 0.113f
C27697 a_2475_13198# a_32082_13174# 0.316f
C27698 a_34090_14178# a_34090_13174# 0.843f
C27699 VDD a_16018_6146# 0.483f
C27700 row_n[3] a_6982_5142# 0.282f
C27701 sample a_1957_12194# 0.345f
C27702 rowon_n[7] a_6890_9158# 0.118f
C27703 a_27974_18194# a_28370_18234# 0.0313f
C27704 VDD a_5374_15544# 0.0779f
C27705 col_n[2] a_5374_4500# 0.0283f
C27706 vcm a_22042_1126# 0.165f
C27707 col_n[12] a_15414_16548# 0.0283f
C27708 col_n[27] a_2475_7174# 0.0531f
C27709 m3_21944_18146# m3_22948_18146# 0.202f
C27710 m2_14784_946# m3_14916_1078# 3.79f
C27711 col[31] a_34090_5142# 0.367f
C27712 a_12914_10162# a_13406_10524# 0.0658f
C27713 a_2275_10186# a_23046_10162# 0.399f
C27714 a_12002_10162# a_12306_10202# 0.0931f
C27715 rowoff_n[15] a_6890_17190# 0.202f
C27716 row_n[14] a_27366_16226# 0.0117f
C27717 rowoff_n[4] a_4974_6146# 0.294f
C27718 a_24050_15182# a_25054_15182# 0.843f
C27719 m2_12776_946# a_13006_2130# 0.843f
C27720 VDD a_31078_10162# 0.483f
C27721 m2_1732_10986# m3_1864_11118# 3.79f
C27722 col[12] a_2475_15206# 0.136f
C27723 col[17] a_2475_4162# 0.136f
C27724 m2_7180_4386# a_6982_4138# 0.165f
C27725 col_n[26] a_29374_5182# 0.084f
C27726 vcm a_2874_4138# 0.1f
C27727 a_8898_7150# a_8990_7150# 0.326f
C27728 rowoff_n[10] a_31078_12170# 0.294f
C27729 rowoff_n[2] a_14010_4138# 0.294f
C27730 a_2475_7174# a_15926_7150# 0.264f
C27731 a_2275_7174# a_13310_7190# 0.144f
C27732 col_n[10] a_13006_16186# 0.251f
C27733 row_n[6] a_27974_8154# 0.0437f
C27734 col_n[7] a_9902_6146# 0.0765f
C27735 m2_1732_3958# sample 0.2f
C27736 rowon_n[10] a_27062_12170# 0.248f
C27737 col_n[17] a_19942_18194# 0.0762f
C27738 col_n[31] rowoff_n[12] 0.0471f
C27739 col_n[24] a_2275_10186# 0.113f
C27740 m2_1732_15002# VDD 0.856f
C27741 m3_1864_6098# a_2966_6146# 0.0302f
C27742 a_15014_17190# a_15014_16186# 0.843f
C27743 VDD a_12002_13174# 0.483f
C27744 rowoff_n[0] a_23046_2130# 0.294f
C27745 a_2275_4162# a_6890_4138# 0.136f
C27746 m3_14916_18146# ctop 0.209f
C27747 col[9] a_2275_18218# 0.0899f
C27748 m2_1732_11990# row_n[10] 0.292f
C27749 vcm a_18026_8154# 0.56f
C27750 a_2275_9182# a_28370_9198# 0.144f
C27751 a_2475_9182# a_30986_9158# 0.264f
C27752 m2_7180_8402# row_n[6] 0.0128f
C27753 col_n[1] a_4370_14540# 0.0283f
C27754 col[14] a_2275_7174# 0.0899f
C27755 m2_13204_4386# row_n[2] 0.0128f
C27756 row_n[10] a_4974_12170# 0.282f
C27757 col[20] a_23046_3134# 0.367f
C27758 a_27974_14178# a_28466_14540# 0.0658f
C27759 a_27062_14178# a_27366_14218# 0.0931f
C27760 rowon_n[14] a_4882_16186# 0.118f
C27761 VDD a_3878_7150# 0.181f
C27762 m2_34864_3958# m3_34996_5094# 0.0341f
C27763 col[30] a_33086_15182# 0.367f
C27764 col[27] a_29982_5142# 0.0682f
C27765 col[29] a_2475_17214# 0.136f
C27766 VDD a_27062_17190# 0.484f
C27767 row_n[0] a_15014_2130# 0.282f
C27768 a_33998_2130# a_34394_2170# 0.0313f
C27769 rowon_n[4] a_14922_6146# 0.118f
C27770 vcm a_8290_2170# 0.155f
C27771 a_2275_6170# a_21950_6146# 0.136f
C27772 vcm a_33086_12170# 0.56f
C27773 row_n[2] a_3878_4138# 0.0437f
C27774 col_n[15] a_18330_3174# 0.084f
C27775 col_n[15] rowoff_n[13] 0.0471f
C27776 a_23958_11166# a_24050_11166# 0.326f
C27777 VDD a_29982_2130# 0.181f
C27778 m2_22240_17438# row_n[15] 0.0128f
C27779 m2_28264_13422# row_n[11] 0.0128f
C27780 rowon_n[6] a_2966_8154# 0.248f
C27781 col_n[0] a_2475_14202# 0.0532f
C27782 col_n[25] a_28370_15222# 0.084f
C27783 m2_34288_9406# row_n[7] 0.0128f
C27784 col_n[4] a_2475_3158# 0.0531f
C27785 col[16] rowoff_n[7] 0.0901f
C27786 col[12] rowoff_n[3] 0.0901f
C27787 col[11] rowoff_n[2] 0.0901f
C27788 col[9] rowoff_n[0] 0.0901f
C27789 col[17] rowoff_n[8] 0.0901f
C27790 col[18] rowoff_n[9] 0.0901f
C27791 col[10] rowoff_n[1] 0.0901f
C27792 col[15] rowoff_n[6] 0.0901f
C27793 col[13] rowoff_n[4] 0.0901f
C27794 col[14] rowoff_n[5] 0.0901f
C27795 col_n[6] a_8898_16186# 0.0765f
C27796 a_2475_3158# a_14010_3134# 0.316f
C27797 a_25054_4138# a_25054_3134# 0.843f
C27798 rowoff_n[8] a_15926_10162# 0.202f
C27799 a_27974_1126# a_2475_1150# 0.264f
C27800 a_25358_1166# a_2275_1150# 0.145f
C27801 row_n[13] a_25966_15182# 0.0437f
C27802 vcm a_23350_6186# 0.155f
C27803 rowoff_n[11] a_19030_13174# 0.294f
C27804 a_18938_8154# a_19334_8194# 0.0313f
C27805 col[31] a_2275_9182# 0.0899f
C27806 vcm a_14010_15182# 0.56f
C27807 VDD a_10906_5142# 0.181f
C27808 row_n[3] a_34394_5182# 0.0117f
C27809 a_24050_1126# VDD 0.035f
C27810 rowon_n[7] a_35094_9158# 0.0141f
C27811 a_7986_17190# a_8290_17230# 0.0931f
C27812 a_2275_17214# a_15014_17190# 0.399f
C27813 a_8898_17190# a_9390_17552# 0.0658f
C27814 rowoff_n[6] a_24962_8154# 0.202f
C27815 col[19] a_22042_13174# 0.367f
C27816 col[16] a_18938_3134# 0.0682f
C27817 m3_22948_18146# a_23046_17190# 0.0303f
C27818 m2_1732_1950# m2_2160_2378# 0.165f
C27819 col_n[1] a_2275_6170# 0.113f
C27820 a_2475_5166# a_29070_5142# 0.316f
C27821 a_15014_5142# a_16018_5142# 0.843f
C27822 col[26] a_28978_15182# 0.0682f
C27823 m3_11904_1078# m3_12908_1078# 0.202f
C27824 col_n[0] rowoff_n[14] 0.0471f
C27825 vcm a_4274_9198# 0.155f
C27826 rowoff_n[15] a_35094_17190# 0.0135f
C27827 rowoff_n[4] a_33998_6146# 0.202f
C27828 ctop a_17022_4138# 4.11f
C27829 m2_23820_946# a_2275_1150# 0.28f
C27830 col[2] rowoff_n[10] 0.0901f
C27831 a_4882_14178# a_4974_14178# 0.326f
C27832 a_3878_14178# a_4274_14218# 0.0313f
C27833 a_2275_14202# a_5278_14218# 0.144f
C27834 a_2475_14202# a_7894_14178# 0.264f
C27835 col_n[16] a_2475_16210# 0.0531f
C27836 row_n[7] a_13006_9158# 0.282f
C27837 col_n[4] a_7286_1166# 0.0839f
C27838 VDD a_25966_9158# 0.181f
C27839 m2_1732_7974# m3_1864_8106# 3.79f
C27840 col_n[21] a_2475_5166# 0.0531f
C27841 col_n[14] a_17326_13214# 0.084f
C27842 rowon_n[11] a_12914_13174# 0.118f
C27843 VDD a_13310_18234# 0.019f
C27844 a_2275_2154# a_20034_2130# 0.399f
C27845 m2_16792_946# VDD 1f
C27846 vcm a_31990_4138# 0.1f
C27847 rowoff_n[9] a_25454_11528# 0.0133f
C27848 a_5978_7150# a_5978_6146# 0.843f
C27849 rowon_n[1] a_22954_3134# 0.118f
C27850 col_n[25] a_28466_7512# 0.0283f
C27851 col[6] a_2475_13198# 0.136f
C27852 vcm a_19334_13214# 0.155f
C27853 VDD a_17422_3496# 0.0779f
C27854 col[11] a_2475_2154# 0.136f
C27855 m2_9764_18014# a_9902_18194# 0.225f
C27856 ctop a_32082_8154# 4.11f
C27857 a_2475_16210# a_22954_16186# 0.264f
C27858 a_2275_16210# a_20338_16226# 0.144f
C27859 VDD a_6890_12170# 0.181f
C27860 rowoff_n[7] a_34490_9520# 0.0133f
C27861 a_2275_4162# a_35094_4138# 0.0924f
C27862 a_18026_4138# a_18330_4178# 0.0931f
C27863 a_18938_4138# a_19430_4500# 0.0658f
C27864 col_n[27] row_n[1] 0.298f
C27865 VDD col[19] 3.83f
C27866 col[8] a_10998_11166# 0.367f
C27867 col_n[28] rowon_n[1] 0.111f
C27868 vcm col[16] 5.46f
C27869 col_n[29] row_n[2] 0.298f
C27870 col_n[26] rowon_n[0] 0.111f
C27871 col_n[8] col[8] 0.489f
C27872 col_n[22] ctop 0.0594f
C27873 col_n[25] row_n[0] 0.298f
C27874 col_n[30] rowon_n[2] 0.111f
C27875 col_n[31] row_n[3] 0.298f
C27876 m2_1732_5966# a_2475_6170# 0.139f
C27877 col[5] a_7894_1126# 0.0682f
C27878 col_n[18] a_2275_8178# 0.113f
C27879 vcm a_12914_7150# 0.1f
C27880 rowoff_n[12] a_6982_14178# 0.294f
C27881 a_30074_9158# a_31078_9158# 0.843f
C27882 col[15] a_17934_13174# 0.0682f
C27883 row_n[10] a_33998_12170# 0.0437f
C27884 vcm a_35398_17230# 0.161f
C27885 rowon_n[14] a_33086_16186# 0.248f
C27886 a_2275_13198# a_13918_13174# 0.136f
C27887 col_n[23] a_26058_7150# 0.251f
C27888 VDD a_32482_7512# 0.0779f
C27889 ctop a_13006_11166# 4.11f
C27890 a_2275_18218# a_2275_17214# 0.0715f
C27891 a_19942_18194# a_20034_18194# 0.0991f
C27892 col_n[30] a_32994_9158# 0.0765f
C27893 VDD a_21950_16186# 0.181f
C27894 col[3] a_2275_16210# 0.0899f
C27895 a_14922_1126# a_15014_1126# 0.0991f
C27896 col[8] a_2275_5166# 0.0899f
C27897 col_n[3] a_6282_11206# 0.084f
C27898 m2_34864_5966# m2_34864_4962# 0.843f
C27899 m2_3164_3382# rowon_n[1] 0.0322f
C27900 m2_27836_946# m2_28840_946# 0.843f
C27901 vcm a_27974_11166# 0.1f
C27902 a_21038_11166# a_21038_10162# 0.843f
C27903 a_3878_10162# a_4370_10524# 0.0658f
C27904 a_2966_10162# a_3270_10202# 0.0931f
C27905 a_2475_10186# a_5978_10162# 0.316f
C27906 row_n[14] a_10998_16186# 0.282f
C27907 m2_30272_17438# a_30074_17190# 0.165f
C27908 col[23] a_2475_15206# 0.136f
C27909 col_n[14] a_17422_5504# 0.0283f
C27910 col[28] a_2475_4162# 0.136f
C27911 a_14922_15182# a_15318_15222# 0.0313f
C27912 a_2275_15206# a_28978_15182# 0.136f
C27913 VDD a_13406_10524# 0.0779f
C27914 col_n[24] a_27462_17552# 0.0283f
C27915 ctop a_28066_15182# 4.11f
C27916 row_n[4] a_21038_6146# 0.282f
C27917 rowon_n[8] a_20946_10162# 0.118f
C27918 rowoff_n[10] a_13406_12532# 0.0133f
C27919 a_33086_8154# a_33390_8194# 0.0931f
C27920 a_33998_8154# a_34490_8516# 0.0658f
C27921 a_31382_1166# vcm 0.16f
C27922 m2_12200_16434# rowon_n[14] 0.0322f
C27923 m2_18224_12418# rowon_n[10] 0.0322f
C27924 row_n[6] a_8290_8194# 0.0117f
C27925 vcm a_8898_14178# 0.1f
C27926 m2_24248_8402# rowon_n[6] 0.0322f
C27927 a_10998_12170# a_12002_12170# 0.843f
C27928 a_2475_12194# a_21038_12170# 0.316f
C27929 m2_30272_4386# rowon_n[2] 0.0322f
C27930 VDD a_4974_4138# 0.483f
C27931 col[4] a_6890_11166# 0.0682f
C27932 VDD a_28466_14540# 0.0779f
C27933 col_n[12] a_15014_5142# 0.251f
C27934 col[20] a_2275_18218# 0.0899f
C27935 col_n[22] a_25054_17190# 0.251f
C27936 rowoff_n[0] a_5374_2492# 0.0133f
C27937 col[25] a_2275_7174# 0.0899f
C27938 col_n[19] a_21950_7150# 0.0765f
C27939 a_29982_5142# a_30074_5142# 0.326f
C27940 rowoff_n[14] a_29470_16548# 0.0133f
C27941 a_2275_9182# a_12002_9158# 0.399f
C27942 m2_21236_15430# a_21038_15182# 0.165f
C27943 rowon_n[2] a_7986_4138# 0.248f
C27944 col_n[0] a_2966_11166# 0.251f
C27945 vcm a_23958_18194# 0.101f
C27946 a_2475_14202# a_2475_13198# 0.0666f
C27947 VDD a_20034_8154# 0.483f
C27948 m2_1732_4962# m3_1864_5094# 3.79f
C27949 col_n[3] a_6378_3496# 0.0283f
C27950 VDD a_9390_17552# 0.0779f
C27951 a_24962_2130# a_25358_2170# 0.0313f
C27952 col_n[13] a_16418_15544# 0.0283f
C27953 m3_13912_1078# VDD 0.0157f
C27954 vcm a_26058_3134# 0.56f
C27955 col_n[26] rowoff_n[13] 0.0471f
C27956 a_2475_6170# a_4882_6146# 0.264f
C27957 a_2275_6170# a_3878_6146# 0.136f
C27958 a_2874_6146# a_3366_6508# 0.0658f
C27959 col_n[10] a_2475_14202# 0.0531f
C27960 rowoff_n[3] a_5978_5142# 0.294f
C27961 a_14922_11166# a_15414_11528# 0.0658f
C27962 a_14010_11166# a_14314_11206# 0.0931f
C27963 col_n[15] a_2475_3158# 0.0531f
C27964 a_2275_11190# a_27062_11166# 0.399f
C27965 col[26] rowoff_n[6] 0.0901f
C27966 col[25] rowoff_n[5] 0.0901f
C27967 col[21] rowoff_n[1] 0.0901f
C27968 col[27] rowoff_n[7] 0.0901f
C27969 col[20] rowoff_n[0] 0.0901f
C27970 col[29] rowoff_n[9] 0.0901f
C27971 col[28] rowoff_n[8] 0.0901f
C27972 col[24] rowoff_n[4] 0.0901f
C27973 col[22] rowoff_n[2] 0.0901f
C27974 col[23] rowoff_n[3] 0.0901f
C27975 m2_28840_18014# a_28978_18194# 0.225f
C27976 m2_5748_18014# a_5978_17190# 0.843f
C27977 row_n[11] a_19030_13174# 0.282f
C27978 a_26058_16186# a_27062_16186# 0.843f
C27979 m2_26832_18014# m3_25960_18146# 0.0341f
C27980 col[6] a_2475_18218# 0.136f
C27981 rowon_n[15] a_18938_17190# 0.118f
C27982 col_n[27] a_30378_4178# 0.084f
C27983 col[0] a_2475_11190# 0.148f
C27984 col_n[1] a_3970_3134# 0.251f
C27985 rowoff_n[1] a_15014_3134# 0.294f
C27986 row_n[1] a_29070_3134# 0.282f
C27987 row_n[13] a_6282_15222# 0.0117f
C27988 col_n[11] a_14010_15182# 0.251f
C27989 vcm a_6982_6146# 0.56f
C27990 rowon_n[5] a_28978_7150# 0.118f
C27991 a_2275_8178# a_17326_8194# 0.144f
C27992 a_2475_8178# a_19942_8154# 0.264f
C27993 col_n[8] a_10906_5142# 0.0765f
C27994 a_10906_8154# a_10998_8154# 0.326f
C27995 m2_12200_13422# a_12002_13174# 0.165f
C27996 col_n[18] a_20946_17190# 0.0765f
C27997 row_n[3] a_16322_5182# 0.0117f
C27998 col_n[7] a_2275_17214# 0.113f
C27999 VDD a_16018_15182# 0.483f
C28000 col_n[12] a_2275_6170# 0.113f
C28001 m2_2160_2378# row_n[0] 0.0194f
C28002 col_n[10] rowoff_n[14] 0.0471f
C28003 a_2275_5166# a_10906_5142# 0.136f
C28004 row_n[5] a_6890_7150# 0.0437f
C28005 a_5886_5142# a_6282_5182# 0.0313f
C28006 col_n[2] a_5374_13536# 0.0283f
C28007 m2_29844_946# m3_30980_1078# 0.0341f
C28008 m3_34996_14130# m3_34996_13126# 0.202f
C28009 m2_31276_9406# a_31078_9158# 0.165f
C28010 rowon_n[9] a_5978_11166# 0.248f
C28011 col[13] rowoff_n[10] 0.0901f
C28012 vcm a_22042_10162# 0.56f
C28013 col[21] a_24050_2130# 0.367f
C28014 a_2475_10186# a_35002_10162# 0.264f
C28015 rowoff_n[15] a_17422_17552# 0.0133f
C28016 col_n[27] a_2475_16210# 0.0531f
C28017 a_2275_10186# a_32386_10202# 0.144f
C28018 col[31] a_34090_14178# 0.367f
C28019 a_29070_15182# a_29374_15222# 0.0931f
C28020 col[2] a_2275_3158# 0.0899f
C28021 a_29982_15182# a_30474_15544# 0.0658f
C28022 col[28] a_30986_4138# 0.0682f
C28023 m2_24824_18014# ctop 0.0422f
C28024 a_1957_2154# a_2275_2154# 0.158f
C28025 a_2475_2154# a_2874_2130# 0.264f
C28026 m2_11196_15430# row_n[13] 0.0128f
C28027 m2_17220_11414# row_n[9] 0.0128f
C28028 m2_23244_7398# row_n[5] 0.0128f
C28029 m2_29268_3382# row_n[1] 0.0128f
C28030 col[17] a_2475_13198# 0.136f
C28031 vcm a_12306_4178# 0.155f
C28032 a_2275_7174# a_25966_7150# 0.136f
C28033 rowoff_n[9] a_7894_11166# 0.202f
C28034 col[22] a_2475_2154# 0.136f
C28035 m2_1732_16006# vcm 0.316f
C28036 col_n[16] a_19334_2170# 0.0839f
C28037 vcm a_2874_13174# 0.1f
C28038 col_n[26] a_29374_14218# 0.084f
C28039 a_25966_12170# a_26058_12170# 0.326f
C28040 VDD a_33998_4138# 0.181f
C28041 col_n[7] a_9902_15182# 0.0765f
C28042 a_2275_16210# a_3970_16186# 0.399f
C28043 row_n[15] ctop 0.183f
C28044 vcm col[27] 5.46f
C28045 VDD col[30] 3.84f
C28046 col_n[13] col[14] 7.13f
C28047 row_n[8] a_27062_10162# 0.282f
C28048 col_n[29] a_2275_8178# 0.113f
C28049 rowoff_n[7] a_16930_9158# 0.202f
C28050 rowon_n[12] a_26970_14178# 0.118f
C28051 a_2475_4162# a_18026_4138# 0.316f
C28052 a_27062_5142# a_27062_4138# 0.843f
C28053 m3_1864_6098# ctop 0.21f
C28054 m2_22240_7398# a_22042_7150# 0.165f
C28055 vcm a_27366_8194# 0.155f
C28056 rowoff_n[13] a_23958_15182# 0.202f
C28057 a_20946_9158# a_21342_9198# 0.0313f
C28058 row_n[10] a_14314_12210# 0.0117f
C28059 ctop a_5978_2130# 4.06f
C28060 vcm a_18026_17190# 0.56f
C28061 col[14] a_2275_16210# 0.0899f
C28062 VDD a_14922_7150# 0.181f
C28063 m2_34864_2954# m3_34996_2082# 0.0341f
C28064 m2_1732_1950# m3_1864_2082# 3.79f
C28065 rowoff_n[5] a_25966_7150# 0.202f
C28066 col[19] a_2275_5166# 0.0899f
C28067 col[20] a_23046_12170# 0.367f
C28068 a_2275_18218# a_19030_18194# 0.0924f
C28069 a_10906_18194# a_11398_18556# 0.0658f
C28070 row_n[0] a_24354_2170# 0.0117f
C28071 col[17] a_19942_2130# 0.0682f
C28072 VDD a_3878_16186# 0.181f
C28073 row_n[12] a_4882_14178# 0.0437f
C28074 a_5886_1126# a_6378_1488# 0.0658f
C28075 a_2275_1150# a_8990_1126# 0.0924f
C28076 col[27] a_29982_14178# 0.0682f
C28077 vcm a_20946_2130# 0.1f
C28078 a_17022_6146# a_18026_6146# 0.843f
C28079 a_2475_6170# a_33086_6146# 0.316f
C28080 m2_8760_946# m2_9188_1374# 0.165f
C28081 rowoff_n[3] a_35002_5142# 0.202f
C28082 row_n[2] a_14922_4138# 0.0437f
C28083 vcm a_8290_11206# 0.155f
C28084 VDD a_6378_1488# 0.0977f
C28085 m2_24824_18014# a_25054_17190# 0.843f
C28086 rowon_n[6] a_14010_8154# 0.248f
C28087 ctop a_21038_6146# 4.11f
C28088 m2_9764_946# col[7] 0.425f
C28089 col_n[15] a_18330_12210# 0.084f
C28090 a_6890_15182# a_6982_15182# 0.326f
C28091 a_2475_15206# a_11910_15182# 0.264f
C28092 a_2275_15206# a_9294_15222# 0.144f
C28093 VDD a_29982_11166# 0.181f
C28094 row_n[4] a_2966_6146# 0.281f
C28095 col_n[4] a_2475_12194# 0.0531f
C28096 a_2275_3158# a_24050_3134# 0.399f
C28097 a_2475_18218# a_17022_18194# 0.0299f
C28098 rowon_n[8] a_2275_10186# 1.79f
C28099 rowoff_n[8] a_26458_10524# 0.0133f
C28100 col_n[9] a_2475_1150# 0.0531f
C28101 m2_13204_5390# a_13006_5142# 0.165f
C28102 col_n[26] a_29470_6508# 0.0283f
C28103 vcm a_34394_6186# 0.155f
C28104 a_7986_8154# a_7986_7150# 0.843f
C28105 vcm a_23350_15222# 0.155f
C28106 a_2475_12194# a_2966_12170# 0.317f
C28107 a_2161_12194# a_2275_12194# 0.183f
C28108 VDD a_21438_5504# 0.0779f
C28109 col[31] a_2275_18218# 0.0899f
C28110 a_35398_1166# VDD 0.0988f
C28111 ctop a_2475_9182# 0.0488f
C28112 row_n[15] a_25054_17190# 0.282f
C28113 a_2475_17214# a_26970_17190# 0.264f
C28114 a_2275_17214# a_24354_17230# 0.144f
C28115 VDD a_10906_14178# 0.181f
C28116 rowoff_n[6] a_35494_8516# 0.0133f
C28117 m2_2736_18014# col[0] 0.347f
C28118 col[9] a_12002_10162# 0.367f
C28119 a_20034_5142# a_20338_5182# 0.0931f
C28120 a_20946_5142# a_21438_5504# 0.0658f
C28121 row_n[5] a_35094_7150# 0.0123f
C28122 col[16] a_18938_12170# 0.0682f
C28123 rowon_n[9] a_35002_11166# 0.118f
C28124 vcm a_16930_9158# 0.1f
C28125 rowoff_n[14] a_11910_16186# 0.202f
C28126 col_n[1] a_2275_15206# 0.113f
C28127 a_32082_10162# a_33086_10162# 0.843f
C28128 col_n[24] a_27062_6146# 0.251f
C28129 col_n[6] a_2275_4162# 0.113f
C28130 vcm a_4274_18234# 0.16f
C28131 a_2275_14202# a_17934_14178# 0.136f
C28132 row_n[7] a_22346_9198# 0.0117f
C28133 VDD a_1957_8178# 0.196f
C28134 col_n[31] a_33998_8154# 0.0765f
C28135 ctop a_17022_13174# 4.11f
C28136 VDD a_25966_18194# 0.343f
C28137 col_n[4] a_7286_10202# 0.084f
C28138 row_n[13] rowoff_n[13] 0.209f
C28139 a_16930_2130# a_17022_2130# 0.326f
C28140 col[0] a_2966_8154# 0.367f
C28141 a_2275_2154# a_29374_2170# 0.144f
C28142 a_2475_2154# a_31990_2130# 0.264f
C28143 col_n[21] a_2475_14202# 0.0531f
C28144 m2_4168_3382# a_3970_3134# 0.165f
C28145 m3_9896_18146# VDD 0.0312f
C28146 row_n[9] a_12914_11166# 0.0437f
C28147 col_n[26] a_2475_3158# 0.0531f
C28148 sample_n rowoff_n[1] 0.14f
C28149 col[31] rowoff_n[0] 0.0901f
C28150 en_bit_n[1] a_2275_1150# 0.0364f
C28151 rowon_n[13] a_12002_15182# 0.248f
C28152 vcm a_31990_13174# 0.1f
C28153 col_n[15] a_18426_4500# 0.0283f
C28154 a_2475_11190# a_9994_11166# 0.316f
C28155 a_23046_12170# a_23046_11166# 0.843f
C28156 col[17] a_2475_18218# 0.136f
C28157 VDD a_28066_3134# 0.483f
C28158 col_n[25] a_28466_16548# 0.0283f
C28159 a_2275_16210# a_32994_16186# 0.136f
C28160 a_16930_16186# a_17326_16226# 0.0313f
C28161 rowon_n[3] a_22042_5142# 0.248f
C28162 VDD a_17422_12532# 0.0779f
C28163 m2_2736_18014# m3_2868_18146# 3.79f
C28164 col[11] a_2475_11190# 0.136f
C28165 m2_1732_13998# rowon_n[12] 0.236f
C28166 ctop a_32082_17190# 4.06f
C28167 m2_7180_10410# rowon_n[8] 0.0322f
C28168 m2_13204_6394# rowon_n[4] 0.0322f
C28169 m2_18224_2378# rowon_n[0] 0.0322f
C28170 col_n[18] a_2275_17214# 0.113f
C28171 m2_18800_18014# col_n[16] 0.243f
C28172 col[5] a_7894_10162# 0.0682f
C28173 vcm a_12914_16186# 0.1f
C28174 a_2475_13198# a_25054_13174# 0.316f
C28175 a_13006_13174# a_14010_13174# 0.843f
C28176 VDD a_8990_6146# 0.483f
C28177 col_n[23] a_2275_6170# 0.113f
C28178 col_n[13] a_16018_4138# 0.251f
C28179 col_n[21] rowoff_n[14] 0.0471f
C28180 col_n[23] a_26058_16186# 0.251f
C28181 VDD a_32482_16548# 0.0779f
C28182 row_n[12] a_33086_14178# 0.282f
C28183 col_n[20] a_22954_6146# 0.0765f
C28184 col_n[30] a_32994_18194# 0.0762f
C28185 col[24] rowoff_n[10] 0.0901f
C28186 vcm a_15014_1126# 0.165f
C28187 m2_28264_15430# rowon_n[13] 0.0322f
C28188 m2_34288_11414# rowon_n[9] 0.0322f
C28189 a_31990_6146# a_32082_6146# 0.326f
C28190 col[8] a_2275_14202# 0.0899f
C28191 m2_5748_946# m3_4876_1078# 0.0341f
C28192 m3_7888_18146# m3_8892_18146# 0.202f
C28193 col[13] a_2275_3158# 0.0899f
C28194 a_2275_10186# a_16018_10162# 0.399f
C28195 rowoff_n[0] VSS 0.63f
C28196 rowoff_n[1] VSS 0.631f
C28197 rowoff_n[2] VSS 0.63f
C28198 rowoff_n[3] VSS 0.63f
C28199 rowoff_n[4] VSS 0.63f
C28200 rowoff_n[5] VSS 0.63f
C28201 rowoff_n[6] VSS 0.63f
C28202 rowoff_n[7] VSS 0.63f
C28203 rowoff_n[8] VSS 0.63f
C28204 rowoff_n[9] VSS 0.63f
C28205 rowoff_n[10] VSS 0.631f
C28206 rowoff_n[11] VSS 0.63f
C28207 rowoff_n[12] VSS 0.63f
C28208 rowoff_n[13] VSS 0.63f
C28209 rowoff_n[14] VSS 0.631f
C28210 rowoff_n[15] VSS 0.714f
C28211 sample_n VSS 11.2f
C28212 col[31] VSS 6.05f
C28213 col[30] VSS 5.99f
C28214 col[29] VSS 6.01f
C28215 col[28] VSS 6.02f
C28216 col[27] VSS 6.02f
C28217 col[26] VSS 6.03f
C28218 col[25] VSS 5.98f
C28219 col[24] VSS 6.02f
C28220 col[23] VSS 6.02f
C28221 col[22] VSS 6.02f
C28222 col[21] VSS 6.02f
C28223 col[20] VSS 6.02f
C28224 col[19] VSS 6.02f
C28225 col[18] VSS 6.02f
C28226 col[17] VSS 5.97f
C28227 col[16] VSS 5.97f
C28228 col[15] VSS 5.97f
C28229 col[14] VSS 6.02f
C28230 col[13] VSS 6.02f
C28231 col[12] VSS 6.02f
C28232 col[11] VSS 6.02f
C28233 col[10] VSS 6.02f
C28234 col[9] VSS 6.02f
C28235 col[8] VSS 6.02f
C28236 col[7] VSS 6.02f
C28237 col[6] VSS 6.02f
C28238 col[5] VSS 6.02f
C28239 col[4] VSS 6.02f
C28240 col[3] VSS 6.02f
C28241 col[2] VSS 6.02f
C28242 col[1] VSS 5.97f
C28243 col[0] VSS 6.18f
C28244 analog_in VSS 0.55f
C28245 en_bit_n[0] VSS 1.01f
C28246 en_bit_n[2] VSS 1f
C28247 en_bit_n[1] VSS 1.01f
C28248 en_C0_n VSS 1.01f
C28249 ctop VSS 19.7f
C28250 sw_n VSS 0.647f
C28251 sw VSS 0.653f
C28252 row_n[0] VSS 7.05f
C28253 rowon_n[0] VSS 5.53f
C28254 row_n[1] VSS 6.98f
C28255 rowon_n[1] VSS 5.47f
C28256 row_n[2] VSS 6.97f
C28257 rowon_n[2] VSS 5.47f
C28258 row_n[3] VSS 6.97f
C28259 rowon_n[3] VSS 5.47f
C28260 row_n[4] VSS 6.97f
C28261 rowon_n[4] VSS 5.47f
C28262 row_n[5] VSS 6.97f
C28263 rowon_n[5] VSS 5.47f
C28264 row_n[6] VSS 6.98f
C28265 rowon_n[6] VSS 5.47f
C28266 row_n[7] VSS 6.97f
C28267 rowon_n[7] VSS 5.47f
C28268 row_n[8] VSS 6.97f
C28269 rowon_n[8] VSS 5.47f
C28270 row_n[9] VSS 6.97f
C28271 rowon_n[9] VSS 5.47f
C28272 row_n[10] VSS 6.98f
C28273 rowon_n[10] VSS 5.47f
C28274 row_n[11] VSS 6.97f
C28275 rowon_n[11] VSS 5.47f
C28276 row_n[12] VSS 6.97f
C28277 rowon_n[12] VSS 5.47f
C28278 row_n[13] VSS 6.97f
C28279 rowon_n[13] VSS 5.47f
C28280 row_n[14] VSS 6.98f
C28281 rowon_n[14] VSS 5.47f
C28282 row_n[15] VSS 6.98f
C28283 rowon_n[15] VSS 5.48f
C28284 col_n[31] VSS 17.1f
C28285 col_n[30] VSS 10.2f
C28286 col_n[29] VSS 10.2f
C28287 col_n[28] VSS 10.3f
C28288 col_n[27] VSS 10.2f
C28289 col_n[26] VSS 10.3f
C28290 col_n[25] VSS 10.2f
C28291 col_n[24] VSS 10f
C28292 col_n[23] VSS 10f
C28293 col_n[22] VSS 10f
C28294 col_n[21] VSS 10f
C28295 col_n[20] VSS 10f
C28296 col_n[19] VSS 10f
C28297 col_n[18] VSS 10f
C28298 col_n[17] VSS 9.62f
C28299 col_n[16] VSS 9.62f
C28300 col_n[15] VSS 9.62f
C28301 col_n[14] VSS 10f
C28302 col_n[13] VSS 10f
C28303 col_n[12] VSS 10f
C28304 col_n[11] VSS 10f
C28305 col_n[10] VSS 10f
C28306 col_n[9] VSS 10f
C28307 col_n[8] VSS 10f
C28308 col_n[7] VSS 10f
C28309 col_n[6] VSS 10f
C28310 col_n[5] VSS 10f
C28311 col_n[4] VSS 10f
C28312 col_n[3] VSS 10f
C28313 col_n[2] VSS 10f
C28314 col_n[1] VSS 9.62f
C28315 vcm VSS 0.444p
C28316 col_n[0] VSS 10f
C28317 sample VSS 15.1f
C28318 VDD VSS 6.19p
C28319 m3_34996_1078# VSS 0.351f
C28320 m3_34568_1078# VSS 0.0609f
C28321 m3_33992_1078# VSS 0.0536f
C28322 m3_32988_1078# VSS 0.155f
C28323 m3_31984_1078# VSS 0.159f
C28324 m3_30980_1078# VSS 0.159f
C28325 m3_29976_1078# VSS 0.159f
C28326 m3_28972_1078# VSS 0.159f
C28327 m3_27968_1078# VSS 0.159f
C28328 m3_26964_1078# VSS 0.162f
C28329 m3_25960_1078# VSS 0.162f
C28330 m3_24956_1078# VSS 0.162f
C28331 m3_23952_1078# VSS 0.162f
C28332 m3_22948_1078# VSS 0.162f
C28333 m3_21944_1078# VSS 0.162f
C28334 m3_20940_1078# VSS 0.162f
C28335 m3_19936_1078# VSS 0.155f
C28336 m3_18932_1078# VSS 0.147f
C28337 m3_17928_1078# VSS 0.151f
C28338 m3_16924_1078# VSS 0.162f
C28339 m3_15920_1078# VSS 0.162f
C28340 m3_14916_1078# VSS 0.162f
C28341 m3_13912_1078# VSS 0.162f
C28342 m3_12908_1078# VSS 0.162f
C28343 m3_11904_1078# VSS 0.162f
C28344 m3_10900_1078# VSS 0.162f
C28345 m3_9896_1078# VSS 0.162f
C28346 m3_8892_1078# VSS 0.162f
C28347 m3_7888_1078# VSS 0.162f
C28348 m3_6884_1078# VSS 0.162f
C28349 m3_5880_1078# VSS 0.162f
C28350 m3_4876_1078# VSS 0.162f
C28351 m3_3872_1078# VSS 0.155f
C28352 m3_2868_1078# VSS 0.161f
C28353 m3_1864_1078# VSS 0.336f
C28354 m3_34996_2082# VSS 0.201f
C28355 m3_2868_2082# VSS 0.0181f
C28356 m3_1864_2082# VSS 0.191f
C28357 m3_34996_3086# VSS 0.201f
C28358 m3_1864_3086# VSS 0.191f
C28359 m3_34996_4090# VSS 0.201f
C28360 m3_1864_4090# VSS 0.191f
C28361 m3_34996_5094# VSS 0.201f
C28362 m3_1864_5094# VSS 0.191f
C28363 m3_34996_6098# VSS 0.201f
C28364 m3_1864_6098# VSS 0.191f
C28365 m3_34996_7102# VSS 0.201f
C28366 m3_1864_7102# VSS 0.191f
C28367 m3_34996_8106# VSS 0.201f
C28368 m3_1864_8106# VSS 0.191f
C28369 m3_34996_9110# VSS 0.201f
C28370 m3_1864_9110# VSS 0.191f
C28371 m3_34996_10114# VSS 0.201f
C28372 m3_1864_10114# VSS 0.191f
C28373 m3_34996_11118# VSS 0.201f
C28374 m3_1864_11118# VSS 0.191f
C28375 m3_34996_12122# VSS 0.201f
C28376 m3_1864_12122# VSS 0.191f
C28377 m3_34996_13126# VSS 0.201f
C28378 m3_1864_13126# VSS 0.191f
C28379 m3_34996_14130# VSS 0.201f
C28380 m3_1864_14130# VSS 0.191f
C28381 m3_34996_15134# VSS 0.201f
C28382 m3_1864_15134# VSS 0.191f
C28383 m3_34996_16138# VSS 0.201f
C28384 m3_1864_16138# VSS 0.191f
C28385 m3_34996_17142# VSS 0.201f
C28386 m3_1864_17142# VSS 0.191f
C28387 m3_34996_18146# VSS 0.271f
C28388 m3_33992_18146# VSS 0.145f
C28389 m3_32988_18146# VSS 0.144f
C28390 m3_31984_18146# VSS 0.122f
C28391 m3_30980_18146# VSS 0.0916f
C28392 m3_29976_18146# VSS 0.144f
C28393 m3_28972_18146# VSS 0.144f
C28394 m3_27968_18146# VSS 0.121f
C28395 m3_26964_18146# VSS 0.0931f
C28396 m3_25960_18146# VSS 0.144f
C28397 m3_24956_18146# VSS 0.144f
C28398 m3_23952_18146# VSS 0.12f
C28399 m3_22948_18146# VSS 0.0947f
C28400 m3_21944_18146# VSS 0.143f
C28401 m3_20940_18146# VSS 0.144f
C28402 m3_19936_18146# VSS 0.119f
C28403 m3_18932_18146# VSS 0.0955f
C28404 m3_17928_18146# VSS 0.143f
C28405 m3_16924_18146# VSS 0.144f
C28406 m3_15920_18146# VSS 0.118f
C28407 m3_14916_18146# VSS 0.0959f
C28408 m3_13912_18146# VSS 0.143f
C28409 m3_12908_18146# VSS 0.144f
C28410 m3_11904_18146# VSS 0.118f
C28411 m3_10900_18146# VSS 0.0963f
C28412 m3_9896_18146# VSS 0.143f
C28413 m3_8892_18146# VSS 0.144f
C28414 m3_7888_18146# VSS 0.118f
C28415 m3_6884_18146# VSS 0.0966f
C28416 m3_5880_18146# VSS 0.143f
C28417 m3_4876_18146# VSS 0.144f
C28418 m3_3872_18146# VSS 0.118f
C28419 m3_2868_18146# VSS 0.0979f
C28420 m3_1864_18146# VSS 0.319f
C28421 m3_1046_19620# VSS 0.645f
C28422 m2_35292_1374# VSS 0.0334f
C28423 m2_34864_946# VSS 1.92f
C28424 m2_33860_946# VSS 0.774f
C28425 m2_33284_1374# VSS 0.0334f
C28426 m2_32856_946# VSS 1.04f
C28427 m2_32280_1374# VSS 0.0334f
C28428 m2_31852_946# VSS 1.07f
C28429 m2_31276_1374# VSS 0.0334f
C28430 m2_30848_946# VSS 1.07f
C28431 m2_30272_1374# VSS 0.0334f
C28432 m2_29844_946# VSS 1.07f
C28433 m2_29268_1374# VSS 0.0334f
C28434 m2_28840_946# VSS 1.07f
C28435 m2_28264_1374# VSS 0.0334f
C28436 m2_27836_946# VSS 1.08f
C28437 m2_27260_1374# VSS 0.0334f
C28438 m2_26832_946# VSS 1.08f
C28439 m2_26256_1374# VSS 0.0334f
C28440 m2_25828_946# VSS 1.08f
C28441 m2_25252_1374# VSS 0.0334f
C28442 m2_24824_946# VSS 1.08f
C28443 m2_24248_1374# VSS 0.0334f
C28444 m2_23820_946# VSS 1.08f
C28445 m2_23244_1374# VSS 0.0334f
C28446 m2_22816_946# VSS 1.08f
C28447 m2_22240_1374# VSS 0.0334f
C28448 m2_21812_946# VSS 1.08f
C28449 m2_21236_1374# VSS 0.0334f
C28450 m2_20808_946# VSS 1.08f
C28451 m2_20232_1374# VSS 0.0272f
C28452 m2_19228_1374# VSS 0.0275f
C28453 m2_18224_1374# VSS 0.0276f
C28454 m2_17220_1374# VSS 0.0334f
C28455 m2_16792_946# VSS 1.08f
C28456 m2_16216_1374# VSS 0.0334f
C28457 m2_15788_946# VSS 1.08f
C28458 m2_15212_1374# VSS 0.0334f
C28459 m2_14784_946# VSS 1.08f
C28460 m2_14208_1374# VSS 0.0334f
C28461 m2_13780_946# VSS 1.08f
C28462 m2_13204_1374# VSS 0.0334f
C28463 m2_12776_946# VSS 1.08f
C28464 m2_12200_1374# VSS 0.0334f
C28465 m2_11772_946# VSS 1.08f
C28466 m2_11196_1374# VSS 0.0334f
C28467 m2_10768_946# VSS 1.08f
C28468 m2_10192_1374# VSS 0.0334f
C28469 m2_9764_946# VSS 1.08f
C28470 m2_9188_1374# VSS 0.0334f
C28471 m2_8760_946# VSS 1.08f
C28472 m2_8184_1374# VSS 0.0334f
C28473 m2_7756_946# VSS 1.08f
C28474 m2_7180_1374# VSS 0.0334f
C28475 m2_6752_946# VSS 1.08f
C28476 m2_6176_1374# VSS 0.0334f
C28477 m2_5748_946# VSS 1.08f
C28478 m2_5172_1374# VSS 0.0334f
C28479 m2_4744_946# VSS 1.08f
C28480 m2_4168_1374# VSS 0.0272f
C28481 m2_3164_1374# VSS 0.0334f
C28482 m2_2736_946# VSS 1.08f
C28483 m2_2160_1374# VSS 0.0222f
C28484 m2_1732_946# VSS 1.8f
C28485 m2_34864_1950# VSS 1.26f
C28486 m2_2736_1950# VSS 0.553f
C28487 m2_1732_1950# VSS 1.21f
C28488 m2_34864_2954# VSS 1.29f
C28489 m2_1732_2954# VSS 1.21f
C28490 m2_34864_3958# VSS 1.28f
C28491 m2_1732_3958# VSS 1.21f
C28492 m2_34864_4962# VSS 1.28f
C28493 m2_1732_4962# VSS 1.21f
C28494 m2_34864_5966# VSS 1.26f
C28495 m2_1732_5966# VSS 1.21f
C28496 m2_34864_6970# VSS 1.28f
C28497 m2_1732_6970# VSS 1.21f
C28498 m2_34864_7974# VSS 1.29f
C28499 m2_1732_7974# VSS 1.21f
C28500 m2_34864_8978# VSS 1.28f
C28501 m2_1732_8978# VSS 1.21f
C28502 m2_34864_9982# VSS 1.26f
C28503 m2_1732_9982# VSS 1.21f
C28504 m2_34864_10986# VSS 1.28f
C28505 m2_1732_10986# VSS 1.21f
C28506 m2_34864_11990# VSS 1.29f
C28507 m2_1732_11990# VSS 1.21f
C28508 m2_34864_12994# VSS 1.28f
C28509 m2_1732_12994# VSS 1.21f
C28510 m2_34864_13998# VSS 1.26f
C28511 m2_1732_13998# VSS 1.21f
C28512 m2_34864_15002# VSS 1.28f
C28513 m2_1732_15002# VSS 1.21f
C28514 m2_34864_16006# VSS 1.29f
C28515 m2_1732_16006# VSS 1.21f
C28516 m2_34864_17010# VSS 1.28f
C28517 m2_1732_17010# VSS 1.21f
C28518 m2_34864_18014# VSS 1.72f
C28519 m2_33860_18014# VSS 1.17f
C28520 m2_32856_18014# VSS 1.18f
C28521 m2_31852_18014# VSS 1.07f
C28522 m2_30848_18014# VSS 1.03f
C28523 m2_29844_18014# VSS 1.16f
C28524 m2_28840_18014# VSS 1.18f
C28525 m2_27836_18014# VSS 1.07f
C28526 m2_26832_18014# VSS 1.03f
C28527 m2_25828_18014# VSS 1.16f
C28528 m2_24824_18014# VSS 1.18f
C28529 m2_23820_18014# VSS 1.07f
C28530 m2_22816_18014# VSS 1.03f
C28531 m2_21812_18014# VSS 1.17f
C28532 m2_20808_18014# VSS 1.18f
C28533 m2_19804_18014# VSS 1.06f
C28534 m2_18800_18014# VSS 1.03f
C28535 m2_17796_18014# VSS 1.17f
C28536 m2_16792_18014# VSS 1.18f
C28537 m2_15788_18014# VSS 1.06f
C28538 m2_14784_18014# VSS 1.04f
C28539 m2_13780_18014# VSS 1.17f
C28540 m2_12776_18014# VSS 1.18f
C28541 m2_11772_18014# VSS 1.06f
C28542 m2_10768_18014# VSS 1.04f
C28543 m2_9764_18014# VSS 1.17f
C28544 m2_8760_18014# VSS 1.18f
C28545 m2_7756_18014# VSS 1.06f
C28546 m2_6752_18014# VSS 1.04f
C28547 m2_5748_18014# VSS 1.17f
C28548 m2_4744_18014# VSS 1.18f
C28549 m2_3740_18014# VSS 1.06f
C28550 m2_2736_18014# VSS 1.04f
C28551 m2_1732_18014# VSS 1.93f
C28552 m2_1046_19620# VSS 0.249f
.ends

.subckt sky130_fd_sc_hd__o21ai_4 VPWR VGND B1 Y A1 A2 VPB VNB
X0 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1 a_115_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2 a_115_297# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3 VPWR A1 a_115_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.14 ps=1.28 w=1 l=0.15
X4 VGND A2 a_32_47# VNB sky130_fd_pr__nfet_01v8 ad=0.104 pd=0.97 as=0.091 ps=0.93 w=0.65 l=0.15
X5 Y B1 a_32_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X6 VGND A1 a_32_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.172 ps=1.83 w=0.65 l=0.15
X7 Y B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X8 a_32_47# B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.185 pd=1.87 as=0.091 ps=0.93 w=0.65 l=0.15
X9 Y B1 a_32_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X10 Y A2 a_115_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X11 a_32_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X12 a_32_47# B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X13 a_32_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X14 a_115_297# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X15 a_32_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.104 ps=0.97 w=0.65 l=0.15
X16 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X17 a_32_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X18 VGND A2 a_32_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X19 Y B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.16 ps=1.32 w=1 l=0.15
X20 VPWR A1 a_115_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X21 Y A2 a_115_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X22 VGND A1 a_32_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X23 a_115_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__o211ai_1 VGND VPWR A1 Y C1 B1 A2 VPB VNB
X0 a_110_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.265 ps=2.53 w=1 l=0.15
X1 VGND A1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.127 pd=1.04 as=0.172 ps=1.83 w=0.65 l=0.15
X2 Y A2 a_110_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.105 ps=1.21 w=1 l=0.15
X3 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.195 ps=1.39 w=1 l=0.15
X4 a_27_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.127 pd=1.04 as=0.127 ps=1.04 w=0.65 l=0.15
X5 a_326_47# B1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.86 as=0.127 ps=1.04 w=0.65 l=0.15
X6 Y C1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.635 pd=3.27 as=0.195 ps=1.39 w=1 l=0.15
X7 Y C1 a_326_47# VNB sky130_fd_pr__nfet_01v8 ad=0.393 pd=2.51 as=0.0683 ps=0.86 w=0.65 l=0.15
.ends

.subckt adc_inverter in out VDD VSS
X0 out in VDD VDD sky130_fd_pr__pfet_01v8 ad=0.118 pd=1.4 as=0.0651 ps=0.73 w=0.42 l=0.15
X1 VDD in out VDD sky130_fd_pr__pfet_01v8 ad=0.0651 pd=0.73 as=0.122 ps=1.42 w=0.42 l=0.15
X2 out in VSS VSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
.ends

.subckt adc_nor a b VSS VDD q
X0 a_312_106# b q VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X1 VSS b q VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2 q a a_120_106# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X3 VDD a a_312_106# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X4 q a VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X5 a_120_106# b VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
.ends

.subckt adc_nor_latch qn q VDD VSS s r
X0 a_806_530# qn VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X1 q r a_806_530# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X2 q r VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X3 a_998_530# qn q VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X4 VSS qn q VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5 VDD r a_998_530# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
X6 a_480_530# q qn VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X7 qn s VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X8 VSS q qn VSS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X9 a_288_530# q VDD VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X10 qn s a_288_530# VDD sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.15
X11 VDD s a_480_530# VDD sky130_fd_pr__pfet_01v8 ad=0.248 pd=2.22 as=0.132 ps=1.13 w=0.8 l=0.15
.ends

.subckt adc_noise_decoup_cell2 nmoscap_bot nmoscap_top pwell mimcap_bot mimcap_top
X0 mimcap_top mimcap_bot sky130_fd_pr__cap_mim_m3_1 l=5.1 w=18.9
X1 nmoscap_top nmoscap_bot pwell sky130_fd_pr__cap_var_lvt w=18.4 l=3.9
.ends

.subckt adc_comp_buffer out in VSS VDD
X0 out a_26_n216# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1 VDD a_26_n216# out VDD sky130_fd_pr__pfet_01v8 ad=0.31 pd=2.62 as=0.165 ps=1.33 w=1 l=0.15
X2 VSS a_26_n216# out VSS sky130_fd_pr__nfet_01v8 ad=0.155 pd=1.62 as=0.0825 ps=0.83 w=0.5 l=0.15
X3 VSS in a_26_n216# VSS sky130_fd_pr__nfet_01v8 ad=0.0825 pd=0.83 as=0.155 ps=1.62 w=0.5 l=0.15
X4 VDD in a_26_n216# VDD sky130_fd_pr__pfet_01v8 ad=0.165 pd=1.33 as=0.31 ps=2.62 w=1 l=0.15
X5 out a_26_n216# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0825 pd=0.83 as=0.0825 ps=0.83 w=0.5 l=0.15
.ends

.subckt adc_comp_circuit bp bn on op VPWR VGND a_30_n1001# a_1611_n1292# adc_comp_buffer_0/out
+ a_470_n1001# a_12_n446# adc_comp_buffer_1/out
Xadc_noise_decoup_cell2_0 VGND op VGND VGND VGND adc_noise_decoup_cell2
Xadc_noise_decoup_cell2_1 VGND on VGND VGND VGND adc_noise_decoup_cell2
Xadc_comp_buffer_0 adc_comp_buffer_0/out bn VGND VPWR adc_comp_buffer
Xadc_comp_buffer_1 adc_comp_buffer_1/out bp VGND VPWR adc_comp_buffer
X0 VPWR a_12_n446# on VPWR sky130_fd_pr__pfet_01v8 ad=0.0775 pd=0.81 as=0.0775 ps=0.81 w=0.5 l=0.15
X1 VGND a_12_n446# a_n28_n1170# VGND sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2 bp a_1611_n1292# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.31 ps=2.31 w=2 l=0.15
X3 a_1090_n348# bn VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.15
X4 VPWR a_12_n446# on VPWR sky130_fd_pr__pfet_01v8 ad=0.0775 pd=0.81 as=0.0775 ps=0.81 w=0.5 l=0.15
X5 a_1877_n348# op a_1877_n348# VPWR sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0 ps=0 w=2 l=0.15
X6 op a_12_n446# VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.0775 pd=0.81 as=0.0775 ps=0.81 w=0.5 l=0.15
X7 VGND bn bp VGND sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.15
X8 a_n28_n1170# a_30_n1001# a_n28_n1170# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.58 pd=4.58 as=0 ps=0 w=2 l=0.15
X9 op a_30_n1001# a_n28_n1170# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.15
X10 on a_470_n1001# a_n28_n1170# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.15
X11 VGND a_12_n446# a_n28_n1170# VGND sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X12 a_n28_n1170# a_12_n446# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X13 on a_470_n1001# a_n28_n1170# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.15
X14 a_n28_n1170# a_470_n1001# a_n28_n1170# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.29 as=0 ps=0 w=2 l=0.15
X15 a_n28_n1170# a_12_n446# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X16 bp on a_1090_n348# VPWR sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.15
X17 a_n28_n1170# a_30_n1001# op VGND sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.15
X18 a_1877_n348# bp VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.15
X19 on a_12_n446# VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.0775 pd=0.81 as=0.0775 ps=0.81 w=0.5 l=0.15
X20 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0 ps=0 w=2 l=0.15
X21 VPWR bn a_1090_n348# VPWR sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.15
X22 a_n28_n1170# a_12_n446# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X23 a_n28_n1170# a_12_n446# a_n28_n1170# VGND sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0 ps=0 w=0.5 l=0.15
X24 bn bp VGND VGND sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.15
X25 a_1877_n348# op bn VPWR sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.15
X26 VPWR a_12_n446# op VPWR sky130_fd_pr__pfet_01v8 ad=0.0775 pd=0.81 as=0.0775 ps=0.81 w=0.5 l=0.15
X27 on a_12_n446# VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.0775 pd=0.81 as=0.0775 ps=0.81 w=0.5 l=0.15
X28 VGND a_12_n446# a_n28_n1170# VGND sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X29 VGND a_1611_n1292# bn VGND sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.31 as=0.33 ps=2.33 w=2 l=0.15
X30 a_1090_n348# bn a_1090_n348# VPWR sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0 ps=0 w=2 l=0.15
X31 a_n28_n1170# a_470_n1001# on VGND sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.15
X32 a_n28_n1170# a_30_n1001# op VGND sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.15
X33 a_n28_n1170# a_470_n1001# on VGND sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.15
X34 VGND a_12_n446# a_n28_n1170# VGND sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X35 a_n28_n1170# a_12_n446# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X36 op a_12_n446# VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.0775 pd=0.81 as=0.0775 ps=0.81 w=0.5 l=0.15
X37 a_1090_n348# on a_1090_n348# VPWR sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0 ps=0 w=2 l=0.15
X38 op a_30_n1001# a_n28_n1170# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.15
X39 VPWR bp a_1877_n348# VPWR sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.15
X40 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.31 as=0 ps=0 w=2 l=0.15
X41 VPWR a_12_n446# VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.155 pd=1.62 as=0 ps=0 w=0.5 l=0.15
X42 VPWR a_12_n446# op VPWR sky130_fd_pr__pfet_01v8 ad=0.0775 pd=0.81 as=0.0775 ps=0.81 w=0.5 l=0.15
X43 VPWR a_12_n446# VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.0775 pd=0.81 as=0 ps=0 w=0.5 l=0.15
X44 a_1877_n348# bp a_1877_n348# VPWR sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0 ps=0 w=2 l=0.15
X45 a_1090_n348# on bp VPWR sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.15
X46 bn op a_1877_n348# VPWR sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.15
X47 a_n28_n1170# a_12_n446# a_n28_n1170# VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.15
.ends

.subckt adc_comp_latch clk inp inn comp_trig latch_qn latch_q VDD VSS
Xadc_inverter_1 adc_inverter_1/in adc_inverter_1/out VDD VSS adc_inverter
Xadc_inverter_2 clk adc_inverter_1/in VDD VSS adc_inverter
Xadc_nor_0 adc_nor_0/a adc_nor_0/b VSS VDD comp_trig adc_nor
Xadc_nor_latch_0 latch_qn latch_q VDD VSS adc_nor_0/b adc_nor_0/a adc_nor_latch
Xadc_comp_circuit_0 adc_comp_circuit_0/bp adc_comp_circuit_0/bn adc_comp_circuit_0/on
+ adc_comp_circuit_0/op VDD VSS inn adc_inverter_1/in adc_nor_0/a inp adc_inverter_1/out
+ adc_nor_0/b adc_comp_circuit
.ends

.subckt sky130_fd_sc_hd__clkbuf_4 VGND VPWR A X VPB VNB
X0 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X1 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0588 ps=0.7 w=0.42 l=0.15
X2 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0703 pd=0.755 as=0.111 ps=1.37 w=0.42 l=0.15
X6 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.14 ps=1.28 w=1 l=0.15
X7 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0703 ps=0.755 w=0.42 l=0.15
X8 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.165 ps=1.33 w=1 l=0.15
X9 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__o211a_1 VGND VPWR X A1 A2 B1 C1 VPB VNB
X0 VGND A1 a_215_47# VNB sky130_fd_pr__nfet_01v8 ad=0.106 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X1 a_510_47# B1 a_215_47# VNB sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.143 ps=1.09 w=0.65 l=0.15
X2 a_79_21# C1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.175 ps=1.35 w=1 l=0.15
X3 VPWR B1 a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.175 pd=1.35 as=0.22 ps=1.44 w=1 l=0.15
X4 a_79_21# A2 a_297_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.22 pd=1.44 as=0.162 ps=1.33 w=1 l=0.15
X5 a_297_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.162 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X6 a_79_21# C1 a_510_47# VNB sky130_fd_pr__nfet_01v8 ad=0.195 pd=1.9 as=0.114 ps=1 w=0.65 l=0.15
X7 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X8 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X9 a_215_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.09 as=0.106 ps=0.975 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__and4b_1 VGND VPWR X D C B A_N VPB VNB
X0 a_297_47# a_27_47# a_193_413# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X1 a_369_47# B a_297_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0735 pd=0.77 as=0.0441 ps=0.63 w=0.42 l=0.15
X2 VPWR D a_193_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.141 pd=1.33 as=0.0662 ps=0.735 w=0.42 l=0.15
X3 X a_193_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.103 ps=1 w=0.65 l=0.15
X4 VPWR A_N a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X5 VGND D a_469_47# VNB sky130_fd_pr__nfet_01v8 ad=0.103 pd=1 as=0.0609 ps=0.71 w=0.42 l=0.15
X6 X a_193_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.141 ps=1.33 w=1 l=0.15
X7 VPWR B a_193_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.128 pd=1.03 as=0.0987 ps=0.89 w=0.42 l=0.15
X8 a_193_413# C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.128 ps=1.03 w=0.42 l=0.15
X9 a_193_413# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0987 pd=0.89 as=0.0567 ps=0.69 w=0.42 l=0.15
X10 a_469_47# C a_369_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.0735 ps=0.77 w=0.42 l=0.15
X11 VGND A_N a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__o21bai_1 VPWR VGND A1 B1_N Y A2 VPB VNB
X0 a_388_297# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.25 as=0.153 ps=1.3 w=1 l=0.15
X1 a_105_352# B1_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X2 a_297_47# a_105_352# Y VNB sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.169 ps=1.82 w=0.65 l=0.15
X3 a_297_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4 VPWR A1 a_388_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.127 ps=1.25 w=1 l=0.15
X5 VGND A2 a_297_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.101 ps=0.96 w=0.65 l=0.15
X6 VPWR B1_N a_105_352# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.178 pd=1.4 as=0.109 ps=1.36 w=0.42 l=0.15
X7 Y a_105_352# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.153 pd=1.3 as=0.178 ps=1.4 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__o22a_2 VGND VPWR A1 A2 B2 B1 X VPB VNB
X0 a_301_47# B2 a_81_21# VNB sky130_fd_pr__nfet_01v8 ad=0.123 pd=1.03 as=0.0878 ps=0.92 w=0.65 l=0.15
X1 VGND A2 a_301_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.123 ps=1.03 w=0.65 l=0.15
X2 a_383_297# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.39 ps=1.78 w=1 l=0.15
X3 VPWR a_81_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.39 pd=1.78 as=0.135 ps=1.27 w=1 l=0.15
X4 a_301_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5 VGND a_81_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6 X a_81_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7 X a_81_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X8 VPWR A1 a_579_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.105 ps=1.21 w=1 l=0.15
X9 a_81_21# B1 a_301_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X10 a_579_297# A2 a_81_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.235 ps=1.47 w=1 l=0.15
X11 a_81_21# B2 a_383_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.235 pd=1.47 as=0.105 ps=1.21 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__o21a_2 VGND VPWR X B1 A2 A1 VPB VNB
X0 VPWR A1 a_470_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.16 ps=1.32 w=1 l=0.15
X1 a_79_21# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.4 ps=1.8 w=1 l=0.15
X2 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.0894 ps=0.925 w=0.65 l=0.15
X3 VGND A2 a_384_47# VNB sky130_fd_pr__nfet_01v8 ad=0.104 pd=0.97 as=0.091 ps=0.93 w=0.65 l=0.15
X4 a_470_297# A2 a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.14 ps=1.28 w=1 l=0.15
X5 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.4 pd=1.8 as=0.138 ps=1.27 w=1 l=0.15
X6 a_384_47# B1 a_79_21# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.172 ps=1.83 w=0.65 l=0.15
X7 a_384_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.104 ps=0.97 w=0.65 l=0.15
X8 X a_79_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.138 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X9 X a_79_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0894 pd=0.925 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__or2_2 VPWR VGND X A B VPB VNB
X0 a_121_297# B a_39_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X1 X a_39_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.107 ps=1 w=0.65 l=0.15
X2 VPWR a_39_297# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3 X a_39_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.156 ps=1.36 w=1 l=0.15
X4 VGND a_39_297# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5 VPWR A a_121_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.156 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X6 VGND A a_39_297# VNB sky130_fd_pr__nfet_01v8 ad=0.107 pd=1 as=0.0567 ps=0.69 w=0.42 l=0.15
X7 a_39_297# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__a221o_2 VPWR VGND C1 B2 B1 A1 A2 X VPB VNB
X0 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.285 pd=2.57 as=0.135 ps=1.27 w=1 l=0.15
X1 a_465_47# A1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X2 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.157 ps=1.32 w=1 l=0.15
X3 a_109_297# B1 a_193_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4 a_193_297# B2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.102 ps=0.965 w=0.65 l=0.15
X6 a_205_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.86 as=0.107 ps=0.98 w=0.65 l=0.15
X7 VPWR A2 a_193_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.157 pd=1.32 as=0.165 ps=1.33 w=1 l=0.15
X8 a_193_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X9 a_27_47# B1 a_205_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0683 ps=0.86 w=0.65 l=0.15
X10 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.185 pd=1.87 as=0.0878 ps=0.92 w=0.65 l=0.15
X11 a_109_297# C1 a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X12 VGND C1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X13 VGND A2 a_465_47# VNB sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.965 as=0.107 ps=0.98 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__o2bb2a_1 VPWR VGND X A1_N A2_N B2 B1 VPB VNB
X0 a_206_369# A1_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.129 pd=1.18 as=0.146 ps=1.34 w=0.42 l=0.15
X1 a_206_369# A2_N a_205_47# VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0662 ps=0.735 w=0.42 l=0.15
X2 VGND B2 a_489_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X3 a_585_369# B2 a_76_199# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0672 ps=0.74 w=0.42 l=0.15
X4 a_489_47# a_206_369# a_76_199# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X5 a_489_47# B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X6 VPWR A2_N a_206_369# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.209 pd=1.35 as=0.129 ps=1.18 w=0.42 l=0.15
X7 a_76_199# a_206_369# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0672 pd=0.74 as=0.209 ps=1.35 w=0.42 l=0.15
X8 a_205_47# A1_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0662 pd=0.735 as=0.0986 ps=0.98 w=0.42 l=0.15
X9 VPWR a_76_199# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.146 pd=1.34 as=0.26 ps=2.52 w=1 l=0.15
X10 VPWR B1 a_585_369# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X11 VGND a_76_199# X VNB sky130_fd_pr__nfet_01v8 ad=0.0986 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__a211o_1 VGND VPWR X C1 A2 A1 B1 VPB VNB
X0 VPWR a_80_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.265 ps=2.53 w=1 l=0.15
X1 a_80_21# C1 a_472_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.155 ps=1.31 w=1 l=0.15
X2 VPWR A2 a_217_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X3 VGND B1 a_80_21# VNB sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.091 ps=0.93 w=0.65 l=0.15
X4 VGND a_80_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.26 pd=1.45 as=0.172 ps=1.83 w=0.65 l=0.15
X5 a_300_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.26 ps=1.45 w=0.65 l=0.15
X6 a_217_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X7 a_80_21# A1 a_300_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X8 a_472_297# B1 a_217_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.14 ps=1.28 w=1 l=0.15
X9 a_80_21# C1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.101 ps=0.96 w=0.65 l=0.15
.ends

.subckt scboundary VSS VDD
X0 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.248 pd=2.1 as=0 ps=0 w=0.69 l=0.71
.ends

.subckt sky130_fd_sc_hd__nand2_4 VGND VPWR B Y A VPB VNB
X0 a_27_47# A Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1 a_27_47# A Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6 a_27_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X7 a_27_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X8 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X9 VGND B a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X10 Y A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X11 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X12 Y A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X13 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X14 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X15 VGND B a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__o31a_1 VGND VPWR X A1 A2 A3 B1 VPB VNB
X0 a_103_199# B1 a_253_47# VNB sky130_fd_pr__nfet_01v8 ad=0.201 pd=1.92 as=0.107 ps=0.98 w=0.65 l=0.15
X1 VPWR a_103_199# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.36 ps=2.72 w=1 l=0.15
X2 a_337_297# A2 a_253_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X3 a_103_199# A3 a_337_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.213 pd=1.42 as=0.165 ps=1.33 w=1 l=0.15
X4 a_253_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.195 ps=1.39 w=1 l=0.15
X5 VPWR B1 a_103_199# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.345 pd=2.69 as=0.213 ps=1.42 w=1 l=0.15
X6 VGND a_103_199# X VNB sky130_fd_pr__nfet_01v8 ad=0.127 pd=1.04 as=0.234 ps=2.02 w=0.65 l=0.15
X7 a_253_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.127 ps=1.04 w=0.65 l=0.15
X8 a_253_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.107 ps=0.98 w=0.65 l=0.15
X9 VGND A2 a_253_47# VNB sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.0878 ps=0.92 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__dfstp_1 VPWR VGND Q SET_B D CLK VPB VNB
X0 VGND a_652_21# a_586_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0882 pd=0.84 as=0.0671 ps=0.75 w=0.42 l=0.15
X1 a_956_413# a_476_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0483 pd=0.65 as=0.0567 ps=0.69 w=0.42 l=0.15
X2 VPWR a_476_47# a_652_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X3 a_586_47# a_193_47# a_476_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.072 ps=0.76 w=0.36 l=0.15
X4 VPWR CLK a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X5 a_476_47# a_27_47# a_381_47# VNB sky130_fd_pr__nfet_01v8 ad=0.072 pd=0.76 as=0.0935 ps=0.965 w=0.36 l=0.15
X6 a_1056_47# a_476_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X7 a_381_47# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.125 pd=1.17 as=0.218 ps=2.2 w=0.84 l=0.15
X8 a_652_21# SET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0798 ps=0.8 w=0.42 l=0.15
X9 a_1224_47# a_27_47# a_1032_413# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X10 a_562_413# a_27_47# a_476_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0567 ps=0.69 w=0.42 l=0.15
X11 VGND a_1032_413# a_1602_47# VNB sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X12 VPWR a_1182_261# a_1140_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X13 Q a_1602_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.149 ps=1.33 w=1 l=0.15
X14 a_1032_413# a_193_47# a_1056_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X15 a_476_47# a_193_47# a_381_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.125 ps=1.17 w=0.42 l=0.15
X16 a_1296_47# a_1182_261# a_1224_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0483 pd=0.65 as=0.0441 ps=0.63 w=0.42 l=0.15
X17 a_193_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X18 VPWR a_652_21# a_562_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.0945 ps=0.87 w=0.42 l=0.15
X19 VPWR SET_B a_1032_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.123 pd=1.17 as=0.109 ps=1.36 w=0.42 l=0.15
X20 a_1032_413# a_27_47# a_956_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0483 ps=0.65 w=0.42 l=0.15
X21 a_1182_261# a_1032_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.218 pd=2.2 as=0.123 ps=1.17 w=0.84 l=0.15
X22 Q a_1602_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X23 a_193_47# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X24 a_1140_413# a_193_47# a_1032_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0819 ps=0.81 w=0.42 l=0.15
X25 VPWR a_1032_413# a_1602_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.166 ps=1.8 w=0.64 l=0.15
X26 a_796_47# SET_B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0882 ps=0.84 w=0.42 l=0.15
X27 a_381_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0935 pd=0.965 as=0.166 ps=1.8 w=0.64 l=0.15
X28 a_1182_261# a_1032_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.6 as=0.114 ps=1.01 w=0.54 l=0.15
X29 a_652_21# a_476_47# a_796_47# VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X30 VGND CLK a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X31 VGND SET_B a_1296_47# VNB sky130_fd_pr__nfet_01v8 ad=0.114 pd=1.01 as=0.0483 ps=0.65 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__a21oi_4 VGND VPWR A2 B1 Y A1 VPB VNB
X0 a_28_297# B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1 a_462_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X2 Y B1 a_28_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.26 ps=2.52 w=1 l=0.15
X3 Y B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X4 a_462_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X5 a_28_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6 a_462_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.104 ps=0.97 w=0.65 l=0.15
X7 Y B1 a_28_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X8 VGND B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.104 pd=0.97 as=0.091 ps=0.93 w=0.65 l=0.15
X9 VGND B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X10 Y A1 a_462_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X11 a_28_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.145 ps=1.29 w=1 l=0.15
X12 VPWR A2 a_28_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X13 Y B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.172 ps=1.83 w=0.65 l=0.15
X14 VGND A2 a_462_47# VNB sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X15 a_28_297# B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.14 ps=1.28 w=1 l=0.15
X16 VPWR A1 a_28_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X17 a_28_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X18 VGND A2 a_462_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X19 VPWR A2 a_28_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.155 ps=1.31 w=1 l=0.15
X20 a_28_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X21 Y A1 a_462_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X22 a_462_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X23 VPWR A1 a_28_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
.ends

.subckt sky130_mm_sc_hd_dlyPoly5ns VPWR VGND in out mid VPB VNB
X0 a_1691_329# out VGND VPB sky130_fd_pr__pfet_01v8_hvt ad=0.24 pd=2.2 as=0.132 ps=1.13 w=0.8 l=0.15
X1 a_1691_329# mid VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.132 pd=1.13 as=0.24 ps=2.2 w=0.8 l=0.15
X2 out mid a_1691_329# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.24 pd=2.2 as=0.132 ps=1.13 w=0.8 l=0.15
X3 VGND out a_1691_329# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.132 pd=1.13 as=0.248 ps=2.22 w=0.8 l=0.15
X4 VGND mid VGND VNB sky130_fd_pr__nfet_01v8 ad=0.399 pd=3.33 as=0 ps=0 w=1.38 l=2.05
X5 a_1632_71# mid VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.126 ps=1.44 w=0.42 l=0.15
X6 VPWR out a_1632_71# VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X7 a_1632_71# out VPWR VNB sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X8 out mid a_1632_71# VNB sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0693 ps=0.75 w=0.42 l=0.15
X9 mid in VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.232 pd=2.18 as=0.232 ps=2.18 w=0.8 l=1.42
X10 mid in VGND VNB sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=3.69
.ends

.subckt sky130_fd_sc_hd__nor2b_1 VGND VPWR B_N A Y VPB VNB
X0 Y a_74_47# a_265_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X1 VPWR B_N a_74_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.157 pd=1.39 as=0.109 ps=1.36 w=0.42 l=0.15
X2 a_265_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.157 ps=1.39 w=1 l=0.15
X3 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.1 ps=0.985 w=0.65 l=0.15
X4 VGND B_N a_74_47# VNB sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.985 as=0.109 ps=1.36 w=0.42 l=0.15
X5 VGND a_74_47# Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__bufbuf_8 VGND VPWR A X VPB VNB
X0 a_318_47# a_206_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1 VPWR a_318_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2 VPWR a_206_47# a_318_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3 X a_318_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4 X a_318_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5 VPWR a_318_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6 X a_318_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7 VGND a_206_47# a_318_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X8 VPWR a_318_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9 X a_318_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X10 a_318_47# a_206_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X11 X a_318_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X12 a_206_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1 ps=0.985 w=0.65 l=0.15
X13 X a_318_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X14 a_206_47# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.154 ps=1.34 w=1 l=0.15
X15 VPWR a_318_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X16 VGND a_206_47# a_318_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X17 VGND a_318_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X18 VGND a_318_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X19 VGND a_318_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X20 X a_318_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X21 VGND a_318_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X22 VPWR a_206_47# a_318_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X23 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.166 ps=1.8 w=0.64 l=0.15
X24 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.985 as=0.109 ps=1.36 w=0.42 l=0.15
X25 X a_318_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
.ends

.subckt adc_clkgen_with_edgedetect VDD clk_comp_out clk_dig_out dlycontrol1_in[0]
+ dlycontrol1_in[1] dlycontrol1_in[2] dlycontrol1_in[3] dlycontrol1_in[4] dlycontrol2_in[0]
+ dlycontrol2_in[1] dlycontrol2_in[2] dlycontrol2_in[3] dlycontrol2_in[4] dlycontrol3_in[0]
+ dlycontrol3_in[1] dlycontrol3_in[2] dlycontrol3_in[3] dlycontrol3_in[4] dlycontrol4_in[0]
+ dlycontrol4_in[1] dlycontrol4_in[2] dlycontrol4_in[3] dlycontrol4_in[4] dlycontrol4_in[5]
+ ena_in enable_dlycontrol_in ndecision_finish_in sample_n_in sample_n_out sample_p_in
+ sample_p_out start_conv_in VSS
XFILLER_10_317 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XFILLER_13_133 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_2.genblk1\[0\].control_invert VDD VSS clkgen.delay_155ns_2.bypass_enable_w\[0\]
+ dlycontrol2_in[0] VDD VSS sky130_fd_sc_hd__inv_2
XFILLER_10_125 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XFILLER_12_10 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XFILLER_12_32 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
Xclkgen.delay_155ns_2.genblk1\[0\].dly_binary.out_mux VSS VDD clkgen.delay_155ns_2.genblk1\[0\].dly_binary.out
+ clkgen.clk_dig_out clkgen.delay_155ns_2.genblk1\[0\].dly_binary.bypass_in clkgen.delay_155ns_2.genblk1\[0\].dly_binary.signal_w\[1\]
+ VDD VSS sky130_fd_sc_hd__mux2_1
Xclkgen.delay_155ns_2.genblk1\[2\].dly_binary.out_mux VSS VDD clkgen.delay_155ns_2.genblk1\[2\].dly_binary.out
+ clkgen.delay_155ns_2.genblk1\[1\].dly_binary.out clkgen.delay_155ns_2.genblk1\[2\].dly_binary.bypass_in
+ clkgen.delay_155ns_2.genblk1\[2\].dly_binary.signal_w\[4\] VDD VSS sky130_fd_sc_hd__mux2_1
Xclkgen.delay_155ns_2.genblk1\[4\].dly_binary.out_mux VSS VDD clkgen.clk_dig_delayed_w
+ clkgen.delay_155ns_2.genblk1\[3\].dly_binary.out clkgen.delay_155ns_2.genblk1\[4\].dly_binary.bypass_in
+ clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[16\] VDD VSS sky130_fd_sc_hd__mux2_1
XFILLER_14_272 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
XANTENNA_clkgen.delay_155ns_1.genblk1\[2\].control_invert_A VSS VDD dlycontrol1_in[2]
+ VDD VSS sky130_fd_sc_hd__diode_2
Xedgedetect.or1 VDD VSS clkgen.enable_loop_in edgedetect.start_conv_edge_w edgedetect.ena_in
+ VDD VSS sky130_fd_sc_hd__or2_1
Xclkgen.delay_155ns_3.genblk1\[0\].dly_binary.genblk1\[0\].delay_unit VDD VSS clkgen.delay_155ns_3.genblk1\[0\].dly_binary.signal_w\[0\]
+ clkgen.delay_155ns_3.genblk1\[0\].dly_binary.signal_w\[1\] clkgen.delay_155ns_3.genblk1\[0\].dly_binary.genblk1\[0\].delay_unit/mid
+ VDD VSS sky130_mm_sc_hd_dlyPoly5ns
XFILLER_16_334 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
XFILLER_4_249 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
Xedgedetect.dly_315ns_1.genblk1\[1\].bypass_enable VDD VSS edgedetect.dly_315ns_1.genblk1\[1\].dly_binary.bypass_in
+ edgedetect.dly_315ns_1.enable_dlycontrol_w edgedetect.dly_315ns_1.bypass_enable_w\[1\]
+ VDD VSS sky130_fd_sc_hd__and2_1
XFILLER_13_3 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XFILLER_3_271 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XFILLER_15_87 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XANTENNA_clkgen.delay_155ns_2.genblk1\[1\].control_invert_A VSS VDD dlycontrol2_in[1]
+ VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_0_241 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
Xclkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[14\].delay_unit VDD VSS clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[14\]
+ clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[15\] clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[14\].delay_unit/mid
+ VDD VSS sky130_mm_sc_hd_dlyPoly5ns
XANTENNA_clkgen.delay_155ns_2.genblk1\[1\].dly_binary.and_bypass_switch_A_N VSS VDD
+ clkgen.delay_155ns_2.genblk1\[1\].dly_binary.bypass_in VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_5_311 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
Xclkgen.delay_155ns_1.genblk1\[2\].bypass_enable VDD VSS clkgen.delay_155ns_1.genblk1\[2\].dly_binary.bypass_in
+ clkgen.delay_155ns_1.enable_dlycontrol_w clkgen.delay_155ns_1.bypass_enable_w\[2\]
+ VDD VSS sky130_fd_sc_hd__and2_1
Xclkgen.delay_155ns_2.genblk1\[3\].bypass_enable VDD VSS clkgen.delay_155ns_2.genblk1\[3\].dly_binary.bypass_in
+ clkgen.delay_155ns_2.enable_dlycontrol_w clkgen.delay_155ns_2.bypass_enable_w\[3\]
+ VDD VSS sky130_fd_sc_hd__and2_1
Xclkgen.delay_155ns_3.genblk1\[4\].bypass_enable VDD VSS clkgen.delay_155ns_3.genblk1\[4\].dly_binary.bypass_in
+ clkgen.delay_155ns_3.enable_dlycontrol_w clkgen.delay_155ns_3.bypass_enable_w\[4\]
+ VDD VSS sky130_fd_sc_hd__and2_1
XFILLER_5_174 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XANTENNA_clkgen.delay_155ns_3.genblk1\[0\].control_invert_A VSS VDD dlycontrol3_in[0]
+ VDD VSS sky130_fd_sc_hd__diode_2
Xedgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[3\].delay_unit VDD VSS edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[3\]
+ edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[4\] edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[3\].delay_unit/mid
+ VDD VSS sky130_mm_sc_hd_dlyPoly5ns
XFILLER_11_276 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XFILLER_18_32 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
Xclkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[1\].delay_unit VDD VSS clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[1\]
+ clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[2\] clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[1\].delay_unit/mid
+ VDD VSS sky130_mm_sc_hd_dlyPoly5ns
Xedgedetect.dly_315ns_1.genblk1\[1\].control_invert VDD VSS edgedetect.dly_315ns_1.bypass_enable_w\[1\]
+ dlycontrol4_in[1] VDD VSS sky130_fd_sc_hd__inv_2
XFILLER_19_151 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XFILLER_3_283 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_6_57 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XFILLER_16_198 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XFILLER_0_253 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
Xedgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[8\].delay_unit VDD VSS edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[8\]
+ edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[9\] edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[8\].delay_unit/mid
+ VDD VSS sky130_mm_sc_hd_dlyPoly5ns
XFILLER_13_113 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XFILLER_5_323 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_2_304 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
Xclkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[12\].delay_unit VDD VSS clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[12\]
+ clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[13\] clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[12\].delay_unit/mid
+ VDD VSS sky130_mm_sc_hd_dlyPoly5ns
XANTENNA_edgedetect.dly_315ns_1.genblk1\[1\].dly_binary.and_bypass_switch_B VSS VDD
+ edgedetect.dly_315ns_1.genblk1\[0\].dly_binary.out VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_5_142 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
Xclkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[6\].delay_unit VDD VSS clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[6\]
+ clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[7\] clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[6\].delay_unit/mid
+ VDD VSS sky130_mm_sc_hd_dlyPoly5ns
XANTENNA_edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.genblk1\[0\].delay_unit_in
+ VSS VDD edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.signal_w\[0\] VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_3_3 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
Xedgedetect.nor1 VSS VDD edgedetect.dly_315ns_1.genblk1\[0\].dly_binary.in edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.out
+ edgedetect.start_conv_edge_w VDD VSS sky130_fd_sc_hd__nor2b_1
Xclkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[0\].delay_unit VDD VSS clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[0\]
+ clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[1\] clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[0\].delay_unit/mid
+ VDD VSS sky130_mm_sc_hd_dlyPoly5ns
XFILLER_11_288 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XFILLER_7_237 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XANTENNA_edgedetect.or1_A VSS VDD edgedetect.start_conv_edge_w VDD VSS sky130_fd_sc_hd__diode_2
Xdelay_sample_p11 VDD VSS sample_p_in sample_p_1 delay_sample_p11/mid VDD VSS sky130_mm_sc_hd_dlyPoly5ns
XFILLER_3_295 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
Xclkgen.delay_155ns_3.genblk1\[1\].control_invert VDD VSS clkgen.delay_155ns_3.bypass_enable_w\[1\]
+ dlycontrol3_in[1] VDD VSS sky130_fd_sc_hd__inv_2
XFILLER_13_306 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XFILLER_0_210 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
XFILLER_0_265 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
Xedgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[3\].delay_unit VDD VSS edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[3\]
+ edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[4\] edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[3\].delay_unit/mid
+ VDD VSS sky130_mm_sc_hd_dlyPoly5ns
Xclkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[5\].delay_unit VDD VSS clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[5\]
+ clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[6\] clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[5\].delay_unit/mid
+ VDD VSS sky130_mm_sc_hd_dlyPoly5ns
XFILLER_5_335 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XFILLER_5_302 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XFILLER_2_316 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
Xclkgen.delay_155ns_3.genblk1\[3\].dly_binary.genblk1\[1\].delay_unit VDD VSS clkgen.delay_155ns_3.genblk1\[3\].dly_binary.signal_w\[1\]
+ clkgen.delay_155ns_3.genblk1\[3\].dly_binary.signal_w\[2\] clkgen.delay_155ns_3.genblk1\[3\].dly_binary.genblk1\[1\].delay_unit/mid
+ VDD VSS sky130_mm_sc_hd_dlyPoly5ns
XFILLER_5_110 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XFILLER_5_121 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
Xedgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[10\].delay_unit VDD VSS edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[10\]
+ edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[11\] edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[10\].delay_unit/mid
+ VDD VSS sky130_mm_sc_hd_dlyPoly5ns
XFILLER_11_256 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[10\].delay_unit VDD VSS clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[10\]
+ clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[11\] clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[10\].delay_unit/mid
+ VDD VSS sky130_mm_sc_hd_dlyPoly5ns
XANTENNA_edgedetect.or1_B VSS VDD edgedetect.ena_in VDD VSS sky130_fd_sc_hd__diode_2
Xedgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[8\].delay_unit VDD VSS edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[8\]
+ edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[9\] edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[8\].delay_unit/mid
+ VDD VSS sky130_mm_sc_hd_dlyPoly5ns
XFILLER_19_120 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_3.genblk1\[3\].dly_binary.genblk1\[6\].delay_unit VDD VSS clkgen.delay_155ns_3.genblk1\[3\].dly_binary.signal_w\[6\]
+ clkgen.delay_155ns_3.genblk1\[3\].dly_binary.signal_w\[7\] clkgen.delay_155ns_3.genblk1\[3\].dly_binary.genblk1\[6\].delay_unit/mid
+ VDD VSS sky130_mm_sc_hd_dlyPoly5ns
Xedgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[11\].delay_unit VDD VSS edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[11\]
+ edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[12\] edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[11\].delay_unit/mid
+ VDD VSS sky130_mm_sc_hd_dlyPoly5ns
XFILLER_16_167 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
XFILLER_11_3 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
Xclkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[4\].delay_unit VDD VSS clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[4\]
+ clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[5\] clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[4\].delay_unit/mid
+ VDD VSS sky130_mm_sc_hd_dlyPoly5ns
Xclkgen.delay_155ns_2.genblk1\[3\].dly_binary.genblk1\[0\].delay_unit VDD VSS clkgen.delay_155ns_2.genblk1\[3\].dly_binary.signal_w\[0\]
+ clkgen.delay_155ns_2.genblk1\[3\].dly_binary.signal_w\[1\] clkgen.delay_155ns_2.genblk1\[3\].dly_binary.genblk1\[0\].delay_unit/mid
+ VDD VSS sky130_mm_sc_hd_dlyPoly5ns
Xedgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[15\].delay_unit VDD VSS edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[15\]
+ edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[16\] edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[15\].delay_unit/mid
+ VDD VSS sky130_mm_sc_hd_dlyPoly5ns
XFILLER_2_328 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
Xclkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[15\].delay_unit VDD VSS clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[15\]
+ clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[16\] clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[15\].delay_unit/mid
+ VDD VSS sky130_mm_sc_hd_dlyPoly5ns
XFILLER_2_125 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
Xclkgen.nor1 VSS VDD clkgen.enable_loop_in clkgen.clk_dig_delayed_w clkgen.delay_155ns_3.genblk1\[0\].dly_binary.in
+ VDD VSS sky130_fd_sc_hd__nor2b_1
XFILLER_11_213 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XFILLER_7_228 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[9\].delay_unit VDD VSS clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[9\]
+ clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[10\] clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[9\].delay_unit/mid
+ VDD VSS sky130_mm_sc_hd_dlyPoly5ns
Xedgedetect.dly_315ns_1.genblk1\[3\].dly_binary.genblk1\[3\].delay_unit VDD VSS edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.signal_w\[3\]
+ edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.signal_w\[4\] edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.genblk1\[3\].delay_unit/mid
+ VDD VSS sky130_mm_sc_hd_dlyPoly5ns
XFILLER_6_272 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
Xclkgen.delay_155ns_2.genblk1\[3\].dly_binary.genblk1\[5\].delay_unit VDD VSS clkgen.delay_155ns_2.genblk1\[3\].dly_binary.signal_w\[5\]
+ clkgen.delay_155ns_2.genblk1\[3\].dly_binary.signal_w\[6\] clkgen.delay_155ns_2.genblk1\[3\].dly_binary.genblk1\[5\].delay_unit/mid
+ VDD VSS sky130_mm_sc_hd_dlyPoly5ns
XANTENNA_clkgen.delay_155ns_1.genblk1\[4\].dly_binary.and_bypass_switch_B VSS VDD
+ clkgen.delay_155ns_1.genblk1\[3\].dly_binary.out VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_3_253 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_3.genblk1\[2\].dly_binary.genblk1\[1\].delay_unit VDD VSS clkgen.delay_155ns_3.genblk1\[2\].dly_binary.signal_w\[1\]
+ clkgen.delay_155ns_3.genblk1\[2\].dly_binary.signal_w\[2\] clkgen.delay_155ns_3.genblk1\[2\].dly_binary.genblk1\[1\].delay_unit/mid
+ VDD VSS sky130_mm_sc_hd_dlyPoly5ns
Xclkgen.delay_155ns_1.genblk1\[2\].control_invert VDD VSS clkgen.delay_155ns_1.bypass_enable_w\[2\]
+ dlycontrol1_in[2] VDD VSS sky130_fd_sc_hd__inv_2
Xedgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[22\].delay_unit VDD VSS edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[22\]
+ edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[23\] edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[22\].delay_unit/mid
+ VDD VSS sky130_mm_sc_hd_dlyPoly5ns
XFILLER_0_223 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XFILLER_8_120 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XANTENNA_edgedetect.dly_315ns_1.enablebuffer_A VSS VDD enable_dlycontrol_in VDD VSS
+ sky130_fd_sc_hd__diode_2
XFILLER_14_244 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
Xedgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[27\].delay_unit VDD VSS edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[27\]
+ edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[28\] edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[27\].delay_unit/mid
+ VDD VSS sky130_mm_sc_hd_dlyPoly5ns
Xclkgen.delay_155ns_1.genblk1\[3\].dly_binary.genblk1\[4\].delay_unit VDD VSS clkgen.delay_155ns_1.genblk1\[3\].dly_binary.signal_w\[4\]
+ clkgen.delay_155ns_1.genblk1\[3\].dly_binary.signal_w\[5\] clkgen.delay_155ns_1.genblk1\[3\].dly_binary.genblk1\[4\].delay_unit/mid
+ VDD VSS sky130_mm_sc_hd_dlyPoly5ns
XANTENNA_clkgen.delay_155ns_1.genblk1\[1\].control_invert_A VSS VDD dlycontrol1_in[1]
+ VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA_clkgen.delay_155ns_2.enablebuffer_A VSS VDD enable_dlycontrol_in VDD VSS
+ sky130_fd_sc_hd__diode_2
XANTENNA_inbuf_3_A VSS VDD ndecision_finish_in VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_1_3 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XFILLER_1_94 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XFILLER_16_306 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_2.genblk1\[2\].dly_binary.genblk1\[0\].delay_unit VDD VSS clkgen.delay_155ns_2.genblk1\[2\].dly_binary.signal_w\[0\]
+ clkgen.delay_155ns_2.genblk1\[2\].dly_binary.signal_w\[1\] clkgen.delay_155ns_2.genblk1\[2\].dly_binary.genblk1\[0\].delay_unit/mid
+ VDD VSS sky130_mm_sc_hd_dlyPoly5ns
XFILLER_3_232 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
Xclkgen.clkdig_inverter VDD VSS clkgen.clk_dig_out clkgen.delay_155ns_1.genblk1\[4\].dly_binary.out
+ VDD VSS sky130_fd_sc_hd__inv_2
XFILLER_3_265 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XFILLER_15_59 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XFILLER_12_320 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XFILLER_16_125 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XFILLER_0_235 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XANTENNA_clkgen.delay_155ns_2.genblk1\[0\].control_invert_A VSS VDD dlycontrol2_in[0]
+ VDD VSS sky130_fd_sc_hd__diode_2
XPHY_0 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XFILLER_17_275 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
Xedgedetect.dly_315ns_1.genblk1\[2\].dly_binary.genblk1\[3\].delay_unit VDD VSS edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.signal_w\[3\]
+ edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.signal_w\[4\] edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.genblk1\[3\].delay_unit/mid
+ VDD VSS sky130_mm_sc_hd_dlyPoly5ns
XFILLER_4_94 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
Xclkgen.delay_155ns_3.genblk1\[1\].dly_binary.genblk1\[1\].delay_unit VDD VSS clkgen.delay_155ns_3.genblk1\[1\].dly_binary.signal_w\[1\]
+ clkgen.delay_155ns_3.genblk1\[1\].dly_binary.signal_w\[2\] clkgen.delay_155ns_3.genblk1\[1\].dly_binary.genblk1\[1\].delay_unit/mid
+ VDD VSS sky130_mm_sc_hd_dlyPoly5ns
XFILLER_19_304 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
XFILLER_19_315 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_3_277 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XFILLER_0_203 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
Xedgedetect.dly_315ns_1.genblk1\[0\].dly_binary.out_mux VSS VDD edgedetect.dly_315ns_1.genblk1\[0\].dly_binary.out
+ edgedetect.dly_315ns_1.genblk1\[0\].dly_binary.in edgedetect.dly_315ns_1.genblk1\[0\].dly_binary.bypass_in
+ edgedetect.dly_315ns_1.genblk1\[0\].dly_binary.signal_w\[1\] VDD VSS sky130_fd_sc_hd__mux2_1
Xdelay_sample_n12 VDD VSS sample_n_in sample_n_1 delay_sample_n12/mid VDD VSS sky130_mm_sc_hd_dlyPoly5ns
XPHY_1 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
Xedgedetect.dly_315ns_1.genblk1\[0\].dly_binary.and_bypass_switch VSS VDD edgedetect.dly_315ns_1.genblk1\[0\].dly_binary.bypass_in
+ edgedetect.dly_315ns_1.genblk1\[0\].dly_binary.signal_w\[0\] edgedetect.dly_315ns_1.genblk1\[0\].dly_binary.in
+ VDD VSS sky130_fd_sc_hd__and2b_1
Xedgedetect.dly_315ns_1.genblk1\[2\].dly_binary.out_mux VSS VDD edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.out
+ edgedetect.dly_315ns_1.genblk1\[1\].dly_binary.out edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.bypass_in
+ edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.signal_w\[4\] VDD VSS sky130_fd_sc_hd__mux2_1
XFILLER_7_94 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
Xinbuf_1 VSS VDD edgedetect.ena_in ena_in VDD VSS sky130_fd_sc_hd__buf_1
XFILLER_8_177 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
Xedgedetect.dly_315ns_1.genblk1\[4\].dly_binary.out_mux VSS VDD edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.out
+ edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.out edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.bypass_in
+ edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[16\] VDD VSS sky130_fd_sc_hd__mux2_1
Xclkgen.delay_155ns_2.genblk1\[1\].dly_binary.genblk1\[0\].delay_unit VDD VSS clkgen.delay_155ns_2.genblk1\[1\].dly_binary.signal_w\[0\]
+ clkgen.delay_155ns_2.genblk1\[1\].dly_binary.signal_w\[1\] clkgen.delay_155ns_2.genblk1\[1\].dly_binary.genblk1\[0\].delay_unit/mid
+ VDD VSS sky130_mm_sc_hd_dlyPoly5ns
XFILLER_14_213 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XFILLER_19_327 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
Xedgedetect.dly_315ns_1.genblk1\[2\].bypass_enable VDD VSS edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.bypass_in
+ edgedetect.dly_315ns_1.enable_dlycontrol_w edgedetect.dly_315ns_1.bypass_enable_w\[2\]
+ VDD VSS sky130_fd_sc_hd__and2_1
Xclkgen.delay_155ns_2.genblk1\[3\].control_invert VDD VSS clkgen.delay_155ns_2.bypass_enable_w\[3\]
+ dlycontrol2_in[3] VDD VSS sky130_fd_sc_hd__inv_2
Xclkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[10\].delay_unit VDD VSS clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[10\]
+ clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[11\] clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[10\].delay_unit/mid
+ VDD VSS sky130_mm_sc_hd_dlyPoly5ns
XFILLER_1_63 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
XFILLER_10_94 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
XANTENNA_clkgen.delay_155ns_2.genblk1\[4\].dly_binary.and_bypass_switch_A_N VSS VDD
+ clkgen.delay_155ns_2.genblk1\[4\].dly_binary.bypass_in VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_3_223 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XFILLER_0_259 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_1.genblk1\[3\].bypass_enable VDD VSS clkgen.delay_155ns_1.genblk1\[3\].dly_binary.bypass_in
+ clkgen.delay_155ns_1.enable_dlycontrol_w clkgen.delay_155ns_1.bypass_enable_w\[3\]
+ VDD VSS sky130_fd_sc_hd__and2_1
XPHY_2 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
Xclkgen.delay_155ns_2.genblk1\[4\].bypass_enable VDD VSS clkgen.delay_155ns_2.genblk1\[4\].dly_binary.bypass_in
+ clkgen.delay_155ns_2.enable_dlycontrol_w clkgen.delay_155ns_2.bypass_enable_w\[4\]
+ VDD VSS sky130_fd_sc_hd__and2_1
Xinbuf_2 VSS VDD edgedetect.dly_315ns_1.genblk1\[0\].dly_binary.in start_conv_in VDD
+ VSS sky130_fd_sc_hd__buf_1
XFILLER_12_152 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XFILLER_8_167 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[15\].delay_unit VDD VSS clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[15\]
+ clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[16\] clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[15\].delay_unit/mid
+ VDD VSS sky130_mm_sc_hd_dlyPoly5ns
XFILLER_4_63 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_1.genblk1\[0\].dly_binary.out_mux VSS VDD clkgen.delay_155ns_1.genblk1\[0\].dly_binary.out
+ clkgen.delay_155ns_1.genblk1\[0\].dly_binary.in clkgen.delay_155ns_1.genblk1\[0\].dly_binary.bypass_in
+ clkgen.delay_155ns_1.genblk1\[0\].dly_binary.signal_w\[1\] VDD VSS sky130_fd_sc_hd__mux2_1
XFILLER_9_19 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_1.genblk1\[2\].dly_binary.out_mux VSS VDD clkgen.delay_155ns_1.genblk1\[2\].dly_binary.out
+ clkgen.delay_155ns_1.genblk1\[1\].dly_binary.out clkgen.delay_155ns_1.genblk1\[2\].dly_binary.bypass_in
+ clkgen.delay_155ns_1.genblk1\[2\].dly_binary.signal_w\[4\] VDD VSS sky130_fd_sc_hd__mux2_1
Xclkgen.delay_155ns_1.genblk1\[4\].dly_binary.out_mux VSS VDD clkgen.delay_155ns_1.genblk1\[4\].dly_binary.out
+ clkgen.delay_155ns_1.genblk1\[3\].dly_binary.out clkgen.delay_155ns_1.genblk1\[4\].dly_binary.bypass_in
+ clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[16\] VDD VSS sky130_fd_sc_hd__mux2_1
Xedgedetect.dly_315ns_1.genblk1\[1\].dly_binary.and_bypass_switch VSS VDD edgedetect.dly_315ns_1.genblk1\[1\].dly_binary.bypass_in
+ edgedetect.dly_315ns_1.genblk1\[1\].dly_binary.signal_w\[0\] edgedetect.dly_315ns_1.genblk1\[0\].dly_binary.out
+ VDD VSS sky130_fd_sc_hd__and2b_1
Xedgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[4\].delay_unit VDD VSS edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[4\]
+ edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[5\] edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[4\].delay_unit/mid
+ VDD VSS sky130_mm_sc_hd_dlyPoly5ns
XFILLER_3_213 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XANTENNA_inbuf_1_A VSS VDD ena_in VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_15_29 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
Xclkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[2\].delay_unit VDD VSS clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[2\]
+ clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[3\] clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[2\].delay_unit/mid
+ VDD VSS sky130_mm_sc_hd_dlyPoly5ns
Xclkgen.delay_155ns_2.genblk1\[0\].dly_binary.genblk1\[0\].delay_unit VDD VSS clkgen.delay_155ns_2.genblk1\[0\].dly_binary.signal_w\[0\]
+ clkgen.delay_155ns_2.genblk1\[0\].dly_binary.signal_w\[1\] clkgen.delay_155ns_2.genblk1\[0\].dly_binary.genblk1\[0\].delay_unit/mid
+ VDD VSS sky130_mm_sc_hd_dlyPoly5ns
XPHY_3 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XFILLER_7_63 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
XFILLER_16_94 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
Xinbuf_3 VSS VDD clkgen.delay_155ns_1.genblk1\[0\].dly_binary.in ndecision_finish_in
+ VDD VSS sky130_fd_sc_hd__buf_1
XFILLER_12_197 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XFILLER_12_164 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XANTENNA_edgedetect.dly_315ns_1.genblk1\[5\].control_invert_A VSS VDD dlycontrol4_in[5]
+ VDD VSS sky130_fd_sc_hd__diode_2
Xedgedetect.dly_315ns_1.genblk1\[4\].control_invert VDD VSS edgedetect.dly_315ns_1.bypass_enable_w\[4\]
+ dlycontrol4_in[4] VDD VSS sky130_fd_sc_hd__inv_2
XFILLER_1_311 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XANTENNA_clkgen.delay_155ns_1.genblk1\[0\].dly_binary.out_mux_S VSS VDD clkgen.delay_155ns_1.genblk1\[0\].dly_binary.bypass_in
+ VDD VSS sky130_fd_sc_hd__diode_2
Xedgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[9\].delay_unit VDD VSS edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[9\]
+ edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[10\] edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[9\].delay_unit/mid
+ VDD VSS sky130_mm_sc_hd_dlyPoly5ns
XFILLER_13_84 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XANTENNA_clkgen.delay_155ns_2.genblk1\[0\].dly_binary.and_bypass_switch_B VSS VDD
+ clkgen.clk_dig_out VDD VSS sky130_fd_sc_hd__diode_2
Xclkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[7\].delay_unit VDD VSS clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[7\]
+ clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[8\] clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[7\].delay_unit/mid
+ VDD VSS sky130_mm_sc_hd_dlyPoly5ns
Xclkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[13\].delay_unit VDD VSS clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[13\]
+ clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[14\] clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[13\].delay_unit/mid
+ VDD VSS sky130_mm_sc_hd_dlyPoly5ns
XFILLER_10_284 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XFILLER_6_244 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XFILLER_1_32 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[1\].delay_unit VDD VSS clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[1\]
+ clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[2\] clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[1\].delay_unit/mid
+ VDD VSS sky130_mm_sc_hd_dlyPoly5ns
XFILLER_2_280 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
Xclkgen.delay_155ns_3.genblk1\[0\].bypass_enable VDD VSS clkgen.delay_155ns_3.genblk1\[0\].dly_binary.bypass_in
+ clkgen.delay_155ns_3.enable_dlycontrol_w clkgen.delay_155ns_3.bypass_enable_w\[0\]
+ VDD VSS sky130_fd_sc_hd__and2_1
XFILLER_12_302 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XFILLER_8_306 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
Xclkgen.delay_155ns_3.genblk1\[1\].dly_binary.out_mux VSS VDD clkgen.delay_155ns_3.genblk1\[1\].dly_binary.out
+ clkgen.delay_155ns_3.genblk1\[0\].dly_binary.out clkgen.delay_155ns_3.genblk1\[1\].dly_binary.bypass_in
+ clkgen.delay_155ns_3.genblk1\[1\].dly_binary.signal_w\[2\] VDD VSS sky130_fd_sc_hd__mux2_1
XPHY_4 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
Xclkgen.delay_155ns_3.genblk1\[3\].dly_binary.out_mux VSS VDD clkgen.delay_155ns_3.genblk1\[3\].dly_binary.out
+ clkgen.delay_155ns_3.genblk1\[2\].dly_binary.out clkgen.delay_155ns_3.genblk1\[3\].dly_binary.bypass_in
+ clkgen.delay_155ns_3.genblk1\[3\].dly_binary.signal_w\[8\] VDD VSS sky130_fd_sc_hd__mux2_1
XFILLER_1_323 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
Xedgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[4\].delay_unit VDD VSS edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[4\]
+ edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[5\] edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[4\].delay_unit/mid
+ VDD VSS sky130_mm_sc_hd_dlyPoly5ns
XFILLER_4_32 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
Xclkgen.delay_155ns_3.genblk1\[4\].control_invert VDD VSS clkgen.delay_155ns_3.bypass_enable_w\[4\]
+ dlycontrol3_in[4] VDD VSS sky130_fd_sc_hd__inv_2
Xclkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[6\].delay_unit VDD VSS clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[6\]
+ clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[7\] clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[6\].delay_unit/mid
+ VDD VSS sky130_mm_sc_hd_dlyPoly5ns
XFILLER_13_74 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XFILLER_9_242 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
XFILLER_9_275 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
Xedgedetect.dly_315ns_1.genblk1\[2\].dly_binary.and_bypass_switch VSS VDD edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.bypass_in
+ edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.signal_w\[0\] edgedetect.dly_315ns_1.genblk1\[1\].dly_binary.out
+ VDD VSS sky130_fd_sc_hd__and2b_1
XFILLER_13_282 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XANTENNA_clkgen.delay_155ns_2.genblk1\[4\].dly_binary.out_mux_S VSS VDD clkgen.delay_155ns_2.genblk1\[4\].dly_binary.bypass_in
+ VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_1_153 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
Xclkgen.delay_155ns_3.genblk1\[3\].dly_binary.genblk1\[2\].delay_unit VDD VSS clkgen.delay_155ns_3.genblk1\[3\].dly_binary.signal_w\[2\]
+ clkgen.delay_155ns_3.genblk1\[3\].dly_binary.signal_w\[3\] clkgen.delay_155ns_3.genblk1\[3\].dly_binary.genblk1\[2\].delay_unit/mid
+ VDD VSS sky130_mm_sc_hd_dlyPoly5ns
XANTENNA_clkgen.delay_155ns_1.genblk1\[0\].control_invert_A VSS VDD dlycontrol1_in[0]
+ VDD VSS sky130_fd_sc_hd__diode_2
Xclkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[0\].delay_unit VDD VSS clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[0\]
+ clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[1\] clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[0\].delay_unit/mid
+ VDD VSS sky130_mm_sc_hd_dlyPoly5ns
XFILLER_3_259 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XFILLER_2_292 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
Xedgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[11\].delay_unit VDD VSS edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[11\]
+ edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[12\] edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[11\].delay_unit/mid
+ VDD VSS sky130_mm_sc_hd_dlyPoly5ns
XFILLER_12_314 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XFILLER_0_229 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[11\].delay_unit VDD VSS clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[11\]
+ clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[12\] clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[11\].delay_unit/mid
+ VDD VSS sky130_mm_sc_hd_dlyPoly5ns
Xedgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[9\].delay_unit VDD VSS edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[9\]
+ edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[10\] edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[9\].delay_unit/mid
+ VDD VSS sky130_mm_sc_hd_dlyPoly5ns
XPHY_5 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XFILLER_7_32 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XFILLER_16_63 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_3.genblk1\[3\].dly_binary.genblk1\[7\].delay_unit VDD VSS clkgen.delay_155ns_3.genblk1\[3\].dly_binary.signal_w\[7\]
+ clkgen.delay_155ns_3.genblk1\[3\].dly_binary.signal_w\[8\] clkgen.delay_155ns_3.genblk1\[3\].dly_binary.genblk1\[7\].delay_unit/mid
+ VDD VSS sky130_mm_sc_hd_dlyPoly5ns
Xedgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[12\].delay_unit VDD VSS edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[12\]
+ edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[13\] edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[12\].delay_unit/mid
+ VDD VSS sky130_mm_sc_hd_dlyPoly5ns
XFILLER_1_335 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
Xclkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[5\].delay_unit VDD VSS clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[5\]
+ clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[6\] clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[5\].delay_unit/mid
+ VDD VSS sky130_mm_sc_hd_dlyPoly5ns
XFILLER_4_173 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_2.genblk1\[3\].dly_binary.genblk1\[1\].delay_unit VDD VSS clkgen.delay_155ns_2.genblk1\[3\].dly_binary.signal_w\[1\]
+ clkgen.delay_155ns_2.genblk1\[3\].dly_binary.signal_w\[2\] clkgen.delay_155ns_2.genblk1\[3\].dly_binary.genblk1\[1\].delay_unit/mid
+ VDD VSS sky130_mm_sc_hd_dlyPoly5ns
XFILLER_13_31 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XFILLER_13_294 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XFILLER_1_187 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
Xedgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[16\].delay_unit VDD VSS edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[16\]
+ edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[17\] edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[16\].delay_unit/mid
+ VDD VSS sky130_mm_sc_hd_dlyPoly5ns
XFILLER_5_290 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_19_63 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XANTENNA_clkgen.delay_155ns_2.genblk1\[2\].dly_binary.out_mux_S VSS VDD clkgen.delay_155ns_2.genblk1\[2\].dly_binary.bypass_in
+ VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_12_326 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
Xclkgen.delay_155ns_1.genblk1\[0\].control_invert VDD VSS clkgen.delay_155ns_1.bypass_enable_w\[0\]
+ dlycontrol1_in[0] VDD VSS sky130_fd_sc_hd__inv_2
Xedgedetect.dly_315ns_1.genblk1\[3\].dly_binary.genblk1\[4\].delay_unit VDD VSS edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.signal_w\[4\]
+ edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.signal_w\[5\] edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.genblk1\[4\].delay_unit/mid
+ VDD VSS sky130_mm_sc_hd_dlyPoly5ns
XPHY_6 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
Xclkgen.delay_155ns_2.genblk1\[3\].dly_binary.genblk1\[6\].delay_unit VDD VSS clkgen.delay_155ns_2.genblk1\[3\].dly_binary.signal_w\[6\]
+ clkgen.delay_155ns_2.genblk1\[3\].dly_binary.signal_w\[7\] clkgen.delay_155ns_2.genblk1\[3\].dly_binary.genblk1\[6\].delay_unit/mid
+ VDD VSS sky130_mm_sc_hd_dlyPoly5ns
XFILLER_12_145 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_3.genblk1\[2\].dly_binary.genblk1\[2\].delay_unit VDD VSS clkgen.delay_155ns_3.genblk1\[2\].dly_binary.signal_w\[2\]
+ clkgen.delay_155ns_3.genblk1\[2\].dly_binary.signal_w\[3\] clkgen.delay_155ns_3.genblk1\[2\].dly_binary.genblk1\[2\].delay_unit/mid
+ VDD VSS sky130_mm_sc_hd_dlyPoly5ns
Xedgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[23\].delay_unit VDD VSS edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[23\]
+ edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[24\] edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[23\].delay_unit/mid
+ VDD VSS sky130_mm_sc_hd_dlyPoly5ns
Xedgedetect.dly_315ns_1.genblk1\[3\].dly_binary.and_bypass_switch VSS VDD edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.bypass_in
+ edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.signal_w\[0\] edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.out
+ VDD VSS sky130_fd_sc_hd__and2b_1
XFILLER_17_237 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_1.genblk1\[3\].dly_binary.genblk1\[0\].delay_unit VDD VSS clkgen.delay_155ns_1.genblk1\[3\].dly_binary.signal_w\[0\]
+ clkgen.delay_155ns_1.genblk1\[3\].dly_binary.signal_w\[1\] clkgen.delay_155ns_1.genblk1\[3\].dly_binary.genblk1\[0\].delay_unit/mid
+ VDD VSS sky130_mm_sc_hd_dlyPoly5ns
XFILLER_9_233 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XFILLER_3_239 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XFILLER_2_261 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_1.genblk1\[3\].dly_binary.genblk1\[5\].delay_unit VDD VSS clkgen.delay_155ns_1.genblk1\[3\].dly_binary.signal_w\[5\]
+ clkgen.delay_155ns_1.genblk1\[3\].dly_binary.signal_w\[6\] clkgen.delay_155ns_1.genblk1\[3\].dly_binary.genblk1\[5\].delay_unit/mid
+ VDD VSS sky130_mm_sc_hd_dlyPoly5ns
Xedgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[28\].delay_unit VDD VSS edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[28\]
+ edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[29\] edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[28\].delay_unit/mid
+ VDD VSS sky130_mm_sc_hd_dlyPoly5ns
XFILLER_15_187 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
Xedgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[30\].delay_unit VDD VSS edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[30\]
+ edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[31\] edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[30\].delay_unit/mid
+ VDD VSS sky130_mm_sc_hd_dlyPoly5ns
XFILLER_12_338 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XPHY_7 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
Xclkgen.delay_155ns_2.genblk1\[2\].dly_binary.genblk1\[1\].delay_unit VDD VSS clkgen.delay_155ns_2.genblk1\[2\].dly_binary.signal_w\[1\]
+ clkgen.delay_155ns_2.genblk1\[2\].dly_binary.signal_w\[2\] clkgen.delay_155ns_2.genblk1\[2\].dly_binary.genblk1\[1\].delay_unit/mid
+ VDD VSS sky130_mm_sc_hd_dlyPoly5ns
XFILLER_16_32 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
XFILLER_17_227 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XFILLER_9_223 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XFILLER_10_244 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XFILLER_19_32 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XFILLER_2_273 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
XFILLER_18_185 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
Xedgedetect.dly_315ns_1.enablebuffer VDD VSS enable_dlycontrol_in edgedetect.dly_315ns_1.enable_dlycontrol_w
+ VDD VSS sky130_fd_sc_hd__buf_4
Xclkgen.delay_155ns_1.genblk1\[2\].dly_binary.genblk1\[0\].delay_unit VDD VSS clkgen.delay_155ns_1.genblk1\[2\].dly_binary.signal_w\[0\]
+ clkgen.delay_155ns_1.genblk1\[2\].dly_binary.signal_w\[1\] clkgen.delay_155ns_1.genblk1\[2\].dly_binary.genblk1\[0\].delay_unit/mid
+ VDD VSS sky130_mm_sc_hd_dlyPoly5ns
Xedgedetect.dly_315ns_1.genblk1\[4\].dly_binary.and_bypass_switch VSS VDD edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.bypass_in
+ edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[0\] edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.out
+ VDD VSS sky130_fd_sc_hd__and2b_1
XPHY_8 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XFILLER_4_302 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_7_195 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XANTENNA_edgedetect.dly_315ns_1.genblk1\[4\].control_invert_A VSS VDD dlycontrol4_in[4]
+ VDD VSS sky130_fd_sc_hd__diode_2
Xclkgen.delay_155ns_1.enablebuffer VDD VSS enable_dlycontrol_in clkgen.delay_155ns_1.enable_dlycontrol_w
+ VDD VSS sky130_fd_sc_hd__buf_4
Xedgedetect.dly_315ns_1.genblk1\[3\].bypass_enable VDD VSS edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.bypass_in
+ edgedetect.dly_315ns_1.enable_dlycontrol_w edgedetect.dly_315ns_1.bypass_enable_w\[3\]
+ VDD VSS sky130_fd_sc_hd__and2_1
XFILLER_13_275 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XFILLER_18_312 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_2.genblk1\[1\].dly_binary.genblk1\[1\].delay_unit VDD VSS clkgen.delay_155ns_2.genblk1\[1\].dly_binary.signal_w\[1\]
+ clkgen.delay_155ns_2.genblk1\[1\].dly_binary.signal_w\[2\] clkgen.delay_155ns_2.genblk1\[1\].dly_binary.genblk1\[1\].delay_unit/mid
+ VDD VSS sky130_mm_sc_hd_dlyPoly5ns
Xclkgen.delay_155ns_2.genblk1\[1\].control_invert VDD VSS clkgen.delay_155ns_2.bypass_enable_w\[1\]
+ dlycontrol2_in[1] VDD VSS sky130_fd_sc_hd__inv_2
XFILLER_15_304 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
XFILLER_15_337 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
XFILLER_2_230 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_1.genblk1\[4\].bypass_enable VDD VSS clkgen.delay_155ns_1.genblk1\[4\].dly_binary.bypass_in
+ clkgen.delay_155ns_1.enable_dlycontrol_w clkgen.delay_155ns_1.bypass_enable_w\[4\]
+ VDD VSS sky130_fd_sc_hd__and2_1
Xclkgen.delay_155ns_3.genblk1\[0\].dly_binary.and_bypass_switch VSS VDD clkgen.delay_155ns_3.genblk1\[0\].dly_binary.bypass_in
+ clkgen.delay_155ns_3.genblk1\[0\].dly_binary.signal_w\[0\] clkgen.delay_155ns_3.genblk1\[0\].dly_binary.in
+ VDD VSS sky130_fd_sc_hd__and2b_1
XFILLER_15_156 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XPHY_9 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
Xclkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[11\].delay_unit VDD VSS clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[11\]
+ clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[12\] clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[11\].delay_unit/mid
+ VDD VSS sky130_mm_sc_hd_dlyPoly5ns
XANTENNA_edgedetect.dly_315ns_1.genblk1\[0\].dly_binary.out_mux_S VSS VDD edgedetect.dly_315ns_1.genblk1\[0\].dly_binary.bypass_in
+ VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_12_104 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XANTENNA_clkgen.delay_155ns_1.enablebuffer_A VSS VDD enable_dlycontrol_in VDD VSS
+ sky130_fd_sc_hd__diode_2
XFILLER_4_314 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_19_292 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XANTENNA_clkgen.delay_155ns_2.genblk1\[2\].dly_binary.and_bypass_switch_A_N VSS VDD
+ clkgen.delay_155ns_2.genblk1\[2\].dly_binary.bypass_in VDD VSS sky130_fd_sc_hd__diode_2
Xedgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[0\].delay_unit VDD VSS edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[0\]
+ edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[1\] edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[0\].delay_unit/mid
+ VDD VSS sky130_mm_sc_hd_dlyPoly5ns
XFILLER_1_125 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_1.genblk1\[1\].dly_binary.genblk1\[0\].delay_unit VDD VSS clkgen.delay_155ns_1.genblk1\[1\].dly_binary.signal_w\[0\]
+ clkgen.delay_155ns_1.genblk1\[1\].dly_binary.signal_w\[1\] clkgen.delay_155ns_1.genblk1\[1\].dly_binary.genblk1\[0\].delay_unit/mid
+ VDD VSS sky130_mm_sc_hd_dlyPoly5ns
XFILLER_18_324 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_10_58 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
Xedgedetect.dly_315ns_1.genblk1\[5\].dly_binary.and_bypass_switch VSS VDD edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.bypass_in
+ edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[0\] edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.out
+ VDD VSS sky130_fd_sc_hd__and2b_1
XFILLER_12_308 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
Xedgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[5\].delay_unit VDD VSS edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[5\]
+ edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[6\] edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[5\].delay_unit/mid
+ VDD VSS sky130_mm_sc_hd_dlyPoly5ns
XANTENNA_clkgen.delay_155ns_1.genblk1\[4\].dly_binary.out_mux_A1 VSS VDD clkgen.delay_155ns_1.genblk1\[3\].dly_binary.out
+ VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_4_326 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
Xclkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[3\].delay_unit VDD VSS clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[3\]
+ clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[4\] clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[3\].delay_unit/mid
+ VDD VSS sky130_mm_sc_hd_dlyPoly5ns
Xedgedetect.dly_315ns_1.genblk1\[2\].control_invert VDD VSS edgedetect.dly_315ns_1.bypass_enable_w\[2\]
+ dlycontrol4_in[2] VDD VSS sky130_fd_sc_hd__inv_2
XFILLER_1_307 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XFILLER_4_167 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XFILLER_13_288 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XFILLER_5_81 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XFILLER_10_214 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XFILLER_18_336 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XFILLER_5_284 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_2.genblk1\[0\].bypass_enable VDD VSS clkgen.delay_155ns_2.genblk1\[0\].dly_binary.bypass_in
+ clkgen.delay_155ns_2.enable_dlycontrol_w clkgen.delay_155ns_2.bypass_enable_w\[0\]
+ VDD VSS sky130_fd_sc_hd__and2_1
XFILLER_5_240 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_3.genblk1\[1\].dly_binary.and_bypass_switch VSS VDD clkgen.delay_155ns_3.genblk1\[1\].dly_binary.bypass_in
+ clkgen.delay_155ns_3.genblk1\[1\].dly_binary.signal_w\[0\] clkgen.delay_155ns_3.genblk1\[0\].dly_binary.out
+ VDD VSS sky130_fd_sc_hd__and2b_1
Xclkgen.delay_155ns_3.genblk1\[1\].bypass_enable VDD VSS clkgen.delay_155ns_3.genblk1\[1\].dly_binary.bypass_in
+ clkgen.delay_155ns_3.enable_dlycontrol_w clkgen.delay_155ns_3.bypass_enable_w\[1\]
+ VDD VSS sky130_fd_sc_hd__and2_1
XFILLER_2_243 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XANTENNA_clkgen.delay_155ns_3.genblk1\[4\].control_invert_A VSS VDD dlycontrol3_in[4]
+ VDD VSS sky130_fd_sc_hd__diode_2
Xclkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[8\].delay_unit VDD VSS clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[8\]
+ clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[9\] clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[8\].delay_unit/mid
+ VDD VSS sky130_mm_sc_hd_dlyPoly5ns
Xclkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[14\].delay_unit VDD VSS clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[14\]
+ clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[15\] clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[14\].delay_unit/mid
+ VDD VSS sky130_mm_sc_hd_dlyPoly5ns
XFILLER_15_125 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
Xclkgen.delay_155ns_2.genblk1\[0\].dly_binary.and_bypass_switch VSS VDD clkgen.delay_155ns_2.genblk1\[0\].dly_binary.bypass_in
+ clkgen.delay_155ns_2.genblk1\[0\].dly_binary.signal_w\[0\] clkgen.clk_dig_out VDD
+ VSS sky130_fd_sc_hd__and2b_1
Xedgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[0\].delay_unit VDD VSS edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[0\]
+ edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[1\] edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[0\].delay_unit/mid
+ VDD VSS sky130_mm_sc_hd_dlyPoly5ns
Xclkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[2\].delay_unit VDD VSS clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[2\]
+ clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[3\] clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[2\].delay_unit/mid
+ VDD VSS sky130_mm_sc_hd_dlyPoly5ns
XFILLER_12_117 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XFILLER_4_338 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
Xclkgen.delay_155ns_1.genblk1\[0\].dly_binary.genblk1\[0\].delay_unit VDD VSS clkgen.delay_155ns_1.genblk1\[0\].dly_binary.signal_w\[0\]
+ clkgen.delay_155ns_1.genblk1\[0\].dly_binary.signal_w\[1\] clkgen.delay_155ns_1.genblk1\[0\].dly_binary.genblk1\[0\].delay_unit/mid
+ VDD VSS sky130_mm_sc_hd_dlyPoly5ns
XANTENNA_clkgen.delay_155ns_1.genblk1\[0\].dly_binary.and_bypass_switch_A_N VSS VDD
+ clkgen.delay_155ns_1.genblk1\[0\].dly_binary.bypass_in VDD VSS sky130_fd_sc_hd__diode_2
Xclkgen.delay_155ns_3.genblk1\[2\].control_invert VDD VSS clkgen.delay_155ns_3.bypass_enable_w\[2\]
+ dlycontrol3_in[2] VDD VSS sky130_fd_sc_hd__inv_2
XFILLER_13_245 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XFILLER_13_59 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XFILLER_0_182 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XANTENNA_clkgen.delay_155ns_2.genblk1\[1\].dly_binary.and_bypass_switch_B VSS VDD
+ clkgen.delay_155ns_2.genblk1\[0\].dly_binary.out VDD VSS sky130_fd_sc_hd__diode_2
Xedgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[5\].delay_unit VDD VSS edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[5\]
+ edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[6\] edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[5\].delay_unit/mid
+ VDD VSS sky130_mm_sc_hd_dlyPoly5ns
Xclkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[7\].delay_unit VDD VSS clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[7\]
+ clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[8\] clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[7\].delay_unit/mid
+ VDD VSS sky130_mm_sc_hd_dlyPoly5ns
XFILLER_10_16 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XFILLER_18_156 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XFILLER_2_255 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_3.genblk1\[3\].dly_binary.genblk1\[3\].delay_unit VDD VSS clkgen.delay_155ns_3.genblk1\[3\].dly_binary.signal_w\[3\]
+ clkgen.delay_155ns_3.genblk1\[3\].dly_binary.signal_w\[4\] clkgen.delay_155ns_3.genblk1\[3\].dly_binary.genblk1\[3\].delay_unit/mid
+ VDD VSS sky130_mm_sc_hd_dlyPoly5ns
XFILLER_2_94 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
XFILLER_7_303 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
Xclkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[1\].delay_unit VDD VSS clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[1\]
+ clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[2\] clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[1\].delay_unit/mid
+ VDD VSS sky130_mm_sc_hd_dlyPoly5ns
XFILLER_11_151 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_2.genblk1\[1\].dly_binary.out_mux VSS VDD clkgen.delay_155ns_2.genblk1\[1\].dly_binary.out
+ clkgen.delay_155ns_2.genblk1\[0\].dly_binary.out clkgen.delay_155ns_2.genblk1\[1\].dly_binary.bypass_in
+ clkgen.delay_155ns_2.genblk1\[1\].dly_binary.signal_w\[2\] VDD VSS sky130_fd_sc_hd__mux2_1
Xedgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[12\].delay_unit VDD VSS edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[12\]
+ edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[13\] edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[12\].delay_unit/mid
+ VDD VSS sky130_mm_sc_hd_dlyPoly5ns
XFILLER_4_125 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[12\].delay_unit VDD VSS clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[12\]
+ clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[13\] clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[12\].delay_unit/mid
+ VDD VSS sky130_mm_sc_hd_dlyPoly5ns
Xclkgen.delay_155ns_2.genblk1\[3\].dly_binary.out_mux VSS VDD clkgen.delay_155ns_2.genblk1\[3\].dly_binary.out
+ clkgen.delay_155ns_2.genblk1\[2\].dly_binary.out clkgen.delay_155ns_2.genblk1\[3\].dly_binary.bypass_in
+ clkgen.delay_155ns_2.genblk1\[3\].dly_binary.signal_w\[8\] VDD VSS sky130_fd_sc_hd__mux2_1
Xclkgen.delay_155ns_3.genblk1\[2\].dly_binary.and_bypass_switch VSS VDD clkgen.delay_155ns_3.genblk1\[2\].dly_binary.bypass_in
+ clkgen.delay_155ns_3.genblk1\[2\].dly_binary.signal_w\[0\] clkgen.delay_155ns_3.genblk1\[1\].dly_binary.out
+ VDD VSS sky130_fd_sc_hd__and2b_1
XFILLER_0_194 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
Xedgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[13\].delay_unit VDD VSS edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[13\]
+ edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[14\] edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[13\].delay_unit/mid
+ VDD VSS sky130_mm_sc_hd_dlyPoly5ns
XFILLER_12_290 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XFILLER_8_272 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
Xclkgen.delay_155ns_2.genblk1\[1\].dly_binary.and_bypass_switch VSS VDD clkgen.delay_155ns_2.genblk1\[1\].dly_binary.bypass_in
+ clkgen.delay_155ns_2.genblk1\[1\].dly_binary.signal_w\[0\] clkgen.delay_155ns_2.genblk1\[0\].dly_binary.out
+ VDD VSS sky130_fd_sc_hd__and2b_1
Xedgedetect.dly_315ns_1.genblk1\[3\].dly_binary.genblk1\[0\].delay_unit VDD VSS edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.signal_w\[0\]
+ edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.signal_w\[1\] edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.genblk1\[0\].delay_unit/mid
+ VDD VSS sky130_mm_sc_hd_dlyPoly5ns
XFILLER_5_231 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[6\].delay_unit VDD VSS clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[6\]
+ clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[7\] clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[6\].delay_unit/mid
+ VDD VSS sky130_mm_sc_hd_dlyPoly5ns
Xclkgen.delay_155ns_2.genblk1\[3\].dly_binary.genblk1\[2\].delay_unit VDD VSS clkgen.delay_155ns_2.genblk1\[3\].dly_binary.signal_w\[2\]
+ clkgen.delay_155ns_2.genblk1\[3\].dly_binary.signal_w\[3\] clkgen.delay_155ns_2.genblk1\[3\].dly_binary.genblk1\[2\].delay_unit/mid
+ VDD VSS sky130_mm_sc_hd_dlyPoly5ns
XFILLER_2_267 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XFILLER_2_223 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
Xedgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[17\].delay_unit VDD VSS edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[17\]
+ edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[18\] edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[17\].delay_unit/mid
+ VDD VSS sky130_mm_sc_hd_dlyPoly5ns
Xclkgen.delay_155ns_1.genblk1\[0\].dly_binary.and_bypass_switch VSS VDD clkgen.delay_155ns_1.genblk1\[0\].dly_binary.bypass_in
+ clkgen.delay_155ns_1.genblk1\[0\].dly_binary.signal_w\[0\] clkgen.delay_155ns_1.genblk1\[0\].dly_binary.in
+ VDD VSS sky130_fd_sc_hd__and2b_1
XFILLER_15_116 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XFILLER_11_300 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XFILLER_7_337 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
XFILLER_7_156 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XFILLER_19_274 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XFILLER_19_285 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
Xedgedetect.dly_315ns_1.genblk1\[3\].dly_binary.genblk1\[5\].delay_unit VDD VSS edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.signal_w\[5\]
+ edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.signal_w\[6\] edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.genblk1\[5\].delay_unit/mid
+ VDD VSS sky130_mm_sc_hd_dlyPoly5ns
XFILLER_16_244 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XFILLER_3_181 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_2.genblk1\[3\].dly_binary.genblk1\[7\].delay_unit VDD VSS clkgen.delay_155ns_2.genblk1\[3\].dly_binary.signal_w\[7\]
+ clkgen.delay_155ns_2.genblk1\[3\].dly_binary.signal_w\[8\] clkgen.delay_155ns_2.genblk1\[3\].dly_binary.genblk1\[7\].delay_unit/mid
+ VDD VSS sky130_mm_sc_hd_dlyPoly5ns
XANTENNA_edgedetect.dly_315ns_1.genblk1\[3\].control_invert_A VSS VDD dlycontrol4_in[3]
+ VDD VSS sky130_fd_sc_hd__diode_2
Xclkgen.delay_155ns_1.genblk1\[3\].control_invert VDD VSS clkgen.delay_155ns_1.bypass_enable_w\[3\]
+ dlycontrol1_in[3] VDD VSS sky130_fd_sc_hd__inv_2
XFILLER_13_236 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_3.genblk1\[2\].dly_binary.genblk1\[3\].delay_unit VDD VSS clkgen.delay_155ns_3.genblk1\[2\].dly_binary.signal_w\[3\]
+ clkgen.delay_155ns_3.genblk1\[2\].dly_binary.signal_w\[4\] clkgen.delay_155ns_3.genblk1\[2\].dly_binary.genblk1\[3\].delay_unit/mid
+ VDD VSS sky130_mm_sc_hd_dlyPoly5ns
Xedgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[24\].delay_unit VDD VSS edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[24\]
+ edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[25\] edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[24\].delay_unit/mid
+ VDD VSS sky130_mm_sc_hd_dlyPoly5ns
Xclkgen.delay_155ns_1.genblk1\[3\].dly_binary.genblk1\[1\].delay_unit VDD VSS clkgen.delay_155ns_1.genblk1\[3\].dly_binary.signal_w\[1\]
+ clkgen.delay_155ns_1.genblk1\[3\].dly_binary.signal_w\[2\] clkgen.delay_155ns_1.genblk1\[3\].dly_binary.genblk1\[1\].delay_unit/mid
+ VDD VSS sky130_mm_sc_hd_dlyPoly5ns
XFILLER_18_125 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XFILLER_2_63 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
Xedgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[29\].delay_unit VDD VSS edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[29\]
+ edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[30\] edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[29\].delay_unit/mid
+ VDD VSS sky130_mm_sc_hd_dlyPoly5ns
Xedgedetect.dly_315ns_1.genblk1\[2\].dly_binary.genblk1\[0\].delay_unit VDD VSS edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.signal_w\[0\]
+ edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.signal_w\[1\] edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.genblk1\[0\].delay_unit/mid
+ VDD VSS sky130_mm_sc_hd_dlyPoly5ns
Xclkgen.delay_155ns_3.genblk1\[3\].dly_binary.and_bypass_switch VSS VDD clkgen.delay_155ns_3.genblk1\[3\].dly_binary.bypass_in
+ clkgen.delay_155ns_3.genblk1\[3\].dly_binary.signal_w\[0\] clkgen.delay_155ns_3.genblk1\[2\].dly_binary.out
+ VDD VSS sky130_fd_sc_hd__and2b_1
Xclkgen.delay_155ns_1.genblk1\[3\].dly_binary.genblk1\[6\].delay_unit VDD VSS clkgen.delay_155ns_1.genblk1\[3\].dly_binary.signal_w\[6\]
+ clkgen.delay_155ns_1.genblk1\[3\].dly_binary.signal_w\[7\] clkgen.delay_155ns_1.genblk1\[3\].dly_binary.genblk1\[6\].delay_unit/mid
+ VDD VSS sky130_mm_sc_hd_dlyPoly5ns
Xedgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[31\].delay_unit VDD VSS edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[31\]
+ edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[32\] edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[31\].delay_unit/mid
+ VDD VSS sky130_mm_sc_hd_dlyPoly5ns
Xclkgen.delay_155ns_2.genblk1\[2\].dly_binary.genblk1\[2\].delay_unit VDD VSS clkgen.delay_155ns_2.genblk1\[2\].dly_binary.signal_w\[2\]
+ clkgen.delay_155ns_2.genblk1\[2\].dly_binary.signal_w\[3\] clkgen.delay_155ns_2.genblk1\[2\].dly_binary.genblk1\[2\].delay_unit/mid
+ VDD VSS sky130_mm_sc_hd_dlyPoly5ns
XFILLER_0_311 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
Xclkgen.delay_155ns_2.genblk1\[2\].dly_binary.and_bypass_switch VSS VDD clkgen.delay_155ns_2.genblk1\[2\].dly_binary.bypass_in
+ clkgen.delay_155ns_2.genblk1\[2\].dly_binary.signal_w\[0\] clkgen.delay_155ns_2.genblk1\[1\].dly_binary.out
+ VDD VSS sky130_fd_sc_hd__and2b_1
XFILLER_10_207 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XFILLER_18_318 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_1.genblk1\[1\].dly_binary.and_bypass_switch VSS VDD clkgen.delay_155ns_1.genblk1\[1\].dly_binary.bypass_in
+ clkgen.delay_155ns_1.genblk1\[1\].dly_binary.signal_w\[0\] clkgen.delay_155ns_1.genblk1\[0\].dly_binary.out
+ VDD VSS sky130_fd_sc_hd__and2b_1
XFILLER_14_94 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
XFILLER_5_222 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XFILLER_19_265 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XFILLER_19_298 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XFILLER_7_125 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
Xclkgen.delay_155ns_1.genblk1\[2\].dly_binary.genblk1\[1\].delay_unit VDD VSS clkgen.delay_155ns_1.genblk1\[2\].dly_binary.signal_w\[1\]
+ clkgen.delay_155ns_1.genblk1\[2\].dly_binary.signal_w\[2\] clkgen.delay_155ns_1.genblk1\[2\].dly_binary.genblk1\[1\].delay_unit/mid
+ VDD VSS sky130_mm_sc_hd_dlyPoly5ns
Xedgedetect.dly_315ns_1.genblk1\[4\].bypass_enable VDD VSS edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.bypass_in
+ edgedetect.dly_315ns_1.enable_dlycontrol_w edgedetect.dly_315ns_1.bypass_enable_w\[4\]
+ VDD VSS sky130_fd_sc_hd__and2_1
XFILLER_17_94 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XFILLER_0_323 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_13_227 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XANTENNA_clkgen.delay_155ns_2.genblk1\[4\].control_invert_A VSS VDD dlycontrol2_in[4]
+ VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_5_278 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_2.enablebuffer VDD VSS enable_dlycontrol_in clkgen.delay_155ns_2.enable_dlycontrol_w
+ VDD VSS sky130_fd_sc_hd__buf_4
XFILLER_2_237 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
Xedgedetect.dly_315ns_1.genblk1\[1\].dly_binary.genblk1\[0\].delay_unit VDD VSS edgedetect.dly_315ns_1.genblk1\[1\].dly_binary.signal_w\[0\]
+ edgedetect.dly_315ns_1.genblk1\[1\].dly_binary.signal_w\[1\] edgedetect.dly_315ns_1.genblk1\[1\].dly_binary.genblk1\[0\].delay_unit/mid
+ VDD VSS sky130_mm_sc_hd_dlyPoly5ns
XFILLER_2_32 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
Xclkgen.delay_155ns_3.genblk1\[4\].dly_binary.and_bypass_switch VSS VDD clkgen.delay_155ns_3.genblk1\[4\].dly_binary.bypass_in
+ clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[0\] clkgen.delay_155ns_3.genblk1\[3\].dly_binary.out
+ VDD VSS sky130_fd_sc_hd__and2b_1
XFILLER_14_185 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XANTENNA_clkgen.delay_155ns_3.genblk1\[3\].control_invert_A VSS VDD dlycontrol3_in[3]
+ VDD VSS sky130_fd_sc_hd__diode_2
Xclkgen.delay_155ns_2.genblk1\[4\].control_invert VDD VSS clkgen.delay_155ns_2.bypass_enable_w\[4\]
+ dlycontrol2_in[4] VDD VSS sky130_fd_sc_hd__inv_2
Xclkgen.delay_155ns_2.genblk1\[3\].dly_binary.and_bypass_switch VSS VDD clkgen.delay_155ns_2.genblk1\[3\].dly_binary.bypass_in
+ clkgen.delay_155ns_2.genblk1\[3\].dly_binary.signal_w\[0\] clkgen.delay_155ns_2.genblk1\[2\].dly_binary.out
+ VDD VSS sky130_fd_sc_hd__and2b_1
XFILLER_19_244 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XFILLER_8_75 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[12\].delay_unit VDD VSS clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[12\]
+ clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[13\] clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[12\].delay_unit/mid
+ VDD VSS sky130_mm_sc_hd_dlyPoly5ns
XFILLER_0_335 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
XANTENNA_clkgen.delay_155ns_2.genblk1\[1\].dly_binary.out_mux_A1 VSS VDD clkgen.delay_155ns_2.genblk1\[0\].dly_binary.out
+ VDD VSS sky130_fd_sc_hd__diode_2
Xclkgen.delay_155ns_1.genblk1\[2\].dly_binary.and_bypass_switch VSS VDD clkgen.delay_155ns_1.genblk1\[2\].dly_binary.bypass_in
+ clkgen.delay_155ns_1.genblk1\[2\].dly_binary.signal_w\[0\] clkgen.delay_155ns_1.genblk1\[1\].dly_binary.out
+ VDD VSS sky130_fd_sc_hd__and2b_1
XFILLER_15_291 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XFILLER_3_151 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
XFILLER_5_32 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XFILLER_14_63 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XFILLER_5_213 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
Xedgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[1\].delay_unit VDD VSS edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[1\]
+ edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[2\] edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[1\].delay_unit/mid
+ VDD VSS sky130_mm_sc_hd_dlyPoly5ns
XFILLER_4_290 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_2_249 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_1.genblk1\[1\].dly_binary.genblk1\[1\].delay_unit VDD VSS clkgen.delay_155ns_1.genblk1\[1\].dly_binary.signal_w\[1\]
+ clkgen.delay_155ns_1.genblk1\[1\].dly_binary.signal_w\[2\] clkgen.delay_155ns_1.genblk1\[1\].dly_binary.genblk1\[1\].delay_unit/mid
+ VDD VSS sky130_mm_sc_hd_dlyPoly5ns
XFILLER_1_271 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_11_315 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_3_311 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_19_256 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XFILLER_8_10 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XFILLER_8_32 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
Xedgedetect.dly_315ns_1.genblk1\[0\].control_invert VDD VSS edgedetect.dly_315ns_1.bypass_enable_w\[0\]
+ dlycontrol4_in[0] VDD VSS sky130_fd_sc_hd__inv_2
Xedgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[6\].delay_unit VDD VSS edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[6\]
+ edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[7\] edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[6\].delay_unit/mid
+ VDD VSS sky130_mm_sc_hd_dlyPoly5ns
XFILLER_17_63 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
Xclkgen.delay_155ns_1.genblk1\[0\].bypass_enable VDD VSS clkgen.delay_155ns_1.genblk1\[0\].dly_binary.bypass_in
+ clkgen.delay_155ns_1.enable_dlycontrol_w clkgen.delay_155ns_1.bypass_enable_w\[0\]
+ VDD VSS sky130_fd_sc_hd__and2_1
Xedgedetect.dly_315ns_1.genblk1\[0\].dly_binary.genblk1\[0\].delay_unit VDD VSS edgedetect.dly_315ns_1.genblk1\[0\].dly_binary.signal_w\[0\]
+ edgedetect.dly_315ns_1.genblk1\[0\].dly_binary.signal_w\[1\] edgedetect.dly_315ns_1.genblk1\[0\].dly_binary.genblk1\[0\].delay_unit/mid
+ VDD VSS sky130_mm_sc_hd_dlyPoly5ns
Xclkgen.delay_155ns_2.genblk1\[1\].bypass_enable VDD VSS clkgen.delay_155ns_2.genblk1\[1\].dly_binary.bypass_in
+ clkgen.delay_155ns_2.enable_dlycontrol_w clkgen.delay_155ns_2.bypass_enable_w\[1\]
+ VDD VSS sky130_fd_sc_hd__and2_1
XFILLER_10_3 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_3.genblk1\[2\].bypass_enable VDD VSS clkgen.delay_155ns_3.genblk1\[2\].dly_binary.bypass_in
+ clkgen.delay_155ns_3.enable_dlycontrol_w clkgen.delay_155ns_3.bypass_enable_w\[2\]
+ VDD VSS sky130_fd_sc_hd__and2_1
XFILLER_12_273 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
XFILLER_12_284 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XFILLER_8_244 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[4\].delay_unit VDD VSS clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[4\]
+ clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[5\] clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[4\].delay_unit/mid
+ VDD VSS sky130_mm_sc_hd_dlyPoly5ns
Xclkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[10\].delay_unit VDD VSS clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[10\]
+ clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[11\] clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[10\].delay_unit/mid
+ VDD VSS sky130_mm_sc_hd_dlyPoly5ns
Xedgedetect.dly_315ns_1.genblk1\[5\].control_invert VDD VSS edgedetect.dly_315ns_1.bypass_enable_w\[5\]
+ dlycontrol4_in[5] VDD VSS sky130_fd_sc_hd__inv_2
XFILLER_2_206 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XPHY_30 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XFILLER_1_283 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
Xclkgen.delay_155ns_2.genblk1\[4\].dly_binary.and_bypass_switch VSS VDD clkgen.delay_155ns_2.genblk1\[4\].dly_binary.bypass_in
+ clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[0\] clkgen.delay_155ns_2.genblk1\[3\].dly_binary.out
+ VDD VSS sky130_fd_sc_hd__and2b_1
XFILLER_11_327 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_11_32 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XANTENNA_clkgen.delay_155ns_1.genblk1\[3\].dly_binary.and_bypass_switch_A_N VSS VDD
+ clkgen.delay_155ns_1.genblk1\[3\].dly_binary.bypass_in VDD VSS sky130_fd_sc_hd__diode_2
Xclkgen.delay_155ns_1.genblk1\[3\].dly_binary.and_bypass_switch VSS VDD clkgen.delay_155ns_1.genblk1\[3\].dly_binary.bypass_in
+ clkgen.delay_155ns_1.genblk1\[3\].dly_binary.signal_w\[0\] clkgen.delay_155ns_1.genblk1\[2\].dly_binary.out
+ VDD VSS sky130_fd_sc_hd__and2b_1
XFILLER_11_179 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
XFILLER_19_213 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XFILLER_8_88 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XFILLER_3_323 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
Xclkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[9\].delay_unit VDD VSS clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[9\]
+ clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[10\] clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[9\].delay_unit/mid
+ VDD VSS sky130_mm_sc_hd_dlyPoly5ns
XFILLER_8_44 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
Xclkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[15\].delay_unit VDD VSS clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[15\]
+ clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[16\] clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[15\].delay_unit/mid
+ VDD VSS sky130_mm_sc_hd_dlyPoly5ns
XANTENNA_edgedetect.dly_315ns_1.genblk1\[1\].dly_binary.out_mux_A1 VSS VDD edgedetect.dly_315ns_1.genblk1\[0\].dly_binary.out
+ VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_0_304 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
Xedgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[1\].delay_unit VDD VSS edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[1\]
+ edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[2\] edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[1\].delay_unit/mid
+ VDD VSS sky130_mm_sc_hd_dlyPoly5ns
Xclkgen.delay_155ns_3.genblk1\[0\].control_invert VDD VSS clkgen.delay_155ns_3.bypass_enable_w\[0\]
+ dlycontrol3_in[0] VDD VSS sky130_fd_sc_hd__inv_2
Xclkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[3\].delay_unit VDD VSS clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[3\]
+ clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[4\] clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[3\].delay_unit/mid
+ VDD VSS sky130_mm_sc_hd_dlyPoly5ns
XANTENNA_clkgen.delay_155ns_1.genblk1\[3\].dly_binary.out_mux_A0 VSS VDD clkgen.delay_155ns_1.genblk1\[3\].dly_binary.signal_w\[8\]
+ VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA_edgedetect.dly_315ns_1.genblk1\[2\].control_invert_A VSS VDD dlycontrol4_in[2]
+ VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_12_296 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XFILLER_14_32 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
XPHY_20 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XPHY_31 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XFILLER_1_295 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_11_306 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XFILLER_11_339 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
Xedgedetect.dly_315ns_1.genblk1\[1\].dly_binary.out_mux VSS VDD edgedetect.dly_315ns_1.genblk1\[1\].dly_binary.out
+ edgedetect.dly_315ns_1.genblk1\[0\].dly_binary.out edgedetect.dly_315ns_1.genblk1\[1\].dly_binary.bypass_in
+ edgedetect.dly_315ns_1.genblk1\[1\].dly_binary.signal_w\[2\] VDD VSS sky130_fd_sc_hd__mux2_1
Xedgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[6\].delay_unit VDD VSS edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[6\]
+ edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[7\] edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[6\].delay_unit/mid
+ VDD VSS sky130_mm_sc_hd_dlyPoly5ns
Xclkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[8\].delay_unit VDD VSS clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[8\]
+ clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[9\] clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[8\].delay_unit/mid
+ VDD VSS sky130_mm_sc_hd_dlyPoly5ns
Xedgedetect.dly_315ns_1.genblk1\[3\].dly_binary.out_mux VSS VDD edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.out
+ edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.out edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.bypass_in
+ edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.signal_w\[8\] VDD VSS sky130_fd_sc_hd__mux2_1
Xclkgen.delay_155ns_3.genblk1\[3\].dly_binary.genblk1\[4\].delay_unit VDD VSS clkgen.delay_155ns_3.genblk1\[3\].dly_binary.signal_w\[4\]
+ clkgen.delay_155ns_3.genblk1\[3\].dly_binary.signal_w\[5\] clkgen.delay_155ns_3.genblk1\[3\].dly_binary.genblk1\[4\].delay_unit/mid
+ VDD VSS sky130_mm_sc_hd_dlyPoly5ns
XANTENNA_inbuf_2_A VSS VDD start_conv_in VDD VSS sky130_fd_sc_hd__diode_2
Xedgedetect.dly_315ns_1.genblk1\[5\].dly_binary.out_mux VSS VDD edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.out
+ edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.out edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.bypass_in
+ edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[32\] VDD VSS sky130_fd_sc_hd__mux2_1
XFILLER_3_335 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XFILLER_17_32 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[2\].delay_unit VDD VSS clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[2\]
+ clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[3\] clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[2\].delay_unit/mid
+ VDD VSS sky130_mm_sc_hd_dlyPoly5ns
XANTENNA_clkgen.delay_155ns_1.genblk1\[3\].dly_binary.out_mux_S VSS VDD clkgen.delay_155ns_1.genblk1\[3\].dly_binary.bypass_in
+ VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_0_146 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
Xedgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[13\].delay_unit VDD VSS edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[13\]
+ edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[14\] edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[13\].delay_unit/mid
+ VDD VSS sky130_mm_sc_hd_dlyPoly5ns
XFILLER_5_13 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XFILLER_5_68 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[13\].delay_unit VDD VSS clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[13\]
+ clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[14\] clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[13\].delay_unit/mid
+ VDD VSS sky130_mm_sc_hd_dlyPoly5ns
XFILLER_5_249 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XPHY_21 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XPHY_32 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XPHY_10 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
Xclkgen.delay_155ns_1.genblk1\[4\].dly_binary.and_bypass_switch VSS VDD clkgen.delay_155ns_1.genblk1\[4\].dly_binary.bypass_in
+ clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[0\] clkgen.delay_155ns_1.genblk1\[3\].dly_binary.out
+ VDD VSS sky130_fd_sc_hd__and2b_1
Xedgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[14\].delay_unit VDD VSS edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[14\]
+ edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[15\] edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[14\].delay_unit/mid
+ VDD VSS sky130_mm_sc_hd_dlyPoly5ns
Xedgedetect.dly_315ns_1.genblk1\[3\].dly_binary.genblk1\[1\].delay_unit VDD VSS edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.signal_w\[1\]
+ edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.signal_w\[2\] edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.genblk1\[1\].delay_unit/mid
+ VDD VSS sky130_mm_sc_hd_dlyPoly5ns
XFILLER_11_89 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
Xclkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[7\].delay_unit VDD VSS clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[7\]
+ clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[8\] clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[7\].delay_unit/mid
+ VDD VSS sky130_mm_sc_hd_dlyPoly5ns
Xoutbuf_1 VSS VDD clkgen.clk_dig_out clk_dig_out VDD VSS sky130_fd_sc_hd__bufbuf_8
XFILLER_14_156 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_2.genblk1\[3\].dly_binary.genblk1\[3\].delay_unit VDD VSS clkgen.delay_155ns_2.genblk1\[3\].dly_binary.signal_w\[3\]
+ clkgen.delay_155ns_2.genblk1\[3\].dly_binary.signal_w\[4\] clkgen.delay_155ns_2.genblk1\[3\].dly_binary.genblk1\[3\].delay_unit/mid
+ VDD VSS sky130_mm_sc_hd_dlyPoly5ns
XANTENNA_edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[0\].delay_unit_in
+ VSS VDD edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[0\] VDD VSS sky130_fd_sc_hd__diode_2
Xedgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[18\].delay_unit VDD VSS edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[18\]
+ edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[19\] edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[18\].delay_unit/mid
+ VDD VSS sky130_mm_sc_hd_dlyPoly5ns
XANTENNA_clkgen.delay_155ns_1.genblk1\[4\].control_invert_A VSS VDD dlycontrol1_in[4]
+ VDD VSS sky130_fd_sc_hd__diode_2
Xedgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[20\].delay_unit VDD VSS edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[20\]
+ edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[21\] edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[20\].delay_unit/mid
+ VDD VSS sky130_mm_sc_hd_dlyPoly5ns
XFILLER_15_284 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_1.genblk1\[1\].control_invert VDD VSS clkgen.delay_155ns_1.bypass_enable_w\[1\]
+ dlycontrol1_in[1] VDD VSS sky130_fd_sc_hd__inv_2
Xclkgen.delay_155ns_1.genblk1\[1\].dly_binary.out_mux VSS VDD clkgen.delay_155ns_1.genblk1\[1\].dly_binary.out
+ clkgen.delay_155ns_1.genblk1\[0\].dly_binary.out clkgen.delay_155ns_1.genblk1\[1\].dly_binary.bypass_in
+ clkgen.delay_155ns_1.genblk1\[1\].dly_binary.signal_w\[2\] VDD VSS sky130_fd_sc_hd__mux2_1
XANTENNA_edgedetect.nor1_B_N VSS VDD edgedetect.dly_315ns_1.genblk1\[0\].dly_binary.in
+ VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_0_136 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_1.genblk1\[3\].dly_binary.out_mux VSS VDD clkgen.delay_155ns_1.genblk1\[3\].dly_binary.out
+ clkgen.delay_155ns_1.genblk1\[2\].dly_binary.out clkgen.delay_155ns_1.genblk1\[3\].dly_binary.bypass_in
+ clkgen.delay_155ns_1.genblk1\[3\].dly_binary.signal_w\[8\] VDD VSS sky130_fd_sc_hd__mux2_1
Xedgedetect.dly_315ns_1.genblk1\[3\].dly_binary.genblk1\[6\].delay_unit VDD VSS edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.signal_w\[6\]
+ edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.signal_w\[7\] edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.genblk1\[6\].delay_unit/mid
+ VDD VSS sky130_mm_sc_hd_dlyPoly5ns
XANTENNA_clkgen.delay_155ns_2.genblk1\[3\].control_invert_A VSS VDD dlycontrol2_in[3]
+ VDD VSS sky130_fd_sc_hd__diode_2
XPHY_33 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XPHY_22 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XPHY_11 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XFILLER_17_198 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XFILLER_1_231 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XFILLER_1_253 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
Xedgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[25\].delay_unit VDD VSS edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[25\]
+ edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[26\] edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[25\].delay_unit/mid
+ VDD VSS sky130_mm_sc_hd_dlyPoly5ns
Xoutbuf_2 VSS VDD clkgen.clk_comp_out clk_comp_out VDD VSS sky130_fd_sc_hd__bufbuf_8
Xclkgen.delay_155ns_1.genblk1\[3\].dly_binary.genblk1\[2\].delay_unit VDD VSS clkgen.delay_155ns_1.genblk1\[3\].dly_binary.signal_w\[2\]
+ clkgen.delay_155ns_1.genblk1\[3\].dly_binary.signal_w\[3\] clkgen.delay_155ns_1.genblk1\[3\].dly_binary.genblk1\[2\].delay_unit/mid
+ VDD VSS sky130_mm_sc_hd_dlyPoly5ns
XFILLER_6_334 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
XANTENNA_clkgen.delay_155ns_3.genblk1\[2\].control_invert_A VSS VDD dlycontrol3_in[2]
+ VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_6_120 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XFILLER_16_208 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XFILLER_12_266 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
Xedgedetect.dly_315ns_1.genblk1\[2\].dly_binary.genblk1\[1\].delay_unit VDD VSS edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.signal_w\[1\]
+ edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.signal_w\[2\] edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.genblk1\[1\].delay_unit/mid
+ VDD VSS sky130_mm_sc_hd_dlyPoly5ns
Xclkgen.delay_155ns_1.genblk1\[3\].dly_binary.genblk1\[7\].delay_unit VDD VSS clkgen.delay_155ns_1.genblk1\[3\].dly_binary.signal_w\[7\]
+ clkgen.delay_155ns_1.genblk1\[3\].dly_binary.signal_w\[8\] clkgen.delay_155ns_1.genblk1\[3\].dly_binary.genblk1\[7\].delay_unit/mid
+ VDD VSS sky130_mm_sc_hd_dlyPoly5ns
XFILLER_17_303 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
Xclkgen.delay_155ns_2.genblk1\[2\].dly_binary.genblk1\[3\].delay_unit VDD VSS clkgen.delay_155ns_2.genblk1\[2\].dly_binary.signal_w\[3\]
+ clkgen.delay_155ns_2.genblk1\[2\].dly_binary.signal_w\[4\] clkgen.delay_155ns_2.genblk1\[2\].dly_binary.genblk1\[3\].delay_unit/mid
+ VDD VSS sky130_mm_sc_hd_dlyPoly5ns
XFILLER_4_284 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XFILLER_4_262 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XPHY_12 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XFILLER_14_306 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XPHY_23 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XPHY_34 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XFILLER_1_243 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
Xoutbuf_3 VSS VDD sample_p_1 sample_p_out VDD VSS sky130_fd_sc_hd__bufbuf_8
XFILLER_14_125 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_3.genblk1\[0\].dly_binary.out_mux VSS VDD clkgen.delay_155ns_3.genblk1\[0\].dly_binary.out
+ clkgen.delay_155ns_3.genblk1\[0\].dly_binary.in clkgen.delay_155ns_3.genblk1\[0\].dly_binary.bypass_in
+ clkgen.delay_155ns_3.genblk1\[0\].dly_binary.signal_w\[1\] VDD VSS sky130_fd_sc_hd__mux2_1
XFILLER_9_151 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XFILLER_9_195 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_3.genblk1\[2\].dly_binary.out_mux VSS VDD clkgen.delay_155ns_3.genblk1\[2\].dly_binary.out
+ clkgen.delay_155ns_3.genblk1\[1\].dly_binary.out clkgen.delay_155ns_3.genblk1\[2\].dly_binary.bypass_in
+ clkgen.delay_155ns_3.genblk1\[2\].dly_binary.signal_w\[4\] VDD VSS sky130_fd_sc_hd__mux2_1
XANTENNA_outbuf_1_A VSS VDD clkgen.clk_dig_out VDD VSS sky130_fd_sc_hd__diode_2
Xedgedetect.dly_315ns_1.genblk1\[5\].bypass_enable VDD VSS edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.bypass_in
+ edgedetect.dly_315ns_1.enable_dlycontrol_w edgedetect.dly_315ns_1.bypass_enable_w\[5\]
+ VDD VSS sky130_fd_sc_hd__and2_1
Xclkgen.delay_155ns_3.genblk1\[4\].dly_binary.out_mux VSS VDD clkgen.clk_comp_out
+ clkgen.delay_155ns_3.genblk1\[3\].dly_binary.out clkgen.delay_155ns_3.genblk1\[4\].dly_binary.bypass_in
+ clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[16\] VDD VSS sky130_fd_sc_hd__mux2_1
XFILLER_6_187 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XFILLER_18_272 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
XFILLER_9_91 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
Xclkgen.delay_155ns_1.genblk1\[2\].dly_binary.genblk1\[2\].delay_unit VDD VSS clkgen.delay_155ns_1.genblk1\[2\].dly_binary.signal_w\[2\]
+ clkgen.delay_155ns_1.genblk1\[2\].dly_binary.signal_w\[3\] clkgen.delay_155ns_1.genblk1\[2\].dly_binary.genblk1\[2\].delay_unit/mid
+ VDD VSS sky130_mm_sc_hd_dlyPoly5ns
XFILLER_17_337 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
XFILLER_4_274 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XFILLER_9_3 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
XPHY_35 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XPHY_24 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XPHY_13 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XFILLER_17_156 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
Xoutbuf_4 VSS VDD sample_n_1 sample_n_out VDD VSS sky130_fd_sc_hd__bufbuf_8
Xclkgen.delay_155ns_3.enablebuffer VDD VSS enable_dlycontrol_in clkgen.delay_155ns_3.enable_dlycontrol_w
+ VDD VSS sky130_fd_sc_hd__buf_4
XANTENNA_clkgen.delay_155ns_2.genblk1\[3\].dly_binary.out_mux_S VSS VDD clkgen.delay_155ns_2.genblk1\[3\].dly_binary.bypass_in
+ VDD VSS sky130_fd_sc_hd__diode_2
Xclkgen.delay_155ns_2.genblk1\[2\].control_invert VDD VSS clkgen.delay_155ns_2.bypass_enable_w\[2\]
+ dlycontrol2_in[2] VDD VSS sky130_fd_sc_hd__inv_2
Xedgedetect.dly_315ns_1.genblk1\[1\].dly_binary.genblk1\[1\].delay_unit VDD VSS edgedetect.dly_315ns_1.genblk1\[1\].dly_binary.signal_w\[1\]
+ edgedetect.dly_315ns_1.genblk1\[1\].dly_binary.signal_w\[2\] edgedetect.dly_315ns_1.genblk1\[1\].dly_binary.genblk1\[1\].delay_unit/mid
+ VDD VSS sky130_mm_sc_hd_dlyPoly5ns
XFILLER_18_284 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XANTENNA_clkgen.delay_155ns_2.genblk1\[4\].dly_binary.out_mux_A0 VSS VDD clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[16\]
+ VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_15_298 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XFILLER_0_94 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XFILLER_12_257 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XFILLER_8_206 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XANTENNA_clkgen.delay_155ns_2.genblk1\[3\].dly_binary.and_bypass_switch_A_N VSS VDD
+ clkgen.delay_155ns_2.genblk1\[3\].dly_binary.bypass_in VDD VSS sky130_fd_sc_hd__diode_2
Xclkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[13\].delay_unit VDD VSS clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[13\]
+ clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[14\] clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[13\].delay_unit/mid
+ VDD VSS sky130_mm_sc_hd_dlyPoly5ns
XANTENNA_edgedetect.dly_315ns_1.genblk1\[1\].control_invert_A VSS VDD dlycontrol4_in[1]
+ VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_4_242 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XPHY_25 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XPHY_36 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XPHY_14 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XANTENNA_delay_sample_n12_in VSS VDD sample_n_in VDD VSS sky130_fd_sc_hd__diode_2
Xedgedetect.dly_315ns_1.genblk1\[0\].bypass_enable VDD VSS edgedetect.dly_315ns_1.genblk1\[0\].dly_binary.bypass_in
+ edgedetect.dly_315ns_1.enable_dlycontrol_w edgedetect.dly_315ns_1.bypass_enable_w\[0\]
+ VDD VSS sky130_fd_sc_hd__and2_1
Xedgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[2\].delay_unit VDD VSS edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[2\]
+ edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[3\] edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[2\].delay_unit/mid
+ VDD VSS sky130_mm_sc_hd_dlyPoly5ns
XANTENNA_edgedetect.dly_315ns_1.genblk1\[0\].dly_binary.and_bypass_switch_B VSS VDD
+ edgedetect.dly_315ns_1.genblk1\[0\].dly_binary.in VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_3_94 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XFILLER_3_307 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XFILLER_10_174 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XFILLER_6_156 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
Xclkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[0\].delay_unit VDD VSS clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[0\]
+ clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[1\] clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[0\].delay_unit/mid
+ VDD VSS sky130_mm_sc_hd_dlyPoly5ns
Xclkgen.delay_155ns_1.genblk1\[1\].bypass_enable VDD VSS clkgen.delay_155ns_1.genblk1\[1\].dly_binary.bypass_in
+ clkgen.delay_155ns_1.enable_dlycontrol_w clkgen.delay_155ns_1.bypass_enable_w\[1\]
+ VDD VSS sky130_fd_sc_hd__and2_1
XANTENNA_clkgen.delay_155ns_2.genblk1\[1\].dly_binary.out_mux_S VSS VDD clkgen.delay_155ns_2.genblk1\[1\].dly_binary.bypass_in
+ VDD VSS sky130_fd_sc_hd__diode_2
Xclkgen.delay_155ns_2.genblk1\[2\].bypass_enable VDD VSS clkgen.delay_155ns_2.genblk1\[2\].dly_binary.bypass_in
+ clkgen.delay_155ns_2.enable_dlycontrol_w clkgen.delay_155ns_2.bypass_enable_w\[2\]
+ VDD VSS sky130_fd_sc_hd__and2_1
Xclkgen.delay_155ns_3.genblk1\[3\].bypass_enable VDD VSS clkgen.delay_155ns_3.genblk1\[3\].dly_binary.bypass_in
+ clkgen.delay_155ns_3.enable_dlycontrol_w clkgen.delay_155ns_3.bypass_enable_w\[3\]
+ VDD VSS sky130_fd_sc_hd__and2_1
XFILLER_17_3 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XFILLER_12_214 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
Xedgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[7\].delay_unit VDD VSS edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[7\]
+ edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[8\] edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[7\].delay_unit/mid
+ VDD VSS sky130_mm_sc_hd_dlyPoly5ns
Xedgedetect.dly_315ns_1.genblk1\[3\].control_invert VDD VSS edgedetect.dly_315ns_1.bypass_enable_w\[3\]
+ dlycontrol4_in[3] VDD VSS sky130_fd_sc_hd__inv_2
XPHY_37 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XPHY_26 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XPHY_15 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XFILLER_17_125 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
Xclkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[5\].delay_unit VDD VSS clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[5\]
+ clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[6\] clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[5\].delay_unit/mid
+ VDD VSS sky130_mm_sc_hd_dlyPoly5ns
Xclkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[11\].delay_unit VDD VSS clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[11\]
+ clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[12\] clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[11\].delay_unit/mid
+ VDD VSS sky130_mm_sc_hd_dlyPoly5ns
XFILLER_10_323 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_13_161 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XFILLER_10_164 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XFILLER_15_256 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XANTENNA_delay_sample_p11_in VSS VDD sample_p_in VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA_clkgen.delay_155ns_1.genblk1\[3\].control_invert_A VSS VDD dlycontrol1_in[3]
+ VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_0_63 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XFILLER_12_226 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
XFILLER_11_270 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XANTENNA_clkgen.delay_155ns_2.genblk1\[0\].dly_binary.out_mux_A1 VSS VDD clkgen.clk_dig_out
+ VDD VSS sky130_fd_sc_hd__diode_2
Xedgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[2\].delay_unit VDD VSS edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[2\]
+ edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[3\] edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[2\].delay_unit/mid
+ VDD VSS sky130_mm_sc_hd_dlyPoly5ns
XFILLER_4_211 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
Xclkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[4\].delay_unit VDD VSS clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[4\]
+ clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[5\] clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[4\].delay_unit/mid
+ VDD VSS sky130_mm_sc_hd_dlyPoly5ns
XPHY_27 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XPHY_38 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XANTENNA_clkgen.delay_155ns_2.genblk1\[2\].control_invert_A VSS VDD dlycontrol2_in[2]
+ VDD VSS sky130_fd_sc_hd__diode_2
XPHY_16 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XFILLER_9_303 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
Xclkgen.delay_155ns_3.genblk1\[3\].control_invert VDD VSS clkgen.delay_155ns_3.bypass_enable_w\[3\]
+ dlycontrol3_in[3] VDD VSS sky130_fd_sc_hd__inv_2
Xclkgen.delay_155ns_3.genblk1\[3\].dly_binary.genblk1\[0\].delay_unit VDD VSS clkgen.delay_155ns_3.genblk1\[3\].dly_binary.signal_w\[0\]
+ clkgen.delay_155ns_3.genblk1\[3\].dly_binary.signal_w\[1\] clkgen.delay_155ns_3.genblk1\[3\].dly_binary.genblk1\[0\].delay_unit/mid
+ VDD VSS sky130_mm_sc_hd_dlyPoly5ns
XFILLER_1_225 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XFILLER_0_280 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_10_335 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
XANTENNA_clkgen.delay_155ns_3.enablebuffer_A VSS VDD enable_dlycontrol_in VDD VSS
+ sky130_fd_sc_hd__diode_2
XFILLER_7_3 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XFILLER_6_306 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XFILLER_13_195 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XFILLER_3_63 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
XFILLER_3_30 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
XANTENNA_clkgen.delay_155ns_3.genblk1\[1\].control_invert_A VSS VDD dlycontrol3_in[1]
+ VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_12_94 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
Xedgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[7\].delay_unit VDD VSS edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[7\]
+ edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[8\] edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[7\].delay_unit/mid
+ VDD VSS sky130_mm_sc_hd_dlyPoly5ns
Xclkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[9\].delay_unit VDD VSS clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[9\]
+ clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[10\] clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[9\].delay_unit/mid
+ VDD VSS sky130_mm_sc_hd_dlyPoly5ns
Xclkgen.delay_155ns_3.genblk1\[3\].dly_binary.genblk1\[5\].delay_unit VDD VSS clkgen.delay_155ns_3.genblk1\[3\].dly_binary.signal_w\[5\]
+ clkgen.delay_155ns_3.genblk1\[3\].dly_binary.signal_w\[6\] clkgen.delay_155ns_3.genblk1\[3\].dly_binary.genblk1\[5\].delay_unit/mid
+ VDD VSS sky130_mm_sc_hd_dlyPoly5ns
Xedgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[10\].delay_unit VDD VSS edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[10\]
+ edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[11\] edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[10\].delay_unit/mid
+ VDD VSS sky130_mm_sc_hd_dlyPoly5ns
XFILLER_11_282 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XFILLER_7_275 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[3\].delay_unit VDD VSS clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[3\]
+ clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[4\] clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[3\].delay_unit/mid
+ VDD VSS sky130_mm_sc_hd_dlyPoly5ns
XFILLER_4_256 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XFILLER_4_201 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XPHY_28 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XFILLER_6_85 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XPHY_17 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XPHY_39 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XFILLER_13_300 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XFILLER_13_311 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
XFILLER_1_237 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XFILLER_1_259 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_9_337 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
Xedgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[14\].delay_unit VDD VSS edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[14\]
+ edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[15\] edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[14\].delay_unit/mid
+ VDD VSS sky130_mm_sc_hd_dlyPoly5ns
XFILLER_0_292 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
Xclkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[14\].delay_unit VDD VSS clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[14\]
+ clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[15\] clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[14\].delay_unit/mid
+ VDD VSS sky130_mm_sc_hd_dlyPoly5ns
XFILLER_11_19 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XFILLER_13_174 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
Xedgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[15\].delay_unit VDD VSS edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[15\]
+ edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[16\] edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[15\].delay_unit/mid
+ VDD VSS sky130_mm_sc_hd_dlyPoly5ns
XFILLER_18_244 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
Xedgedetect.dly_315ns_1.genblk1\[3\].dly_binary.genblk1\[2\].delay_unit VDD VSS edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.signal_w\[2\]
+ edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.signal_w\[3\] edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.genblk1\[2\].delay_unit/mid
+ VDD VSS sky130_mm_sc_hd_dlyPoly5ns
Xclkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[8\].delay_unit VDD VSS clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[8\]
+ clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[9\] clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[8\].delay_unit/mid
+ VDD VSS sky130_mm_sc_hd_dlyPoly5ns
XANTENNA_edgedetect.dly_315ns_1.genblk1\[0\].dly_binary.and_bypass_switch_A_N VSS
+ VDD edgedetect.dly_315ns_1.genblk1\[0\].dly_binary.bypass_in VDD VSS sky130_fd_sc_hd__diode_2
Xclkgen.delay_155ns_2.genblk1\[3\].dly_binary.genblk1\[4\].delay_unit VDD VSS clkgen.delay_155ns_2.genblk1\[3\].dly_binary.signal_w\[4\]
+ clkgen.delay_155ns_2.genblk1\[3\].dly_binary.signal_w\[5\] clkgen.delay_155ns_2.genblk1\[3\].dly_binary.genblk1\[4\].delay_unit/mid
+ VDD VSS sky130_mm_sc_hd_dlyPoly5ns
XFILLER_0_32 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XFILLER_9_63 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_3.genblk1\[2\].dly_binary.genblk1\[0\].delay_unit VDD VSS clkgen.delay_155ns_3.genblk1\[2\].dly_binary.signal_w\[0\]
+ clkgen.delay_155ns_3.genblk1\[2\].dly_binary.signal_w\[1\] clkgen.delay_155ns_3.genblk1\[2\].dly_binary.genblk1\[0\].delay_unit/mid
+ VDD VSS sky130_mm_sc_hd_dlyPoly5ns
Xedgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[19\].delay_unit VDD VSS edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[19\]
+ edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[20\] edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[19\].delay_unit/mid
+ VDD VSS sky130_mm_sc_hd_dlyPoly5ns
XFILLER_11_294 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XFILLER_18_94 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
Xedgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[21\].delay_unit VDD VSS edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[21\]
+ edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[22\] edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[21\].delay_unit/mid
+ VDD VSS sky130_mm_sc_hd_dlyPoly5ns
XANTENNA_edgedetect.dly_315ns_1.genblk1\[0\].dly_binary.out_mux_A1 VSS VDD edgedetect.dly_315ns_1.genblk1\[0\].dly_binary.in
+ VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_4_268 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XFILLER_4_235 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XPHY_18 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XPHY_29 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
Xedgedetect.dly_315ns_1.genblk1\[3\].dly_binary.genblk1\[7\].delay_unit VDD VSS edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.signal_w\[7\]
+ edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.signal_w\[8\] edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.genblk1\[7\].delay_unit/mid
+ VDD VSS sky130_mm_sc_hd_dlyPoly5ns
Xclkgen.delay_155ns_1.genblk1\[4\].control_invert VDD VSS clkgen.delay_155ns_1.bypass_enable_w\[4\]
+ dlycontrol1_in[4] VDD VSS sky130_fd_sc_hd__inv_2
XFILLER_12_63 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
Xedgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[26\].delay_unit VDD VSS edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[26\]
+ edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[27\] edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[26\].delay_unit/mid
+ VDD VSS sky130_mm_sc_hd_dlyPoly5ns
Xclkgen.delay_155ns_1.genblk1\[3\].dly_binary.genblk1\[3\].delay_unit VDD VSS clkgen.delay_155ns_1.genblk1\[3\].dly_binary.signal_w\[3\]
+ clkgen.delay_155ns_1.genblk1\[3\].dly_binary.signal_w\[4\] clkgen.delay_155ns_1.genblk1\[3\].dly_binary.genblk1\[3\].delay_unit/mid
+ VDD VSS sky130_mm_sc_hd_dlyPoly5ns
XFILLER_2_174 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XFILLER_12_207 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XANTENNA_edgedetect.dly_315ns_1.genblk1\[0\].control_invert_A VSS VDD dlycontrol4_in[0]
+ VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_6_43 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XPHY_19 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
Xedgedetect.dly_315ns_1.genblk1\[2\].dly_binary.genblk1\[2\].delay_unit VDD VSS edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.signal_w\[2\]
+ edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.signal_w\[3\] edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.genblk1\[2\].delay_unit/mid
+ VDD VSS sky130_mm_sc_hd_dlyPoly5ns
XFILLER_15_74 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_3.genblk1\[1\].dly_binary.genblk1\[0\].delay_unit VDD VSS clkgen.delay_155ns_3.genblk1\[1\].dly_binary.signal_w\[0\]
+ clkgen.delay_155ns_3.genblk1\[1\].dly_binary.signal_w\[1\] clkgen.delay_155ns_3.genblk1\[1\].dly_binary.genblk1\[0\].delay_unit/mid
+ VDD VSS sky130_mm_sc_hd_dlyPoly5ns
XFILLER_18_213 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XFILLER_5_3 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XFILLER_15_216 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
XFILLER_2_164 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XFILLER_9_32 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XFILLER_18_63 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XFILLER_11_241 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
XFILLER_11_263 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XFILLER_4_226 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XFILLER_19_182 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_1.genblk1\[2\].dly_binary.genblk1\[3\].delay_unit VDD VSS clkgen.delay_155ns_1.genblk1\[2\].dly_binary.signal_w\[3\]
+ clkgen.delay_155ns_1.genblk1\[2\].dly_binary.signal_w\[4\] clkgen.delay_155ns_1.genblk1\[2\].dly_binary.genblk1\[3\].delay_unit/mid
+ VDD VSS sky130_mm_sc_hd_dlyPoly5ns
XFILLER_1_218 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
.ends

.subckt sky130_fd_sc_hd__dfstp_2 VPWR VGND Q SET_B D CLK VPB VNB
X0 VGND a_652_21# a_586_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0882 pd=0.84 as=0.0671 ps=0.75 w=0.42 l=0.15
X1 a_956_413# a_476_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0567 ps=0.69 w=0.42 l=0.15
X2 a_1136_413# a_193_47# a_1028_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0819 ps=0.81 w=0.42 l=0.15
X3 VPWR a_476_47# a_652_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X4 a_586_47# a_193_47# a_476_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.072 ps=0.76 w=0.36 l=0.15
X5 a_1228_47# a_27_47# a_1028_413# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0735 ps=0.77 w=0.42 l=0.15
X6 VPWR CLK a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X7 a_476_47# a_27_47# a_381_47# VNB sky130_fd_pr__nfet_01v8 ad=0.072 pd=0.76 as=0.0935 ps=0.965 w=0.36 l=0.15
X8 a_1056_47# a_476_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X9 a_381_47# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.125 pd=1.17 as=0.218 ps=2.2 w=0.84 l=0.15
X10 a_652_21# SET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0798 ps=0.8 w=0.42 l=0.15
X11 VPWR a_1602_47# Q VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X12 a_562_413# a_27_47# a_476_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0567 ps=0.69 w=0.42 l=0.15
X13 VGND a_1028_413# a_1602_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X14 VGND a_1602_47# Q VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X15 Q a_1602_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X16 a_1028_413# a_193_47# a_1056_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0735 pd=0.77 as=0.0441 ps=0.63 w=0.42 l=0.15
X17 a_476_47# a_193_47# a_381_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.125 ps=1.17 w=0.42 l=0.15
X18 a_193_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X19 VPWR a_1028_413# a_1602_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X20 VPWR a_652_21# a_562_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.0945 ps=0.87 w=0.42 l=0.15
X21 Q a_1602_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X22 a_1028_413# a_27_47# a_956_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0441 ps=0.63 w=0.42 l=0.15
X23 VPWR a_1178_261# a_1136_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X24 a_193_47# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X25 a_1178_261# a_1028_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.223 pd=2.21 as=0.121 ps=1.16 w=0.84 l=0.15
X26 a_796_47# SET_B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0882 ps=0.84 w=0.42 l=0.15
X27 a_1300_47# a_1178_261# a_1228_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X28 a_381_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0935 pd=0.965 as=0.166 ps=1.8 w=0.64 l=0.15
X29 a_1178_261# a_1028_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.6 as=0.114 ps=1.01 w=0.54 l=0.15
X30 a_652_21# a_476_47# a_796_47# VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X31 VPWR SET_B a_1028_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.121 pd=1.16 as=0.109 ps=1.36 w=0.42 l=0.15
X32 VGND CLK a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X33 VGND SET_B a_1300_47# VNB sky130_fd_pr__nfet_01v8 ad=0.114 pd=1.01 as=0.0441 ps=0.63 w=0.42 l=0.15
.ends

.subckt adc_top VDD VSS inp_analog inn_analog rst_n clk_vcm start_conversion_in 
+ conversion_finished_out conversion_finished_osr_out
+ config_1_in[15] config_1_in[14] config_1_in[13] config_1_in[12] config_1_in[11] config_1_in[10]
+ config_1_in[9] config_1_in[8] config_1_in[7] config_1_in[6] config_1_in[5] config_1_in[4]
+ config_1_in[3] config_1_in[2] config_1_in[1] config_1_in[0]
+ config_2_in[15] config_2_in[14] config_2_in[13] config_2_in[12] config_2_in[11] config_2_in[10]
+ config_2_in[9] config_2_in[8] config_2_in[7] config_2_in[6] config_2_in[5] config_2_in[4]
+ config_2_in[3] config_2_in[2] config_2_in[1] config_2_in[0]
+ result_out[15] result_out[14] result_out[13] result_out[12] result_out[11] result_out[10]
+ result_out[9] result_out[8] result_out[7] result_out[6] result_out[5] result_out[4]
+ result_out[3] result_out[2] result_out[1] result_out[0]
X_3155_ VSS VDD net59 _0045_ net71 net40 VDD VSS sky130_fd_sc_hd__dfrtp_1
X_3086_ VDD VSS _1342_ _0971_ _0799_ VDD VSS sky130_fd_sc_hd__xor2_1
X_2106_ VDD VSS _1125_ _0068_ core.pdc.col_out\[27\] _0070_ _1102_ _0160_ VDD VSS
+ sky130_fd_sc_hd__a221o_1
X_2037_ VDD VSS _0120_ _0098_ VDD VSS sky130_fd_sc_hd__inv_2
X_2939_ VSS VDD _0830_ _0831_ VDD VSS sky130_fd_sc_hd__clkbuf_2
XANTENNA__1534__A VSS VDD net15 VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__3132__CLK VSS VDD clknet_2_0__leaf_clk_dig_dummy VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_92_309 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
XFILLER_93_25 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XFILLER_26_41 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XFILLER_26_85 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
XANTENNA__2084__B VSS VDD _0113_ VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_3_45 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XFILLER_83_309 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XANTENNA__1987__A2 VSS VDD _1053_ VDD VSS sky130_fd_sc_hd__diode_2
X_2724_ VSS VDD _0620_ _0622_ _0621_ VDD VSS sky130_fd_sc_hd__nand2_1
X_2655_ VSS VDD _0288_ _0560_ _0530_ VDD VSS sky130_fd_sc_hd__nand2_1
X_1606_ VDD VSS _1154_ _1153_ VDD VSS sky130_fd_sc_hd__inv_2
X_2586_ VSS VDD _1300_ _0501_ _0502_ VDD VSS sky130_fd_sc_hd__nor2_1
X_1537_ VSS VDD _1075_ _1084_ _1070_ _1064_ core.ndc.col_out_n\[1\] _1094_ VDD VSS
+ sky130_fd_sc_hd__o221a_2
X_1468_ VSS VDD _1028_ _1030_ _1029_ VDD VSS sky130_fd_sc_hd__nand2_1
X_3138_ VSS VDD clknet_2_0__leaf_clk_dig_dummy _0028_ net85 core.cnb.result_out\[6\]
+ VDD VSS sky130_fd_sc_hd__dfrtp_1
X_3069_ VDD VSS _0955_ _0954_ VDD VSS sky130_fd_sc_hd__inv_2
XFILLER_88_25 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XFILLER_77_103 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XANTENNA__2095__A VSS VDD _0065_ VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1439__A VSS VDD _1002_ VDD VSS sky130_fd_sc_hd__diode_2
Xgenblk2\[3\].buf_p_rown VSS VDD pmatrix_row_core_n_buffered\[3\] core.pdc.row_out_n\[3\]
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
XANTENNA__3178__CLK VSS VDD net58 VDD VSS sky130_fd_sc_hd__diode_2
X_2440_ VSS VDD _1332_ core.pdc.rowon_bottotop_n\[5\] _1342_ VDD VSS sky130_fd_sc_hd__nor2_2
X_2371_ VSS VDD _0384_ core.osr.result_r\[18\] _0387_ VDD VSS sky130_fd_sc_hd__nand2b_1
XFILLER_56_309 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_83_128 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XANTENNA__1902__A VSS VDD core.pdc.rowoff_out_n\[5\] VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__2082__A1 VSS VDD _1284_ VDD VSS sky130_fd_sc_hd__diode_2
X_2707_ VSS VDD _0376_ _0605_ _0606_ _0517_ VDD VSS sky130_fd_sc_hd__o21ai_1
X_2638_ VSS VDD core.osr.next_result_w\[7\] _0545_ _0535_ VDD VSS sky130_fd_sc_hd__nand2_1
X_2569_ VSS VDD _1395_ _0483_ _0490_ VDD VSS sky130_fd_sc_hd__nor2_1
XFILLER_59_136 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XANTENNA__2908__A VSS VDD _0799_ VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_87_489 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XFILLER_130_11 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
XFILLER_23_31 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XANTENNA__2362__B VSS VDD _0241_ VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_139_53 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XFILLER_139_97 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_136_141 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_99_35 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XFILLER_99_57 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_48_72 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_0_24 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XFILLER_0_57 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_9_22 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
X_1940_ VSS VDD _1396_ _1395_ _1394_ _1079_ _1085_ VDD VSS sky130_fd_sc_hd__a211o_2
X_1871_ VSS VDD core.ndc.rowoff_out_n\[8\] _1321_ _1352_ VDD VSS sky130_fd_sc_hd__nor2_1
X_2423_ VSS VDD _1356_ _1352_ core.ndc.row_out_n\[4\] VDD VSS sky130_fd_sc_hd__nor2_1
X_2354_ VSS VDD _0371_ _0373_ _0372_ VDD VSS sky130_fd_sc_hd__nand2_1
X_2285_ VSS VDD _0309_ _0311_ _0307_ VDD VSS sky130_fd_sc_hd__nand2_1
XANTENNA__2447__B VSS VDD core.pdc.rowon_out_n\[15\] VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_52_301 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
Xgenblk2\[0\].buf_n_rown VSS VDD nmatrix_row_core_n_buffered\[0\] core.ndc.row_out_n\[0\]
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
XFILLER_100_25 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XANTENNA__2182__B VSS VDD _0220_ VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1802__A1 VSS VDD _1126_ VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1802__B2 VSS VDD _1296_ VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_60_29 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_118_141 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_118_130 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XFILLER_109_23 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
XANTENNA__1807__A VSS VDD core.cnb.data_register_r\[8\] VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_47_128 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XFILLER_55_161 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XFILLER_55_183 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_34_85 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XANTENNA__2267__B VSS VDD core.cnb.result_out\[6\] VDD VSS sky130_fd_sc_hd__diode_2
X_2070_ VDD VSS core.pdc.col_out_n\[18\] core.pdc.col_out\[18\] VDD VSS sky130_fd_sc_hd__clkinv_2
XANTENNA__1598__S VSS VDD _1077_ VDD VSS sky130_fd_sc_hd__diode_2
X_2972_ VSS VDD _0054_ _0757_ _0863_ _0861_ _1055_ _0688_ VDD VSS sky130_fd_sc_hd__a32o_1
X_1923_ VSS VDD _1362_ core.ndc.rowoff_out_n\[5\] _1384_ VDD VSS sky130_fd_sc_hd__nor2_1
X_1854_ VSS VDD _1340_ _1026_ _1341_ _1300_ VDD VSS sky130_fd_sc_hd__o21ai_1
XANTENNA__1627__A VSS VDD _1032_ VDD VSS sky130_fd_sc_hd__diode_2
X_1785_ VSS VDD _1124_ _1291_ _1275_ VDD VSS sky130_fd_sc_hd__nand2_1
X_2406_ VDD VSS _0414_ core.osr.is_last_sample _0412_ _0415_ VDD VSS sky130_fd_sc_hd__or3_1
X_2337_ VDD VSS _0358_ _0357_ VDD VSS sky130_fd_sc_hd__inv_2
X_2268_ VSS VDD _0296_ _0294_ _0255_ _0293_ _0295_ VDD VSS sky130_fd_sc_hd__a31o_1
Xgenblk2\[4\].buf_p_rowonn VSS VDD pmatrix_rowon_core_n_buffered\[4\] core.pdc.rowon_out_n\[4\]
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
X_2199_ VSS VDD core.cnb.next_average_sum_w\[3\] _0234_ VDD VSS sky130_fd_sc_hd__clkbuf_1
XANTENNA_nmat_col_n[8] VSS VDD nmatrix_col_core_n_buffered\[8\] VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_52_197 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_112_5 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XFILLER_20_76 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XFILLER_136_65 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_96_47 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XANTENNA__1711__A0 VSS VDD _1242_ VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA_input18_A VSS VDD config_2_in[0] VDD VSS sky130_fd_sc_hd__diode_2
X_1570_ VSS VDD _1058_ _1037_ _1122_ VDD VSS sky130_fd_sc_hd__nor2_1
X_3171_ VSS VDD net61 core.osr.next_result_w\[11\] net73 core.osr.result_r\[11\] VDD
+ VSS sky130_fd_sc_hd__dfrtp_1
X_2122_ VSS VDD _1396_ _0171_ _1188_ VDD VSS sky130_fd_sc_hd__nand2_1
XFILLER_19_150 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
XFILLER_47_481 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
X_2053_ VDD VSS _0131_ _0132_ VDD VSS sky130_fd_sc_hd__clkinv_2
XFILLER_34_153 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
X_2955_ VDD VSS _0847_ _0471_ VDD VSS sky130_fd_sc_hd__inv_2
X_1906_ VDD VSS _1376_ _1375_ VDD VSS sky130_fd_sc_hd__inv_2
X_2886_ VDD VSS _0780_ _0777_ _0779_ VDD VSS sky130_fd_sc_hd__or2_1
X_1837_ VSS VDD core.cnb.data_register_r\[10\] _1326_ VDD VSS sky130_fd_sc_hd__clkbuf_2
X_1768_ VSS VDD _1176_ _1280_ _1279_ VDD VSS sky130_fd_sc_hd__nand2_1
X_1699_ VDD VSS _1232_ _1233_ VDD VSS sky130_fd_sc_hd__clkinv_2
XFILLER_85_510 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_122_23 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XANTENNA__2249__A1 VSS VDD core.cnb.result_out\[4\] VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1820__A VSS VDD _1312_ VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_40_101 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_25_153 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XANTENNA__3160__RESET_B VSS VDD net81 VDD VSS sky130_fd_sc_hd__diode_2
Xgenblk2\[8\].buf_p_rown VSS VDD pmatrix_row_core_n_buffered\[8\] core.pdc.row_out_n\[8\]
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xoutput42 VDD VSS result_out[13] net42 VDD VSS sky130_fd_sc_hd__buf_2
Xoutput53 VDD VSS result_out[9] net53 VDD VSS sky130_fd_sc_hd__buf_2
XANTENNA__2098__A VSS VDD _0065_ VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1999__B1 VSS VDD _1259_ VDD VSS sky130_fd_sc_hd__diode_2
X_2740_ VSS VDD _0206_ _0636_ _0635_ VDD VSS sky130_fd_sc_hd__nand2_1
XANTENNA__2561__A VSS VDD _0482_ VDD VSS sky130_fd_sc_hd__diode_2
X_2671_ VSS VDD _0347_ _1002_ _0574_ _0348_ VDD VSS sky130_fd_sc_hd__nand3_1
XFILLER_75_5 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
X_1622_ VDD VSS _1167_ _1168_ VDD VSS sky130_fd_sc_hd__clkinv_2
X_1553_ VDD VSS core.ndc.col_out_n\[2\] core.ndc.col_out\[2\] VDD VSS sky130_fd_sc_hd__inv_2
XANTENNA__2500__S VSS VDD _0220_ VDD VSS sky130_fd_sc_hd__diode_2
X_1484_ VDD VSS _1044_ core.cnb.data_register_r\[5\] VDD VSS sky130_fd_sc_hd__buf_2
XANTENNA__1624__B VSS VDD _1045_ VDD VSS sky130_fd_sc_hd__diode_2
X_3154_ VSS VDD net59 _0044_ net71 net39 VDD VSS sky130_fd_sc_hd__dfrtp_1
XANTENNA__1640__A VSS VDD _1039_ VDD VSS sky130_fd_sc_hd__diode_2
X_3085_ VSS VDD _0966_ _0970_ _0969_ VDD VSS sky130_fd_sc_hd__nand2_1
X_2105_ VDD VSS _0160_ _0103_ _1092_ VDD VSS sky130_fd_sc_hd__and2_1
X_2036_ VSS VDD _0118_ _0119_ _1235_ VDD VSS sky130_fd_sc_hd__nand2_1
X_2938_ VSS VDD _0820_ _0829_ _0830_ _0753_ VDD VSS sky130_fd_sc_hd__nand3_1
XANTENNA__2471__A VSS VDD core.pdc.row_out_n\[2\] VDD VSS sky130_fd_sc_hd__diode_2
X_2869_ VSS VDD _0649_ _0701_ _0763_ _0762_ VDD VSS sky130_fd_sc_hd__nand3_1
Xgenblk1\[3\].buf_p_coln VSS VDD pmatrix_col_core_n_buffered\[3\] core.pdc.col_out_n\[3\]
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
XANTENNA__1914__B1 VSS VDD core.ndc.rowon_bottotop_n\[5\] VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_9_105 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
XFILLER_42_41 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XANTENNA__2381__A VSS VDD _0394_ VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1709__B VSS VDD _1213_ VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_47_9 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XFILLER_67_82 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_83_81 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
Xgenblk2\[5\].buf_n_rown VSS VDD nmatrix_row_core_n_buffered\[5\] core.ndc.row_bottotop_n\[5\]
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
X_2723_ VDD VSS _0530_ _0356_ _1018_ _0621_ VDD VSS sky130_fd_sc_hd__a21oi_1
X_2654_ VSS VDD _0557_ _0559_ _0558_ VDD VSS sky130_fd_sc_hd__nand2_1
X_1605_ VSS VDD _1105_ _1078_ _1153_ _1135_ VDD VSS sky130_fd_sc_hd__a21oi_2
X_2585_ VSS VDD _0488_ _0501_ _1067_ VDD VSS sky130_fd_sc_hd__nand2_1
XANTENNA__1635__A VSS VDD core.ndc.col_out_n\[7\] VDD VSS sky130_fd_sc_hd__diode_2
X_1536_ VSS VDD _1091_ _1094_ _1093_ VDD VSS sky130_fd_sc_hd__nand2_1
X_1467_ VSS VDD core.cnb.data_register_r\[11\] _1029_ core.cnb.data_register_r\[10\]
+ VDD VSS sky130_fd_sc_hd__nor2_2
X_3137_ VSS VDD clknet_2_0__leaf_clk_dig_dummy _0027_ net79 core.cnb.result_out\[5\]
+ VDD VSS sky130_fd_sc_hd__dfrtp_2
X_3068_ VDD VSS _1326_ _0954_ _0799_ VDD VSS sky130_fd_sc_hd__xor2_1
X_2019_ VSS VDD _0107_ _0108_ _1135_ VDD VSS sky130_fd_sc_hd__nand2_1
XFILLER_50_273 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
XFILLER_10_148 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XANTENNA__1545__A VSS VDD _1032_ VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_92_107 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XFILLER_92_129 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XANTENNA__2823__B VSS VDD core.cnb.data_register_r\[1\] VDD VSS sky130_fd_sc_hd__diode_2
Xgenblk1\[0\].buf_n_coln VDD VSS core.ndc.col_out_n\[0\] nmatrix_col_core_n_buffered\[0\]
+ VDD VSS sky130_fd_sc_hd__buf_6
X_2370_ VSS VDD core.osr.next_result_w\[17\] _0386_ VDD VSS sky130_fd_sc_hd__clkbuf_1
XFILLER_68_137 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XANTENNA__1902__B VSS VDD _1325_ VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__3122__CLK VSS VDD clknet_2_2__leaf_clk_dig_dummy VDD VSS sky130_fd_sc_hd__diode_2
X_2706_ VSS VDD _0381_ _0385_ _0605_ _0517_ VDD VSS sky130_fd_sc_hd__nand3_1
X_2637_ VSS VDD core.osr.next_result_w\[9\] _0544_ _0533_ VDD VSS sky130_fd_sc_hd__nand2_1
XFILLER_58_29 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
X_2568_ VDD VSS _0489_ _0488_ VDD VSS sky130_fd_sc_hd__dlymetal6s2s_1
X_2499_ VSS VDD _0004_ _0440_ VDD VSS sky130_fd_sc_hd__clkbuf_1
X_1519_ VDD VSS _1077_ _1041_ VDD VSS sky130_fd_sc_hd__buf_2
XFILLER_114_35 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XFILLER_114_79 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XFILLER_130_56 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_23_43 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XFILLER_99_14 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_136_153 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XFILLER_99_69 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XFILLER_93_405 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XANTENNA__1722__B VSS VDD _1102_ VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_93_449 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_0_69 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
X_1870_ VDD VSS core.ndc.rowoff_out_n\[8\] _1351_ VDD VSS sky130_fd_sc_hd__inv_2
XFILLER_80_93 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
X_2422_ VSS VDD _1350_ _1354_ core.ndc.row_out_n\[3\] VDD VSS sky130_fd_sc_hd__nor2_1
X_2353_ VSS VDD _0352_ _0372_ _0370_ VDD VSS sky130_fd_sc_hd__or2b_1
X_2284_ VDD VSS _0310_ _0307_ _0309_ VDD VSS sky130_fd_sc_hd__or2_1
XANTENNA__1632__B VSS VDD _1177_ VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_61_891 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
X_1999_ VSS VDD _1259_ _0090_ _0088_ _1224_ core.pdc.col_out_n\[7\] _0093_ VDD VSS
+ sky130_fd_sc_hd__o221a_1
XFILLER_118_153 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XFILLER_109_57 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XANTENNA__3185__RESET_B VSS VDD net87 VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__3168__CLK VSS VDD net66 VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_55_195 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XFILLER_34_97 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_34_75 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XFILLER_50_85 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_59_94 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_93_213 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XFILLER_46_151 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
X_2971_ VSS VDD _0862_ _0790_ _0863_ _0805_ VDD VSS sky130_fd_sc_hd__nand3_1
X_1922_ VSS VDD _1372_ _1369_ _1378_ core.pdc.rowon_out_n\[12\] VDD VSS sky130_fd_sc_hd__a21o_2
X_1853_ VSS VDD _1340_ _1339_ _1303_ VDD VSS sky130_fd_sc_hd__nand2_2
XANTENNA__1796__A1 VSS VDD _1091_ VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1796__B2 VSS VDD _1296_ VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1908__A VSS VDD _1377_ VDD VSS sky130_fd_sc_hd__diode_2
X_1784_ VDD VSS _1289_ _1290_ VDD VSS sky130_fd_sc_hd__clkinv_2
XFILLER_115_134 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
Xgenblk1\[8\].buf_p_coln VSS VDD pmatrix_col_core_n_buffered\[8\] core.pdc.col_out_n\[8\]
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
X_2405_ VDD VSS _0414_ _0413_ VDD VSS sky130_fd_sc_hd__inv_2
XANTENNA__2458__B VSS VDD core.ndc.rowon_out_n\[3\] VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_29_118 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
X_2336_ VSS VDD core.osr.result_r\[12\] _0357_ core.osr.result_r\[13\] VDD VSS sky130_fd_sc_hd__nand2_1
X_2267_ VDD VSS _0295_ _0251_ core.cnb.result_out\[6\] VDD VSS sky130_fd_sc_hd__and2_1
X_2198_ VSS VDD _0234_ _0233_ _0232_ _0209_ VDD VSS sky130_fd_sc_hd__and3_1
XANTENNA_nmat_col_n[7] VSS VDD nmatrix_col_core_n_buffered\[7\] VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_52_187 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XFILLER_136_77 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
XANTENNA__1553__A VSS VDD core.ndc.col_out\[2\] VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__2368__B VSS VDD _0255_ VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1711__A1 VSS VDD _1202_ VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_48_416 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XFILLER_45_74 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XFILLER_83_290 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XFILLER_45_85 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XANTENNA__1778__A1 VSS VDD _1284_ VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1728__A VSS VDD core.ndc.col_out_n\[16\] VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1463__A VSS VDD net14 VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_112_126 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
X_3170_ VSS VDD net61 core.osr.next_result_w\[10\] net73 core.osr.result_r\[10\] VDD
+ VSS sky130_fd_sc_hd__dfrtp_1
X_2121_ VSS VDD _1401_ _0170_ _1096_ VDD VSS sky130_fd_sc_hd__nand2_1
X_2052_ VSS VDD _1227_ _0094_ _0131_ VDD VSS sky130_fd_sc_hd__nor2_1
XANTENNA__1910__B VSS VDD _1342_ VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_47_493 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
X_2954_ VSS VDD _0845_ _0846_ _0475_ VDD VSS sky130_fd_sc_hd__nand2_1
X_1905_ VSS VDD _1038_ _1339_ _1375_ VDD VSS sky130_fd_sc_hd__nor2_1
XANTENNA__2741__B VSS VDD net54 VDD VSS sky130_fd_sc_hd__diode_2
X_2885_ VSS VDD _0778_ _0779_ _0718_ VDD VSS sky130_fd_sc_hd__nand2_1
X_1836_ VDD VSS _1325_ _1324_ VDD VSS sky130_fd_sc_hd__buf_2
X_1767_ VDD VSS _1279_ _1032_ VDD VSS sky130_fd_sc_hd__buf_2
X_1698_ VSS VDD _1227_ _1231_ _1232_ VDD VSS sky130_fd_sc_hd__nor2_1
XANTENNA__2497__A2 VSS VDD _0220_ VDD VSS sky130_fd_sc_hd__diode_2
X_2319_ VDD VSS _0342_ _0341_ VDD VSS sky130_fd_sc_hd__inv_2
XFILLER_66_29 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_85_522 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
XANTENNA__1820__B VSS VDD _1022_ VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_40_113 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
Xgenblk1\[5\].buf_n_coln VDD VSS core.ndc.col_out_n\[5\] nmatrix_col_core_n_buffered\[5\]
+ VDD VSS sky130_fd_sc_hd__buf_6
Xoutput43 VDD VSS result_out[14] net43 VDD VSS sky130_fd_sc_hd__buf_2
XANTENNA__2098__B VSS VDD _0115_ VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1696__A0 VSS VDD _1229_ VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA_input30_A VSS VDD config_2_in[6] VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1730__B VSS VDD _1213_ VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1999__A1 VSS VDD _1224_ VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_31_113 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
X_2670_ VDD VSS _1008_ _0363_ _0524_ _0573_ VDD VSS sky130_fd_sc_hd__a21oi_1
X_1621_ VSS VDD _1131_ _1166_ _1167_ VDD VSS sky130_fd_sc_hd__nor2_1
X_1552_ VDD VSS _1096_ core.ndc.col_out\[2\] _1091_ _1107_ _1100_ _1102_ VDD VSS sky130_fd_sc_hd__a221o_4
X_1483_ VSS VDD _1042_ _1043_ VDD VSS sky130_fd_sc_hd__clkbuf_2
X_3153_ VSS VDD net59 _0043_ net71 net53 VDD VSS sky130_fd_sc_hd__dfrtp_1
XFILLER_100_118 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XANTENNA__1921__A VSS VDD _1383_ VDD VSS sky130_fd_sc_hd__diode_2
X_2104_ VDD VSS core.pdc.col_out\[26\] core.pdc.col_out_n\[26\] VDD VSS sky130_fd_sc_hd__clkinv_2
X_3084_ VDD VSS _0918_ _0912_ _1022_ _0969_ VDD VSS sky130_fd_sc_hd__or3_1
XFILLER_47_290 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
X_2035_ VDD VSS _0118_ _0074_ VDD VSS sky130_fd_sc_hd__inv_2
XFILLER_22_146 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XFILLER_50_477 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
X_2937_ VSS VDD _0828_ _0809_ _0806_ _0829_ VDD VSS sky130_fd_sc_hd__nor3_1
XANTENNA__2471__B VSS VDD core.pdc.rowon_out_n\[2\] VDD VSS sky130_fd_sc_hd__diode_2
X_2868_ VSS VDD core.cnb.shift_register_r\[12\] _0698_ _0762_ VDD VSS sky130_fd_sc_hd__nor2_1
X_1819_ VSS VDD _1071_ _1312_ VDD VSS sky130_fd_sc_hd__clkbuf_2
X_2799_ VDD VSS _0694_ _0678_ core.cnb.shift_register_r\[15\] VDD VSS sky130_fd_sc_hd__and2_1
XFILLER_133_67 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XFILLER_85_374 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XFILLER_93_49 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
XFILLER_13_113 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_42_53 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XANTENNA__1725__B VSS VDD _1177_ VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1669__A0 VSS VDD _1208_ VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_95_116 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
XANTENNA__1741__A VSS VDD _1033_ VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_95_149 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XFILLER_67_94 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XANTENNA__1460__B VSS VDD core.cnb.data_register_r\[8\] VDD VSS sky130_fd_sc_hd__diode_2
Xgenblk2\[13\].buf_n_rowonn VSS VDD nmatrix_rowon_core_n_buffered\[13\] core.ndc.rowon_out_n\[13\]
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
X_2722_ VSS VDD _0618_ _0619_ _0620_ _0528_ VDD VSS sky130_fd_sc_hd__nand3_1
X_2653_ VSS VDD core.osr.next_result_w\[11\] _0558_ _0533_ VDD VSS sky130_fd_sc_hd__nand2_1
X_2584_ VSS VDD core.cnb.result_out\[7\] _0461_ _0500_ _0029_ VDD VSS sky130_fd_sc_hd__o21a_1
X_1604_ VDD VSS _1152_ _1092_ VDD VSS sky130_fd_sc_hd__buf_2
X_1535_ VDD VSS _1093_ _1092_ VDD VSS sky130_fd_sc_hd__buf_2
X_1466_ VSS VDD core.cnb.data_register_r\[9\] core.cnb.data_register_r\[8\] _1028_
+ VDD VSS sky130_fd_sc_hd__nor2_1
X_3136_ VSS VDD clknet_2_0__leaf_clk_dig_dummy _0026_ net78 core.cnb.result_out\[4\]
+ VDD VSS sky130_fd_sc_hd__dfrtp_2
XFILLER_55_525 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
X_3067_ VSS VDD _0952_ _0059_ _0953_ VDD VSS sky130_fd_sc_hd__nand2_1
X_2018_ VSS VDD _1390_ _0107_ _1122_ VDD VSS sky130_fd_sc_hd__nand2_1
XANTENNA__2482__A VSS VDD core.pdc.row_out_n\[15\] VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA_fanout80_A VSS VDD net81 VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__2657__A VSS VDD _0983_ VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1561__A VSS VDD _1114_ VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_37_53 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XANTENNA__1736__A VSS VDD _1124_ VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1471__A VSS VDD core.ndc.rowoff_out_n\[0\] VDD VSS sky130_fd_sc_hd__diode_2
X_2705_ VSS VDD _0602_ _0046_ _0604_ VDD VSS sky130_fd_sc_hd__nand2_1
X_2636_ VSS VDD _0038_ _0541_ _0540_ _0539_ _0543_ VDD VSS sky130_fd_sc_hd__a31o_1
XANTENNA__1593__A2 VSS VDD _1141_ VDD VSS sky130_fd_sc_hd__diode_2
X_2567_ VSS VDD _0487_ _0473_ _0488_ VDD VSS sky130_fd_sc_hd__nor2_1
X_2498_ VSS VDD _0440_ core.cnb.shift_register_r\[3\] _0203_ core.cnb.shift_register_r\[2\]
+ VDD VSS sky130_fd_sc_hd__mux2_1
X_1518_ VDD VSS _1076_ core.cnb.data_register_r\[3\] VDD VSS sky130_fd_sc_hd__buf_2
X_1449_ VDD VSS _1013_ core.osr.sample_count_r\[7\] VDD VSS sky130_fd_sc_hd__inv_2
Xvcm net1 vcm/phi2 vcm/phi1_n vcm/phi1 vcm/phi2_n vcm/vcm VDD vcm/mimtop1 vcm/mimtop2
+ vcm/mimbot1 VSS adc_vcm_generator
XFILLER_55_311 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XFILLER_55_333 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
X_3119_ VSS VDD clknet_2_0__leaf_clk_dig_dummy _0019_ net84 core.cnb.sampled_avg_control_r\[0\]
+ VDD VSS sky130_fd_sc_hd__dfrtp_4
XFILLER_82_141 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
XFILLER_130_68 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XFILLER_139_11 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_136_121 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_99_26 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XANTENNA__1556__A VSS VDD _1039_ VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_93_417 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XFILLER_104_91 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XFILLER_9_57 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_80_50 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
X_2421_ VSS VDD _1331_ _1329_ core.ndc.row_out_n\[2\] _1357_ VDD VSS sky130_fd_sc_hd__a21oi_2
XFILLER_89_81 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
X_2352_ VSS VDD _0309_ _0351_ _0371_ _0370_ VDD VSS sky130_fd_sc_hd__nand3_1
X_2283_ VSS VDD _0308_ _0300_ _0309_ _0294_ VDD VSS sky130_fd_sc_hd__o21ai_2
XFILLER_52_358 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
XFILLER_100_49 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
X_1998_ VSS VDD _0092_ _0093_ _1155_ VDD VSS sky130_fd_sc_hd__nand2_1
XFILLER_133_113 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_109_69 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
X_2619_ VSS VDD _1011_ _0528_ VDD VSS sky130_fd_sc_hd__clkbuf_2
XFILLER_87_200 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_125_57 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XFILLER_125_79 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_87_277 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XFILLER_83_461 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XANTENNA__2373__C VSS VDD _0240_ VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__2451__B1 VSS VDD _1328_ VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_51_380 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_126_1 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_50_97 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XFILLER_38_108 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XANTENNA__3112__CLK VSS VDD clknet_2_3__leaf_clk_dig_dummy VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_93_225 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XFILLER_46_163 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XFILLER_75_94 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
X_2970_ VSS VDD _0792_ _0862_ _0789_ VDD VSS sky130_fd_sc_hd__nand2_1
X_1921_ VSS VDD core.pdc.rowon_out_n\[11\] _1383_ VDD VSS sky130_fd_sc_hd__clkbuf_1
XFILLER_98_5 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_91_71 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
X_1852_ VDD VSS _1339_ _1338_ VDD VSS sky130_fd_sc_hd__inv_2
XANTENNA__1796__A2 VSS VDD _1279_ VDD VSS sky130_fd_sc_hd__diode_2
X_1783_ VSS VDD _1131_ _1194_ _1289_ VDD VSS sky130_fd_sc_hd__nor2_1
X_2404_ VSS VDD _0410_ _0413_ core.osr.sample_count_r\[5\] VDD VSS sky130_fd_sc_hd__nand2_1
X_2335_ VDD VSS _0356_ core.osr.next_result_w\[12\] VDD VSS sky130_fd_sc_hd__clkinv_2
X_2266_ VSS VDD _0292_ _0294_ _0291_ VDD VSS sky130_fd_sc_hd__nand2_1
X_2197_ VSS VDD _0227_ _0233_ core.cnb.average_sum_r\[3\] VDD VSS sky130_fd_sc_hd__nand2_1
XANTENNA_nmat_col_n[6] VSS VDD nmatrix_col_core_n_buffered\[6\] VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_52_144 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XANTENNA__1834__A VSS VDD _1323_ VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__3135__CLK VSS VDD clknet_2_0__leaf_clk_dig_dummy VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_29_43 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
XANTENNA__2665__A VSS VDD core.osr.next_result_w\[8\] VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_56_461 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_45_97 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_6_25 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XFILLER_61_96 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
X_2120_ VDD VSS core.pdc.col_out_n\[29\] core.pdc.col_out\[29\] VDD VSS sky130_fd_sc_hd__clkinv_2
XFILLER_86_93 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
X_2051_ VSS VDD _1396_ _0130_ _1152_ VDD VSS sky130_fd_sc_hd__nand2_1
XFILLER_47_461 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XFILLER_34_133 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
X_2953_ VSS VDD _0844_ _0845_ _0834_ VDD VSS sky130_fd_sc_hd__nand2_1
X_1904_ VDD VSS _1374_ _1026_ _1373_ VDD VSS sky130_fd_sc_hd__or2_1
XANTENNA__1638__B VSS VDD _1053_ VDD VSS sky130_fd_sc_hd__diode_2
X_2884_ VSS VDD _0718_ _0720_ _0778_ _0719_ VDD VSS sky130_fd_sc_hd__nand3_1
X_1835_ VSS VDD net14 _1324_ _1308_ VDD VSS sky130_fd_sc_hd__nand2_1
X_1766_ VDD VSS core.ndc.col_out\[23\] core.ndc.col_out_n\[23\] VDD VSS sky130_fd_sc_hd__inv_2
X_1697_ VDD VSS _1231_ _1230_ VDD VSS sky130_fd_sc_hd__inv_2
XFILLER_106_37 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
X_2318_ VSS VDD core.osr.result_r\[11\] _0341_ core.cnb.result_out\[11\] VDD VSS sky130_fd_sc_hd__nand2_1
X_2249_ VSS VDD _0278_ core.cnb.result_out\[4\] _0279_ _0271_ VDD VSS sky130_fd_sc_hd__o21ai_2
XFILLER_82_18 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XFILLER_40_125 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XFILLER_15_89 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XANTENNA__1829__A VSS VDD _1022_ VDD VSS sky130_fd_sc_hd__diode_2
Xgenblk2\[0\].buf_p_rowonn VSS VDD pmatrix_rowon_core_n_buffered\[0\] core.pdc.rowon_out_n\[0\]
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xoutput44 VDD VSS result_out[15] net44 VDD VSS sky130_fd_sc_hd__buf_2
XANTENNA__1696__A1 VSS VDD _1161_ VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA_input23_A VSS VDD config_2_in[14] VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_91_515 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_56_85 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XFILLER_31_125 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XANTENNA__1739__A VSS VDD core.ndc.col_out_n\[18\] VDD VSS sky130_fd_sc_hd__diode_2
X_1620_ VDD VSS _1166_ _1165_ VDD VSS sky130_fd_sc_hd__inv_2
X_1551_ VDD VSS _1107_ _1106_ _1092_ VDD VSS sky130_fd_sc_hd__and2_1
XANTENNA__1474__A VSS VDD _1033_ VDD VSS sky130_fd_sc_hd__diode_2
X_1482_ VDD VSS _1042_ _1041_ VDD VSS sky130_fd_sc_hd__inv_2
XFILLER_97_92 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_86_309 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
X_3152_ VSS VDD net57 _0042_ net69 net52 VDD VSS sky130_fd_sc_hd__dfrtp_1
X_2103_ VDD VSS _1152_ _0146_ core.pdc.col_out\[26\] _0118_ _1102_ _0159_ VDD VSS
+ sky130_fd_sc_hd__a221o_1
X_3083_ VSS VDD _0967_ _0968_ _0060_ _0758_ VDD VSS sky130_fd_sc_hd__o21ai_1
X_2034_ VDD VSS _0116_ _0117_ VDD VSS sky130_fd_sc_hd__clkinv_2
XFILLER_50_423 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XFILLER_50_445 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XFILLER_50_489 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
X_2936_ VSS VDD _0825_ _0726_ _0828_ _0827_ VDD VSS sky130_fd_sc_hd__nand3_1
X_2867_ VSS VDD _0471_ _0761_ _0760_ VDD VSS sky130_fd_sc_hd__nand2_1
X_1818_ VDD VSS _1310_ _1311_ VDD VSS sky130_fd_sc_hd__clkinv_2
X_2798_ VSS VDD _0640_ _0660_ _0693_ _0454_ VDD VSS sky130_fd_sc_hd__nand3_1
XFILLER_117_25 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
X_1749_ VSS VDD _1212_ _1269_ _1177_ VDD VSS sky130_fd_sc_hd__nand2_1
XFILLER_133_13 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XFILLER_93_17 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XFILLER_26_66 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XFILLER_13_125 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_49_501 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XFILLER_49_512 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XANTENNA__1669__A1 VSS VDD _1197_ VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA_genblk2\[14\].buf_p_rowonn_A VSS VDD core.pdc.rowon_out_n\[14\] VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__3014__A VSS VDD _1312_ VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1469__A VSS VDD net14 VDD VSS sky130_fd_sc_hd__diode_2
X_2721_ VSS VDD core.osr.next_result_w\[18\] _0619_ _0533_ VDD VSS sky130_fd_sc_hd__nand2_1
X_2652_ VDD VSS core.osr.next_result_w\[9\] _0535_ _0556_ _0557_ VDD VSS sky130_fd_sc_hd__a21oi_1
X_1603_ VDD VSS core.ndc.col_out_n\[5\] core.ndc.col_out\[5\] VDD VSS sky130_fd_sc_hd__inv_2
X_2583_ VDD VSS _0489_ _1067_ _0500_ _0498_ _1117_ _0439_ VDD VSS sky130_fd_sc_hd__a221o_1
X_1534_ VSS VDD net15 _1092_ VDD VSS sky130_fd_sc_hd__clkbuf_2
X_1465_ VSS VDD core.ndc.rowoff_out_n\[0\] _1025_ _1027_ VDD VSS sky130_fd_sc_hd__nand2_2
X_3204_ VSS VDD net65 core.osr.is_last_sample net84 core.osr.data_valid_r VDD VSS
+ sky130_fd_sc_hd__dfrtp_1
X_3135_ VSS VDD clknet_2_0__leaf_clk_dig_dummy _0025_ net78 core.cnb.result_out\[3\]
+ VDD VSS sky130_fd_sc_hd__dfrtp_1
X_3066_ VSS VDD _0758_ _0953_ _1303_ VDD VSS sky130_fd_sc_hd__nand2_1
X_2017_ VSS VDD _0106_ _1133_ _1390_ _1137_ VDD VSS sky130_fd_sc_hd__mux2_1
XANTENNA__2482__B VSS VDD core.pdc.rowon_out_n\[15\] VDD VSS sky130_fd_sc_hd__diode_2
X_2919_ VSS VDD _0810_ _0730_ _0811_ _0731_ VDD VSS sky130_fd_sc_hd__nand3_1
XFILLER_128_24 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XFILLER_128_79 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XFILLER_88_17 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XANTENNA_fanout73_A VSS VDD net83 VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1561__B VSS VDD _1037_ VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_139_141 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_68_117 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XANTENNA__1471__B VSS VDD core.ndc.rowon_out_n\[0\] VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_83_109 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XANTENNA__1927__A VSS VDD core.ndc.rowon_out_n\[0\] VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_71_1 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
X_2704_ VDD VSS _0604_ _0603_ VDD VSS sky130_fd_sc_hd__inv_2
X_2635_ VDD VSS _0394_ core.cnb.result_out\[0\] _0542_ _0543_ net48 VDD VSS sky130_fd_sc_hd__a22o_1
X_2566_ VDD VSS core.cnb.data_register_r\[0\] _0482_ _1076_ core.cnb.data_register_r\[1\]
+ _0487_ VDD VSS sky130_fd_sc_hd__or4_1
X_1517_ VDD VSS _1075_ _1074_ VDD VSS sky130_fd_sc_hd__buf_2
XFILLER_59_106 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
X_2497_ VSS VDD _0220_ _0439_ _0003_ _0437_ VDD VSS sky130_fd_sc_hd__o21ai_1
XANTENNA__2477__B VSS VDD core.pdc.row_out_n\[10\] VDD VSS sky130_fd_sc_hd__diode_2
X_1448_ VSS VDD _1011_ _1012_ _0985_ VDD VSS sky130_fd_sc_hd__nand2_1
X_3118_ VSS VDD clknet_2_2__leaf_clk_dig_dummy _0018_ net86 core.cnb.shift_register_r\[16\]
+ VDD VSS sky130_fd_sc_hd__dfrtp_1
XFILLER_130_25 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
X_3049_ VSS VDD _0882_ _0868_ _0937_ _0906_ VDD VSS sky130_fd_sc_hd__nand3_1
XFILLER_90_29 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
XFILLER_139_23 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XFILLER_136_133 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
XANTENNA_nmat_rowoff_n[1] VSS VDD core.ndc.rowoff_out_n\[1\] VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_64_74 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XFILLER_9_69 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
Xfanout90 VSS VDD net92 net90 VDD VSS sky130_fd_sc_hd__clkbuf_2
XANTENNA__1747__A VSS VDD _1187_ VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1466__B VSS VDD core.cnb.data_register_r\[8\] VDD VSS sky130_fd_sc_hd__diode_2
X_2420_ VSS VDD _1344_ _1359_ core.ndc.row_out_n\[1\] VDD VSS sky130_fd_sc_hd__nor2_1
XANTENNA__1980__B1 VSS VDD _1259_ VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__3191__CLK VSS VDD clknet_2_1__leaf_clk_dig_dummy VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_89_93 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
X_2351_ VSS VDD _0370_ core.osr.result_r\[15\] core.osr.result_r\[14\] _0358_ VDD
+ VSS sky130_fd_sc_hd__and3_1
X_2282_ VSS VDD _0290_ _0297_ _0298_ _0308_ VDD VSS sky130_fd_sc_hd__o21a_1
XFILLER_92_440 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XFILLER_92_473 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
X_1997_ VDD VSS _0092_ _0091_ VDD VSS sky130_fd_sc_hd__inv_2
XFILLER_133_125 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
X_2618_ VSS VDD _0519_ core.osr.next_result_w\[3\] _0527_ core.osr.next_result_w\[7\]
+ _0526_ _0524_ VDD VSS sky130_fd_sc_hd__o221ai_1
X_2549_ VSS VDD _0472_ _0438_ _0473_ VDD VSS sky130_fd_sc_hd__nor2_1
XFILLER_87_212 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_18_56 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_115_91 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_46_175 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
X_1920_ VDD VSS _1383_ _1382_ _1373_ VDD VSS sky130_fd_sc_hd__or2_1
XFILLER_91_83 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XANTENNA__2861__A VSS VDD _0691_ VDD VSS sky130_fd_sc_hd__diode_2
X_1851_ VSS VDD _1338_ _1326_ core.cnb.data_register_r\[11\] VDD VSS sky130_fd_sc_hd__nand2_2
X_1782_ VDD VSS core.ndc.col_out_n\[26\] core.ndc.col_out\[26\] VDD VSS sky130_fd_sc_hd__clkinv_2
XFILLER_115_103 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
X_2403_ VSS VDD core.osr.sample_count_r\[5\] _0410_ _0412_ VDD VSS sky130_fd_sc_hd__nor2_1
X_2334_ VSS VDD _0355_ _0354_ _0356_ _0241_ VDD VSS sky130_fd_sc_hd__nand3_2
X_2265_ VDD VSS _0293_ _0291_ _0292_ VDD VSS sky130_fd_sc_hd__or2_1
X_2196_ VSS VDD _0228_ _0232_ _0231_ VDD VSS sky130_fd_sc_hd__nand2_1
XFILLER_52_123 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XFILLER_111_38 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XANTENNA_nmat_col_n[5] VSS VDD nmatrix_col_core_n_buffered\[5\] VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_20_57 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XANTENNA_genblk1\[7\].buf_n_coln_A VSS VDD core.ndc.col_out_n\[7\] VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__2011__A VSS VDD _0101_ VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_56_473 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XANTENNA__1760__A VSS VDD _1131_ VDD VSS sky130_fd_sc_hd__diode_2
X_2050_ VDD VSS core.pdc.col_out_n\[14\] core.pdc.col_out\[14\] VDD VSS sky130_fd_sc_hd__clkinv_2
XANTENNA_genblk2\[12\].buf_p_rown_A VSS VDD core.pdc.row_out_n\[12\] VDD VSS sky130_fd_sc_hd__diode_2
X_2952_ VSS VDD _0842_ _0844_ _0843_ VDD VSS sky130_fd_sc_hd__nand2_1
X_1903_ VSS VDD _1342_ _1327_ _1373_ VDD VSS sky130_fd_sc_hd__nor2_1
X_2883_ VDD VSS _0777_ _0776_ VDD VSS sky130_fd_sc_hd__inv_2
X_1834_ VDD VSS core.pdc.row_out_n\[3\] _1323_ VDD VSS sky130_fd_sc_hd__inv_2
X_1765_ VSS VDD core.ndc.col_out_n\[23\] _1278_ VDD VSS sky130_fd_sc_hd__clkbuf_1
XANTENNA__2530__S VSS VDD net54 VDD VSS sky130_fd_sc_hd__diode_2
X_1696_ VSS VDD _1230_ _1161_ _1041_ _1229_ VDD VSS sky130_fd_sc_hd__mux2_1
X_2317_ VSS VDD core.osr.result_r\[11\] core.cnb.result_out\[11\] _0340_ VDD VSS sky130_fd_sc_hd__nor2_1
X_2248_ VDD VSS _0277_ _0276_ _0252_ _0278_ VDD VSS sky130_fd_sc_hd__a21o_1
XANTENNA__1670__A VSS VDD _1033_ VDD VSS sky130_fd_sc_hd__diode_2
X_2179_ VDD VSS _0218_ core.cnb.average_sum_r\[0\] VDD VSS sky130_fd_sc_hd__inv_2
XFILLER_25_145 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XFILLER_15_57 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XFILLER_31_23 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XANTENNA__3102__CLK VSS VDD clknet_2_0__leaf_clk_dig_dummy VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1564__B VSS VDD _1117_ VDD VSS sky130_fd_sc_hd__diode_2
Xoutput45 VDD VSS result_out[1] net45 VDD VSS sky130_fd_sc_hd__buf_2
XANTENNA__2676__A VSS VDD _0395_ VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1580__A VSS VDD core.ndc.col_out\[4\] VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_48_248 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XANTENNA_input16_A VSS VDD config_1_in[8] VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_56_42 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XFILLER_56_281 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
X_1550_ VSS VDD _1106_ _1105_ _1104_ _1103_ _1088_ VDD VSS sky130_fd_sc_hd__a31o_1
XANTENNA_pmat_col[31] VSS VDD core.pdc.col_out\[31\] VDD VSS sky130_fd_sc_hd__diode_2
X_1481_ VSS VDD _1041_ core.ndc.rowon_out_n\[0\] _1040_ VDD VSS sky130_fd_sc_hd__nand2_2
X_3151_ VSS VDD net57 _0041_ net71 net51 VDD VSS sky130_fd_sc_hd__dfrtp_1
X_2102_ VDD VSS _0159_ _0158_ VDD VSS sky130_fd_sc_hd__inv_2
X_3082_ VSS VDD _0758_ _0968_ _1326_ VDD VSS sky130_fd_sc_hd__nand2_1
X_2033_ VSS VDD _1033_ _0115_ _0116_ VDD VSS sky130_fd_sc_hd__nor2_1
XANTENNA__3125__CLK VSS VDD clknet_2_3__leaf_clk_dig_dummy VDD VSS sky130_fd_sc_hd__diode_2
X_2935_ VSS VDD _0826_ _0731_ _0827_ _0725_ VDD VSS sky130_fd_sc_hd__nand3_1
X_2866_ VDD VSS _0760_ _0759_ VDD VSS sky130_fd_sc_hd__inv_2
X_1817_ VSS VDD _1309_ _1038_ _1310_ VDD VSS sky130_fd_sc_hd__nor2_1
XANTENNA__1665__A VSS VDD core.ndc.col_out_n\[9\] VDD VSS sky130_fd_sc_hd__diode_2
X_2797_ VSS VDD _0471_ _0692_ _0686_ VDD VSS sky130_fd_sc_hd__nand2_1
X_1748_ VSS VDD _1221_ _1268_ _1173_ VDD VSS sky130_fd_sc_hd__nand2_1
XFILLER_89_104 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XFILLER_117_37 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
X_1679_ VDD VSS _1217_ _1198_ VDD VSS sky130_fd_sc_hd__inv_2
XANTENNA_input8_A VSS VDD config_1_in[15] VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__2496__A VSS VDD _0438_ VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_93_29 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XFILLER_13_137 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
XANTENNA__1850__A2 VSS VDD _1312_ VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_42_88 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XANTENNA__1575__A VSS VDD _1053_ VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_101_1 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
Xgenblk2\[11\].buf_p_rown VSS VDD pmatrix_row_core_n_buffered\[11\] core.pdc.row_out_n\[11\]
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
XFILLER_49_524 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
X_2720_ VDD VSS _0568_ core.osr.next_result_w\[14\] _0617_ _0618_ VDD VSS sky130_fd_sc_hd__a21oi_1
XFILLER_80_6 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
X_2651_ VDD VSS _1001_ core.osr.next_result_w\[7\] _0530_ _0556_ VDD VSS sky130_fd_sc_hd__a21o_1
X_1602_ VSS VDD _1151_ core.ndc.col_out\[5\] VDD VSS sky130_fd_sc_hd__clkbuf_2
X_2582_ VDD VSS core.cnb.result_out\[6\] _0439_ _0028_ _0497_ _1104_ _0499_ VDD VSS
+ sky130_fd_sc_hd__a221o_1
X_1533_ VSS VDD _1078_ _1090_ _1086_ _1091_ VDD VSS sky130_fd_sc_hd__mux2_2
X_1464_ VSS VDD _1026_ _1027_ VDD VSS sky130_fd_sc_hd__clkbuf_2
X_3203_ VSS VDD net65 _0064_ net78 core.osr.osr_mode_r\[2\] VDD VSS sky130_fd_sc_hd__dfrtp_1
X_3134_ VSS VDD clknet_2_0__leaf_clk_dig_dummy _0024_ net78 core.cnb.result_out\[2\]
+ VDD VSS sky130_fd_sc_hd__dfrtp_1
XFILLER_55_505 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
X_3065_ VSS VDD _0950_ _0781_ _0952_ _0951_ VDD VSS sky130_fd_sc_hd__nand3_1
X_2016_ VDD VSS core.pdc.col_out_n\[9\] core.pdc.col_out\[9\] VDD VSS sky130_fd_sc_hd__clkinv_2
XFILLER_50_221 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XFILLER_10_107 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
X_2918_ VSS VDD _0638_ _0706_ _0810_ VDD VSS sky130_fd_sc_hd__nor2_1
X_2849_ VSS VDD _0744_ _0645_ _0644_ _0654_ _0650_ VDD VSS sky130_fd_sc_hd__and4_1
XANTENNA_nmat_sample_n VSS VDD _0001_ VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA_fanout66_A VSS VDD net67 VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_139_153 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XFILLER_68_129 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XFILLER_73_891 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
X_2703_ VDD VSS core.osr.next_result_w\[8\] net41 _1020_ _0603_ _0562_ VDD VSS sky130_fd_sc_hd__a22o_1
X_2634_ VSS VDD _0983_ _0542_ VDD VSS sky130_fd_sc_hd__clkbuf_2
X_2565_ VSS VDD _0024_ _0486_ VDD VSS sky130_fd_sc_hd__clkbuf_1
X_1516_ VSS VDD _1073_ _1074_ VDD VSS sky130_fd_sc_hd__clkbuf_2
X_2496_ VSS VDD _0438_ _0439_ VDD VSS sky130_fd_sc_hd__clkbuf_2
X_1447_ VDD VSS _1011_ _1009_ VDD VSS sky130_fd_sc_hd__inv_2
X_3117_ VSS VDD clknet_2_2__leaf_clk_dig_dummy _0017_ net93 core.cnb.shift_register_r\[15\]
+ VDD VSS sky130_fd_sc_hd__dfrtp_1
XANTENNA__2774__A VSS VDD _0637_ VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_55_368 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
X_3048_ VSS VDD _0909_ _0922_ _0936_ _0935_ VDD VSS sky130_fd_sc_hd__nand3_1
XFILLER_64_891 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XFILLER_90_19 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XFILLER_23_57 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XFILLER_139_57 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_2_114 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XANTENNA_nmat_rowoff_n[0] VSS VDD core.ndc.rowoff_out_n\[0\] VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_9_15 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XFILLER_70_883 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
Xfanout91 VDD VSS net91 net92 VDD VSS sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout80 VDD VSS net80 net81 VDD VSS sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__2221__A2 VSS VDD _0240_ VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1747__B VSS VDD _1152_ VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1980__A1 VSS VDD _1224_ VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__2859__A VSS VDD core.cnb.pswitch_out\[0\] VDD VSS sky130_fd_sc_hd__diode_2
X_2350_ VSS VDD _0366_ _0369_ _0368_ VDD VSS sky130_fd_sc_hd__nand2_1
X_2281_ VSS VDD _0305_ _0307_ _0306_ VDD VSS sky130_fd_sc_hd__and2b_1
XANTENNA__1799__B2 VSS VDD _1296_ VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1799__A1 VSS VDD _1121_ VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_61_883 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
X_1996_ VSS VDD _1045_ _1169_ _0091_ _1409_ VDD VSS sky130_fd_sc_hd__o21ai_2
XFILLER_133_137 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
X_2617_ VSS VDD _0288_ _0526_ _1002_ VDD VSS sky130_fd_sc_hd__nand2_1
XANTENNA__1673__A VSS VDD _1092_ VDD VSS sky130_fd_sc_hd__diode_2
X_2548_ VDD VSS _0471_ _0472_ VDD VSS sky130_fd_sc_hd__buf_6
Xgenblk1\[12\].buf_p_coln VSS VDD pmatrix_col_core_n_buffered\[12\] core.pdc.col_out_n\[12\]
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
X_2479_ VSS VDD core.pdc.rowon_out_n\[12\] core.pdc.rowoff_out_n\[12\] core.pdc.row_out_n\[12\]
+ VDD VSS sky130_fd_sc_hd__nand2_1
XFILLER_18_13 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_18_68 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
XFILLER_34_23 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XANTENNA__1848__A VSS VDD _1335_ VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_75_41 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XFILLER_61_113 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_131_91 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XANTENNA__2861__B VSS VDD _0208_ VDD VSS sky130_fd_sc_hd__diode_2
X_1850_ VSS VDD _1337_ _1309_ _1312_ _1332_ _1336_ VDD VSS sky130_fd_sc_hd__a31o_1
X_1781_ VSS VDD _1035_ _1143_ _1220_ _1259_ core.ndc.col_out_n\[26\] _1288_ VDD VSS
+ sky130_fd_sc_hd__o221a_1
X_2402_ VDD VSS _0411_ core.osr.next_sample_count_w\[4\] VDD VSS sky130_fd_sc_hd__clkinv_2
X_2333_ VSS VDD _0353_ _0355_ core.osr.result_r\[12\] VDD VSS sky130_fd_sc_hd__nand2_1
XANTENNA__2902__B1 VSS VDD _1076_ VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__2101__B VSS VDD _1072_ VDD VSS sky130_fd_sc_hd__diode_2
X_2264_ VSS VDD _0286_ _0292_ _0282_ VDD VSS sky130_fd_sc_hd__nand2_1
X_2195_ VDD VSS _0231_ core.cnb.average_sum_r\[3\] VDD VSS sky130_fd_sc_hd__inv_2
XFILLER_52_102 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XANTENNA_nmat_col_n[4] VSS VDD nmatrix_col_core_n_buffered\[4\] VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_52_179 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XANTENNA__1668__A VSS VDD _1206_ VDD VSS sky130_fd_sc_hd__diode_2
X_1979_ VSS VDD _0077_ _0078_ _1155_ VDD VSS sky130_fd_sc_hd__nand2_1
XFILLER_121_118 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
Xgenblk2\[6\].buf_n_rowonn VSS VDD nmatrix_rowon_core_n_buffered\[6\] core.ndc.rowon_out_n\[6\]
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
XANTENNA__2011__B VSS VDD _1275_ VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_45_11 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_43_113 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XFILLER_43_124 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XANTENNA__3181__CLK VSS VDD clknet_2_1__leaf_clk_dig_dummy VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1578__A VSS VDD _1126_ VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1760__B VSS VDD _1243_ VDD VSS sky130_fd_sc_hd__diode_2
X_2951_ VSS VDD _0753_ _0843_ VDD VSS sky130_fd_sc_hd__clkinvlp_2
X_1902_ VSS VDD core.pdc.rowoff_out_n\[5\] core.pdc.rowon_out_n\[4\] _1325_ VDD VSS
+ sky130_fd_sc_hd__nand2_1
X_2882_ VSS VDD _0774_ _0776_ _0775_ VDD VSS sky130_fd_sc_hd__nand2_1
X_1833_ VSS VDD _1322_ core.pdc.rowoff_out_n\[8\] _1323_ _1321_ VDD VSS sky130_fd_sc_hd__o21ai_2
X_1764_ VSS VDD _1278_ _1277_ _1276_ _1274_ VDD VSS sky130_fd_sc_hd__and3_1
X_1695_ VSS VDD _1136_ _1229_ _1228_ VDD VSS sky130_fd_sc_hd__nand2_1
X_2316_ VSS VDD _0338_ _0339_ _0328_ VDD VSS sky130_fd_sc_hd__nand2_1
X_2247_ VSS VDD _0275_ _0277_ _0274_ VDD VSS sky130_fd_sc_hd__nand2_1
XFILLER_122_38 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XANTENNA__2103__A1 VSS VDD _1152_ VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__2103__B2 VSS VDD _1102_ VDD VSS sky130_fd_sc_hd__diode_2
X_2178_ VSS VDD core.cnb.next_average_counter_w\[4\] _0217_ VDD VSS sky130_fd_sc_hd__clkbuf_1
XFILLER_53_466 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XFILLER_40_149 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XFILLER_31_68 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_31_57 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
XFILLER_31_46 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XANTENNA__1917__A1 VSS VDD core.ndc.rowoff_out_n\[5\] VDD VSS sky130_fd_sc_hd__diode_2
Xoutput46 VDD VSS result_out[2] net46 VDD VSS sky130_fd_sc_hd__buf_2
XFILLER_56_32 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
XFILLER_56_293 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XANTENNA__1605__B1 VSS VDD _1135_ VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__2030__B1 VSS VDD _1259_ VDD VSS sky130_fd_sc_hd__diode_2
Xgenblk2\[13\].buf_n_rown VSS VDD nmatrix_row_core_n_buffered\[13\] core.ndc.row_out_n\[13\]
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
X_1480_ VSS VDD _1040_ _1038_ _1039_ VDD VSS sky130_fd_sc_hd__nand2_2
XFILLER_98_116 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
X_3150_ VSS VDD net57 _0040_ net69 net50 VDD VSS sky130_fd_sc_hd__dfrtp_1
X_3081_ VSS VDD _0965_ _0691_ _0967_ _0966_ VDD VSS sky130_fd_sc_hd__nand3_1
X_2101_ VSS VDD _0077_ _0158_ _1072_ VDD VSS sky130_fd_sc_hd__nand2_1
X_2032_ VSS VDD _1389_ _1201_ _1199_ _0115_ VDD VSS sky130_fd_sc_hd__mux2_2
X_2934_ VSS VDD _0826_ _0762_ _0645_ _0722_ VDD VSS sky130_fd_sc_hd__and3_1
X_2865_ VSS VDD _0677_ _0713_ _0759_ VDD VSS sky130_fd_sc_hd__nor2_1
X_1816_ VDD VSS _1309_ _1308_ VDD VSS sky130_fd_sc_hd__buf_2
X_2796_ VSS VDD core.cnb.data_register_r\[0\] _0690_ _0687_ _0210_ _0050_ _0691_ VDD
+ VSS sky130_fd_sc_hd__o221a_1
XANTENNA__2021__B1 VSS VDD _1064_ VDD VSS sky130_fd_sc_hd__diode_2
X_1747_ VSS VDD _1187_ _1267_ _1152_ VDD VSS sky130_fd_sc_hd__nand2_1
X_1678_ VDD VSS core.ndc.col_out\[10\] core.ndc.col_out_n\[10\] VDD VSS sky130_fd_sc_hd__inv_2
XANTENNA__2012__A0 VSS VDD _1186_ VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_107_93 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XANTENNA__2618__A2 VSS VDD core.osr.next_result_w\[3\] VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__2079__B1 VSS VDD _1125_ VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_83_85 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
X_2650_ VDD VSS _0554_ _0553_ _0555_ _0040_ VDD VSS sky130_fd_sc_hd__a21o_1
X_1601_ VSS VDD _1144_ _1150_ _1140_ _1151_ VDD VSS sky130_fd_sc_hd__or3b_1
X_2581_ VSS VDD _0439_ _0498_ _0499_ VDD VSS sky130_fd_sc_hd__nor2_1
X_1532_ VSS VDD _1036_ _1089_ _1090_ VDD VSS sky130_fd_sc_hd__nor2_1
X_1463_ VDD VSS _1026_ net14 VDD VSS sky130_fd_sc_hd__dlymetal6s2s_1
X_3202_ VSS VDD net64 _0063_ net78 core.osr.osr_mode_r\[1\] VDD VSS sky130_fd_sc_hd__dfrtp_1
Xgenblk1\[17\].buf_p_coln VSS VDD pmatrix_col_core_n_buffered\[17\] core.pdc.col_out_n\[17\]
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
XFILLER_55_517 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
X_3133_ VSS VDD clknet_2_0__leaf_clk_dig_dummy _0023_ net84 core.cnb.result_out\[1\]
+ VDD VSS sky130_fd_sc_hd__dfrtp_2
XFILLER_94_141 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
X_3064_ VSS VDD _0942_ _0902_ _0951_ _0948_ VDD VSS sky130_fd_sc_hd__nand3_1
X_2015_ VDD VSS core.pdc.col_out_n\[9\] _0105_ VDD VSS sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_90_380 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_10_119 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
X_2917_ VSS VDD _0454_ _0808_ _0809_ VDD VSS sky130_fd_sc_hd__nor2_1
XFILLER_12_59 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
X_2848_ VSS VDD _0738_ _0742_ _0743_ VDD VSS sky130_fd_sc_hd__nor2_1
X_2779_ VSS VDD _0672_ _0675_ _0674_ VDD VSS sky130_fd_sc_hd__nand2_1
XANTENNA__3188__RESET_B VSS VDD net87 VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_37_45 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XFILLER_46_517 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XANTENNA_fanout59_A VSS VDD net61 VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1586__A VSS VDD _1135_ VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_78_63 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_78_85 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XANTENNA__3115__CLK VSS VDD clknet_2_2__leaf_clk_dig_dummy VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_76_141 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XFILLER_91_122 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
X_2702_ VSS VDD _0599_ _0602_ _0601_ VDD VSS sky130_fd_sc_hd__nand2_1
X_2633_ VDD VSS _0541_ _0537_ core.osr.next_result_w\[2\] VDD VSS sky130_fd_sc_hd__or2_1
XFILLER_57_1 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
X_2564_ VSS VDD _0486_ core.cnb.result_out\[2\] _0480_ _0485_ VDD VSS sky130_fd_sc_hd__mux2_1
X_1515_ VDD VSS _1073_ _1072_ VDD VSS sky130_fd_sc_hd__inv_2
X_2495_ VSS VDD _0438_ _0208_ core.cnb.shift_register_r\[2\] VDD VSS sky130_fd_sc_hd__nand2_2
X_1446_ VSS VDD _1009_ _1010_ core.osr.sample_count_r\[2\] VDD VSS sky130_fd_sc_hd__nand2_1
XANTENNA_clkbuf_2_3__f_clk_dig_dummy_A VSS VDD clknet_0_clk_dig_dummy VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_67_130 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_55_325 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
X_3116_ VSS VDD clknet_2_2__leaf_clk_dig_dummy _0016_ net93 core.cnb.shift_register_r\[14\]
+ VDD VSS sky130_fd_sc_hd__dfrtp_1
XFILLER_82_122 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
X_3047_ VSS VDD _0934_ _0935_ _0906_ VDD VSS sky130_fd_sc_hd__nand2_1
XFILLER_130_38 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XANTENNA__3097__S VSS VDD _0241_ VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_139_69 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
Xgenblk1\[14\].buf_n_coln VDD VSS core.ndc.col_out_n\[14\] nmatrix_col_core_n_buffered\[14\]
+ VDD VSS sky130_fd_sc_hd__buf_6
XANTENNA__2949__B VSS VDD _0482_ VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__3138__CLK VSS VDD clknet_2_0__leaf_clk_dig_dummy VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_48_11 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XFILLER_58_141 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
XFILLER_46_314 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_73_100 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_0_29 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
Xgenblk2\[14\].buf_p_rowonn VSS VDD pmatrix_rowon_core_n_buffered\[14\] core.pdc.rowon_out_n\[14\]
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
XFILLER_54_380 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
XFILLER_120_60 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_80_31 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
Xfanout92 VDD VSS net92 net94 VDD VSS sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout70 VSS VDD net83 net70 VDD VSS sky130_fd_sc_hd__clkbuf_2
Xfanout81 VDD VSS net81 net82 VDD VSS sky130_fd_sc_hd__buf_2
XFILLER_127_113 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XANTENNA__2205__A VSS VDD core.cnb.result_out\[0\] VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1763__B VSS VDD _1188_ VDD VSS sky130_fd_sc_hd__diode_2
X_2280_ VSS VDD core.osr.result_r\[8\] _0306_ core.cnb.result_out\[8\] VDD VSS sky130_fd_sc_hd__nand2_1
XFILLER_29_5 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_92_453 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_52_339 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
X_1995_ VDD VSS _0090_ _0089_ VDD VSS sky130_fd_sc_hd__inv_2
X_2616_ VDD VSS _0523_ net46 _0395_ _0036_ _0525_ VDD VSS sky130_fd_sc_hd__a22o_1
XANTENNA__1954__A VSS VDD _1272_ VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_133_149 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
X_2547_ VDD VSS _0470_ _0471_ VDD VSS sky130_fd_sc_hd__buf_6
X_2478_ VSS VDD core.pdc.row_out_n\[11\] core.pdc.rowoff_out_n\[11\] core.pdc.rowon_out_n\[11\]
+ VDD VSS sky130_fd_sc_hd__nand2_1
X_1429_ VSS VDD core.osr.osr_mode_r\[2\] _0989_ _0993_ VDD VSS sky130_fd_sc_hd__nor2_1
XFILLER_18_25 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XFILLER_51_361 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XANTENNA__2025__A VSS VDD _0101_ VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_109_124 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
XFILLER_50_78 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
XFILLER_93_206 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XFILLER_75_53 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XFILLER_46_199 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XFILLER_131_81 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
Xnmat_sample_buf VSS VDD nmat_sample_switch_buffered net55 VDD VSS sky130_fd_sc_hd__clkbuf_1
XFILLER_91_63 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
X_1780_ VSS VDD _1149_ _1288_ _1284_ VDD VSS sky130_fd_sc_hd__nand2_1
XANTENNA__1774__A VSS VDD _1095_ VDD VSS sky130_fd_sc_hd__diode_2
X_2401_ VDD VSS _0410_ core.osr.is_last_sample _0409_ _0411_ VDD VSS sky130_fd_sc_hd__or3_1
X_2332_ VDD VSS _0354_ core.osr.result_r\[12\] _0353_ VDD VSS sky130_fd_sc_hd__or2_1
X_2263_ VDD VSS _0291_ _0289_ _0290_ VDD VSS sky130_fd_sc_hd__and2_1
XFILLER_84_228 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
X_2194_ VSS VDD core.cnb.next_average_sum_w\[2\] _0230_ VDD VSS sky130_fd_sc_hd__clkbuf_1
XFILLER_92_261 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
XANTENNA_nmat_col_n[3] VSS VDD nmatrix_col_core_n_buffered\[3\] VDD VSS sky130_fd_sc_hd__diode_2
X_1978_ VSS VDD _0077_ _1146_ _1400_ _1147_ VDD VSS sky130_fd_sc_hd__mux2_1
XFILLER_121_108 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XANTENNA_nmat_col[19] VSS VDD core.ndc.col_out\[19\] VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_48_409 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XFILLER_29_57 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_28_144 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XFILLER_90_209 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XFILLER_83_272 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
XANTENNA__1859__A VSS VDD _1325_ VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1578__B VSS VDD _1129_ VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_101_84 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_6_17 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XANTENNA__1594__A VSS VDD _1074_ VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_120_141 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XANTENNA__1533__S VSS VDD _1078_ VDD VSS sky130_fd_sc_hd__diode_2
X_2950_ VSS VDD _0832_ _0842_ _0833_ VDD VSS sky130_fd_sc_hd__nand2_1
XANTENNA__1488__B VSS VDD _1047_ VDD VSS sky130_fd_sc_hd__diode_2
X_1901_ VSS VDD core.pdc.rowoff_out_n\[5\] _1372_ _1309_ VDD VSS sky130_fd_sc_hd__nand2_2
X_2881_ VSS VDD _0771_ _0772_ _0775_ _0482_ VDD VSS sky130_fd_sc_hd__nand3_1
X_1832_ VDD VSS _1308_ _1304_ _1038_ _1300_ _1322_ VDD VSS sky130_fd_sc_hd__or4_1
X_1763_ VSS VDD _1180_ _1277_ _1188_ VDD VSS sky130_fd_sc_hd__nand2_1
X_1694_ VDD VSS _1228_ _1105_ VDD VSS sky130_fd_sc_hd__inv_2
XFILLER_106_29 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
X_2315_ VSS VDD _0326_ _0338_ _0330_ VDD VSS sky130_fd_sc_hd__nand2_1
X_2246_ VDD VSS _0276_ _0274_ _0275_ VDD VSS sky130_fd_sc_hd__or2_1
X_2177_ VSS VDD _0217_ _0216_ _0215_ _0210_ VDD VSS sky130_fd_sc_hd__and3_1
XFILLER_25_103 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
Xclkbuf_2_1__f_clk_dig_dummy VSS VDD clknet_0_clk_dig_dummy clknet_2_1__leaf_clk_dig_dummy
+ VDD VSS sky130_fd_sc_hd__clkbuf_16
Xgenblk1\[24\].buf_p_coln VSS VDD pmatrix_col_core_n_buffered\[24\] core.pdc.col_out_n\[24\]
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xoutput47 VDD VSS result_out[3] net47 VDD VSS sky130_fd_sc_hd__buf_2
Xoutput36 VDD VSS conversion_finished_osr_out net36 VDD VSS sky130_fd_sc_hd__buf_2
XANTENNA__2957__B VSS VDD core.cnb.data_register_r\[1\] VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1550__B1 VSS VDD _1088_ VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_56_77 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
XFILLER_56_99 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_56_272 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XFILLER_16_147 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XANTENNA__1589__A VSS VDD _1138_ VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA_genblk1\[3\].buf_n_coln_A VSS VDD core.ndc.col_out_n\[3\] VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1605__A1 VSS VDD _1078_ VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__2030__A1 VSS VDD _1074_ VDD VSS sky130_fd_sc_hd__diode_2
X_3080_ VSS VDD _0964_ _0966_ _0955_ VDD VSS sky130_fd_sc_hd__nand2_1
X_2100_ VDD VSS core.pdc.col_out_n\[25\] core.pdc.col_out\[25\] VDD VSS sky130_fd_sc_hd__inv_2
X_2031_ VDD VSS core.pdc.col_out_n\[12\] core.pdc.col_out\[12\] VDD VSS sky130_fd_sc_hd__clkinv_2
XFILLER_22_106 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
X_2933_ VSS VDD _0821_ _0824_ _0825_ VDD VSS sky130_fd_sc_hd__nor2_1
XFILLER_87_1 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
X_2864_ VSS VDD _0051_ _0757_ _0755_ _0721_ core.cnb.data_register_r\[1\] _0758_ VDD
+ VSS sky130_fd_sc_hd__a32o_1
X_1815_ VSS VDD core.cnb.data_register_r\[11\] _1308_ VDD VSS sky130_fd_sc_hd__clkbuf_2
X_2795_ VSS VDD _0460_ _0691_ _0670_ VDD VSS sky130_fd_sc_hd__nor2_2
XANTENNA__1946__B VSS VDD _1155_ VDD VSS sky130_fd_sc_hd__diode_2
X_1746_ VDD VSS core.ndc.col_out\[19\] core.ndc.col_out_n\[19\] VDD VSS sky130_fd_sc_hd__inv_2
XANTENNA__2021__A1 VSS VDD _1224_ VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__2123__A VSS VDD _1039_ VDD VSS sky130_fd_sc_hd__diode_2
X_1677_ VSS VDD _1216_ core.ndc.col_out_n\[10\] VDD VSS sky130_fd_sc_hd__clkbuf_2
XANTENNA__3171__CLK VSS VDD net61 VDD VSS sky130_fd_sc_hd__diode_2
Xgenblk1\[19\].buf_n_coln VDD VSS core.ndc.col_out_n\[19\] nmatrix_col_core_n_buffered\[19\]
+ VDD VSS sky130_fd_sc_hd__buf_6
XANTENNA__1681__B VSS VDD _1173_ VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_85_312 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
X_2229_ VSS VDD _0259_ _0261_ _0258_ VDD VSS sky130_fd_sc_hd__nand2_1
XFILLER_26_25 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XANTENNA__2796__C1 VSS VDD _0691_ VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__2012__A1 VSS VDD _1197_ VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__2033__A VSS VDD _1033_ VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_107_50 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
XFILLER_107_72 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_67_65 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XANTENNA_input21_A VSS VDD config_2_in[12] VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__2079__A1 VSS VDD _1102_ VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_83_53 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XFILLER_91_337 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XANTENNA__2208__A VSS VDD _0241_ VDD VSS sky130_fd_sc_hd__diode_2
Xgenblk1\[21\].buf_n_coln VDD VSS core.ndc.col_out_n\[21\] nmatrix_col_core_n_buffered\[21\]
+ VDD VSS sky130_fd_sc_hd__buf_6
XFILLER_83_97 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_8_110 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
X_1600_ VSS VDD _1149_ _1150_ _1032_ VDD VSS sky130_fd_sc_hd__nand2_1
X_2580_ VSS VDD _0489_ _0498_ _1160_ VDD VSS sky130_fd_sc_hd__nand2_1
X_1531_ VDD VSS _1089_ _1088_ VDD VSS sky130_fd_sc_hd__inv_2
X_1462_ VSS VDD _1024_ _1025_ core.cnb.data_register_r\[11\] VDD VSS sky130_fd_sc_hd__nand2_1
X_3201_ VSS VDD net65 _0062_ net78 core.osr.osr_mode_r\[0\] VDD VSS sky130_fd_sc_hd__dfrtp_2
X_3132_ VSS VDD clknet_2_0__leaf_clk_dig_dummy _0022_ net84 core.cnb.result_out\[0\]
+ VDD VSS sky130_fd_sc_hd__dfrtp_2
X_3063_ VSS VDD _0944_ _0950_ _0949_ VDD VSS sky130_fd_sc_hd__nand2_1
X_2014_ VSS VDD _0105_ _0104_ _0102_ _0100_ VDD VSS sky130_fd_sc_hd__and3_1
XFILLER_90_392 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
X_2916_ VSS VDD _0807_ _0808_ _0725_ VDD VSS sky130_fd_sc_hd__nand2_1
X_2847_ VSS VDD _0742_ _0649_ _0724_ _0741_ VDD VSS sky130_fd_sc_hd__and3_1
X_2778_ VSS VDD _0674_ _0640_ _0652_ _0673_ VDD VSS sky130_fd_sc_hd__nand3b_1
XANTENNA__1692__A VSS VDD core.ndc.col_out_n\[12\] VDD VSS sky130_fd_sc_hd__diode_2
X_1729_ VDD VSS _1255_ _1074_ _1243_ VDD VSS sky130_fd_sc_hd__or2_1
XFILLER_37_13 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_46_507 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XFILLER_37_57 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XANTENNA__1992__B1 VSS VDD _1082_ VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_78_75 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XFILLER_78_97 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XFILLER_76_131 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XFILLER_91_134 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XANTENNA__2880__B VSS VDD core.cnb.pswitch_out\[2\] VDD VSS sky130_fd_sc_hd__diode_2
X_2701_ VDD VSS _0601_ _0600_ VDD VSS sky130_fd_sc_hd__inv_2
X_2632_ VSS VDD _1019_ _0540_ VDD VSS sky130_fd_sc_hd__clkbuf_2
X_2563_ VSS VDD _0483_ _0485_ _0484_ VDD VSS sky130_fd_sc_hd__or2b_1
X_1514_ VSS VDD _1071_ _1072_ net15 VDD VSS sky130_fd_sc_hd__nor2_2
X_2494_ VDD VSS _0437_ core.cnb.is_holding_result_w VDD VSS sky130_fd_sc_hd__inv_2
X_1445_ VSS VDD _1008_ _1009_ core.osr.osr_mode_r\[1\] VDD VSS sky130_fd_sc_hd__nor2_2
XFILLER_67_142 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
X_3115_ VSS VDD clknet_2_2__leaf_clk_dig_dummy _0015_ net93 core.cnb.shift_register_r\[13\]
+ VDD VSS sky130_fd_sc_hd__dfrtp_1
XFILLER_55_337 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
X_3046_ VSS VDD _0928_ _0933_ _0934_ _0870_ VDD VSS sky130_fd_sc_hd__o21ai_1
XFILLER_82_134 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
XANTENNA_fanout71_A VSS VDD net73 VDD VSS sky130_fd_sc_hd__diode_2
Xfanout60 VSS VDD net60 net61 VDD VSS sky130_fd_sc_hd__clkbuf_1
Xfanout71 VSS VDD net73 net71 VDD VSS sky130_fd_sc_hd__clkbuf_2
Xfanout82 VDD VSS net82 net83 VDD VSS sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_80_65 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XFILLER_127_103 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XANTENNA__1965__B1 VSS VDD _1125_ VDD VSS sky130_fd_sc_hd__diode_2
Xfanout93 VDD VSS net93 net94 VDD VSS sky130_fd_sc_hd__buf_2
XFILLER_127_125 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_49_197 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XFILLER_92_465 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
X_1994_ VSS VDD _1394_ _1242_ _1202_ _0089_ VDD VSS sky130_fd_sc_hd__mux2_2
XANTENNA__2115__B VSS VDD _1096_ VDD VSS sky130_fd_sc_hd__diode_2
Xgenblk1\[29\].buf_p_coln VSS VDD pmatrix_col_core_n_buffered\[29\] core.pdc.col_out_n\[29\]
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
X_2615_ VDD VSS _0525_ _0524_ core.osr.next_result_w\[6\] VDD VSS sky130_fd_sc_hd__or2_1
XANTENNA__2131__A VSS VDD core.cnb.data_register_r\[2\] VDD VSS sky130_fd_sc_hd__diode_2
X_2546_ VDD VSS _0469_ _0468_ _0470_ _0203_ VDD VSS sky130_fd_sc_hd__a21boi_2
XFILLER_125_28 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
X_2477_ VSS VDD core.pdc.rowon_out_n\[10\] core.pdc.rowoff_out_n\[10\] core.pdc.row_out_n\[10\]
+ VDD VSS sky130_fd_sc_hd__nand2_1
X_1428_ VDD VSS _0992_ _0991_ VDD VSS sky130_fd_sc_hd__inv_2
XFILLER_18_37 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XFILLER_55_101 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XFILLER_83_421 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
X_3029_ VDD VSS _0916_ _0830_ _0856_ _0917_ VDD VSS sky130_fd_sc_hd__a21o_1
XFILLER_51_373 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XANTENNA__3105__CLK VSS VDD clknet_2_2__leaf_clk_dig_dummy VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_50_24 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XANTENNA__2025__B VSS VDD _1093_ VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_50_35 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XANTENNA__1947__B1 VSS VDD _1259_ VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_124_128 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XFILLER_59_77 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
Xgenblk1\[31\].buf_p_coln VSS VDD pmatrix_col_core_n_buffered\[31\] core.pdc.col_out_n\[31\]
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
XFILLER_61_137 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XANTENNA_genblk2\[1\].buf_n_rown_A VSS VDD core.ndc.row_out_n\[1\] VDD VSS sky130_fd_sc_hd__diode_2
X_2400_ VSS VDD _0999_ _0406_ _0410_ VDD VSS sky130_fd_sc_hd__nor2_1
X_2331_ VSS VDD _0353_ _0351_ _0309_ _0352_ VDD VSS sky130_fd_sc_hd__a21bo_1
X_2262_ VSS VDD core.cnb.result_out\[6\] _0290_ core.osr.result_r\[6\] VDD VSS sky130_fd_sc_hd__nand2_1
X_2193_ VSS VDD _0230_ _0229_ _0228_ _0209_ VDD VSS sky130_fd_sc_hd__and3_1
XANTENNA_nmat_col_n[2] VSS VDD nmatrix_col_core_n_buffered\[2\] VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA_genblk2\[0\].buf_p_rowonn_A VSS VDD core.pdc.rowon_out_n\[0\] VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__3128__CLK VSS VDD clknet_2_3__leaf_clk_dig_dummy VDD VSS sky130_fd_sc_hd__diode_2
X_1977_ VDD VSS _0076_ _0075_ VDD VSS sky130_fd_sc_hd__inv_2
XANTENNA__1684__B VSS VDD _1177_ VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA_genblk2\[1\].buf_n_rowonn_A VSS VDD core.ndc.rowon_out_n\[1\] VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA_nmat_col[18] VSS VDD core.ndc.col_out\[18\] VDD VSS sky130_fd_sc_hd__diode_2
X_2529_ VSS VDD _0018_ _0456_ VDD VSS sky130_fd_sc_hd__clkbuf_1
XFILLER_29_69 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_56_421 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_45_57 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_43_148 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XFILLER_101_41 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_51_181 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
Xgenblk1\[26\].buf_n_coln VSS VDD nmatrix_col_core_n_buffered\[26\] core.ndc.col_out_n\[26\]
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
XFILLER_101_96 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_6_29 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_10_93 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XFILLER_86_64 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_86_53 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XFILLER_47_421 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XANTENNA__1769__B VSS VDD _1213_ VDD VSS sky130_fd_sc_hd__diode_2
X_1900_ VSS VDD _1023_ _1372_ _1022_ VDD VSS sky130_fd_sc_hd__nand2_1
X_2880_ VSS VDD _0773_ _0774_ core.cnb.pswitch_out\[2\] VDD VSS sky130_fd_sc_hd__nand2_1
X_1831_ VSS VDD _1321_ _1318_ core.pdc.rowoff_out_n\[8\] _1311_ core.pdc.row_out_n\[2\]
+ VDD VSS sky130_fd_sc_hd__o22a_1
XANTENNA__1785__A VSS VDD _1124_ VDD VSS sky130_fd_sc_hd__diode_2
X_1762_ VSS VDD _1187_ _1276_ _1275_ VDD VSS sky130_fd_sc_hd__nand2_1
X_1693_ VDD VSS _1227_ _1073_ VDD VSS sky130_fd_sc_hd__buf_2
XFILLER_103_109 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XFILLER_106_19 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
X_2314_ VDD VSS _0337_ core.osr.next_result_w\[10\] VDD VSS sky130_fd_sc_hd__buf_6
X_2245_ VSS VDD _0267_ _0275_ _0265_ VDD VSS sky130_fd_sc_hd__nand2_1
X_2176_ VSS VDD _0214_ _0216_ core.cnb.average_counter_r\[4\] VDD VSS sky130_fd_sc_hd__nand2_1
Xoutput48 VDD VSS result_out[4] net48 VDD VSS sky130_fd_sc_hd__buf_2
Xoutput37 VDD VSS conversion_finished_out net65 VDD VSS sky130_fd_sc_hd__buf_2
XANTENNA_genblk1\[18\].buf_n_coln_A VSS VDD core.ndc.col_out_n\[18\] VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_88_398 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XANTENNA__1605__A2 VSS VDD _1105_ VDD VSS sky130_fd_sc_hd__diode_2
Xgenblk2\[2\].buf_n_rowonn VSS VDD nmatrix_rowon_core_n_buffered\[2\] core.ndc.rowon_out_n\[2\]
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
XANTENNA_pmat_col[4] VSS VDD core.pdc.col_out\[4\] VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__2030__A2 VSS VDD _0113_ VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_137_81 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
X_2030_ VSS VDD _1259_ _0088_ _0113_ _1074_ core.pdc.col_out_n\[12\] _0114_ VDD VSS
+ sky130_fd_sc_hd__o221a_1
XFILLER_22_118 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
X_2932_ VSS VDD _0737_ _0813_ _0824_ _0823_ VDD VSS sky130_fd_sc_hd__nand3_1
XFILLER_94_3 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
X_2863_ VSS VDD _0688_ _0758_ VDD VSS sky130_fd_sc_hd__clkbuf_2
X_1814_ VSS VDD _1300_ _1306_ _1307_ VDD VSS sky130_fd_sc_hd__nor2_1
X_2794_ VDD VSS _0690_ _0689_ _0686_ VDD VSS sky130_fd_sc_hd__and2_1
X_1745_ VSS VDD _1266_ core.ndc.col_out_n\[19\] VDD VSS sky130_fd_sc_hd__clkbuf_2
XFILLER_7_94 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
X_1676_ VSS VDD _1216_ _1215_ _1214_ _1211_ VDD VSS sky130_fd_sc_hd__and3_1
XFILLER_85_302 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
X_2228_ VDD VSS _0260_ _0258_ _0259_ VDD VSS sky130_fd_sc_hd__or2_1
X_2159_ VSS VDD _0203_ _0189_ _0202_ VDD VSS sky130_fd_sc_hd__nand2_2
XANTENNA__2796__B1 VSS VDD core.cnb.data_register_r\[0\] VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_42_69 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XANTENNA__2033__B VSS VDD _0115_ VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA_pmat_analog_in VSS VDD ANTENNA_pmat_analog_in/DIODE VDD VSS sky130_fd_sc_hd__diode_2
Xpmat_95 VSS VDD net95 pmat_95/HI VDD VSS sky130_fd_sc_hd__conb_1
XFILLER_107_84 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XFILLER_91_305 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XANTENNA_input14_A VSS VDD config_1_in[6] VDD VSS sky130_fd_sc_hd__diode_2
X_1530_ VSS VDD _1088_ _1085_ _1087_ VDD VSS sky130_fd_sc_hd__nor2_4
X_1461_ VSS VDD _1022_ _1023_ _1024_ VDD VSS sky130_fd_sc_hd__nor2_1
X_3200_ VSS VDD net64 core.osr.next_sample_count_w\[8\] net77 core.osr.sample_count_r\[8\]
+ VDD VSS sky130_fd_sc_hd__dfrtp_1
X_3131_ VSS VDD clknet_2_3__leaf_clk_dig_dummy core.cnb.next_average_sum_w\[4\] net91
+ core.cnb.average_sum_r\[4\] VDD VSS sky130_fd_sc_hd__dfrtp_1
XANTENNA_genblk2\[5\].buf_p_rowonn_A VSS VDD core.pdc.rowon_bottotop_n\[5\] VDD VSS
+ sky130_fd_sc_hd__diode_2
XANTENNA_nmat_col_n[19] VSS VDD nmatrix_col_core_n_buffered\[19\] VDD VSS sky130_fd_sc_hd__diode_2
X_3062_ VDD VSS _0949_ _0948_ VDD VSS sky130_fd_sc_hd__inv_2
X_2013_ VSS VDD _0103_ _0104_ _1101_ VDD VSS sky130_fd_sc_hd__nand2_1
XFILLER_76_891 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
X_2915_ VSS VDD _0807_ _0694_ _0644_ _0722_ VDD VSS sky130_fd_sc_hd__and3_1
XFILLER_12_17 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
X_2846_ VSS VDD _0646_ _0634_ _0740_ _0741_ VDD VSS sky130_fd_sc_hd__nor3_1
X_2777_ VSS VDD _0653_ _0673_ core.cnb.shift_register_r\[11\] VDD VSS sky130_fd_sc_hd__nand2_1
X_1728_ VDD VSS core.ndc.col_out\[16\] core.ndc.col_out_n\[16\] VDD VSS sky130_fd_sc_hd__inv_2
X_1659_ VSS VDD _1059_ _1052_ _1201_ _1200_ VDD VSS sky130_fd_sc_hd__o21ai_1
XANTENNA_input6_A VSS VDD config_1_in[13] VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_37_25 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_37_69 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_67_891 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XFILLER_53_24 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_53_57 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XANTENNA__1992__A1 VSS VDD _1114_ VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_5_136 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XFILLER_94_53 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XFILLER_91_146 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_73_883 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
X_2700_ VSS VDD core.osr.next_result_w\[10\] _1019_ _0600_ _1011_ VDD VSS sky130_fd_sc_hd__o21ai_1
XANTENNA__1793__A VSS VDD core.ndc.col_out\[28\] VDD VSS sky130_fd_sc_hd__diode_2
X_2631_ VSS VDD _0534_ _0536_ _0539_ _0538_ VDD VSS sky130_fd_sc_hd__nand3_1
X_2562_ VSS VDD _0478_ _0484_ _0482_ VDD VSS sky130_fd_sc_hd__nand2_1
X_1513_ VDD VSS _1071_ core.cnb.data_register_r\[8\] VDD VSS sky130_fd_sc_hd__inv_2
XFILLER_4_40 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
X_2493_ VSS VDD _0220_ _0434_ _0002_ core.cnb.enable_loop_out VDD VSS sky130_fd_sc_hd__o21ai_1
X_1444_ VDD VSS _0993_ _1008_ VDD VSS sky130_fd_sc_hd__clkinv_2
X_3114_ VSS VDD clknet_2_2__leaf_clk_dig_dummy _0014_ net93 core.cnb.shift_register_r\[12\]
+ VDD VSS sky130_fd_sc_hd__dfrtp_2
X_3045_ VSS VDD _0931_ _1114_ _0933_ _0932_ VDD VSS sky130_fd_sc_hd__nand3_1
XFILLER_64_883 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
X_2829_ VSS VDD _0642_ _0724_ VDD VSS sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout64_A VSS VDD net66 VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_64_45 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XANTENNA__3184__CLK VSS VDD clknet_2_1__leaf_clk_dig_dummy VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_64_89 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XFILLER_54_393 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
Xfanout61 VSS VDD net67 net61 VDD VSS sky130_fd_sc_hd__clkbuf_2
Xfanout72 VDD VSS net72 net73 VDD VSS sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout83 VSS VDD net34 net83 VDD VSS sky130_fd_sc_hd__clkbuf_2
Xfanout94 VDD VSS net94 net34 VDD VSS sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__1965__A1 VSS VDD _1121_ VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_127_137 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XANTENNA__1965__B2 VSS VDD _1413_ VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_64_113 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
XFILLER_92_477 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
X_1993_ VDD VSS _0088_ _0087_ VDD VSS sky130_fd_sc_hd__inv_2
X_2614_ VSS VDD _0994_ _0524_ VDD VSS sky130_fd_sc_hd__clkbuf_2
X_2545_ VDD VSS _0469_ _0222_ _0207_ VDD VSS sky130_fd_sc_hd__or2_1
X_2476_ VSS VDD core.pdc.row_out_n\[9\] core.pdc.rowoff_out_n\[9\] core.pdc.rowon_out_n\[9\]
+ VDD VSS sky130_fd_sc_hd__nand2_1
X_1427_ VSS VDD _0991_ core.osr.osr_mode_r\[2\] _0990_ _0989_ VDD VSS sky130_fd_sc_hd__and3_1
XFILLER_83_400 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
XFILLER_83_433 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
X_3028_ VSS VDD _0916_ _0818_ _0751_ _0910_ VDD VSS sky130_fd_sc_hd__and3_1
XFILLER_83_477 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XANTENNA__1698__A VSS VDD _1227_ VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_133_7 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XANTENNA__1947__A1 VSS VDD _1224_ VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_50_47 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_109_137 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
Xgenblk2\[4\].buf_p_rown VSS VDD pmatrix_row_core_n_buffered\[4\] core.pdc.row_out_n\[4\]
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
XFILLER_93_219 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
Xgenblk2\[10\].buf_p_rowonn VSS VDD pmatrix_rowon_core_n_buffered\[10\] core.pdc.rowon_out_n\[10\]
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
X_2330_ VSS VDD _0352_ _0350_ _0342_ _0329_ _0343_ _0324_ VDD VSS sky130_fd_sc_hd__a221oi_1
X_2261_ VDD VSS _0289_ core.cnb.result_out\[6\] core.osr.result_r\[6\] VDD VSS sky130_fd_sc_hd__or2_1
XFILLER_34_5 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
X_2192_ VSS VDD _0223_ _0229_ _0226_ VDD VSS sky130_fd_sc_hd__nand2_1
XFILLER_37_113 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_92_241 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XANTENNA_nmat_col_n[1] VSS VDD nmatrix_col_core_n_buffered\[1\] VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_92_296 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
X_1976_ VSS VDD _0075_ _1208_ _1394_ _1197_ VDD VSS sky130_fd_sc_hd__mux2_1
XANTENNA__2142__A VSS VDD core.cnb.sampled_avg_control_r\[0\] VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_106_107 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XANTENNA_nmat_col[17] VSS VDD core.ndc.col_out\[17\] VDD VSS sky130_fd_sc_hd__diode_2
X_2528_ VSS VDD _0456_ net54 _0219_ _0454_ VDD VSS sky130_fd_sc_hd__mux2_1
X_2459_ VSS VDD core.ndc.rowon_out_n\[4\] core.ndc.rowoff_out_n\[4\] core.ndc.row_out_n\[4\]
+ VDD VSS sky130_fd_sc_hd__nand2_1
XANTENNA__2106__B2 VSS VDD _1102_ VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__2106__A1 VSS VDD _1125_ VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_56_433 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_56_477 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_61_24 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_101_53 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XANTENNA__2036__B VSS VDD _1235_ VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_51_193 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_61_57 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XANTENNA__2052__A VSS VDD _1227_ VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_126_50 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_19_113 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XFILLER_86_76 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XFILLER_19_124 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_34_116 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
X_1830_ VDD VSS _1321_ _1320_ VDD VSS sky130_fd_sc_hd__inv_2
XFILLER_89_6 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XANTENNA__1785__B VSS VDD _1275_ VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__2584__A1 VSS VDD core.cnb.result_out\[7\] VDD VSS sky130_fd_sc_hd__diode_2
X_1761_ VDD VSS _1275_ _1072_ VDD VSS sky130_fd_sc_hd__buf_2
X_1692_ VDD VSS core.ndc.col_out\[12\] core.ndc.col_out_n\[12\] VDD VSS sky130_fd_sc_hd__inv_2
Xgenblk2\[1\].buf_n_rown VSS VDD nmatrix_row_core_n_buffered\[1\] core.ndc.row_out_n\[1\]
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
X_2313_ VDD VSS _0337_ _0334_ _0336_ VDD VSS sky130_fd_sc_hd__and2_1
XFILLER_25_1 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
X_2244_ VDD VSS _0274_ _0272_ _0273_ VDD VSS sky130_fd_sc_hd__and2_1
X_2175_ VDD VSS _0215_ core.cnb.average_counter_r\[4\] _0214_ VDD VSS sky130_fd_sc_hd__or2_1
XANTENNA_cgen_dlycontrol4_in[5] VSS VDD net8 VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__2024__B1 VSS VDD _1208_ VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__2575__A1 VSS VDD core.cnb.result_out\[4\] VDD VSS sky130_fd_sc_hd__diode_2
X_1959_ VDD VSS _1411_ _1410_ VDD VSS sky130_fd_sc_hd__inv_2
Xoutput49 VDD VSS result_out[5] net49 VDD VSS sky130_fd_sc_hd__buf_2
Xoutput38 VDD VSS result_out[0] net38 VDD VSS sky130_fd_sc_hd__buf_2
XANTENNA__2600__A VSS VDD _1328_ VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_88_355 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XANTENNA__1550__A2 VSS VDD _1104_ VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_16_116 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XANTENNA__2047__A VSS VDD _1413_ VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_112_85 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XANTENNA_pmat_col[3] VSS VDD core.pdc.col_out\[3\] VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_137_93 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XANTENNA__3118__CLK VSS VDD clknet_2_2__leaf_clk_dig_dummy VDD VSS sky130_fd_sc_hd__diode_2
X_2931_ VSS VDD _0822_ _0730_ _0823_ _0731_ VDD VSS sky130_fd_sc_hd__nand3_1
XFILLER_30_141 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
X_2862_ VDD VSS _0757_ _0756_ VDD VSS sky130_fd_sc_hd__inv_2
X_1813_ VSS VDD _1302_ _1306_ _1305_ VDD VSS sky130_fd_sc_hd__nand2_1
X_2793_ VDD VSS _0688_ _0689_ VDD VSS sky130_fd_sc_hd__clkinv_4
X_1744_ VSS VDD _1266_ _1265_ _1264_ _1262_ VDD VSS sky130_fd_sc_hd__and3_1
Xgenblk2\[7\].buf_p_rowonn VSS VDD pmatrix_rowon_core_n_buffered\[7\] core.pdc.rowon_out_n\[7\]
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
X_1675_ VSS VDD _1138_ _1215_ _1177_ VDD VSS sky130_fd_sc_hd__nand2_1
X_2227_ VSS VDD _0249_ _0259_ _0247_ VDD VSS sky130_fd_sc_hd__nand2_1
X_2158_ VSS VDD _0200_ _0202_ _0201_ VDD VSS sky130_fd_sc_hd__nand2_1
X_2089_ VDD VSS _0151_ _0152_ VDD VSS sky130_fd_sc_hd__clkinv_2
XANTENNA__2796__A1 VSS VDD _0210_ VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_88_141 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XFILLER_91_317 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XFILLER_83_33 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_91_328 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XFILLER_16_60 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XFILLER_8_145 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
X_1460_ VSS VDD core.cnb.data_register_r\[9\] _1023_ core.cnb.data_register_r\[8\]
+ VDD VSS sky130_fd_sc_hd__nand2_1
XFILLER_79_141 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
X_3130_ VSS VDD clknet_2_3__leaf_clk_dig_dummy core.cnb.next_average_sum_w\[3\] net91
+ core.cnb.average_sum_r\[3\] VDD VSS sky130_fd_sc_hd__dfrtp_1
XFILLER_94_100 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XANTENNA_nmat_col_n[18] VSS VDD nmatrix_col_core_n_buffered\[18\] VDD VSS sky130_fd_sc_hd__diode_2
X_3061_ VSS VDD _0946_ _0948_ _0947_ VDD VSS sky130_fd_sc_hd__nand2_1
X_2012_ VSS VDD _0103_ _1197_ _1394_ _1186_ VDD VSS sky130_fd_sc_hd__mux2_1
X_2914_ VSS VDD _0806_ _0454_ _0730_ _0725_ VDD VSS sky130_fd_sc_hd__and3_1
XANTENNA__2134__B VSS VDD core.cnb.sampled_avg_control_r\[0\] VDD VSS sky130_fd_sc_hd__diode_2
X_2845_ VSS VDD _0653_ _0740_ _0739_ VDD VSS sky130_fd_sc_hd__nand2_1
XFILLER_12_29 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XFILLER_128_29 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
X_2776_ VSS VDD _0669_ _0660_ _0672_ _0671_ VDD VSS sky130_fd_sc_hd__nand3_1
X_1727_ VDD VSS core.ndc.col_out_n\[16\] _1254_ VDD VSS sky130_fd_sc_hd__buf_2
X_1658_ VDD VSS _1200_ _1055_ VDD VSS sky130_fd_sc_hd__inv_2
X_1589_ VDD VSS _1139_ _1138_ VDD VSS sky130_fd_sc_hd__inv_2
Xgenblk2\[9\].buf_p_rown VSS VDD pmatrix_row_core_n_buffered\[9\] core.pdc.row_out_n\[9\]
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
XFILLER_85_133 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XFILLER_37_37 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XFILLER_53_36 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_139_113 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XANTENNA__2325__A VSS VDD core.cnb.result_out\[11\] VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_89_461 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_91_158 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XFILLER_91_169 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
X_2630_ VSS VDD _0519_ _0279_ _0537_ _0538_ VDD VSS sky130_fd_sc_hd__o21a_1
XANTENNA__3066__A VSS VDD _0758_ VDD VSS sky130_fd_sc_hd__diode_2
X_2561_ VSS VDD _0482_ _0478_ _0483_ VDD VSS sky130_fd_sc_hd__nor2_1
X_2492_ VSS VDD _2492_/X _0436_ VDD VSS sky130_fd_sc_hd__buf_1
X_1512_ VSS VDD _1070_ _1069_ _1054_ _1067_ VDD VSS sky130_fd_sc_hd__mux2_1
X_1443_ VDD VSS _0999_ _0994_ core.osr.sample_count_r\[6\] _1007_ VDD VSS sky130_fd_sc_hd__a21o_1
XFILLER_4_52 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_4_85 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
X_3113_ VSS VDD clknet_2_3__leaf_clk_dig_dummy _0013_ net93 core.cnb.shift_register_r\[11\]
+ VDD VSS sky130_fd_sc_hd__dfrtp_2
XANTENNA__2448__B1 VSS VDD core.pdc.rowon_bottotop_n\[5\] VDD VSS sky130_fd_sc_hd__diode_2
X_3044_ VSS VDD _0930_ _0932_ _0918_ VDD VSS sky130_fd_sc_hd__nand2_1
Xgenblk1\[4\].buf_p_coln VSS VDD pmatrix_col_core_n_buffered\[4\] core.pdc.col_out_n\[4\]
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
X_2828_ VSS VDD _0723_ _0644_ _0679_ _0722_ VDD VSS sky130_fd_sc_hd__and3_1
X_2759_ VSS VDD _0649_ _0652_ _0655_ _0654_ VDD VSS sky130_fd_sc_hd__nand3_1
XFILLER_86_464 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
XFILLER_46_328 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
XFILLER_46_339 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
XFILLER_86_486 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XANTENNA_fanout57_A VSS VDD net58 VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_64_57 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XANTENNA__1662__A1 VSS VDD _1199_ VDD VSS sky130_fd_sc_hd__diode_2
Xfanout73 VSS VDD net83 net73 VDD VSS sky130_fd_sc_hd__clkbuf_2
Xfanout62 VDD VSS net62 net63 VDD VSS sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout84 VSS VDD net85 net84 VDD VSS sky130_fd_sc_hd__clkbuf_2
XFILLER_80_78 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
XFILLER_13_61 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
Xgenblk2\[6\].buf_n_rown VSS VDD nmatrix_row_core_n_buffered\[6\] core.ndc.row_out_n\[6\]
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
XFILLER_49_100 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_49_122 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_92_412 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XFILLER_52_309 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_92_489 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
X_1992_ VSS VDD _1082_ _1114_ _0087_ _1412_ VDD VSS sky130_fd_sc_hd__o21ai_2
X_2613_ VSS VDD _0519_ core.osr.next_result_w\[2\] core.osr.next_result_w\[4\] _1003_
+ _0523_ _0520_ VDD VSS sky130_fd_sc_hd__o221a_1
XFILLER_133_108 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
X_2544_ VDD VSS _0466_ _0465_ _0467_ _0468_ VDD VSS sky130_fd_sc_hd__a21oi_1
X_2475_ VSS VDD core.pdc.row_out_n\[7\] core.pdc.rowoff_out_n\[7\] core.pdc.rowon_out_n\[7\]
+ VDD VSS sky130_fd_sc_hd__nand2_1
X_1426_ VDD VSS _0990_ core.osr.osr_mode_r\[1\] VDD VSS sky130_fd_sc_hd__inv_2
XFILLER_83_445 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XFILLER_83_467 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
X_3027_ VDD VSS _0915_ _0914_ VDD VSS sky130_fd_sc_hd__inv_2
XFILLER_83_489 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_50_59 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XFILLER_132_141 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
Xgenblk1\[1\].buf_n_coln VDD VSS core.ndc.col_out_n\[1\] nmatrix_col_core_n_buffered\[1\]
+ VDD VSS sky130_fd_sc_hd__buf_6
XFILLER_115_52 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XFILLER_46_169 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XANTENNA__3181__RESET_B VSS VDD net86 VDD VSS sky130_fd_sc_hd__diode_2
X_2260_ VDD VSS core.osr.next_result_w\[5\] _0288_ VDD VSS sky130_fd_sc_hd__inv_2
X_2191_ VDD VSS _0228_ _0227_ VDD VSS sky130_fd_sc_hd__inv_2
XFILLER_37_136 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XFILLER_37_125 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
XFILLER_1_53 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XANTENNA_nmat_col_n[0] VSS VDD nmatrix_col_core_n_buffered\[0\] VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_92_253 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XFILLER_92_275 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XFILLER_92_286 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
X_1975_ VSS VDD _0074_ _1141_ _1389_ _1111_ VDD VSS sky130_fd_sc_hd__mux2_1
Xpmat pmatrix_row_core_n_buffered\[0\] pmatrix_row_core_n_buffered\[1\] pmatrix_row_core_n_buffered\[2\]
+ pmatrix_row_core_n_buffered\[3\] pmatrix_row_core_n_buffered\[4\] pmatrix_row_core_n_buffered\[5\]
+ pmatrix_row_core_n_buffered\[6\] pmatrix_row_core_n_buffered\[7\] pmatrix_row_core_n_buffered\[8\]
+ pmatrix_row_core_n_buffered\[9\] pmatrix_row_core_n_buffered\[10\] pmatrix_row_core_n_buffered\[11\]
+ pmatrix_row_core_n_buffered\[12\] pmatrix_row_core_n_buffered\[13\] pmatrix_row_core_n_buffered\[14\]
+ pmatrix_row_core_n_buffered\[15\] pmatrix_rowon_core_n_buffered\[0\] pmatrix_rowon_core_n_buffered\[1\]
+ pmatrix_rowon_core_n_buffered\[2\] pmatrix_rowon_core_n_buffered\[3\] pmatrix_rowon_core_n_buffered\[4\]
+ pmatrix_rowon_core_n_buffered\[5\] pmatrix_rowon_core_n_buffered\[6\] pmatrix_rowon_core_n_buffered\[7\]
+ pmatrix_rowon_core_n_buffered\[8\] pmatrix_rowon_core_n_buffered\[9\] pmatrix_rowon_core_n_buffered\[10\]
+ pmatrix_rowon_core_n_buffered\[11\] pmatrix_rowon_core_n_buffered\[12\] pmatrix_rowon_core_n_buffered\[13\]
+ pmatrix_rowon_core_n_buffered\[14\] pmatrix_rowon_core_n_buffered\[15\] core.pdc.rowoff_out_n\[0\]
+ core.pdc.rowoff_out_n\[1\] core.pdc.rowoff_out_n\[2\] core.pdc.rowoff_out_n\[3\]
+ core.pdc.rowoff_out_n\[4\] core.pdc.rowoff_out_n\[5\] core.pdc.rowoff_out_n\[6\]
+ core.pdc.rowoff_out_n\[7\] core.pdc.rowoff_out_n\[8\] core.pdc.rowoff_out_n\[9\]
+ core.pdc.rowoff_out_n\[10\] core.pdc.rowoff_out_n\[11\] core.pdc.rowoff_out_n\[12\]
+ core.pdc.rowoff_out_n\[13\] core.pdc.rowoff_out_n\[14\] core.pdc.rowoff_out_n\[15\]
+ vcm/vcm sample_pmatrix_cgen _0000_ pmatrix_col_core_n_buffered\[31\] pmatrix_col_core_n_buffered\[30\]
+ pmatrix_col_core_n_buffered\[29\] pmatrix_col_core_n_buffered\[28\] pmatrix_col_core_n_buffered\[27\]
+ pmatrix_col_core_n_buffered\[26\] pmatrix_col_core_n_buffered\[25\] pmatrix_col_core_n_buffered\[24\]
+ pmatrix_col_core_n_buffered\[23\] pmatrix_col_core_n_buffered\[22\] pmatrix_col_core_n_buffered\[21\]
+ pmatrix_col_core_n_buffered\[20\] pmatrix_col_core_n_buffered\[19\] pmatrix_col_core_n_buffered\[18\]
+ pmatrix_col_core_n_buffered\[17\] pmatrix_col_core_n_buffered\[16\] pmatrix_col_core_n_buffered\[15\]
+ pmatrix_col_core_n_buffered\[14\] pmatrix_col_core_n_buffered\[13\] pmatrix_col_core_n_buffered\[12\]
+ pmatrix_col_core_n_buffered\[11\] pmatrix_col_core_n_buffered\[10\] pmatrix_col_core_n_buffered\[9\]
+ pmatrix_col_core_n_buffered\[8\] pmatrix_col_core_n_buffered\[7\] pmatrix_col_core_n_buffered\[6\]
+ pmatrix_col_core_n_buffered\[5\] pmatrix_col_core_n_buffered\[4\] pmatrix_col_core_n_buffered\[3\]
+ pmatrix_col_core_n_buffered\[2\] pmatrix_col_core_n_buffered\[1\] pmatrix_col_core_n_buffered\[0\]
+ core.cnb.data_register_r\[2\] core.cnb.data_register_r\[1\] core.cnb.data_register_r\[0\]
+ net95 pmat_sample_switch_buffered pmat_sample_switch_n_buffered inp_analog core.pdc.col_out\[0\]
+ core.pdc.col_out\[1\] core.pdc.col_out\[2\] core.pdc.col_out\[3\] core.pdc.col_out\[4\]
+ core.pdc.col_out\[5\] core.pdc.col_out\[6\] core.pdc.col_out\[7\] core.pdc.col_out\[8\]
+ core.pdc.col_out\[9\] core.pdc.col_out\[10\] core.pdc.col_out\[11\] core.pdc.col_out\[12\]
+ core.pdc.col_out\[13\] core.pdc.col_out\[14\] core.pdc.col_out\[15\] core.pdc.col_out\[16\]
+ core.pdc.col_out\[17\] core.pdc.col_out\[18\] core.pdc.col_out\[19\] core.pdc.col_out\[20\]
+ core.pdc.col_out\[21\] core.pdc.col_out\[22\] core.pdc.col_out\[23\] core.pdc.col_out\[24\]
+ core.pdc.col_out\[25\] core.pdc.col_out\[26\] core.pdc.col_out\[27\] core.pdc.col_out\[28\]
+ core.pdc.col_out\[29\] core.pdc.col_out\[30\] core.pdc.col_out\[31\] VDD VSS ctop_pmatrix_analog
+ adc_array_matrix_12bit
XFILLER_20_29 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_106_119 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_136_29 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XANTENNA__3174__CLK VSS VDD net58 VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_114_152 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XANTENNA_nmat_col[16] VSS VDD core.ndc.col_out\[16\] VDD VSS sky130_fd_sc_hd__diode_2
X_2527_ VSS VDD _0017_ _0455_ VDD VSS sky130_fd_sc_hd__clkbuf_1
XFILLER_88_515 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
X_2458_ VSS VDD core.ndc.row_out_n\[3\] core.ndc.rowoff_out_n\[3\] core.ndc.rowon_out_n\[3\]
+ VDD VSS sky130_fd_sc_hd__nand2_1
X_2389_ VSS VDD _0985_ _0397_ _0401_ VDD VSS sky130_fd_sc_hd__nor2_1
XFILLER_28_136 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XFILLER_56_445 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XFILLER_56_489 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_83_253 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
XANTENNA__1502__A VSS VDD _1053_ VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__2317__B VSS VDD core.cnb.result_out\[11\] VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_61_36 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XFILLER_61_69 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_126_62 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_120_122 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_19_136 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XANTENNA__2243__A VSS VDD core.cnb.result_out\[4\] VDD VSS sky130_fd_sc_hd__diode_2
X_1760_ VDD VSS _1274_ _1131_ _1243_ VDD VSS sky130_fd_sc_hd__or2_1
X_1691_ VSS VDD _1035_ _1225_ _1153_ _1224_ core.ndc.col_out_n\[12\] _1226_ VDD VSS
+ sky130_fd_sc_hd__o221a_2
X_2312_ VSS VDD _0251_ _0336_ _0335_ VDD VSS sky130_fd_sc_hd__nand2_1
XFILLER_111_100 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
X_2243_ VSS VDD core.cnb.result_out\[4\] _0273_ core.osr.result_r\[4\] VDD VSS sky130_fd_sc_hd__nand2_1
X_2174_ VDD VSS _0214_ _0193_ VDD VSS sky130_fd_sc_hd__inv_2
XANTENNA_cgen_dlycontrol4_in[4] VSS VDD net7 VDD VSS sky130_fd_sc_hd__diode_2
X_1958_ VSS VDD _1047_ _1057_ _1410_ _1409_ VDD VSS sky130_fd_sc_hd__o21ai_2
X_1889_ VSS VDD _1306_ _1362_ core.pdc.rowon_out_n\[1\] _1364_ VDD VSS sky130_fd_sc_hd__o21ai_2
Xoutput39 VDD VSS result_out[10] net39 VDD VSS sky130_fd_sc_hd__buf_2
XFILLER_102_111 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XANTENNA__1550__A3 VSS VDD _1105_ VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_56_14 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
XFILLER_56_220 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XFILLER_16_128 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_112_42 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XANTENNA__2047__B VSS VDD _1235_ VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA_pmat_col[2] VSS VDD core.pdc.col_out\[2\] VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_97_43 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
Xgenblk1\[9\].buf_p_coln VSS VDD pmatrix_col_core_n_buffered\[9\] core.pdc.col_out_n\[9\]
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
XFILLER_90_510 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
X_2930_ VSS VDD _0638_ _0766_ _0822_ VDD VSS sky130_fd_sc_hd__nor2_1
XFILLER_15_150 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
X_2861_ VSS VDD _0691_ _0756_ _0208_ VDD VSS sky130_fd_sc_hd__nand2_1
X_1812_ VDD VSS _1305_ _1304_ VDD VSS sky130_fd_sc_hd__inv_2
X_2792_ VSS VDD _0208_ _0688_ _0670_ VDD VSS sky130_fd_sc_hd__nor2_2
X_1743_ VDD VSS _1265_ _1227_ _1225_ VDD VSS sky130_fd_sc_hd__or2_1
X_1674_ VSS VDD _1212_ _1214_ _1213_ VDD VSS sky130_fd_sc_hd__nand2_1
XFILLER_97_131 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
X_2226_ VDD VSS _0258_ _0256_ _0257_ VDD VSS sky130_fd_sc_hd__and2_1
X_2157_ VDD VSS _0201_ core.cnb.average_counter_r\[4\] _0187_ VDD VSS sky130_fd_sc_hd__or2_1
XFILLER_26_17 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XANTENNA__2493__A1 VSS VDD core.cnb.enable_loop_out VDD VSS sky130_fd_sc_hd__diode_2
X_2088_ VSS VDD _1227_ _0072_ _0151_ VDD VSS sky130_fd_sc_hd__nor2_1
XFILLER_13_109 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XANTENNA_fanout87_A VSS VDD net94 VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_107_42 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XFILLER_67_57 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XFILLER_67_46 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XFILLER_123_96 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
XFILLER_83_45 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XANTENNA_genblk1\[14\].buf_n_coln_A VSS VDD core.ndc.col_out_n\[14\] VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA_nmat_col_n[17] VSS VDD nmatrix_col_core_n_buffered\[17\] VDD VSS sky130_fd_sc_hd__diode_2
X_3060_ VSS VDD _0945_ _0947_ _0507_ VDD VSS sky130_fd_sc_hd__nand2_1
X_2011_ VSS VDD _0101_ _0102_ _1275_ VDD VSS sky130_fd_sc_hd__nand2_1
XFILLER_90_340 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XFILLER_50_237 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
X_2913_ VDD VSS _0805_ _0804_ VDD VSS sky130_fd_sc_hd__inv_2
X_2844_ VDD VSS _0739_ core.cnb.shift_register_r\[11\] VDD VSS sky130_fd_sc_hd__inv_2
XANTENNA__1738__B1 VSS VDD _1035_ VDD VSS sky130_fd_sc_hd__diode_2
X_2775_ VSS VDD core.cnb.shift_register_r\[16\] _0670_ _0671_ VDD VSS sky130_fd_sc_hd__nor2_1
X_1726_ VSS VDD _1254_ _1253_ _1252_ _1250_ VDD VSS sky130_fd_sc_hd__and3_1
X_1657_ VDD VSS _1052_ _1199_ _1059_ _1036_ VDD VSS sky130_fd_sc_hd__o21ai_4
X_1588_ VSS VDD _1138_ _1137_ _1077_ _1133_ VDD VSS sky130_fd_sc_hd__mux2_1
Xgenblk1\[6\].buf_n_coln VDD VSS core.ndc.col_out_n\[6\] nmatrix_col_core_n_buffered\[6\]
+ VDD VSS sky130_fd_sc_hd__buf_6
X_2209_ VDD VSS _0239_ core.osr.next_result_w\[0\] _0242_ VDD VSS sky130_fd_sc_hd__xor2_1
X_3189_ VSS VDD clknet_2_1__leaf_clk_dig_dummy _0059_ net81 core.cnb.data_register_r\[9\]
+ VDD VSS sky130_fd_sc_hd__dfrtp_2
XANTENNA__3108__CLK VSS VDD clknet_2_3__leaf_clk_dig_dummy VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_53_48 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XANTENNA__1510__A VSS VDD _1047_ VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__2325__B VSS VDD _0255_ VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_139_125 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_118_41 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_118_85 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_78_45 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XFILLER_89_440 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XFILLER_89_473 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_91_104 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XFILLER_94_88 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XANTENNA__1968__B1 VSS VDD _1088_ VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_64_6 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XANTENNA__2251__A VSS VDD core.cnb.result_out\[5\] VDD VSS sky130_fd_sc_hd__diode_2
X_2560_ VSS VDD core.cnb.data_register_r\[2\] _0482_ VDD VSS sky130_fd_sc_hd__clkbuf_2
X_2491_ VDD VSS net17 _1040_ net16 _0436_ VDD VSS sky130_fd_sc_hd__or3_1
X_1511_ VSS VDD _1068_ _1069_ _1037_ VDD VSS sky130_fd_sc_hd__nor2_2
X_1442_ VSS VDD _1006_ _1005_ _0998_ _0997_ _0988_ VDD VSS sky130_fd_sc_hd__and4_1
XFILLER_4_97 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XANTENNA__3082__A VSS VDD _0758_ VDD VSS sky130_fd_sc_hd__diode_2
X_3112_ VSS VDD clknet_2_3__leaf_clk_dig_dummy _0012_ net93 core.cnb.shift_register_r\[10\]
+ VDD VSS sky130_fd_sc_hd__dfrtp_1
X_3043_ VDD VSS _0831_ _0930_ _0856_ _0931_ VDD VSS sky130_fd_sc_hd__a21o_1
XFILLER_139_29 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
X_2827_ VDD VSS _0722_ _0659_ VDD VSS sky130_fd_sc_hd__inv_2
X_2758_ VSS VDD core.cnb.shift_register_r\[11\] _0653_ _0654_ VDD VSS sky130_fd_sc_hd__nor2_1
X_1709_ VSS VDD _1240_ _1241_ _1213_ VDD VSS sky130_fd_sc_hd__nand2_1
X_2689_ VSS VDD core.osr.next_result_w\[13\] _0590_ _0535_ VDD VSS sky130_fd_sc_hd__nand2_1
XANTENNA__1505__A VSS VDD core.ndc.col_out_n\[0\] VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_86_498 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XFILLER_64_14 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
Xfanout74 VDD VSS net74 net76 VDD VSS sky130_fd_sc_hd__buf_2
Xfanout63 VDD VSS net63 net66 VDD VSS sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout85 VDD VSS net85 net87 VDD VSS sky130_fd_sc_hd__buf_2
XFILLER_13_73 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
XFILLER_89_33 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XANTENNA__2071__A VSS VDD _0081_ VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_89_44 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_89_281 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XFILLER_49_134 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XFILLER_38_81 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XFILLER_49_178 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
X_1991_ VDD VSS core.pdc.col_out_n\[6\] core.pdc.col_out\[6\] VDD VSS sky130_fd_sc_hd__clkinv_2
XANTENNA__2602__A1 VSS VDD core.cnb.result_out\[11\] VDD VSS sky130_fd_sc_hd__diode_2
X_2612_ VDD VSS _0521_ net45 _0395_ _0035_ _0522_ VDD VSS sky130_fd_sc_hd__a22o_1
X_2543_ VSS VDD _0181_ _0207_ _0467_ core.cnb.average_sum_r\[1\] VDD VSS sky130_fd_sc_hd__o21ai_1
X_2474_ VSS VDD core.pdc.rowon_out_n\[6\] core.pdc.rowoff_out_n\[6\] core.pdc.row_out_n\[6\]
+ VDD VSS sky130_fd_sc_hd__nand2_1
X_1425_ VDD VSS _0989_ core.osr.osr_mode_r\[0\] VDD VSS sky130_fd_sc_hd__inv_2
XFILLER_18_29 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XANTENNA__1979__B VSS VDD _1155_ VDD VSS sky130_fd_sc_hd__diode_2
X_3026_ VSS VDD _0475_ _0914_ _0913_ _1117_ _0911_ VDD VSS sky130_fd_sc_hd__o211ai_1
XFILLER_34_17 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XFILLER_51_310 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
XFILLER_91_490 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
XFILLER_51_398 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
Xnmat_sample_buf_n VSS VDD nmat_sample_switch_n_buffered core.cnb.enable_loop_out
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
XANTENNA__1995__A VSS VDD _0089_ VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_59_25 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XFILLER_132_153 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XFILLER_132_131 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XFILLER_75_68 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
XFILLER_75_57 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XFILLER_131_30 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
X_2190_ VSS VDD _0226_ _0223_ _0227_ VDD VSS sky130_fd_sc_hd__nor2_1
XFILLER_1_21 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
X_1974_ VDD VSS core.pdc.col_out\[4\] core.pdc.col_out_n\[4\] VDD VSS sky130_fd_sc_hd__clkinv_2
XFILLER_136_19 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XFILLER_114_131 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
XANTENNA_nmat_col[15] VSS VDD core.ndc.col_out\[15\] VDD VSS sky130_fd_sc_hd__diode_2
X_2526_ VSS VDD _0455_ _0454_ _0219_ core.cnb.shift_register_r\[15\] VDD VSS sky130_fd_sc_hd__mux2_1
X_2457_ VSS VDD core.ndc.row_out_n\[2\] core.ndc.rowoff_out_n\[2\] core.ndc.rowon_out_n\[2\]
+ VDD VSS sky130_fd_sc_hd__nand2_1
XFILLER_29_17 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
X_2388_ VSS VDD core.osr.sample_count_r\[2\] _0398_ _0400_ VDD VSS sky130_fd_sc_hd__nor2_1
XFILLER_45_38 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
X_3009_ VSS VDD _0884_ _0877_ _0898_ _0895_ VDD VSS sky130_fd_sc_hd__nand3_1
XFILLER_10_41 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XFILLER_10_52 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XFILLER_126_85 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XFILLER_126_74 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XFILLER_120_134 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
XANTENNA__3058__A1 VSS VDD _0799_ VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_35_82 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
X_1690_ VSS VDD _1172_ _1226_ _1093_ VDD VSS sky130_fd_sc_hd__nand2_1
XANTENNA__1792__B2 VSS VDD _1125_ VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__2897__C VSS VDD _1395_ VDD VSS sky130_fd_sc_hd__diode_2
X_2311_ VDD VSS _0335_ core.cnb.result_out\[10\] VDD VSS sky130_fd_sc_hd__inv_2
X_2242_ VDD VSS _0272_ core.cnb.result_out\[4\] core.osr.result_r\[4\] VDD VSS sky130_fd_sc_hd__or2_1
X_2173_ VSS VDD core.cnb.next_average_counter_w\[3\] _0213_ VDD VSS sky130_fd_sc_hd__clkbuf_1
XANTENNA__1603__A VSS VDD core.ndc.col_out\[5\] VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__2137__C VSS VDD core.cnb.sampled_avg_control_r\[0\] VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA_cgen_dlycontrol4_in[3] VSS VDD net6 VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__3141__CLK VSS VDD clknet_2_0__leaf_clk_dig_dummy VDD VSS sky130_fd_sc_hd__diode_2
X_1957_ VDD VSS _1409_ _1400_ VDD VSS sky130_fd_sc_hd__buf_2
X_1888_ VSS VDD _1363_ _1364_ _1303_ VDD VSS sky130_fd_sc_hd__nor2_2
X_2509_ VSS VDD _0446_ core.cnb.shift_register_r\[8\] _0444_ core.cnb.shift_register_r\[7\]
+ VDD VSS sky130_fd_sc_hd__mux2_1
XFILLER_102_123 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XANTENNA__1513__A VSS VDD core.cnb.data_register_r\[8\] VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA_genblk2\[2\].buf_p_rown_A VSS VDD core.pdc.row_out_n\[2\] VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_112_54 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_112_98 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_90_522 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
X_2860_ VSS VDD _0718_ _0754_ _0755_ _0719_ VDD VSS sky130_fd_sc_hd__nand3_1
X_1811_ VSS VDD _1303_ _1304_ core.cnb.data_register_r\[10\] VDD VSS sky130_fd_sc_hd__nand2_1
X_2791_ VSS VDD _0686_ _0687_ core.cnb.data_register_r\[0\] VDD VSS sky130_fd_sc_hd__nand2_1
X_1742_ VDD VSS _1263_ _1264_ VDD VSS sky130_fd_sc_hd__clkinv_2
X_1673_ VDD VSS _1213_ _1092_ VDD VSS sky130_fd_sc_hd__buf_2
XFILLER_97_143 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
X_2225_ VSS VDD core.cnb.result_out\[2\] _0257_ core.osr.result_r\[2\] VDD VSS sky130_fd_sc_hd__nand2_1
XANTENNA__2429__A VSS VDD _1342_ VDD VSS sky130_fd_sc_hd__diode_2
X_2156_ VSS VDD _0193_ _0196_ _0200_ _0199_ VDD VSS sky130_fd_sc_hd__nand3_1
XFILLER_26_29 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XANTENNA__2493__A2 VSS VDD _0220_ VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_53_235 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XFILLER_53_246 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XFILLER_93_393 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
X_2087_ VDD VSS core.pdc.col_out\[22\] core.pdc.col_out_n\[22\] VDD VSS sky130_fd_sc_hd__clkinv_2
XANTENNA_nmat_sample_buf_A VSS VDD net55 VDD VSS sky130_fd_sc_hd__diode_2
X_2989_ VSS VDD _0877_ _0879_ _0878_ VDD VSS sky130_fd_sc_hd__nand2_1
XFILLER_123_42 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
XANTENNA__3187__CLK VSS VDD clknet_2_1__leaf_clk_dig_dummy VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_83_57 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XANTENNA_genblk2\[12\].buf_p_rowonn_A VSS VDD core.pdc.rowon_out_n\[12\] VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA_cgen_dlycontrol3_in[4] VSS VDD net23 VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA_nmat_col_n[16] VSS VDD nmatrix_col_core_n_buffered\[16\] VDD VSS sky130_fd_sc_hd__diode_2
X_2010_ VSS VDD _0101_ _1085_ _1395_ _1390_ _1132_ VDD VSS sky130_fd_sc_hd__a31o_1
XFILLER_76_883 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XANTENNA__1600__B VSS VDD _1032_ VDD VSS sky130_fd_sc_hd__diode_2
X_2912_ VSS VDD _0802_ _0804_ _0803_ VDD VSS sky130_fd_sc_hd__nand2_1
X_2843_ VSS VDD _0732_ _0734_ _0738_ _0737_ VDD VSS sky130_fd_sc_hd__nand3_1
X_2774_ VSS VDD _0637_ _0670_ VDD VSS sky130_fd_sc_hd__inv_1
XANTENNA__1738__A1 VSS VDD _1259_ VDD VSS sky130_fd_sc_hd__diode_2
X_1725_ VSS VDD _1182_ _1253_ _1177_ VDD VSS sky130_fd_sc_hd__nand2_1
X_1656_ VSS VDD _1198_ _1186_ _1054_ _1197_ VDD VSS sky130_fd_sc_hd__mux2_1
X_1587_ VSS VDD _1122_ _1137_ _1136_ VDD VSS sky130_fd_sc_hd__nor2_2
XFILLER_85_113 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
X_2208_ VSS VDD _0241_ _0242_ core.osr.result_r\[0\] VDD VSS sky130_fd_sc_hd__nand2_1
XFILLER_67_883 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
X_3188_ VSS VDD clknet_2_1__leaf_clk_dig_dummy _0058_ net87 core.cnb.data_register_r\[8\]
+ VDD VSS sky130_fd_sc_hd__dfrtp_4
X_2139_ VSS VDD _0181_ _0183_ _0182_ VDD VSS sky130_fd_sc_hd__nand2_1
Xgenblk2\[3\].buf_p_rowonn VSS VDD pmatrix_rowon_core_n_buffered\[3\] core.pdc.rowon_out_n\[3\]
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
XFILLER_139_137 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XFILLER_118_53 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_118_97 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_134_52 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
XFILLER_89_485 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_134_85 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_94_45 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XANTENNA_input12_A VSS VDD config_1_in[4] VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1701__A VSS VDD net15 VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_43_93 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
X_2490_ VDD VSS net36 _0435_ VDD VSS sky130_fd_sc_hd__inv_2
X_1510_ VDD VSS _1068_ _1047_ VDD VSS sky130_fd_sc_hd__inv_2
X_1441_ VSS VDD core.osr.sample_count_r\[6\] _1003_ _1001_ _0999_ _1005_ _1004_ VDD
+ VSS sky130_fd_sc_hd__o221a_1
X_3111_ VSS VDD clknet_2_3__leaf_clk_dig_dummy _0011_ net90 core.cnb.shift_register_r\[9\]
+ VDD VSS sky130_fd_sc_hd__dfrtp_2
XFILLER_67_113 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
X_3042_ VSS VDD _0930_ _0910_ _0833_ _0726_ _0929_ VDD VSS sky130_fd_sc_hd__and4_1
XANTENNA__1656__A0 VSS VDD _1197_ VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_48_382 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XFILLER_51_525 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XFILLER_90_182 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XFILLER_23_19 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XANTENNA_pmat_sample_buf_n_A VSS VDD core.cnb.enable_loop_out VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__2442__A VSS VDD core.ndc.rowoff_out_n\[5\] VDD VSS sky130_fd_sc_hd__diode_2
X_2826_ VDD VSS _0719_ _0718_ _0720_ _0721_ VDD VSS sky130_fd_sc_hd__a21o_1
X_2757_ VDD VSS _0653_ core.cnb.shift_register_r\[10\] VDD VSS sky130_fd_sc_hd__inv_2
XFILLER_2_109 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
X_2688_ VSS VDD _0347_ _0568_ _0589_ _0348_ VDD VSS sky130_fd_sc_hd__nand3_1
X_1708_ VDD VSS _1240_ _1108_ VDD VSS sky130_fd_sc_hd__inv_2
X_1639_ VDD VSS _1183_ _1182_ VDD VSS sky130_fd_sc_hd__inv_2
XANTENNA_input4_A VSS VDD config_1_in[11] VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_86_411 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
XFILLER_86_444 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XFILLER_73_116 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XFILLER_104_77 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
Xfanout64 VSS VDD net66 net64 VDD VSS sky130_fd_sc_hd__clkbuf_2
Xfanout75 VDD VSS net75 net76 VDD VSS sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout86 VDD VSS net86 net87 VDD VSS sky130_fd_sc_hd__buf_2
XANTENNA__2071__B VSS VDD _1213_ VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_8_1 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_2_2__f_clk_dig_dummy_A VSS VDD clknet_0_clk_dig_dummy VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_64_127 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
X_1990_ VSS VDD _0086_ core.pdc.col_out_n\[6\] VDD VSS sky130_fd_sc_hd__clkbuf_2
XANTENNA__2262__A VSS VDD core.cnb.result_out\[6\] VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_118_118 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
X_2611_ VSS VDD _0288_ _0522_ _0517_ VDD VSS sky130_fd_sc_hd__nand2_1
X_2542_ VDD VSS core.cnb.average_sum_r\[2\] _0195_ _0198_ _0466_ VDD VSS sky130_fd_sc_hd__a21oi_1
XANTENNA_nmat_col[31] VSS VDD core.ndc.col_out\[31\] VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__3093__A VSS VDD _0758_ VDD VSS sky130_fd_sc_hd__diode_2
X_2473_ VSS VDD core.pdc.row_out_n\[4\] core.pdc.rowoff_out_n\[4\] core.pdc.rowon_out_n\[4\]
+ VDD VSS sky130_fd_sc_hd__nand2_1
X_1424_ VSS VDD _0987_ _0988_ _0983_ VDD VSS sky130_fd_sc_hd__nor2_2
XFILLER_83_414 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XANTENNA__1629__B1 VSS VDD _1118_ VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_55_127 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
X_3025_ VSS VDD _0912_ _0472_ _0913_ _0911_ VDD VSS sky130_fd_sc_hd__o21ai_1
XANTENNA__2172__A VSS VDD _0210_ VDD VSS sky130_fd_sc_hd__diode_2
X_2809_ VDD VSS _0704_ _0703_ VDD VSS sky130_fd_sc_hd__inv_2
XFILLER_117_151 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XFILLER_115_76 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
XFILLER_131_42 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_61_108 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XFILLER_54_160 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XFILLER_54_193 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XFILLER_91_57 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XFILLER_24_51 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XFILLER_40_72 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XFILLER_40_94 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
Xnmat_96 VSS VDD nmat_96/LO net96 VDD VSS sky130_fd_sc_hd__conb_1
XANTENNA__3190__RESET_B VSS VDD net81 VDD VSS sky130_fd_sc_hd__diode_2
Xcomp comp/clk ctop_pmatrix_analog ctop_nmatrix_analog decision_finish_comp_n comp/latch_qn
+ core.cnb.comparator_in VDD VSS adc_comp_latch
XFILLER_37_105 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
XFILLER_92_200 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
XFILLER_1_33 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
X_1973_ VDD VSS _1121_ _0068_ core.pdc.col_out\[4\] _0070_ _1296_ _0073_ VDD VSS sky130_fd_sc_hd__a221o_1
XFILLER_60_1 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XANTENNA_nmat_col[14] VSS VDD core.ndc.col_out\[14\] VDD VSS sky130_fd_sc_hd__diode_2
X_2525_ VSS VDD core.cnb.shift_register_r\[16\] _0454_ VDD VSS sky130_fd_sc_hd__clkbuf_2
X_2456_ VSS VDD core.ndc.rowon_out_n\[1\] core.ndc.rowoff_out_n\[1\] core.ndc.row_out_n\[1\]
+ VDD VSS sky130_fd_sc_hd__nand2_1
XFILLER_29_29 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
X_2387_ VDD VSS core.osr.next_sample_count_w\[1\] _0399_ VDD VSS sky130_fd_sc_hd__inv_2
XFILLER_83_211 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XANTENNA__2167__A VSS VDD _0210_ VDD VSS sky130_fd_sc_hd__diode_2
X_3008_ VSS VDD _0887_ _0897_ _0896_ VDD VSS sky130_fd_sc_hd__nand2_1
XFILLER_83_299 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XFILLER_10_64 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XFILLER_86_35 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XFILLER_19_73 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XANTENNA__3191__SET_B VSS VDD net82 VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_47_469 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_55_491 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_42_141 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_51_60 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XANTENNA__1792__A2 VSS VDD _1279_ VDD VSS sky130_fd_sc_hd__diode_2
X_2310_ VSS VDD _0331_ _0255_ _0334_ _0333_ VDD VSS sky130_fd_sc_hd__nand3_1
X_2241_ VSS VDD _0988_ _0271_ VDD VSS sky130_fd_sc_hd__clkbuf_2
XFILLER_111_113 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
X_2172_ VSS VDD _0213_ _0193_ _0194_ _0210_ VDD VSS sky130_fd_sc_hd__and3_1
XFILLER_46_491 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XANTENNA_cgen_dlycontrol4_in[2] VSS VDD net5 VDD VSS sky130_fd_sc_hd__diode_2
X_1956_ VDD VSS core.pdc.col_out_n\[2\] core.pdc.col_out\[2\] VDD VSS sky130_fd_sc_hd__inv_2
X_1887_ VDD VSS _1363_ _1029_ VDD VSS sky130_fd_sc_hd__inv_2
X_2508_ VSS VDD _0008_ _0445_ VDD VSS sky130_fd_sc_hd__clkbuf_1
XFILLER_102_135 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XANTENNA__1940__C1 VSS VDD _1085_ VDD VSS sky130_fd_sc_hd__diode_2
X_2439_ VSS VDD _1376_ core.ndc.rowon_out_n\[2\] _1385_ VDD VSS sky130_fd_sc_hd__nand2_1
XFILLER_56_255 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XFILLER_112_66 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_24_130 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XFILLER_24_141 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_21_63 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
XFILLER_21_85 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_47_277 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XFILLER_30_122 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_62_81 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
X_1810_ VSS VDD core.cnb.data_register_r\[9\] _1303_ VDD VSS sky130_fd_sc_hd__clkbuf_2
XFILLER_7_21 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
X_2790_ VSS VDD _0677_ _0685_ _0686_ VDD VSS sky130_fd_sc_hd__nand2b_1
X_1741_ VSS VDD _1033_ _1153_ _1263_ VDD VSS sky130_fd_sc_hd__nor2_1
XANTENNA__2270__A VSS VDD core.cnb.result_out\[7\] VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_7_65 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
X_1672_ VDD VSS _1207_ _1103_ _1206_ _1212_ VDD VSS sky130_fd_sc_hd__a21o_1
X_2224_ VDD VSS _0256_ core.cnb.result_out\[2\] core.osr.result_r\[2\] VDD VSS sky130_fd_sc_hd__or2_1
X_2155_ VSS VDD _0197_ _0198_ _0199_ core.cnb.average_counter_r\[3\] VDD VSS sky130_fd_sc_hd__o21ai_1
XFILLER_93_361 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
X_2086_ VDD VSS _0101_ _1173_ core.pdc.col_out\[22\] _0103_ _1096_ _0150_ VDD VSS
+ sky130_fd_sc_hd__a221o_1
XFILLER_42_29 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
X_2988_ VSS VDD _0874_ _1113_ _0878_ _0875_ VDD VSS sky130_fd_sc_hd__nand3_1
X_1939_ VDD VSS core.cnb.data_register_r\[3\] _1395_ VDD VSS sky130_fd_sc_hd__clkinv_2
XANTENNA__2180__A VSS VDD _0208_ VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_83_25 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XFILLER_83_69 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_16_85 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XANTENNA_genblk2\[15\].buf_p_rown_A VSS VDD core.pdc.row_out_n\[15\] VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA_cgen_dlycontrol3_in[3] VSS VDD net22 VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__3131__CLK VSS VDD clknet_2_3__leaf_clk_dig_dummy VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA_nmat_col_n[15] VSS VDD nmatrix_col_core_n_buffered\[15\] VDD VSS sky130_fd_sc_hd__diode_2
X_2911_ VSS VDD _0798_ _1200_ _0803_ _0800_ VDD VSS sky130_fd_sc_hd__nand3_1
X_2842_ VSS VDD _0736_ _0725_ _0737_ _0724_ VDD VSS sky130_fd_sc_hd__nand3_1
X_2773_ VSS VDD _0669_ _0635_ _0206_ _0668_ VDD VSS sky130_fd_sc_hd__and3_1
X_1724_ VSS VDD _1251_ _1252_ _1213_ VDD VSS sky130_fd_sc_hd__nand2_1
X_1655_ VDD VSS _1196_ _1197_ VDD VSS sky130_fd_sc_hd__clkinv_2
X_1586_ VDD VSS _1136_ _1135_ VDD VSS sky130_fd_sc_hd__inv_2
XFILLER_85_125 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
X_2207_ VSS VDD _0240_ _0241_ VDD VSS sky130_fd_sc_hd__clkbuf_4
X_3187_ VSS VDD clknet_2_1__leaf_clk_dig_dummy _0057_ net85 core.cnb.data_register_r\[7\]
+ VDD VSS sky130_fd_sc_hd__dfrtp_4
X_2138_ VDD VSS _0182_ core.cnb.average_counter_r\[1\] core.cnb.average_counter_r\[0\]
+ VDD VSS sky130_fd_sc_hd__or2_1
XANTENNA__1998__B VSS VDD _1155_ VDD VSS sky130_fd_sc_hd__diode_2
X_2069_ VSS VDD _1075_ _0115_ _0069_ _1126_ core.pdc.col_out_n\[18\] _0141_ VDD VSS
+ sky130_fd_sc_hd__o221a_1
XFILLER_118_65 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XANTENNA_fanout92_A VSS VDD net94 VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_89_497 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
XFILLER_94_13 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_134_97 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_94_57 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_94_79 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XFILLER_27_84 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XANTENNA__1968__A2 VSS VDD _1104_ VDD VSS sky130_fd_sc_hd__diode_2
X_1440_ VDD VSS _1004_ core.osr.sample_count_r\[8\] _0992_ VDD VSS sky130_fd_sc_hd__or2_1
X_3110_ VSS VDD clknet_2_3__leaf_clk_dig_dummy _0010_ net90 core.cnb.shift_register_r\[8\]
+ VDD VSS sky130_fd_sc_hd__dfrtp_1
XANTENNA_genblk1\[10\].buf_n_coln_A VSS VDD core.ndc.col_out_n\[10\] VDD VSS sky130_fd_sc_hd__diode_2
X_3041_ VSS VDD _0929_ _0818_ _0827_ _0745_ VDD VSS sky130_fd_sc_hd__and3_1
XANTENNA__1656__A1 VSS VDD _1186_ VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__2605__B1 VSS VDD _0395_ VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_90_1 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
X_2825_ VDD VSS _0720_ _0687_ VDD VSS sky130_fd_sc_hd__inv_2
X_2756_ VSS VDD _0651_ _0646_ _0652_ VDD VSS sky130_fd_sc_hd__nor2_1
X_2687_ VDD VSS _1008_ _0376_ _0524_ _0588_ VDD VSS sky130_fd_sc_hd__a21oi_1
X_1707_ VDD VSS _1238_ _1239_ VDD VSS sky130_fd_sc_hd__clkinv_2
X_1638_ VSS VDD _1061_ _1182_ _1053_ VDD VSS sky130_fd_sc_hd__nand2_1
X_1569_ VDD VSS _1121_ _1101_ VDD VSS sky130_fd_sc_hd__buf_2
XFILLER_46_309 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XFILLER_104_23 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XFILLER_104_34 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XFILLER_104_45 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
Xgenblk2\[12\].buf_p_rown VSS VDD pmatrix_row_core_n_buffered\[12\] core.pdc.row_out_n\[12\]
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
XANTENNA__2617__B VSS VDD _1002_ VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_120_88 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
Xfanout65 VSS VDD net65 net66 VDD VSS sky130_fd_sc_hd__clkbuf_1
Xfanout54 VDD VSS net54 net55 VDD VSS sky130_fd_sc_hd__buf_2
XANTENNA_cgen_dlycontrol2_in[4] VSS VDD net33 VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_13_42 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
Xfanout76 VSS VDD net82 net76 VDD VSS sky130_fd_sc_hd__clkbuf_2
Xfanout87 VDD VSS net87 net94 VDD VSS sky130_fd_sc_hd__buf_2
XFILLER_80_59 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XFILLER_13_86 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_89_24 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
XFILLER_89_57 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_89_261 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XFILLER_89_272 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XFILLER_49_158 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XFILLER_92_404 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XANTENNA__1712__A VSS VDD _1034_ VDD VSS sky130_fd_sc_hd__diode_2
X_2610_ VSS VDD _0521_ _0517_ core.osr.next_result_w\[3\] _0519_ _0520_ VDD VSS sky130_fd_sc_hd__o211a_1
X_2541_ VSS VDD _0462_ _0463_ _0465_ _0464_ VDD VSS sky130_fd_sc_hd__nand3_1
XFILLER_126_141 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
X_2472_ VSS VDD core.pdc.row_out_n\[3\] core.pdc.rowoff_out_n\[3\] core.pdc.rowon_out_n\[3\]
+ VDD VSS sky130_fd_sc_hd__nand2_1
X_1423_ VSS VDD _0987_ _0986_ _0985_ core.osr.sample_count_r\[0\] _0984_ VDD VSS sky130_fd_sc_hd__and4b_1
XANTENNA__1629__A1 VSS VDD _1085_ VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_55_139 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
X_3024_ VSS VDD _0835_ _0834_ _0912_ VDD VSS sky130_fd_sc_hd__nor2_1
XANTENNA__2437__B VSS VDD core.pdc.rowon_out_n\[0\] VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_70_109 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
X_2808_ VSS VDD _0674_ _0703_ _0702_ VDD VSS sky130_fd_sc_hd__nand2_1
X_2739_ VSS VDD core.cnb.shift_register_r\[6\] core.cnb.shift_register_r\[7\] _0635_
+ VDD VSS sky130_fd_sc_hd__nor2_1
XANTENNA__1565__A0 VSS VDD _1112_ VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_115_66 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
XFILLER_86_253 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_46_128 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XANTENNA__2347__B VSS VDD _0240_ VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_91_25 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_24_85 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_108_141 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_1_45 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XANTENNA__1588__S VSS VDD _1077_ VDD VSS sky130_fd_sc_hd__diode_2
X_1972_ VSS VDD _0065_ _0072_ _0073_ VDD VSS sky130_fd_sc_hd__nor2_1
Xgenblk2\[12\].buf_n_rowonn VSS VDD nmatrix_rowon_core_n_buffered\[12\] core.ndc.rowon_out_n\[12\]
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
XANTENNA_nmat_col[13] VSS VDD core.ndc.col_out\[13\] VDD VSS sky130_fd_sc_hd__diode_2
X_2524_ VSS VDD _0016_ _0453_ VDD VSS sky130_fd_sc_hd__clkbuf_1
X_2455_ VSS VDD core.pdc.rowon_out_n\[0\] _1362_ core.ndc.rowon_out_n\[14\] _1365_
+ VDD VSS sky130_fd_sc_hd__o21ai_2
X_2386_ VDD VSS _0398_ core.osr.is_last_sample _0396_ _0399_ VDD VSS sky130_fd_sc_hd__or3_1
XFILLER_28_106 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_45_29 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
X_3007_ VSS VDD _0895_ _0896_ VDD VSS sky130_fd_sc_hd__clkinvlp_2
XANTENNA__2183__A VSS VDD core.cnb.comparator_in VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_51_164 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XFILLER_101_57 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
XFILLER_124_7 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_105_144 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_19_85 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_42_153 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
X_2240_ VSS VDD _0270_ core.osr.next_result_w\[3\] VDD VSS sky130_fd_sc_hd__clkbuf_2
X_2171_ VSS VDD core.cnb.next_average_counter_w\[2\] _0212_ VDD VSS sky130_fd_sc_hd__clkbuf_1
XANTENNA_cgen_dlycontrol4_in[1] VSS VDD net4 VDD VSS sky130_fd_sc_hd__diode_2
Xgenblk1\[13\].buf_p_coln VSS VDD pmatrix_col_core_n_buffered\[13\] core.pdc.col_out_n\[13\]
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
X_1955_ VDD VSS _1398_ _1279_ core.pdc.col_out\[2\] _1406_ _1296_ _1408_ VDD VSS sky130_fd_sc_hd__a221o_1
X_1886_ VSS VDD _1038_ _1362_ VDD VSS sky130_fd_sc_hd__clkbuf_2
X_2507_ VSS VDD _0445_ core.cnb.shift_register_r\[7\] _0444_ core.cnb.shift_register_r\[6\]
+ VDD VSS sky130_fd_sc_hd__mux2_1
XANTENNA__1940__B1 VSS VDD _1079_ VDD VSS sky130_fd_sc_hd__diode_2
X_2438_ VDD VSS _1340_ _1027_ _1364_ core.ndc.rowon_out_n\[1\] VDD VSS sky130_fd_sc_hd__a21o_1
X_2369_ VDD VSS _0386_ _0381_ _0385_ VDD VSS sky130_fd_sc_hd__and2_1
XFILLER_112_23 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XFILLER_112_78 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
XFILLER_115_3 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_97_24 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XANTENNA_nmat_col_n[31] VSS VDD nmatrix_col_core_n_buffered\[31\] VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_97_57 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
XANTENNA_input35_A VSS VDD start_conversion_in VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__2088__A VSS VDD _1227_ VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1720__A VSS VDD core.ndc.col_out_n\[15\] VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_46_72 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XFILLER_30_134 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
XFILLER_62_71 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
X_1740_ VSS VDD _1157_ _1262_ _1152_ VDD VSS sky130_fd_sc_hd__nand2_1
XFILLER_7_77 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
X_1671_ VDD VSS _1210_ _1211_ VDD VSS sky130_fd_sc_hd__clkinv_2
X_2223_ VSS VDD _0988_ _0255_ VDD VSS sky130_fd_sc_hd__clkbuf_2
X_2154_ VDD VSS _0198_ _0181_ VDD VSS sky130_fd_sc_hd__inv_2
XFILLER_16_1 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XANTENNA__1630__A VSS VDD _1175_ VDD VSS sky130_fd_sc_hd__diode_2
X_2085_ VDD VSS _0150_ _0149_ VDD VSS sky130_fd_sc_hd__inv_2
Xgenblk2\[9\].buf_n_rowonn VSS VDD nmatrix_rowon_core_n_buffered\[9\] core.ndc.rowon_out_n\[9\]
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
X_2987_ VSS VDD _0876_ _0877_ _1058_ VDD VSS sky130_fd_sc_hd__nand2_1
XANTENNA__2461__A VSS VDD core.ndc.row_out_n\[7\] VDD VSS sky130_fd_sc_hd__diode_2
X_1938_ VDD VSS _1394_ _1388_ VDD VSS sky130_fd_sc_hd__buf_2
X_1869_ VSS VDD net14 _1308_ _1351_ VDD VSS sky130_fd_sc_hd__nor2_1
XFILLER_123_11 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_123_66 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
Xgenblk1\[10\].buf_n_coln VDD VSS core.ndc.col_out_n\[10\] nmatrix_col_core_n_buffered\[10\]
+ VDD VSS sky130_fd_sc_hd__buf_6
XANTENNA__1540__A VSS VDD _1095_ VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_16_97 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_52_281 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_32_52 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XANTENNA__2090__B VSS VDD _1235_ VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1715__A VSS VDD core.ndc.col_out_n\[14\] VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA_cgen_dlycontrol3_in[2] VSS VDD net21 VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA_nmat_col_n[14] VSS VDD nmatrix_col_core_n_buffered\[14\] VDD VSS sky130_fd_sc_hd__diode_2
X_2910_ VSS VDD _0801_ _0802_ _1055_ VDD VSS sky130_fd_sc_hd__nand2_1
X_2841_ VSS VDD _0646_ _0735_ _0736_ VDD VSS sky130_fd_sc_hd__nor2_1
X_2772_ VSS VDD core.cnb.shift_register_r\[2\] _0667_ _0668_ VDD VSS sky130_fd_sc_hd__nor2_1
X_1723_ VDD VSS _1251_ _1049_ VDD VSS sky130_fd_sc_hd__inv_2
X_1654_ VSS VDD _1195_ _1196_ _1051_ VDD VSS sky130_fd_sc_hd__nand2_1
X_1585_ VSS VDD _1135_ _1134_ _1050_ VDD VSS sky130_fd_sc_hd__nor2_4
X_2206_ VDD VSS _0240_ _0988_ VDD VSS sky130_fd_sc_hd__buf_2
XFILLER_54_502 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
X_3186_ VSS VDD clknet_2_1__leaf_clk_dig_dummy _0056_ net85 core.cnb.data_register_r\[6\]
+ VDD VSS sky130_fd_sc_hd__dfrtp_2
X_2137_ VSS VDD _0176_ _0180_ _0181_ core.cnb.sampled_avg_control_r\[0\] VDD VSS sky130_fd_sc_hd__nand3_1
XANTENNA__2456__A VSS VDD core.ndc.rowon_out_n\[1\] VDD VSS sky130_fd_sc_hd__diode_2
X_2068_ VSS VDD _0120_ _0141_ _1155_ VDD VSS sky130_fd_sc_hd__nand2_1
XFILLER_5_108 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XFILLER_118_77 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
XANTENNA__1535__A VSS VDD _1092_ VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_134_32 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XANTENNA_fanout85_A VSS VDD net87 VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_94_25 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XFILLER_94_69 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
Xgenblk2\[14\].buf_n_rown VSS VDD nmatrix_row_core_n_buffered\[14\] core.ndc.row_out_n\[14\]
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
XFILLER_27_63 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_27_41 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XFILLER_27_96 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XANTENNA__1968__A3 VSS VDD _1105_ VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__3184__RESET_B VSS VDD net87 VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_4_67 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
X_3040_ VSS VDD _0926_ _1055_ _0928_ _0927_ VDD VSS sky130_fd_sc_hd__nand3_1
XFILLER_51_505 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_83_1 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
X_2824_ VSS VDD _0714_ _0716_ _0719_ core.cnb.pswitch_out\[1\] VDD VSS sky130_fd_sc_hd__nand3_1
XFILLER_136_109 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
X_2755_ VSS VDD _0650_ _0651_ _0642_ VDD VSS sky130_fd_sc_hd__nand2_1
X_2686_ VSS VDD _0585_ _0044_ _0587_ VDD VSS sky130_fd_sc_hd__nand2_1
X_1706_ VSS VDD _1227_ _1166_ _1238_ VDD VSS sky130_fd_sc_hd__nor2_1
X_1637_ VSS VDD _1180_ _1181_ _1096_ VDD VSS sky130_fd_sc_hd__nand2_1
X_1568_ VDD VSS core.ndc.col_out\[3\] core.ndc.col_out_n\[3\] VDD VSS sky130_fd_sc_hd__inv_2
XFILLER_48_18 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XFILLER_48_29 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XFILLER_86_424 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_58_137 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
X_1499_ VSS VDD _1059_ _1058_ _1044_ VDD VSS sky130_fd_sc_hd__nand2_2
X_3169_ VSS VDD net66 core.osr.next_result_w\[9\] net76 core.osr.result_r\[9\] VDD
+ VSS sky130_fd_sc_hd__dfrtp_1
XFILLER_104_57 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_54_398 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
XFILLER_120_78 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
XANTENNA__2633__B VSS VDD core.osr.next_result_w\[2\] VDD VSS sky130_fd_sc_hd__diode_2
Xfanout55 VSS VDD core.cnb.is_sampling_w net55 VDD VSS sky130_fd_sc_hd__clkbuf_4
XFILLER_80_38 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XANTENNA_cgen_dlycontrol2_in[3] VSS VDD net32 VDD VSS sky130_fd_sc_hd__diode_2
Xfanout88 VSS VDD net92 net88 VDD VSS sky130_fd_sc_hd__clkbuf_2
Xfanout77 VDD VSS net77 net80 VDD VSS sky130_fd_sc_hd__buf_2
Xfanout66 VSS VDD net67 net66 VDD VSS sky130_fd_sc_hd__clkbuf_2
XANTENNA__3121__CLK VSS VDD clknet_2_2__leaf_clk_dig_dummy VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_129_76 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_13_98 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
XANTENNA__2532__A0 VSS VDD core.cnb.sampled_avg_control_r\[1\] VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_89_295 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XFILLER_38_62 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XANTENNA__1712__B VSS VDD _1243_ VDD VSS sky130_fd_sc_hd__diode_2
Xgenblk1\[18\].buf_p_coln VSS VDD pmatrix_col_core_n_buffered\[18\] core.pdc.col_out_n\[18\]
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
XFILLER_118_109 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
X_2540_ VSS VDD _0231_ _0177_ _0464_ _0186_ VDD VSS sky130_fd_sc_hd__o21ai_1
X_2471_ VSS VDD core.pdc.row_out_n\[2\] core.pdc.rowoff_out_n\[2\] core.pdc.rowon_out_n\[2\]
+ VDD VSS sky130_fd_sc_hd__nand2_1
X_1422_ VSS VDD core.osr.sample_count_r\[5\] core.osr.sample_count_r\[3\] core.osr.sample_count_r\[1\]
+ _0986_ VDD VSS sky130_fd_sc_hd__nor3_1
XANTENNA__1903__A VSS VDD _1342_ VDD VSS sky130_fd_sc_hd__diode_2
X_3023_ VSS VDD _0910_ _0911_ _0827_ VDD VSS sky130_fd_sc_hd__nand2_1
XFILLER_83_449 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_51_346 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XFILLER_60_891 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
X_2807_ VSS VDD _0702_ _0639_ _0701_ _0699_ VDD VSS sky130_fd_sc_hd__nand3b_1
X_2738_ VSS VDD _0633_ _0634_ core.cnb.shift_register_r\[9\] VDD VSS sky130_fd_sc_hd__nand2_1
XANTENNA__1565__A1 VSS VDD _1118_ VDD VSS sky130_fd_sc_hd__diode_2
X_2669_ VDD VSS _0565_ _0572_ _0042_ _0571_ VDD VSS sky130_fd_sc_hd__o21bai_1
Xgenblk1\[20\].buf_p_coln VSS VDD pmatrix_col_core_n_buffered\[20\] core.pdc.col_out_n\[20\]
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
XFILLER_86_265 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_46_107 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XANTENNA__2644__A VSS VDD core.osr.next_result_w\[8\] VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_91_37 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_24_64 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_24_97 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_40_85 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XFILLER_108_153 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XFILLER_49_72 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
XFILLER_1_57 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XANTENNA__3167__CLK VSS VDD net61 VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_65_71 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XANTENNA__2554__A VSS VDD core.cnb.pswitch_out\[1\] VDD VSS sky130_fd_sc_hd__diode_2
X_1971_ VDD VSS _0072_ _0071_ VDD VSS sky130_fd_sc_hd__inv_2
XANTENNA_nmat_col[12] VSS VDD core.ndc.col_out\[12\] VDD VSS sky130_fd_sc_hd__diode_2
X_2523_ VSS VDD _0453_ core.cnb.shift_register_r\[15\] _0219_ core.cnb.shift_register_r\[14\]
+ VDD VSS sky130_fd_sc_hd__mux2_1
XFILLER_46_1 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
X_2454_ VDD VSS core.ndc.rowon_out_n\[13\] _0431_ VDD VSS sky130_fd_sc_hd__inv_2
X_2385_ VDD VSS _0398_ _0397_ VDD VSS sky130_fd_sc_hd__inv_2
XANTENNA_cgen_dlycontrol1_in[4] VSS VDD net28 VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_28_118 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
Xinput1 VSS VDD net1 clk_vcm VDD VSS sky130_fd_sc_hd__clkbuf_1
XFILLER_56_449 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
Xgenblk1\[15\].buf_n_coln VDD VSS core.ndc.col_out_n\[15\] nmatrix_col_core_n_buffered\[15\]
+ VDD VSS sky130_fd_sc_hd__buf_6
X_3006_ VSS VDD _0893_ _0895_ _0894_ VDD VSS sky130_fd_sc_hd__nand2_1
XFILLER_10_77 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
XFILLER_19_53 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XFILLER_19_97 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_47_449 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_35_41 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_111_126 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
X_2170_ VSS VDD _0212_ _0197_ _0192_ _0210_ VDD VSS sky130_fd_sc_hd__and3_1
XANTENNA__1900__B VSS VDD _1022_ VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA_cgen_dlycontrol4_in[0] VSS VDD net3 VDD VSS sky130_fd_sc_hd__diode_2
X_1954_ VSS VDD _1272_ _1407_ _1408_ VDD VSS sky130_fd_sc_hd__nor2_1
X_1885_ VSS VDD core.pdc.row_out_n\[15\] _1361_ core.ndc.rowon_out_n\[0\] VDD VSS
+ sky130_fd_sc_hd__nand2_2
X_2506_ VSS VDD _0208_ _0444_ VDD VSS sky130_fd_sc_hd__clkbuf_2
XFILLER_88_316 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
X_2437_ VSS VDD _1341_ core.ndc.row_out_n\[15\] core.pdc.rowon_out_n\[0\] VDD VSS
+ sky130_fd_sc_hd__nand2_1
X_2368_ VDD VSS _0385_ _0384_ _0255_ VDD VSS sky130_fd_sc_hd__and2_1
X_2299_ VSS VDD _0309_ _0307_ _0323_ _0317_ VDD VSS sky130_fd_sc_hd__nand3_1
XFILLER_24_121 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XANTENNA__1538__A VSS VDD core.ndc.col_out_n\[1\] VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__2641__B VSS VDD core.osr.next_result_w\[3\] VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__2088__B VSS VDD _0072_ VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__3138__RESET_B VSS VDD net85 VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA_input28_A VSS VDD config_2_in[4] VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_46_95 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_7_34 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
X_1670_ VSS VDD _1033_ _1209_ _1210_ VDD VSS sky130_fd_sc_hd__nor2_1
X_2222_ VDD VSS core.osr.next_result_w\[1\] _0254_ VDD VSS sky130_fd_sc_hd__inv_2
X_2153_ VSS VDD _0191_ _0197_ _0184_ VDD VSS sky130_fd_sc_hd__nand2_1
XFILLER_53_216 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
X_2084_ VDD VSS _0149_ _1039_ _0113_ VDD VSS sky130_fd_sc_hd__or2_1
XFILLER_21_102 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XFILLER_21_113 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XFILLER_21_124 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
X_2986_ VSS VDD _0874_ _0876_ _0875_ VDD VSS sky130_fd_sc_hd__nand2_1
X_1937_ VDD VSS core.pdc.col_out_n\[0\] core.pdc.col_out\[0\] VDD VSS sky130_fd_sc_hd__inv_2
X_1868_ VSS VDD _1324_ _1333_ _1350_ VDD VSS sky130_fd_sc_hd__nor2_1
X_1799_ VDD VSS _1121_ _1083_ core.ndc.col_out\[30\] _1247_ _1296_ _1298_ VDD VSS
+ sky130_fd_sc_hd__a221o_1
XFILLER_107_57 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XFILLER_88_168 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XFILLER_123_23 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_84_396 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XFILLER_52_293 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XFILLER_12_146 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XFILLER_32_64 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XFILLER_79_113 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XANTENNA_cgen_dlycontrol3_in[1] VSS VDD net20 VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA_nmat_col_n[13] VSS VDD nmatrix_col_core_n_buffered\[13\] VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_94_149 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
XFILLER_87_190 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
XFILLER_90_300 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XFILLER_50_208 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
X_2840_ VSS VDD _0663_ _0735_ _0641_ VDD VSS sky130_fd_sc_hd__nand2_1
X_2771_ VDD VSS _0667_ core.cnb.shift_register_r\[3\] VDD VSS sky130_fd_sc_hd__inv_2
X_1722_ VSS VDD _1249_ _1250_ _1102_ VDD VSS sky130_fd_sc_hd__nand2_1
X_1653_ VSS VDD _1066_ _1195_ _1104_ VDD VSS sky130_fd_sc_hd__nand2_1
X_1584_ VSS VDD core.cnb.data_register_r\[6\] core.cnb.data_register_r\[5\] _1134_
+ VDD VSS sky130_fd_sc_hd__nor2_1
Xgenblk1\[25\].buf_p_coln VSS VDD pmatrix_col_core_n_buffered\[25\] core.pdc.col_out_n\[25\]
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
X_2205_ VDD VSS _0239_ core.cnb.result_out\[0\] VDD VSS sky130_fd_sc_hd__inv_2
X_3185_ VSS VDD clknet_2_1__leaf_clk_dig_dummy _0055_ net87 core.cnb.data_register_r\[5\]
+ VDD VSS sky130_fd_sc_hd__dfrtp_1
X_2136_ VDD VSS _0180_ core.cnb.sampled_avg_control_r\[2\] VDD VSS sky130_fd_sc_hd__inv_2
XANTENNA__2456__B VSS VDD core.ndc.row_out_n\[1\] VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_54_514 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_93_193 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
X_2067_ VDD VSS core.pdc.col_out\[17\] core.pdc.col_out_n\[17\] VDD VSS sky130_fd_sc_hd__clkinv_2
X_2969_ VDD VSS _0861_ _0805_ _0860_ VDD VSS sky130_fd_sc_hd__or2_1
XANTENNA__1551__A VSS VDD _1106_ VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_84_182 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XANTENNA__2382__A VSS VDD _0395_ VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA_pmat_rowoff_n[8] VSS VDD core.pdc.rowoff_out_n\[8\] VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_4_79 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XANTENNA__1461__A VSS VDD _1022_ VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__2557__A VSS VDD _0438_ VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_48_374 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XFILLER_90_141 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_51_517 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XFILLER_90_163 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XFILLER_90_174 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XANTENNA__2066__B1 VSS VDD _0089_ VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__2605__A2 VSS VDD _0995_ VDD VSS sky130_fd_sc_hd__diode_2
X_2823_ VSS VDD _0717_ _0718_ core.cnb.data_register_r\[1\] VDD VSS sky130_fd_sc_hd__nand2_1
XFILLER_76_1 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
X_2754_ VSS VDD core.cnb.shift_register_r\[8\] core.cnb.shift_register_r\[9\] _0650_
+ VDD VSS sky130_fd_sc_hd__nor2_1
X_1705_ VDD VSS core.ndc.col_out\[13\] core.ndc.col_out_n\[13\] VDD VSS sky130_fd_sc_hd__inv_2
X_2685_ VDD VSS _0587_ _0586_ VDD VSS sky130_fd_sc_hd__inv_2
XANTENNA__1636__A VSS VDD _1129_ VDD VSS sky130_fd_sc_hd__diode_2
X_1636_ VDD VSS _1180_ _1129_ VDD VSS sky130_fd_sc_hd__inv_2
X_1567_ VSS VDD _1075_ _1109_ _1108_ _1064_ core.ndc.col_out_n\[3\] _1120_ VDD VSS
+ sky130_fd_sc_hd__o221a_2
X_1498_ VSS VDD core.cnb.data_register_r\[6\] _1058_ VDD VSS sky130_fd_sc_hd__clkbuf_2
XFILLER_86_436 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
X_3168_ VSS VDD net66 core.osr.next_result_w\[8\] net76 core.osr.result_r\[8\] VDD
+ VSS sky130_fd_sc_hd__dfrtp_1
XFILLER_104_69 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XFILLER_64_29 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
X_2119_ VSS VDD core.pdc.col_out_n\[29\] _0169_ VDD VSS sky130_fd_sc_hd__clkbuf_1
X_3099_ VSS VDD _0981_ core.osr.osr_mode_r\[2\] _0241_ net13 VDD VSS sky130_fd_sc_hd__mux2_1
Xfanout56 VDD VSS net56 net57 VDD VSS sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_cgen_dlycontrol2_in[2] VSS VDD net31 VDD VSS sky130_fd_sc_hd__diode_2
Xfanout89 VDD VSS net89 net92 VDD VSS sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout78 VDD VSS net78 net80 VDD VSS sky130_fd_sc_hd__buf_2
Xfanout67 VSS VDD net37 net67 VDD VSS sky130_fd_sc_hd__clkbuf_2
XFILLER_129_88 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XANTENNA__1546__A VSS VDD _1101_ VDD VSS sky130_fd_sc_hd__diode_2
Xgenblk1\[22\].buf_n_coln VDD VSS core.ndc.col_out_n\[22\] nmatrix_col_core_n_buffered\[22\]
+ VDD VSS sky130_fd_sc_hd__buf_6
XFILLER_49_116 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XFILLER_38_85 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_92_428 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XANTENNA_input10_A VSS VDD config_1_in[2] VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_70_61 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XANTENNA__1456__A VSS VDD _0983_ VDD VSS sky130_fd_sc_hd__diode_2
X_2470_ VSS VDD core.pdc.row_out_n\[1\] core.pdc.rowoff_out_n\[1\] core.pdc.rowon_out_n\[1\]
+ VDD VSS sky130_fd_sc_hd__nand2_1
X_1421_ VDD VSS _0985_ core.osr.sample_count_r\[2\] VDD VSS sky130_fd_sc_hd__inv_2
X_3022_ VDD VSS _0910_ _0809_ VDD VSS sky130_fd_sc_hd__inv_2
XFILLER_63_141 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
X_2806_ VSS VDD _0700_ _0659_ _0701_ VDD VSS sky130_fd_sc_hd__nor2_1
X_2737_ VDD VSS _0633_ core.cnb.shift_register_r\[8\] VDD VSS sky130_fd_sc_hd__inv_2
X_2668_ VDD VSS _0394_ core.osr.next_result_w\[4\] _0542_ _0572_ net52 VDD VSS sky130_fd_sc_hd__a22o_1
X_1619_ VSS VDD _1165_ _1164_ _1041_ _1161_ VDD VSS sky130_fd_sc_hd__mux2_1
XFILLER_59_29 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
X_2599_ VDD VSS _0439_ _0335_ _0512_ _0032_ VDD VSS sky130_fd_sc_hd__a21oi_1
XFILLER_115_57 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
XANTENNA_input2_A VSS VDD config_1_in[0] VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_75_17 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_86_277 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XANTENNA__2644__B VSS VDD _1002_ VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_91_16 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
XFILLER_24_76 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XFILLER_24_43 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XFILLER_138_3 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_40_64 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XFILLER_123_113 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_1_69 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XFILLER_45_141 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
X_1970_ VSS VDD _0071_ _1115_ _1052_ _1389_ _1045_ VDD VSS sky130_fd_sc_hd__a31o_1
X_2522_ VSS VDD _0015_ _0452_ VDD VSS sky130_fd_sc_hd__clkbuf_1
X_2453_ VSS VDD _1380_ _0431_ _1306_ VDD VSS sky130_fd_sc_hd__nand2_1
XANTENNA_cgen_sample_p_in VSS VDD net55 VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_39_1 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
X_2384_ VSS VDD core.osr.sample_count_r\[0\] _0397_ core.osr.sample_count_r\[1\] VDD
+ VSS sky130_fd_sc_hd__nand2_1
XANTENNA_cgen_dlycontrol1_in[3] VSS VDD net27 VDD VSS sky130_fd_sc_hd__diode_2
Xinput2 VSS VDD net2 config_1_in[0] VDD VSS sky130_fd_sc_hd__clkbuf_1
XANTENNA__3111__CLK VSS VDD clknet_2_3__leaf_clk_dig_dummy VDD VSS sky130_fd_sc_hd__diode_2
X_3005_ VSS VDD _0890_ _1051_ _0894_ _0891_ VDD VSS sky130_fd_sc_hd__nand3_1
XFILLER_36_141 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_51_144 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XANTENNA__2480__A VSS VDD core.pdc.rowon_out_n\[13\] VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_105_113 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_19_21 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XANTENNA_fanout60_A VSS VDD net61 VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_47_439 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XFILLER_42_122 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_35_53 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XANTENNA__1718__B VSS VDD _1093_ VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1734__A VSS VDD core.ndc.col_out_n\[17\] VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__3134__CLK VSS VDD clknet_2_0__leaf_clk_dig_dummy VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__2549__B VSS VDD _0438_ VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_93_501 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XFILLER_18_152 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
X_1953_ VSS VDD _1123_ _1403_ _1068_ _1407_ VDD VSS sky130_fd_sc_hd__o21a_1
XANTENNA__2504__S VSS VDD _0220_ VDD VSS sky130_fd_sc_hd__diode_2
X_1884_ VSS VDD _1358_ _1361_ _1026_ VDD VSS sky130_fd_sc_hd__nand2_1
XANTENNA__1909__A VSS VDD _1340_ VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1628__B VSS VDD _1173_ VDD VSS sky130_fd_sc_hd__diode_2
X_2505_ VSS VDD _0007_ _0443_ VDD VSS sky130_fd_sc_hd__clkbuf_1
X_2436_ VDD VSS _1331_ _1320_ _1307_ core.ndc.row_out_n\[14\] VDD VSS sky130_fd_sc_hd__a21oi_1
XANTENNA__1644__A VSS VDD _1032_ VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1940__A2 VSS VDD _1395_ VDD VSS sky130_fd_sc_hd__diode_2
X_2367_ VSS VDD _0377_ _0384_ _0383_ VDD VSS sky130_fd_sc_hd__nand2_1
X_2298_ VSS VDD core.osr.next_result_w\[9\] _0321_ _0322_ VDD VSS sky130_fd_sc_hd__nand2_2
XFILLER_56_225 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XANTENNA__2475__A VSS VDD core.pdc.row_out_n\[7\] VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_72_29 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_21_11 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XFILLER_21_77 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XFILLER_47_225 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XFILLER_47_247 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_47_269 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XFILLER_46_85 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
XANTENNA__1729__A VSS VDD _1074_ VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_7_46 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XANTENNA_pmat_en_bit_n[2] VSS VDD core.cnb.data_register_r\[2\] VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_30_5 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
X_2221_ VSS VDD _0253_ core.cnb.result_out\[1\] _0254_ _0240_ VDD VSS sky130_fd_sc_hd__o21ai_2
XFILLER_87_81 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
X_2152_ VSS VDD _0194_ _0196_ _0195_ VDD VSS sky130_fd_sc_hd__nand2_1
X_2083_ VDD VSS core.pdc.col_out_n\[21\] core.pdc.col_out\[21\] VDD VSS sky130_fd_sc_hd__clkinv_2
XANTENNA__2635__B1 VSS VDD _0394_ VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__2742__B VSS VDD _0637_ VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_21_136 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
X_2985_ VSS VDD _0799_ _0875_ _0873_ VDD VSS sky130_fd_sc_hd__nand2_1
X_1936_ VDD VSS _1284_ _1391_ _1393_ core.pdc.col_out\[0\] VDD VSS sky130_fd_sc_hd__a21o_1
X_1867_ VSS VDD _1349_ _1325_ core.ndc.row_bottotop_n\[5\] _1027_ core.pdc.row_out_n\[10\]
+ VDD VSS sky130_fd_sc_hd__o22a_2
X_1798_ VSS VDD _1272_ _1109_ _1298_ VDD VSS sky130_fd_sc_hd__nor2_1
Xgenblk1\[27\].buf_n_coln VSS VDD nmatrix_col_core_n_buffered\[27\] core.ndc.col_out_n\[27\]
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
XFILLER_88_158 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
X_2419_ VDD VSS _0424_ core.osr.next_sample_count_w\[8\] VDD VSS sky130_fd_sc_hd__clkinv_2
XFILLER_123_35 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XFILLER_84_320 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
XFILLER_83_17 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XFILLER_84_386 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XFILLER_16_77 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
XFILLER_120_3 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XANTENNA_cgen_dlycontrol3_in[0] VSS VDD net19 VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_79_125 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XANTENNA_nmat_col_n[12] VSS VDD nmatrix_col_core_n_buffered\[12\] VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_94_117 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XANTENNA__1731__B VSS VDD _1188_ VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__2562__B VSS VDD _0482_ VDD VSS sky130_fd_sc_hd__diode_2
X_2770_ VSS VDD _0656_ _0665_ _0666_ VDD VSS sky130_fd_sc_hd__nor2_1
X_1721_ VDD VSS _1249_ _1246_ VDD VSS sky130_fd_sc_hd__inv_2
X_1652_ VDD VSS _1194_ _1193_ VDD VSS sky130_fd_sc_hd__inv_2
X_1583_ VDD VSS _1133_ _1132_ VDD VSS sky130_fd_sc_hd__inv_2
X_2204_ VSS VDD core.cnb.next_average_sum_w\[4\] _0238_ VDD VSS sky130_fd_sc_hd__clkbuf_1
X_3184_ VSS VDD clknet_2_1__leaf_clk_dig_dummy _0054_ net87 core.cnb.data_register_r\[4\]
+ VDD VSS sky130_fd_sc_hd__dfrtp_2
X_2135_ VDD VSS core.cnb.average_counter_r\[3\] _0178_ core.cnb.average_counter_r\[4\]
+ _0179_ VDD VSS sky130_fd_sc_hd__a21o_1
X_2066_ VDD VSS _0139_ _1173_ core.pdc.col_out\[17\] _0089_ _1296_ _0140_ VDD VSS
+ sky130_fd_sc_hd__a221o_1
XANTENNA__1831__A1 VSS VDD core.pdc.rowoff_out_n\[8\] VDD VSS sky130_fd_sc_hd__diode_2
X_2968_ VSS VDD _0841_ _0852_ _0860_ _0859_ VDD VSS sky130_fd_sc_hd__nand3_1
X_1919_ VSS VDD _1026_ _1029_ _1382_ VDD VSS sky130_fd_sc_hd__nor2_1
XFILLER_118_13 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
X_2899_ VDD VSS _0792_ _0782_ _0775_ VDD VSS sky130_fd_sc_hd__and2_1
XFILLER_134_23 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
Xgenblk2\[5\].buf_n_rowonn VSS VDD nmatrix_rowon_core_n_buffered\[5\] core.ndc.rowon_bottotop_n\[5\]
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
XANTENNA__1551__B VSS VDD _1092_ VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_27_21 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
Xgenblk2\[0\].buf_p_rown VSS VDD pmatrix_row_core_n_buffered\[0\] core.pdc.row_out_n\[0\]
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
XFILLER_43_31 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XFILLER_138_141 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XANTENNA__2602__S VSS VDD _0438_ VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_67_106 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
XFILLER_90_197 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XANTENNA__2066__B2 VSS VDD _1296_ VDD VSS sky130_fd_sc_hd__diode_2
X_2822_ VSS VDD _0714_ _0717_ _0716_ VDD VSS sky130_fd_sc_hd__nand2_1
X_2753_ VDD VSS _0639_ _0649_ VDD VSS sky130_fd_sc_hd__buf_6
X_1704_ VSS VDD _1237_ core.ndc.col_out_n\[13\] VDD VSS sky130_fd_sc_hd__clkbuf_2
XANTENNA__1577__B1 VSS VDD _1082_ VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_69_1 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
X_2684_ VDD VSS net39 core.osr.next_result_w\[6\] _0562_ _0586_ _0393_ VDD VSS sky130_fd_sc_hd__a22o_1
X_1635_ VDD VSS core.ndc.col_out\[7\] core.ndc.col_out_n\[7\] VDD VSS sky130_fd_sc_hd__inv_2
X_1566_ VDD VSS _1120_ _1110_ _1119_ VDD VSS sky130_fd_sc_hd__or2_1
XANTENNA__1652__A VSS VDD _1193_ VDD VSS sky130_fd_sc_hd__diode_2
X_1497_ VSS VDD _1056_ _1057_ VDD VSS sky130_fd_sc_hd__clkbuf_4
X_3167_ VSS VDD net61 core.osr.next_result_w\[7\] net73 core.osr.result_r\[7\] VDD
+ VSS sky130_fd_sc_hd__dfrtp_1
X_3098_ VSS VDD _0063_ _0980_ VDD VSS sky130_fd_sc_hd__clkbuf_1
X_2118_ VSS VDD _0169_ _0168_ _0167_ _0166_ VDD VSS sky130_fd_sc_hd__and3_1
XFILLER_120_14 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
X_2049_ VSS VDD core.pdc.col_out_n\[14\] _0129_ VDD VSS sky130_fd_sc_hd__clkbuf_1
XFILLER_120_36 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XANTENNA_cgen_dlycontrol2_in[1] VSS VDD net30 VDD VSS sky130_fd_sc_hd__diode_2
Xfanout57 VDD VSS net57 net58 VDD VSS sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout68 VSS VDD net69 net68 VDD VSS sky130_fd_sc_hd__clkbuf_2
Xfanout79 VDD VSS net79 net80 VDD VSS sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__1562__A VSS VDD _1113_ VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__2377__B VSS VDD _0240_ VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_38_97 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
XFILLER_54_52 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XANTENNA__2824__C VSS VDD core.cnb.pswitch_out\[1\] VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_54_85 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XANTENNA__2599__A2 VSS VDD _0439_ VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_126_111 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XANTENNA__1737__A VSS VDD _1074_ VDD VSS sky130_fd_sc_hd__diode_2
X_1420_ VDD VSS core.osr.sample_count_r\[6\] core.osr.sample_count_r\[8\] core.osr.sample_count_r\[7\]
+ core.osr.sample_count_r\[4\] _0984_ VDD VSS sky130_fd_sc_hd__or4_1
XANTENNA__1472__A VSS VDD net15 VDD VSS sky130_fd_sc_hd__diode_2
X_3021_ VSS VDD _0860_ _0909_ _0908_ VDD VSS sky130_fd_sc_hd__nand2_1
X_2805_ VSS VDD _0645_ _0700_ _0642_ VDD VSS sky130_fd_sc_hd__nand2_1
XANTENNA__1647__A VSS VDD _1190_ VDD VSS sky130_fd_sc_hd__diode_2
X_2736_ VSS VDD _0630_ _0049_ _0632_ VDD VSS sky130_fd_sc_hd__nand2_1
X_2667_ VSS VDD _0566_ _0570_ _0571_ VDD VSS sky130_fd_sc_hd__nor2_1
X_1618_ VDD VSS _1164_ _1163_ VDD VSS sky130_fd_sc_hd__inv_2
XANTENNA__1970__B1 VSS VDD _1045_ VDD VSS sky130_fd_sc_hd__diode_2
X_2598_ VSS VDD _1022_ _0509_ _0501_ _1328_ _0512_ _0461_ VDD VSS sky130_fd_sc_hd__o221a_1
XANTENNA__3190__CLK VSS VDD clknet_2_1__leaf_clk_dig_dummy VDD VSS sky130_fd_sc_hd__diode_2
X_1549_ VSS VDD _1105_ _1056_ _1050_ VDD VSS sky130_fd_sc_hd__nor2_4
XFILLER_75_29 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_131_57 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_54_197 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XANTENNA__1557__A VSS VDD _1085_ VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_123_125 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XANTENNA_genblk2\[8\].buf_p_rowonn_A VSS VDD core.pdc.rowon_out_n\[8\] VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_92_215 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
XFILLER_92_248 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XANTENNA__3012__A VSS VDD _0799_ VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA_genblk2\[9\].buf_n_rowonn_A VSS VDD core.ndc.rowon_out_n\[9\] VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA_nmat_col[10] VSS VDD core.ndc.col_out\[10\] VDD VSS sky130_fd_sc_hd__diode_2
X_2521_ VSS VDD _0452_ core.cnb.shift_register_r\[14\] _0219_ core.cnb.shift_register_r\[13\]
+ VDD VSS sky130_fd_sc_hd__mux2_1
X_2452_ VDD VSS core.ndc.rowon_out_n\[12\] _0430_ VDD VSS sky130_fd_sc_hd__inv_2
X_2383_ VSS VDD core.osr.sample_count_r\[0\] core.osr.sample_count_r\[1\] _0396_ VDD
+ VSS sky130_fd_sc_hd__nor2_1
XANTENNA_cgen_dlycontrol1_in[2] VSS VDD net26 VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_83_204 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
Xinput3 VSS VDD config_1_in[10] net3 VDD VSS sky130_fd_sc_hd__clkbuf_2
XANTENNA__1930__A VSS VDD core.pdc.rowon_out_n\[0\] VDD VSS sky130_fd_sc_hd__diode_2
X_3004_ VSS VDD _0892_ _0893_ _1117_ VDD VSS sky130_fd_sc_hd__nand2_1
XFILLER_83_248 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XFILLER_91_281 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_101_27 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XANTENNA__2480__B VSS VDD core.pdc.row_out_n\[13\] VDD VSS sky130_fd_sc_hd__diode_2
X_2719_ VSS VDD _0517_ _0380_ _0617_ VDD VSS sky130_fd_sc_hd__nor2_1
XFILLER_126_13 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_105_125 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_120_106 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
XFILLER_87_521 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
XFILLER_19_109 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XFILLER_19_33 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_42_134 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
XFILLER_92_60 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XANTENNA__2581__A VSS VDD _0439_ VDD VSS sky130_fd_sc_hd__diode_2
X_1952_ VDD VSS _1406_ _1405_ VDD VSS sky130_fd_sc_hd__inv_2
X_1883_ VSS VDD _1360_ core.pdc.row_out_n\[14\] _1359_ VDD VSS sky130_fd_sc_hd__nor2_2
XANTENNA__1909__B VSS VDD core.pdc.rowoff_out_n\[8\] VDD VSS sky130_fd_sc_hd__diode_2
X_2504_ VSS VDD _0443_ core.cnb.shift_register_r\[6\] _0220_ core.cnb.shift_register_r\[5\]
+ VDD VSS sky130_fd_sc_hd__mux2_1
X_2435_ VSS VDD core.ndc.row_bottotop_n\[10\] _1318_ core.pdc.rowoff_out_n\[8\] _1369_
+ core.ndc.row_out_n\[13\] VDD VSS sky130_fd_sc_hd__o22a_1
X_2366_ VDD VSS _0383_ _0382_ VDD VSS sky130_fd_sc_hd__inv_2
X_2297_ VSS VDD _0252_ _0322_ core.cnb.result_out\[9\] VDD VSS sky130_fd_sc_hd__nand2_1
XFILLER_56_237 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
Xgenblk2\[5\].buf_p_rown VSS VDD pmatrix_row_core_n_buffered\[5\] core.ndc.row_bottotop_n\[10\]
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
XANTENNA__1835__A VSS VDD net14 VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_47_204 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_46_20 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XFILLER_47_259 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
XFILLER_15_101 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XFILLER_46_53 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
Xgenblk2\[13\].buf_p_rowonn VSS VDD pmatrix_rowon_core_n_buffered\[13\] core.pdc.rowon_out_n\[13\]
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
XANTENNA__1729__B VSS VDD _1243_ VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__3101__CLK VSS VDD clknet_2_0__leaf_clk_dig_dummy VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA_pmat_en_bit_n[1] VSS VDD core.cnb.data_register_r\[1\] VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_97_104 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
X_2220_ VDD VSS _0250_ _0249_ _0252_ _0253_ VDD VSS sky130_fd_sc_hd__a21o_1
Xpmat_sample_buf VSS VDD pmat_sample_switch_buffered net55 VDD VSS sky130_fd_sc_hd__clkbuf_1
XFILLER_23_5 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
X_2151_ VDD VSS _0195_ _0177_ _0186_ VDD VSS sky130_fd_sc_hd__and2_1
XFILLER_93_321 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
X_2082_ VSS VDD _1284_ _0106_ _0148_ core.pdc.col_out_n\[21\] VDD VSS sky130_fd_sc_hd__o21a_1
XFILLER_93_376 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XFILLER_93_387 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XANTENNA__2635__A1 VSS VDD core.cnb.result_out\[0\] VDD VSS sky130_fd_sc_hd__diode_2
X_2984_ VDD VSS _0874_ _0873_ _0784_ VDD VSS sky130_fd_sc_hd__or2_1
Xgenblk1\[0\].buf_p_coln VSS VDD pmatrix_col_core_n_buffered\[0\] core.pdc.col_out_n\[0\]
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
X_1935_ VDD VSS _1393_ _1392_ VDD VSS sky130_fd_sc_hd__inv_2
X_1866_ VDD VSS _1349_ _1329_ VDD VSS sky130_fd_sc_hd__inv_2
X_1797_ VDD VSS core.ndc.col_out_n\[29\] core.ndc.col_out\[29\] VDD VSS sky130_fd_sc_hd__inv_2
X_2418_ VDD VSS _0423_ core.osr.is_last_sample _0422_ _0424_ VDD VSS sky130_fd_sc_hd__or3_1
XANTENNA__2486__A VSS VDD sample_nmatrix_cgen VDD VSS sky130_fd_sc_hd__diode_2
X_2349_ VDD VSS _0368_ core.osr.result_r\[15\] VDD VSS sky130_fd_sc_hd__inv_2
XFILLER_84_332 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XANTENNA__3124__CLK VSS VDD clknet_2_2__leaf_clk_dig_dummy VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_32_99 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_79_137 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XANTENNA__2396__A VSS VDD _0394_ VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_94_129 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XANTENNA_input33_A VSS VDD config_2_in[9] VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_57_85 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
Xgenblk2\[2\].buf_n_rown VSS VDD nmatrix_row_core_n_buffered\[2\] core.ndc.row_out_n\[2\]
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
XANTENNA__3004__B VSS VDD _1117_ VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_90_368 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
X_1720_ VDD VSS core.ndc.col_out\[15\] core.ndc.col_out_n\[15\] VDD VSS sky130_fd_sc_hd__inv_2
X_1651_ VSS VDD _1193_ _1192_ _1191_ _1077_ VDD VSS sky130_fd_sc_hd__o21a_2
XANTENNA__1475__A VSS VDD _1034_ VDD VSS sky130_fd_sc_hd__diode_2
X_1582_ VDD VSS _1113_ _1079_ _1051_ _1132_ VDD VSS sky130_fd_sc_hd__a21o_1
X_2203_ VSS VDD _0238_ _0237_ _0236_ _0209_ VDD VSS sky130_fd_sc_hd__and3_1
X_3183_ VSS VDD clknet_2_1__leaf_clk_dig_dummy _0053_ net86 core.cnb.data_register_r\[3\]
+ VDD VSS sky130_fd_sc_hd__dfrtp_2
X_2134_ VSS VDD _0177_ _0178_ core.cnb.sampled_avg_control_r\[0\] VDD VSS sky130_fd_sc_hd__nand2_1
XFILLER_93_173 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
X_2065_ VSS VDD _0065_ _1405_ _0140_ VDD VSS sky130_fd_sc_hd__nor2_1
XFILLER_139_109 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
X_2967_ VSS VDD _0857_ _1076_ _0859_ _0858_ VDD VSS sky130_fd_sc_hd__nand3_1
X_1918_ VSS VDD core.pdc.rowon_out_n\[10\] _1381_ VDD VSS sky130_fd_sc_hd__clkbuf_1
X_2898_ VSS VDD _0789_ _0791_ _0790_ VDD VSS sky130_fd_sc_hd__nand2_1
X_1849_ VDD VSS _1336_ _1026_ VDD VSS sky130_fd_sc_hd__buf_2
XFILLER_118_25 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XFILLER_76_107 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XFILLER_138_153 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XANTENNA__2066__A2 VSS VDD _1173_ VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_72_891 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
X_2821_ VSS VDD _0471_ _0686_ _0716_ _0715_ VDD VSS sky130_fd_sc_hd__nand3_1
X_2752_ VSS VDD _0648_ _0640_ _0647_ _0634_ VDD VSS sky130_fd_sc_hd__nand3b_1
X_1703_ VSS VDD _1237_ _1236_ _1234_ _1233_ VDD VSS sky130_fd_sc_hd__and3_1
X_2683_ VDD VSS _0581_ _0584_ _0585_ _0583_ VDD VSS sky130_fd_sc_hd__o21bai_1
X_1634_ VSS VDD _1179_ core.ndc.col_out_n\[7\] VDD VSS sky130_fd_sc_hd__clkbuf_2
X_1565_ VSS VDD _1119_ _1118_ _1077_ _1112_ VDD VSS sky130_fd_sc_hd__mux2_1
XANTENNA__1933__A VSS VDD _1057_ VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_86_405 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XFILLER_58_107 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XFILLER_58_129 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
X_1496_ VSS VDD _1055_ _1056_ core.cnb.data_register_r\[3\] VDD VSS sky130_fd_sc_hd__nand2_1
X_3166_ VSS VDD net60 core.osr.next_result_w\[6\] net72 core.osr.result_r\[6\] VDD
+ VSS sky130_fd_sc_hd__dfrtp_1
X_3097_ VSS VDD _0980_ core.osr.osr_mode_r\[1\] _0241_ net12 VDD VSS sky130_fd_sc_hd__mux2_1
X_2117_ VSS VDD _0077_ _0168_ _1235_ VDD VSS sky130_fd_sc_hd__nand2_1
X_2048_ VSS VDD _0129_ _0128_ _0127_ _0123_ VDD VSS sky130_fd_sc_hd__and3_1
XFILLER_120_48 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XANTENNA_cgen_dlycontrol2_in[0] VSS VDD net29 VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_63_891 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
Xfanout58 VSS VDD net67 net58 VDD VSS sky130_fd_sc_hd__clkbuf_2
Xfanout69 VSS VDD net70 net69 VDD VSS sky130_fd_sc_hd__clkbuf_2
XFILLER_13_13 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_129_13 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_129_57 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XFILLER_38_21 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
XFILLER_54_64 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_126_101 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XFILLER_70_85 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_79_94 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XANTENNA__1472__B VSS VDD core.cnb.data_register_r\[8\] VDD VSS sky130_fd_sc_hd__diode_2
X_3020_ VDD VSS _0908_ _0906_ _0907_ VDD VSS sky130_fd_sc_hd__and2_1
XFILLER_95_93 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XFILLER_60_883 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
X_2804_ VSS VDD _0698_ _0699_ core.cnb.shift_register_r\[12\] VDD VSS sky130_fd_sc_hd__nand2_1
XFILLER_117_123 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
X_2735_ VDD VSS _0632_ _0631_ VDD VSS sky130_fd_sc_hd__inv_2
X_2666_ VSS VDD _0567_ _0570_ _0569_ VDD VSS sky130_fd_sc_hd__nand2_1
XANTENNA_clkbuf_2_1__f_clk_dig_dummy_A VSS VDD clknet_0_clk_dig_dummy VDD VSS sky130_fd_sc_hd__diode_2
X_1617_ VDD VSS _1163_ _1050_ _1162_ VDD VSS sky130_fd_sc_hd__or2_2
X_2597_ VSS VDD _0031_ _0511_ VDD VSS sky130_fd_sc_hd__clkbuf_1
XFILLER_115_15 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
X_1548_ VSS VDD _1058_ _1104_ VDD VSS sky130_fd_sc_hd__clkbuf_4
X_1479_ VDD VSS _1039_ net15 VDD VSS sky130_fd_sc_hd__inv_2
XFILLER_86_235 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
X_3149_ VSS VDD net59 _0039_ net71 net49 VDD VSS sky130_fd_sc_hd__dfrtp_1
XFILLER_54_121 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XFILLER_131_69 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_50_360 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XANTENNA__1573__A VSS VDD _1095_ VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_85_290 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
Xgenblk1\[5\].buf_p_coln VSS VDD pmatrix_col_core_n_buffered\[5\] core.pdc.col_out_n\[5\]
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
X_2520_ VSS VDD _0014_ _0451_ VDD VSS sky130_fd_sc_hd__clkbuf_1
X_2451_ VDD VSS _1328_ _1369_ _1365_ _0430_ _1331_ VDD VSS sky130_fd_sc_hd__a22o_1
X_2382_ VSS VDD _0395_ core.osr.next_sample_count_w\[0\] core.osr.sample_count_r\[0\]
+ VDD VSS sky130_fd_sc_hd__nand2_1
XANTENNA_cgen_dlycontrol1_in[1] VSS VDD net25 VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_56_408 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
Xinput4 VSS VDD config_1_in[11] net4 VDD VSS sky130_fd_sc_hd__clkbuf_2
XANTENNA__1930__B VSS VDD _1040_ VDD VSS sky130_fd_sc_hd__diode_2
X_3003_ VSS VDD _0890_ _0892_ _0891_ VDD VSS sky130_fd_sc_hd__nand2_1
XFILLER_51_124 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XFILLER_91_293 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
X_2718_ VDD VSS _0616_ _0615_ VDD VSS sky130_fd_sc_hd__inv_2
XFILLER_10_25 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
X_2649_ VDD VSS _0394_ core.osr.next_result_w\[2\] _0542_ _0555_ net50 VDD VSS sky130_fd_sc_hd__a22o_1
XFILLER_86_18 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XFILLER_19_45 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
Xgenblk2\[7\].buf_n_rown VSS VDD nmatrix_row_core_n_buffered\[7\] core.ndc.row_out_n\[7\]
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
XANTENNA__1568__A VSS VDD core.ndc.col_out_n\[3\] VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__2671__B VSS VDD _1002_ VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_129_1 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_76_95 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_33_113 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XANTENNA__3180__CLK VSS VDD clknet_2_3__leaf_clk_dig_dummy VDD VSS sky130_fd_sc_hd__diode_2
X_1951_ VSS VDD _1405_ _1403_ _1090_ _1404_ VDD VSS sky130_fd_sc_hd__a21bo_1
X_1882_ VSS VDD _1311_ _1349_ _1360_ VDD VSS sky130_fd_sc_hd__nor2_1
X_2503_ VSS VDD _0006_ _0442_ VDD VSS sky130_fd_sc_hd__clkbuf_1
X_2434_ VSS VDD _1325_ _1321_ core.pdc.rowoff_out_n\[8\] _1328_ core.ndc.row_out_n\[12\]
+ VDD VSS sky130_fd_sc_hd__o22a_1
X_2365_ VSS VDD core.osr.result_r\[16\] _0382_ core.osr.result_r\[17\] VDD VSS sky130_fd_sc_hd__nand2_1
XANTENNA__1689__B1 VSS VDD _1199_ VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1941__A VSS VDD _1396_ VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_84_503 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
X_2296_ VSS VDD _0319_ _0271_ _0321_ _0320_ VDD VSS sky130_fd_sc_hd__nand3_1
XFILLER_2_81 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
Xgenblk1\[2\].buf_n_coln VDD VSS core.ndc.col_out_n\[2\] nmatrix_col_core_n_buffered\[2\]
+ VDD VSS sky130_fd_sc_hd__buf_6
XFILLER_52_488 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_137_13 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_137_57 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_47_216 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XANTENNA__1570__B VSS VDD _1037_ VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_15_113 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_102_71 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XANTENNA_pmat_en_bit_n[0] VSS VDD core.cnb.data_register_r\[0\] VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__3187__RESET_B VSS VDD net85 VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1761__A VSS VDD _1072_ VDD VSS sky130_fd_sc_hd__diode_2
X_2150_ VSS VDD _0192_ _0194_ _0190_ VDD VSS sky130_fd_sc_hd__nand2_1
XANTENNA__1480__B VSS VDD _1039_ VDD VSS sky130_fd_sc_hd__diode_2
X_2081_ VSS VDD _0075_ _0148_ _1284_ VDD VSS sky130_fd_sc_hd__nand2_1
XFILLER_93_333 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
X_2983_ VSS VDD _0704_ _0873_ _0695_ VDD VSS sky130_fd_sc_hd__nand2_1
XFILLER_21_149 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
X_1934_ VSS VDD _1390_ _1392_ _1069_ VDD VSS sky130_fd_sc_hd__nand2_1
X_1865_ VDD VSS core.ndc.row_bottotop_n\[5\] _1348_ VDD VSS sky130_fd_sc_hd__inv_2
X_1796_ VDD VSS _1297_ _1296_ _1100_ _1091_ _1279_ core.ndc.col_out\[29\] VDD VSS
+ sky130_fd_sc_hd__a221o_2
XANTENNA__2571__A1 VSS VDD _0439_ VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_107_27 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
X_2417_ VDD VSS _0423_ _0419_ core.osr.sample_count_r\[8\] VDD VSS sky130_fd_sc_hd__and2_1
X_2348_ VDD VSS core.osr.next_result_w\[14\] _0367_ VDD VSS sky130_fd_sc_hd__inv_2
X_2279_ VSS VDD core.osr.result_r\[8\] core.cnb.result_out\[8\] _0305_ VDD VSS sky130_fd_sc_hd__nor2_1
XFILLER_16_68 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XANTENNA_nmat_col_n[10] VSS VDD nmatrix_col_core_n_buffered\[10\] VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1581__A VSS VDD _1039_ VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA_input26_A VSS VDD config_2_in[2] VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_57_97 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XFILLER_90_347 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
X_1650_ VSS VDD _1077_ _1192_ _1132_ VDD VSS sky130_fd_sc_hd__nand2_1
X_1581_ VSS VDD _1039_ _1131_ VDD VSS sky130_fd_sc_hd__clkbuf_2
XANTENNA__2553__A1 VSS VDD core.cnb.result_out\[0\] VDD VSS sky130_fd_sc_hd__diode_2
X_2202_ VDD VSS _0237_ _0235_ _0233_ VDD VSS sky130_fd_sc_hd__or2_1
XFILLER_85_108 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
X_3182_ VSS VDD clknet_2_1__leaf_clk_dig_dummy _0052_ net86 core.cnb.data_register_r\[2\]
+ VDD VSS sky130_fd_sc_hd__dfrtp_1
X_2133_ VSS VDD core.cnb.sampled_avg_control_r\[2\] _0176_ _0177_ VDD VSS sky130_fd_sc_hd__nor2_1
XFILLER_93_185 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XANTENNA__2069__B1 VSS VDD _1075_ VDD VSS sky130_fd_sc_hd__diode_2
X_2064_ VDD VSS _0139_ _0125_ VDD VSS sky130_fd_sc_hd__inv_2
X_2966_ VSS VDD _0855_ _0858_ _0856_ VDD VSS sky130_fd_sc_hd__nand2_1
X_1917_ VSS VDD _1381_ _1362_ core.ndc.rowoff_out_n\[5\] _1380_ VDD VSS sky130_fd_sc_hd__a21bo_1
X_2897_ VSS VDD _0786_ _0787_ _0790_ _1395_ VDD VSS sky130_fd_sc_hd__nand3_1
X_1848_ VDD VSS core.pdc.row_out_n\[6\] _1335_ VDD VSS sky130_fd_sc_hd__inv_2
X_1779_ VDD VSS core.ndc.col_out_n\[25\] core.ndc.col_out\[25\] VDD VSS sky130_fd_sc_hd__inv_2
XFILLER_76_119 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_94_29 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XFILLER_138_121 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XANTENNA_pmat_rowoff_n[5] VSS VDD core.pdc.rowoff_out_n\[5\] VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_108_92 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
XANTENNA__3015__B VSS VDD _1312_ VDD VSS sky130_fd_sc_hd__diode_2
X_2820_ VSS VDD _0713_ _0715_ VDD VSS sky130_fd_sc_hd__clkinvlp_2
XFILLER_129_143 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
X_2751_ VSS VDD _0643_ _0646_ _0647_ VDD VSS sky130_fd_sc_hd__nor2_1
X_2682_ VSS VDD core.osr.next_result_w\[8\] _0540_ _0584_ _0528_ VDD VSS sky130_fd_sc_hd__o21ai_1
X_1702_ VSS VDD _1149_ _1236_ _1235_ VDD VSS sky130_fd_sc_hd__nand2_1
XANTENNA__1577__A2 VSS VDD _1128_ VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1486__A VSS VDD _1045_ VDD VSS sky130_fd_sc_hd__diode_2
X_1633_ VSS VDD _1179_ _1178_ _1174_ _1168_ VDD VSS sky130_fd_sc_hd__and3_1
X_1564_ VSS VDD _1116_ _1118_ _1117_ VDD VSS sky130_fd_sc_hd__nand2_1
X_1495_ VDD VSS core.cnb.data_register_r\[4\] _1055_ VDD VSS sky130_fd_sc_hd__buf_4
XANTENNA__3114__CLK VSS VDD clknet_2_2__leaf_clk_dig_dummy VDD VSS sky130_fd_sc_hd__diode_2
X_3165_ VSS VDD net60 core.osr.next_result_w\[5\] net72 core.osr.result_r\[5\] VDD
+ VSS sky130_fd_sc_hd__dfrtp_1
XFILLER_66_141 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
X_3096_ VSS VDD _0062_ _0979_ VDD VSS sky130_fd_sc_hd__clkbuf_1
X_2116_ VSS VDD _1406_ _0167_ _1188_ VDD VSS sky130_fd_sc_hd__nand2_1
X_2047_ VSS VDD _1413_ _0128_ _1235_ VDD VSS sky130_fd_sc_hd__nand2_1
Xfanout59 VDD VSS net59 net61 VDD VSS sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_13_25 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
X_2949_ VSS VDD _0839_ _0482_ _0841_ _0840_ VDD VSS sky130_fd_sc_hd__nand3_1
XFILLER_129_25 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_135_113 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XANTENNA__2004__B VSS VDD _1284_ VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA_genblk1\[17\].buf_n_coln_A VSS VDD core.ndc.col_out_n\[17\] VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA_fanout76_A VSS VDD net82 VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_54_32 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_54_76 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XFILLER_110_60 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
Xgenblk2\[1\].buf_n_rowonn VSS VDD nmatrix_rowon_core_n_buffered\[1\] core.ndc.rowon_out_n\[1\]
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
XFILLER_70_97 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XANTENNA__3137__CLK VSS VDD clknet_2_0__leaf_clk_dig_dummy VDD VSS sky130_fd_sc_hd__diode_2
Xgenblk1\[7\].buf_n_coln VDD VSS core.ndc.col_out_n\[7\] nmatrix_col_core_n_buffered\[7\]
+ VDD VSS sky130_fd_sc_hd__buf_6
X_2803_ VDD VSS _0698_ core.cnb.shift_register_r\[13\] VDD VSS sky130_fd_sc_hd__inv_2
X_2734_ VDD VSS _0393_ core.cnb.result_out\[11\] _0562_ _0631_ net44 VDD VSS sky130_fd_sc_hd__a22o_1
X_2665_ VSS VDD core.osr.next_result_w\[8\] _0569_ _0568_ VDD VSS sky130_fd_sc_hd__nand2_1
X_2596_ VSS VDD _0511_ core.cnb.result_out\[9\] _0480_ _0510_ VDD VSS sky130_fd_sc_hd__mux2_1
X_1616_ VDD VSS _1162_ _1036_ _1134_ VDD VSS sky130_fd_sc_hd__and2_1
XFILLER_115_27 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
X_1547_ VSS VDD _1078_ _1103_ VDD VSS sky130_fd_sc_hd__clkbuf_2
X_1478_ VSS VDD _1031_ _1038_ VDD VSS sky130_fd_sc_hd__clkbuf_2
X_3148_ VSS VDD net56 _0038_ net68 net48 VDD VSS sky130_fd_sc_hd__dfrtp_1
X_3079_ VDD VSS _0965_ _0955_ _0964_ VDD VSS sky130_fd_sc_hd__or2_1
XFILLER_24_35 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XFILLER_108_102 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XANTENNA__1748__B VSS VDD _1173_ VDD VSS sky130_fd_sc_hd__diode_2
X_2450_ VSS VDD _1378_ core.ndc.rowon_out_n\[11\] _1370_ VDD VSS sky130_fd_sc_hd__nand2_1
X_2381_ VDD VSS _0394_ _0395_ VDD VSS sky130_fd_sc_hd__buf_4
XANTENNA_cgen_dlycontrol1_in[0] VSS VDD net18 VDD VSS sky130_fd_sc_hd__diode_2
Xinput5 VSS VDD config_1_in[12] net5 VDD VSS sky130_fd_sc_hd__clkbuf_2
X_3002_ VSS VDD _0847_ _0891_ _0888_ VDD VSS sky130_fd_sc_hd__nand2_1
XFILLER_91_261 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_51_169 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XANTENNA__2534__S VSS VDD net54 VDD VSS sky130_fd_sc_hd__diode_2
X_2717_ VDD VSS core.osr.next_result_w\[10\] net43 _0393_ _0615_ _0562_ VDD VSS sky130_fd_sc_hd__a22o_1
X_2648_ VDD VSS _0554_ _0516_ _0520_ VDD VSS sky130_fd_sc_hd__or2_1
X_2579_ VDD VSS _0027_ _0496_ _0497_ _0461_ core.cnb.result_out\[5\] VDD VSS sky130_fd_sc_hd__o2bb2a_1
XFILLER_47_409 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_19_57 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XFILLER_76_85 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XFILLER_46_453 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_33_136 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_33_125 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XFILLER_92_95 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
X_1950_ VSS VDD _1400_ _1404_ _1086_ VDD VSS sky130_fd_sc_hd__nand2_1
X_1881_ VSS VDD _1336_ _1358_ _1359_ VDD VSS sky130_fd_sc_hd__nor2_1
X_2502_ VSS VDD _0442_ core.cnb.shift_register_r\[5\] _0203_ core.cnb.shift_register_r\[4\]
+ VDD VSS sky130_fd_sc_hd__mux2_1
XANTENNA__2583__C1 VSS VDD _0439_ VDD VSS sky130_fd_sc_hd__diode_2
X_2433_ VDD VSS core.ndc.row_out_n\[11\] _0427_ VDD VSS sky130_fd_sc_hd__inv_2
X_2364_ VDD VSS core.osr.result_r\[16\] _0377_ core.osr.result_r\[17\] _0381_ VDD
+ VSS sky130_fd_sc_hd__a21o_1
XFILLER_110_141 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
X_2295_ VSS VDD _0318_ _0320_ _0317_ VDD VSS sky130_fd_sc_hd__nand2_1
XFILLER_84_515 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_52_445 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
XANTENNA__2491__C VSS VDD _1040_ VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_137_25 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XANTENNA__3095__S VSS VDD _0241_ VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_137_69 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_87_342 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XFILLER_15_125 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_11_80 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XFILLER_127_91 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_87_51 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
X_2080_ VDD VSS core.pdc.col_out_n\[20\] core.pdc.col_out\[20\] VDD VSS sky130_fd_sc_hd__inv_2
XFILLER_93_367 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
XANTENNA__2096__B2 VSS VDD _1102_ VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1489__A VSS VDD _1037_ VDD VSS sky130_fd_sc_hd__diode_2
X_2982_ VSS VDD _0055_ _0757_ _0872_ _0871_ _1114_ _0688_ VDD VSS sky130_fd_sc_hd__a32o_1
X_1933_ VDD VSS _1089_ _1390_ _1057_ _1391_ VDD VSS sky130_fd_sc_hd__or3_1
X_1864_ VSS VDD _1308_ _1318_ _1348_ VDD VSS sky130_fd_sc_hd__nor2_1
Xinput30 VDD VSS net30 config_2_in[6] VDD VSS sky130_fd_sc_hd__dlymetal6s2s_1
X_1795_ VSS VDD _1272_ _1143_ _1297_ VDD VSS sky130_fd_sc_hd__nor2_1
X_2416_ VSS VDD core.osr.sample_count_r\[8\] _0419_ _0422_ VDD VSS sky130_fd_sc_hd__nor2_1
X_2347_ VSS VDD _0365_ _0240_ _0367_ _0366_ VDD VSS sky130_fd_sc_hd__nand3_1
X_2278_ VSS VDD _0304_ core.osr.next_result_w\[7\] VDD VSS sky130_fd_sc_hd__clkbuf_2
XFILLER_16_47 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XFILLER_79_106 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
XANTENNA__3170__CLK VSS VDD net61 VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_57_32 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XANTENNA__2693__A VSS VDD _0395_ VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA_input19_A VSS VDD config_2_in[10] VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_90_359 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
X_1580_ VDD VSS core.ndc.col_out_n\[4\] core.ndc.col_out\[4\] VDD VSS sky130_fd_sc_hd__inv_2
XANTENNA__2002__A1 VSS VDD _1082_ VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_98_72 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
X_2201_ VSS VDD _0233_ _0236_ _0235_ VDD VSS sky130_fd_sc_hd__nand2_1
X_3181_ VSS VDD clknet_2_1__leaf_clk_dig_dummy _0051_ net86 core.cnb.data_register_r\[1\]
+ VDD VSS sky130_fd_sc_hd__dfrtp_4
X_2132_ VDD VSS _0176_ core.cnb.sampled_avg_control_r\[1\] VDD VSS sky130_fd_sc_hd__inv_2
XANTENNA__2069__A1 VSS VDD _1126_ VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_93_197 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XANTENNA__2069__B2 VSS VDD _0115_ VDD VSS sky130_fd_sc_hd__diode_2
X_2063_ VDD VSS core.pdc.col_out_n\[16\] core.pdc.col_out\[16\] VDD VSS sky130_fd_sc_hd__clkinv_2
XANTENNA__2108__A VSS VDD _1131_ VDD VSS sky130_fd_sc_hd__diode_2
X_2965_ VDD VSS _0855_ _0831_ _0856_ _0857_ VDD VSS sky130_fd_sc_hd__a21o_1
X_1916_ VSS VDD _1372_ _1380_ _1331_ VDD VSS sky130_fd_sc_hd__nand2_1
X_2896_ VSS VDD _0788_ _0789_ _1076_ VDD VSS sky130_fd_sc_hd__nand2_1
X_1847_ VDD VSS _1331_ _1320_ _1334_ _1335_ VDD VSS sky130_fd_sc_hd__a21o_1
X_1778_ VSS VDD core.ndc.col_out\[25\] _1157_ _1284_ _1285_ _1287_ VDD VSS sky130_fd_sc_hd__a211o_2
XANTENNA_genblk2\[5\].buf_p_rown_A VSS VDD core.ndc.row_bottotop_n\[10\] VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_138_133 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
XANTENNA__1576__B VSS VDD _1057_ VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_104_1 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
XFILLER_84_41 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_84_85 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XANTENNA__1767__A VSS VDD _1032_ VDD VSS sky130_fd_sc_hd__diode_2
X_2750_ VSS VDD _0646_ _0644_ _0645_ VDD VSS sky130_fd_sc_hd__nand2_2
X_2681_ VSS VDD _0356_ _0582_ _0583_ _0517_ VDD VSS sky130_fd_sc_hd__o21ai_1
X_1701_ VDD VSS _1235_ net15 VDD VSS sky130_fd_sc_hd__buf_2
X_1632_ VSS VDD _1176_ _1178_ _1177_ VDD VSS sky130_fd_sc_hd__nand2_1
XANTENNA__3171__RESET_B VSS VDD net73 VDD VSS sky130_fd_sc_hd__diode_2
X_1563_ VDD VSS _1117_ core.cnb.data_register_r\[7\] VDD VSS sky130_fd_sc_hd__buf_2
X_1494_ VSS VDD _1041_ _1054_ VDD VSS sky130_fd_sc_hd__clkbuf_2
XANTENNA__2110__B VSS VDD _1177_ VDD VSS sky130_fd_sc_hd__diode_2
X_3164_ VSS VDD net62 core.osr.next_result_w\[4\] net74 core.osr.result_r\[4\] VDD
+ VSS sky130_fd_sc_hd__dfrtp_1
X_3095_ VSS VDD _0979_ core.osr.osr_mode_r\[0\] _0241_ net11 VDD VSS sky130_fd_sc_hd__mux2_1
X_2115_ VSS VDD _1398_ _0166_ _1096_ VDD VSS sky130_fd_sc_hd__nand2_1
X_2046_ VDD VSS _0126_ _0127_ VDD VSS sky130_fd_sc_hd__clkinv_2
XANTENNA__1677__A VSS VDD _1216_ VDD VSS sky130_fd_sc_hd__diode_2
X_2948_ VDD VSS _0840_ _0791_ VDD VSS sky130_fd_sc_hd__inv_2
XFILLER_129_37 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
XFILLER_135_125 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
X_2879_ VSS VDD _0771_ _0773_ _0772_ VDD VSS sky130_fd_sc_hd__nand2_1
XANTENNA__2020__B VSS VDD _1093_ VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_57_131 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XFILLER_85_462 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XFILLER_85_495 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XFILLER_110_50 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XFILLER_70_21 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XFILLER_110_72 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_79_85 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
X_2802_ VSS VDD _0684_ _0696_ _0697_ VDD VSS sky130_fd_sc_hd__nor2_1
X_2733_ VSS VDD _0628_ _0630_ _0629_ VDD VSS sky130_fd_sc_hd__nand2_1
XANTENNA__2105__B VSS VDD _1092_ VDD VSS sky130_fd_sc_hd__diode_2
X_2664_ VSS VDD _1001_ _0568_ VDD VSS sky130_fd_sc_hd__clkbuf_2
X_2595_ VDD VSS _0510_ _0508_ _0509_ VDD VSS sky130_fd_sc_hd__or2_1
X_1615_ VSS VDD _1160_ _1161_ _1051_ VDD VSS sky130_fd_sc_hd__nor2_2
Xgenblk2\[6\].buf_p_rowonn VSS VDD pmatrix_rowon_core_n_buffered\[6\] core.pdc.rowon_out_n\[6\]
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
XANTENNA_cgen_enable_dlycontrol_in VSS VDD net24 VDD VSS sky130_fd_sc_hd__diode_2
X_1546_ VDD VSS _1102_ _1101_ VDD VSS sky130_fd_sc_hd__buf_2
X_1477_ VDD VSS _1037_ _1036_ VDD VSS sky130_fd_sc_hd__inv_2
X_3147_ VSS VDD net56 _0037_ net68 net47 VDD VSS sky130_fd_sc_hd__dfrtp_1
X_3078_ VSS VDD _0957_ _0964_ _0963_ VDD VSS sky130_fd_sc_hd__nand2_1
XANTENNA__2435__A1 VSS VDD core.pdc.rowoff_out_n\[8\] VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__2435__B2 VSS VDD core.ndc.row_bottotop_n\[10\] VDD VSS sky130_fd_sc_hd__diode_2
X_2029_ VSS VDD _0084_ _0114_ _1155_ VDD VSS sky130_fd_sc_hd__nand2_1
XANTENNA_genblk2\[15\].buf_p_rowonn_A VSS VDD core.pdc.rowon_out_n\[15\] VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_40_79 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XFILLER_6_5 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_49_88 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_105_94 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XANTENNA__3104__CLK VSS VDD clknet_2_2__leaf_clk_dig_dummy VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_81_97 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
X_2380_ VSS VDD _0393_ _0394_ VDD VSS sky130_fd_sc_hd__clkbuf_2
Xinput6 VSS VDD config_1_in[13] net6 VDD VSS sky130_fd_sc_hd__clkbuf_2
X_3001_ VSS VDD _0795_ _0890_ _0889_ VDD VSS sky130_fd_sc_hd__nand2_1
XFILLER_83_229 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
XFILLER_101_19 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XFILLER_91_273 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
XFILLER_51_159 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
X_2716_ VSS VDD _0612_ _0047_ _0614_ VDD VSS sky130_fd_sc_hd__nand2_1
X_2647_ VDD VSS _1000_ core.osr.next_result_w\[10\] _0552_ _0553_ VDD VSS sky130_fd_sc_hd__a21o_1
XANTENNA__1674__B VSS VDD _1213_ VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_126_38 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
X_2578_ VDD VSS _1065_ _0489_ _0480_ _0497_ VDD VSS sky130_fd_sc_hd__a21oi_1
X_1529_ VDD VSS _1087_ _1044_ VDD VSS sky130_fd_sc_hd__inv_2
XANTENNA__3127__CLK VSS VDD clknet_2_3__leaf_clk_dig_dummy VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_51_67 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_51_89 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XANTENNA_nmat_row_n[1] VSS VDD nmatrix_row_core_n_buffered\[1\] VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_104_150 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
XFILLER_76_31 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XFILLER_93_505 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_18_112 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
XFILLER_33_148 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
X_1880_ VSS VDD _1317_ _1358_ _1029_ VDD VSS sky130_fd_sc_hd__nand2_1
XANTENNA__1775__A VSS VDD _1126_ VDD VSS sky130_fd_sc_hd__diode_2
X_2501_ VSS VDD _0005_ _0441_ VDD VSS sky130_fd_sc_hd__clkbuf_1
X_2432_ VSS VDD _1322_ _0427_ _1330_ VDD VSS sky130_fd_sc_hd__nand2_1
X_2363_ VDD VSS core.osr.next_result_w\[16\] _0380_ VDD VSS sky130_fd_sc_hd__inv_2
XANTENNA__1689__A2 VSS VDD _1206_ VDD VSS sky130_fd_sc_hd__diode_2
X_2294_ VDD VSS _0319_ _0317_ _0318_ VDD VSS sky130_fd_sc_hd__or2_1
XFILLER_112_29 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XFILLER_137_37 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_55_295 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_15_137 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XANTENNA__1595__A VSS VDD _1045_ VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__2096__A2 VSS VDD _1275_ VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_46_262 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
XFILLER_46_273 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
XFILLER_46_295 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
X_2981_ VSS VDD _0863_ _0802_ _0872_ _0870_ VDD VSS sky130_fd_sc_hd__nand3_1
X_1932_ VDD VSS _1390_ _1389_ VDD VSS sky130_fd_sc_hd__dlymetal6s2s_1
X_1863_ VDD VSS core.pdc.row_out_n\[9\] _1347_ VDD VSS sky130_fd_sc_hd__inv_2
Xinput31 VDD VSS net31 config_2_in[7] VDD VSS sky130_fd_sc_hd__dlymetal6s2s_1
Xinput20 VDD VSS net20 config_2_in[11] VDD VSS sky130_fd_sc_hd__dlymetal6s2s_1
X_1794_ VDD VSS _1296_ _1095_ VDD VSS sky130_fd_sc_hd__buf_2
X_2415_ VDD VSS core.osr.next_sample_count_w\[7\] _0421_ VDD VSS sky130_fd_sc_hd__inv_2
X_2346_ VSS VDD _0353_ core.osr.result_r\[14\] _0366_ _0358_ VDD VSS sky130_fd_sc_hd__nand3_1
X_2277_ VSS VDD core.cnb.result_out\[7\] _0271_ _0303_ _0304_ VDD VSS sky130_fd_sc_hd__o21a_1
XFILLER_12_118 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_20_151 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XFILLER_90_316 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_113_50 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
XFILLER_73_76 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
X_2200_ VDD VSS _0235_ core.cnb.average_sum_r\[4\] VDD VSS sky130_fd_sc_hd__inv_2
X_3180_ VSS VDD clknet_2_3__leaf_clk_dig_dummy _0050_ net86 core.cnb.data_register_r\[0\]
+ VDD VSS sky130_fd_sc_hd__dfrtp_4
X_2131_ VDD VSS core.cnb.data_register_r\[2\] core.cnb.pswitch_out\[2\] VDD VSS sky130_fd_sc_hd__clkinv_2
X_2062_ VSS VDD _1075_ _0135_ _0094_ _1064_ core.pdc.col_out_n\[16\] _0138_ VDD VSS
+ sky130_fd_sc_hd__o221a_1
XFILLER_75_891 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XANTENNA__2108__B VSS VDD _0091_ VDD VSS sky130_fd_sc_hd__diode_2
X_2964_ VSS VDD _0847_ _0856_ VDD VSS sky130_fd_sc_hd__clkbuf_2
X_1915_ VSS VDD core.ndc.rowoff_out_n\[5\] core.ndc.row_bottotop_n\[5\] core.ndc.rowon_bottotop_n\[5\]
+ VDD VSS sky130_fd_sc_hd__nand2_2
X_2895_ VSS VDD _0786_ _0788_ _0787_ VDD VSS sky130_fd_sc_hd__nand2_1
X_1846_ VSS VDD _1333_ _1316_ _1334_ VDD VSS sky130_fd_sc_hd__nor2_1
X_1777_ VDD VSS _1287_ _1286_ VDD VSS sky130_fd_sc_hd__inv_2
XFILLER_89_449 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XANTENNA__1504__A1 VSS VDD _1035_ VDD VSS sky130_fd_sc_hd__diode_2
X_2329_ VSS VDD _0351_ _0317_ _0307_ _0350_ VDD VSS sky130_fd_sc_hd__and3_1
XFILLER_66_891 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XFILLER_43_13 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XANTENNA__1873__A VSS VDD _1353_ VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1592__B VSS VDD _1112_ VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_68_87 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XANTENNA_input31_A VSS VDD config_2_in[7] VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_84_53 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XFILLER_90_102 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XFILLER_84_75 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XFILLER_72_883 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
X_2680_ VSS VDD core.osr.next_result_w\[10\] _0582_ _0568_ VDD VSS sky130_fd_sc_hd__nand2_1
X_1700_ VDD VSS _1234_ _1034_ _1204_ VDD VSS sky130_fd_sc_hd__or2_1
X_1631_ VDD VSS _1177_ _1072_ VDD VSS sky130_fd_sc_hd__buf_2
XANTENNA__1783__A VSS VDD _1131_ VDD VSS sky130_fd_sc_hd__diode_2
X_1562_ VSS VDD _1113_ _1115_ _1116_ VDD VSS sky130_fd_sc_hd__nor2_1
X_1493_ VSS VDD _1052_ _1053_ VDD VSS sky130_fd_sc_hd__clkbuf_4
X_3163_ VSS VDD net63 core.osr.next_result_w\[3\] net74 core.osr.result_r\[3\] VDD
+ VSS sky130_fd_sc_hd__dfrtp_1
XANTENNA__3140__RESET_B VSS VDD net81 VDD VSS sky130_fd_sc_hd__diode_2
X_2114_ VDD VSS core.pdc.col_out_n\[28\] core.pdc.col_out\[28\] VDD VSS sky130_fd_sc_hd__clkinv_2
X_3094_ VSS VDD _0977_ _0061_ _0978_ VDD VSS sky130_fd_sc_hd__nand2_1
XFILLER_81_113 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
X_2045_ VSS VDD _1227_ _0125_ _0126_ VDD VSS sky130_fd_sc_hd__nor2_1
XFILLER_63_883 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
X_2947_ VDD VSS _0475_ _0837_ _0838_ _0839_ VDD VSS sky130_fd_sc_hd__a21oi_1
XFILLER_129_49 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
X_2878_ VSS VDD _0772_ _0471_ _0760_ _0770_ VDD VSS sky130_fd_sc_hd__nand3b_1
XANTENNA__1973__B2 VSS VDD _1296_ VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1973__A1 VSS VDD _1121_ VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_135_137 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
X_1829_ VSS VDD _1022_ _1319_ _1320_ VDD VSS sky130_fd_sc_hd__nor2_1
XFILLER_79_75 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XFILLER_135_81 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_63_113 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XANTENNA__3183__CLK VSS VDD clknet_2_1__leaf_clk_dig_dummy VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_91_477 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
X_2801_ VSS VDD _0693_ _0696_ _0695_ VDD VSS sky130_fd_sc_hd__nand2_1
X_2732_ VDD VSS _0530_ _0363_ _1018_ _0629_ VDD VSS sky130_fd_sc_hd__a21oi_1
XANTENNA__1955__B2 VSS VDD _1296_ VDD VSS sky130_fd_sc_hd__diode_2
X_2663_ VSS VDD core.osr.next_result_w\[10\] _0567_ _0535_ VDD VSS sky130_fd_sc_hd__nand2_1
X_2594_ VSS VDD _1303_ _0503_ _0509_ VDD VSS sky130_fd_sc_hd__nor2_1
X_1614_ VSS VDD _1058_ _1066_ _1160_ VDD VSS sky130_fd_sc_hd__nor2_1
X_1545_ VSS VDD _1032_ _1101_ VDD VSS sky130_fd_sc_hd__clkbuf_2
XANTENNA__2121__B VSS VDD _1096_ VDD VSS sky130_fd_sc_hd__diode_2
X_1476_ VSS VDD _1036_ core.cnb.data_register_r\[3\] core.cnb.data_register_r\[4\]
+ VDD VSS sky130_fd_sc_hd__nor2_4
XFILLER_86_249 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
X_3146_ VSS VDD net56 _0036_ net68 net46 VDD VSS sky130_fd_sc_hd__dfrtp_1
XFILLER_54_113 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
X_3077_ VSS VDD _0948_ _0960_ _0962_ _0963_ VDD VSS sky130_fd_sc_hd__o21a_1
X_2028_ VSS VDD _1136_ _1228_ _0113_ _1394_ VDD VSS sky130_fd_sc_hd__o21ai_2
XANTENNA__1688__A VSS VDD _1074_ VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__2791__B VSS VDD core.cnb.data_register_r\[0\] VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1643__B1 VSS VDD _1186_ VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA_fanout81_A VSS VDD net82 VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_45_113 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_81_32 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XFILLER_81_76 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XANTENNA_genblk1\[13\].buf_n_coln_A VSS VDD core.ndc.col_out_n\[13\] VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_114_107 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XANTENNA__2222__A VSS VDD _0254_ VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1780__B VSS VDD _1284_ VDD VSS sky130_fd_sc_hd__diode_2
Xinput7 VSS VDD config_1_in[14] net7 VDD VSS sky130_fd_sc_hd__clkbuf_2
X_3000_ VDD VSS _0889_ _0888_ VDD VSS sky130_fd_sc_hd__inv_2
XANTENNA__2116__B VSS VDD _1188_ VDD VSS sky130_fd_sc_hd__diode_2
Xgenblk2\[13\].buf_p_rown VSS VDD pmatrix_row_core_n_buffered\[13\] core.pdc.row_out_n\[13\]
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
X_2715_ VDD VSS _0614_ _0613_ VDD VSS sky130_fd_sc_hd__inv_2
XANTENNA__2132__A VSS VDD core.cnb.sampled_avg_control_r\[1\] VDD VSS sky130_fd_sc_hd__diode_2
X_2646_ VSS VDD _0550_ _0552_ _0551_ VDD VSS sky130_fd_sc_hd__nand2_1
X_2577_ VSS VDD _0493_ _0496_ _1114_ VDD VSS sky130_fd_sc_hd__nand2_1
XANTENNA__1690__B VSS VDD _1093_ VDD VSS sky130_fd_sc_hd__diode_2
X_1528_ VSS VDD _1079_ _1085_ _1086_ VDD VSS sky130_fd_sc_hd__nor2_1
X_1459_ VDD VSS core.cnb.data_register_r\[10\] _1022_ VDD VSS sky130_fd_sc_hd__clkinv_2
XFILLER_27_113 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_55_433 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
X_3129_ VSS VDD clknet_2_3__leaf_clk_dig_dummy core.cnb.next_average_sum_w\[2\] net91
+ core.cnb.average_sum_r\[2\] VDD VSS sky130_fd_sc_hd__dfrtp_1
XFILLER_55_455 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
XFILLER_50_160 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_51_46 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XANTENNA__2042__A VSS VDD _0089_ VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA_nmat_row_n[0] VSS VDD nmatrix_row_core_n_buffered\[0\] VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_93_517 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
XANTENNA__2032__A0 VSS VDD _1199_ VDD VSS sky130_fd_sc_hd__diode_2
X_2500_ VSS VDD _0441_ core.cnb.shift_register_r\[4\] _0220_ core.cnb.shift_register_r\[3\]
+ VDD VSS sky130_fd_sc_hd__mux2_1
XANTENNA__2583__B2 VSS VDD _1117_ VDD VSS sky130_fd_sc_hd__diode_2
X_2431_ VSS VDD core.ndc.row_bottotop_n\[10\] _1321_ _1311_ _1027_ core.ndc.row_out_n\[10\]
+ VDD VSS sky130_fd_sc_hd__o22a_1
XANTENNA__1791__A VSS VDD _1272_ VDD VSS sky130_fd_sc_hd__diode_2
X_2362_ VSS VDD _0378_ _0241_ _0380_ _0379_ VDD VSS sky130_fd_sc_hd__nand3_1
X_2293_ VSS VDD _0311_ _0318_ _0306_ VDD VSS sky130_fd_sc_hd__nand2_1
XFILLER_56_208 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XANTENNA_nmat_sample_buf_n_A VSS VDD core.cnb.enable_loop_out VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1966__A VSS VDD core.pdc.col_out\[3\] VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_137_49 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
X_2629_ VDD VSS _0537_ _1011_ VDD VSS sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_46_57 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
XFILLER_46_79 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XFILLER_102_41 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XANTENNA__2037__A VSS VDD _0098_ VDD VSS sky130_fd_sc_hd__diode_2
Xgenblk2\[10\].buf_n_rown VSS VDD nmatrix_row_core_n_buffered\[10\] core.ndc.row_out_n\[10\]
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
XANTENNA__1595__B VSS VDD _1079_ VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_97_119 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XANTENNA__1525__C1 VSS VDD _1082_ VDD VSS sky130_fd_sc_hd__diode_2
Xgenblk2\[15\].buf_n_rowonn VSS VDD nmatrix_rowon_core_n_buffered\[15\] core.ndc.rowon_out_n\[15\]
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
XFILLER_46_230 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
XFILLER_46_241 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
X_2980_ VDD VSS _0802_ _0863_ _0870_ _0871_ VDD VSS sky130_fd_sc_hd__a21o_1
XANTENNA__1786__A VSS VDD _1106_ VDD VSS sky130_fd_sc_hd__diode_2
X_1931_ VSS VDD _1388_ _1389_ VDD VSS sky130_fd_sc_hd__clkbuf_2
X_1862_ VDD VSS _1347_ _1344_ _1346_ VDD VSS sky130_fd_sc_hd__or2_2
Xinput21 VDD VSS net21 config_2_in[12] VDD VSS sky130_fd_sc_hd__dlymetal6s2s_1
Xinput10 VSS VDD net10 config_1_in[2] VDD VSS sky130_fd_sc_hd__clkbuf_1
XANTENNA__2005__B1 VSS VDD _1035_ VDD VSS sky130_fd_sc_hd__diode_2
X_1793_ VDD VSS core.ndc.col_out_n\[28\] core.ndc.col_out\[28\] VDD VSS sky130_fd_sc_hd__inv_2
Xinput32 VDD VSS net32 config_2_in[8] VDD VSS sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_107_19 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
X_2414_ VSS VDD _1021_ _0420_ _0419_ _0421_ VDD VSS sky130_fd_sc_hd__or3b_1
XANTENNA__3117__CLK VSS VDD clknet_2_2__leaf_clk_dig_dummy VDD VSS sky130_fd_sc_hd__diode_2
X_2345_ VSS VDD _0359_ _0365_ _0364_ VDD VSS sky130_fd_sc_hd__nand2_1
X_2276_ VSS VDD _0302_ _0255_ _0303_ _0301_ VDD VSS sky130_fd_sc_hd__o21ai_1
XFILLER_84_369 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_48_506 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_90_328 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_73_88 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_22_92 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
XFILLER_98_41 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
Xgenblk1\[14\].buf_p_coln VSS VDD pmatrix_col_core_n_buffered\[14\] core.pdc.col_out_n\[14\]
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
XANTENNA__2230__A VSS VDD _0255_ VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_98_85 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XANTENNA__3045__B VSS VDD _1114_ VDD VSS sky130_fd_sc_hd__diode_2
X_2130_ VDD VSS core.pdc.col_out\[31\] core.pdc.col_out_n\[31\] VDD VSS sky130_fd_sc_hd__clkinv_2
XFILLER_14_5 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
X_2061_ VSS VDD _1391_ _0138_ _1093_ VDD VSS sky130_fd_sc_hd__nand2_1
X_2963_ VSS VDD _0855_ _0818_ _0745_ _0854_ VDD VSS sky130_fd_sc_hd__and3_1
X_1914_ VSS VDD _1336_ _1366_ core.pdc.rowon_out_n\[9\] core.ndc.rowon_bottotop_n\[5\]
+ VDD VSS sky130_fd_sc_hd__a21oi_2
X_2894_ VSS VDD _0787_ _0783_ _0472_ _0785_ VDD VSS sky130_fd_sc_hd__nand3b_1
X_1845_ VSS VDD _1332_ _1333_ _1300_ VDD VSS sky130_fd_sc_hd__nand2_1
X_1776_ VDD VSS _1286_ _1033_ _1119_ VDD VSS sky130_fd_sc_hd__or2_1
X_2328_ VSS VDD _0332_ _0344_ _0350_ VDD VSS sky130_fd_sc_hd__nor2_1
XFILLER_84_111 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
X_2259_ VSS VDD _0288_ _0287_ _0240_ _0280_ VDD VSS sky130_fd_sc_hd__o21a_2
XFILLER_43_25 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XANTENNA__2985__A VSS VDD _0799_ VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_68_99 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
XFILLER_88_494 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XANTENNA_input24_A VSS VDD config_2_in[15] VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_84_21 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
XFILLER_90_125 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
X_1630_ VDD VSS _1176_ _1175_ VDD VSS sky130_fd_sc_hd__inv_2
X_1561_ VSS VDD _1114_ _1037_ _1115_ VDD VSS sky130_fd_sc_hd__nor2_1
X_1492_ VSS VDD _1051_ _1052_ VDD VSS sky130_fd_sc_hd__clkbuf_2
X_3162_ VSS VDD net63 core.osr.next_result_w\[2\] net75 core.osr.result_r\[2\] VDD
+ VSS sky130_fd_sc_hd__dfrtp_1
X_2113_ VSS VDD core.pdc.col_out_n\[28\] _0165_ VDD VSS sky130_fd_sc_hd__clkbuf_1
X_3093_ VSS VDD _0758_ _0978_ _1309_ VDD VSS sky130_fd_sc_hd__nand2_1
XANTENNA__3180__RESET_B VSS VDD net86 VDD VSS sky130_fd_sc_hd__diode_2
X_2044_ VSS VDD _1161_ _1403_ _0124_ _0125_ VDD VSS sky130_fd_sc_hd__o21a_1
XFILLER_50_501 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
X_2946_ VSS VDD _0475_ _0835_ _0838_ VDD VSS sky130_fd_sc_hd__nor2_1
Xgenblk1\[11\].buf_n_coln VSS VDD nmatrix_col_core_n_buffered\[11\] core.ndc.col_out_n\[11\]
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
X_2877_ VSS VDD _0761_ _0771_ _0770_ VDD VSS sky130_fd_sc_hd__nand2_1
XFILLER_135_105 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
X_1828_ VDD VSS _1319_ _1028_ VDD VSS sky130_fd_sc_hd__inv_2
XANTENNA__1974__A VSS VDD core.pdc.col_out\[4\] VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_135_149 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
X_1759_ VDD VSS core.ndc.col_out_n\[22\] core.ndc.col_out\[22\] VDD VSS sky130_fd_sc_hd__inv_2
XANTENNA_nmat_col[9] VSS VDD core.ndc.col_out\[9\] VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__2029__B VSS VDD _1155_ VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA_genblk2\[1\].buf_p_rown_A VSS VDD core.pdc.row_out_n\[1\] VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__2045__A VSS VDD _1227_ VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_110_85 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_135_93 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_48_144 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_63_125 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XANTENNA__2881__C VSS VDD _0482_ VDD VSS sky130_fd_sc_hd__diode_2
X_2800_ VSS VDD _0640_ _0682_ _0695_ _0694_ VDD VSS sky130_fd_sc_hd__nand3_1
X_2731_ VSS VDD _0623_ _0628_ _0627_ VDD VSS sky130_fd_sc_hd__nand2_1
XANTENNA__1794__A VSS VDD _1095_ VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1955__A2 VSS VDD _1279_ VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_117_138 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
X_2662_ VDD VSS _1008_ _0356_ _0524_ _0566_ VDD VSS sky130_fd_sc_hd__a21oi_1
X_1613_ VDD VSS core.ndc.col_out_n\[6\] core.ndc.col_out\[6\] VDD VSS sky130_fd_sc_hd__inv_2
X_2593_ VSS VDD _0507_ _0502_ _0508_ VDD VSS sky130_fd_sc_hd__nor2_1
XFILLER_132_119 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
X_1544_ VDD VSS _1100_ _1099_ VDD VSS sky130_fd_sc_hd__inv_2
XFILLER_5_84 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
X_1475_ VDD VSS _1035_ _1034_ VDD VSS sky130_fd_sc_hd__buf_2
XANTENNA__2668__B1 VSS VDD _0394_ VDD VSS sky130_fd_sc_hd__diode_2
X_3145_ VSS VDD net56 _0035_ net68 net45 VDD VSS sky130_fd_sc_hd__dfrtp_1
X_3076_ VSS VDD _0962_ _0961_ _0833_ _0918_ _0507_ VDD VSS sky130_fd_sc_hd__a211o_1
X_2027_ VDD VSS core.pdc.col_out_n\[11\] core.pdc.col_out\[11\] VDD VSS sky130_fd_sc_hd__clkinv_2
XFILLER_50_331 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
XANTENNA__1643__A1 VSS VDD _1113_ VDD VSS sky130_fd_sc_hd__diode_2
X_2929_ VDD VSS _0821_ _0818_ VDD VSS sky130_fd_sc_hd__inv_2
Xgenblk2\[15\].buf_n_rown VSS VDD nmatrix_row_core_n_buffered\[15\] core.ndc.row_out_n\[15\]
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
XFILLER_108_116 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_40_37 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_123_108 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XFILLER_49_35 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_49_57 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XFILLER_105_74 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_45_125 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XFILLER_60_128 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_81_88 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
XFILLER_114_119 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_122_141 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
Xinput8 VSS VDD config_1_in[15] net8 VDD VSS sky130_fd_sc_hd__clkbuf_2
XFILLER_51_117 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
X_2714_ VDD VSS core.osr.next_result_w\[9\] net42 _1020_ _0613_ _0562_ VDD VSS sky130_fd_sc_hd__a22o_1
X_2645_ VDD VSS _1001_ core.osr.next_result_w\[6\] _1009_ _0551_ VDD VSS sky130_fd_sc_hd__a21oi_1
XFILLER_10_29 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
X_2576_ VSS VDD _0026_ _0495_ VDD VSS sky130_fd_sc_hd__clkbuf_1
XANTENNA__2889__B1 VSS VDD _0482_ VDD VSS sky130_fd_sc_hd__diode_2
X_1527_ VDD VSS _1085_ _1081_ VDD VSS sky130_fd_sc_hd__buf_2
X_1458_ VSS VDD _1021_ core.osr.is_last_sample VDD VSS sky130_fd_sc_hd__clkbuf_2
X_3128_ VSS VDD clknet_2_3__leaf_clk_dig_dummy core.cnb.next_average_sum_w\[1\] net90
+ core.cnb.average_sum_r\[1\] VDD VSS sky130_fd_sc_hd__dfrtp_1
XFILLER_27_125 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_55_423 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XFILLER_55_445 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
X_3059_ VDD VSS _0946_ _0507_ _0945_ VDD VSS sky130_fd_sc_hd__or2_1
Xgenblk2\[2\].buf_p_rowonn VSS VDD pmatrix_rowon_core_n_buffered\[2\] core.pdc.rowon_out_n\[2\]
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
XFILLER_51_36 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XANTENNA__2042__B VSS VDD _1279_ VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__3173__CLK VSS VDD net61 VDD VSS sky130_fd_sc_hd__diode_2
Xgenblk1\[19\].buf_p_coln VSS VDD pmatrix_col_core_n_buffered\[19\] core.pdc.col_out_n\[19\]
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
XFILLER_18_103 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XFILLER_46_412 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XFILLER_46_434 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_41_150 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XFILLER_25_81 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XANTENNA__2583__A2 VSS VDD _1067_ VDD VSS sky130_fd_sc_hd__diode_2
X_2430_ VDD VSS _0426_ core.ndc.row_bottotop_n\[10\] VDD VSS sky130_fd_sc_hd__clkinv_2
XANTENNA__1791__B VSS VDD _1175_ VDD VSS sky130_fd_sc_hd__diode_2
X_2361_ VSS VDD _0377_ _0379_ core.osr.result_r\[16\] VDD VSS sky130_fd_sc_hd__nand2_1
X_2292_ VSS VDD _0314_ _0316_ _0317_ VDD VSS sky130_fd_sc_hd__nor2_1
XANTENNA__2099__A1 VSS VDD _0081_ VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_2_85 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XANTENNA__2099__B2 VSS VDD _1096_ VDD VSS sky130_fd_sc_hd__diode_2
Xgenblk1\[21\].buf_p_coln VSS VDD pmatrix_col_core_n_buffered\[21\] core.pdc.col_out_n\[21\]
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
XFILLER_52_437 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
X_2628_ VSS VDD core.osr.next_result_w\[6\] _0536_ _0535_ VDD VSS sky130_fd_sc_hd__nand2_1
X_2559_ VSS VDD _0023_ _0481_ VDD VSS sky130_fd_sc_hd__clkbuf_1
XFILLER_46_36 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_102_97 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XFILLER_11_50 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
XFILLER_2_1 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_93_337 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_46_253 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XFILLER_46_286 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
X_1930_ VSS VDD core.pdc.rowon_out_n\[0\] _1388_ _1040_ VDD VSS sky130_fd_sc_hd__nand2_1
X_1861_ VDD VSS _1346_ _1345_ VDD VSS sky130_fd_sc_hd__inv_2
XANTENNA__1786__B VSS VDD _1188_ VDD VSS sky130_fd_sc_hd__diode_2
Xinput22 VDD VSS net22 config_2_in[13] VDD VSS sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_52_90 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
Xinput11 VSS VDD net11 config_1_in[3] VDD VSS sky130_fd_sc_hd__clkbuf_1
XANTENNA__2005__B2 VSS VDD _0072_ VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__2005__A1 VSS VDD _1126_ VDD VSS sky130_fd_sc_hd__diode_2
Xgenblk1\[16\].buf_n_coln VDD VSS core.ndc.col_out_n\[16\] nmatrix_col_core_n_buffered\[16\]
+ VDD VSS sky130_fd_sc_hd__buf_6
X_1792_ VDD VSS _1295_ _1125_ _1240_ _1294_ _1279_ core.ndc.col_out\[28\] VDD VSS
+ sky130_fd_sc_hd__a221o_2
Xinput33 VDD VSS net33 config_2_in[9] VDD VSS sky130_fd_sc_hd__dlymetal6s2s_1
X_2413_ VSS VDD _0417_ _0420_ _1013_ VDD VSS sky130_fd_sc_hd__nand2_1
XFILLER_88_109 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
X_2344_ VDD VSS _0364_ core.osr.result_r\[14\] VDD VSS sky130_fd_sc_hd__inv_2
XFILLER_96_120 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
X_2275_ VSS VDD _0302_ _0300_ _0290_ _0294_ VDD VSS sky130_fd_sc_hd__and3_1
XFILLER_92_392 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_32_38 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XFILLER_57_13 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_48_518 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XFILLER_57_57 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XFILLER_73_67 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XFILLER_7_113 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XANTENNA__1994__A0 VSS VDD _1202_ VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_98_53 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_98_97 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
X_2060_ VDD VSS core.pdc.col_out_n\[15\] core.pdc.col_out\[15\] VDD VSS sky130_fd_sc_hd__clkinv_2
XANTENNA__1797__A VSS VDD core.ndc.col_out\[29\] VDD VSS sky130_fd_sc_hd__diode_2
X_2962_ VSS VDD _0854_ _0737_ _0734_ _0853_ VDD VSS sky130_fd_sc_hd__and3_1
X_1913_ VSS VDD core.pdc.rowon_out_n\[8\] _1379_ core.ndc.rowon_out_n\[15\] VDD VSS
+ sky130_fd_sc_hd__nand2_2
X_2893_ VSS VDD _0784_ _0786_ _0785_ VDD VSS sky130_fd_sc_hd__nand2_1
XFILLER_8_62 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
X_1844_ VSS VDD _1303_ _1326_ _1332_ VDD VSS sky130_fd_sc_hd__nor2_1
X_1775_ VSS VDD _1126_ _1231_ _1285_ VDD VSS sky130_fd_sc_hd__nor2_1
Xnmat nmatrix_row_core_n_buffered\[0\] nmatrix_row_core_n_buffered\[1\] nmatrix_row_core_n_buffered\[2\]
+ nmatrix_row_core_n_buffered\[3\] nmatrix_row_core_n_buffered\[4\] nmatrix_row_core_n_buffered\[5\]
+ nmatrix_row_core_n_buffered\[6\] nmatrix_row_core_n_buffered\[7\] nmatrix_row_core_n_buffered\[8\]
+ nmatrix_row_core_n_buffered\[9\] nmatrix_row_core_n_buffered\[10\] nmatrix_row_core_n_buffered\[11\]
+ nmatrix_row_core_n_buffered\[12\] nmatrix_row_core_n_buffered\[13\] nmatrix_row_core_n_buffered\[14\]
+ nmatrix_row_core_n_buffered\[15\] nmatrix_rowon_core_n_buffered\[0\] nmatrix_rowon_core_n_buffered\[1\]
+ nmatrix_rowon_core_n_buffered\[2\] nmatrix_rowon_core_n_buffered\[3\] nmatrix_rowon_core_n_buffered\[4\]
+ nmatrix_rowon_core_n_buffered\[5\] nmatrix_rowon_core_n_buffered\[6\] nmatrix_rowon_core_n_buffered\[7\]
+ nmatrix_rowon_core_n_buffered\[8\] nmatrix_rowon_core_n_buffered\[9\] nmatrix_rowon_core_n_buffered\[10\]
+ nmatrix_rowon_core_n_buffered\[11\] nmatrix_rowon_core_n_buffered\[12\] nmatrix_rowon_core_n_buffered\[13\]
+ nmatrix_rowon_core_n_buffered\[14\] nmatrix_rowon_core_n_buffered\[15\] core.ndc.rowoff_out_n\[0\]
+ core.ndc.rowoff_out_n\[1\] core.ndc.rowoff_out_n\[2\] core.ndc.rowoff_out_n\[3\]
+ core.ndc.rowoff_out_n\[4\] core.ndc.rowoff_out_n\[5\] core.ndc.rowoff_out_n\[6\]
+ core.ndc.rowoff_out_n\[7\] core.ndc.rowoff_out_n\[8\] core.ndc.rowoff_out_n\[9\]
+ core.ndc.rowoff_out_n\[10\] core.ndc.rowoff_out_n\[11\] core.ndc.rowoff_out_n\[12\]
+ core.ndc.rowoff_out_n\[13\] core.ndc.rowoff_out_n\[14\] core.ndc.rowoff_out_n\[15\]
+ vcm/vcm sample_nmatrix_cgen _0001_ nmatrix_col_core_n_buffered\[31\] nmatrix_col_core_n_buffered\[30\]
+ nmatrix_col_core_n_buffered\[29\] nmatrix_col_core_n_buffered\[28\] nmatrix_col_core_n_buffered\[27\]
+ nmatrix_col_core_n_buffered\[26\] nmatrix_col_core_n_buffered\[25\] nmatrix_col_core_n_buffered\[24\]
+ nmatrix_col_core_n_buffered\[23\] nmatrix_col_core_n_buffered\[22\] nmatrix_col_core_n_buffered\[21\]
+ nmatrix_col_core_n_buffered\[20\] nmatrix_col_core_n_buffered\[19\] nmatrix_col_core_n_buffered\[18\]
+ nmatrix_col_core_n_buffered\[17\] nmatrix_col_core_n_buffered\[16\] nmatrix_col_core_n_buffered\[15\]
+ nmatrix_col_core_n_buffered\[14\] nmatrix_col_core_n_buffered\[13\] nmatrix_col_core_n_buffered\[12\]
+ nmatrix_col_core_n_buffered\[11\] nmatrix_col_core_n_buffered\[10\] nmatrix_col_core_n_buffered\[9\]
+ nmatrix_col_core_n_buffered\[8\] nmatrix_col_core_n_buffered\[7\] nmatrix_col_core_n_buffered\[6\]
+ nmatrix_col_core_n_buffered\[5\] nmatrix_col_core_n_buffered\[4\] nmatrix_col_core_n_buffered\[3\]
+ nmatrix_col_core_n_buffered\[2\] nmatrix_col_core_n_buffered\[1\] nmatrix_col_core_n_buffered\[0\]
+ core.cnb.pswitch_out\[2\] core.cnb.pswitch_out\[1\] core.cnb.pswitch_out\[0\] net96
+ nmat_sample_switch_buffered nmat_sample_switch_n_buffered inn_analog core.ndc.col_out\[0\]
+ core.ndc.col_out\[1\] core.ndc.col_out\[2\] core.ndc.col_out\[3\] core.ndc.col_out\[4\]
+ core.ndc.col_out\[5\] core.ndc.col_out\[6\] core.ndc.col_out\[7\] core.ndc.col_out\[8\]
+ core.ndc.col_out\[9\] core.ndc.col_out\[10\] core.ndc.col_out\[11\] core.ndc.col_out\[12\]
+ core.ndc.col_out\[13\] core.ndc.col_out\[14\] core.ndc.col_out\[15\] core.ndc.col_out\[16\]
+ core.ndc.col_out\[17\] core.ndc.col_out\[18\] core.ndc.col_out\[19\] core.ndc.col_out\[20\]
+ core.ndc.col_out\[21\] core.ndc.col_out\[22\] core.ndc.col_out\[23\] core.ndc.col_out\[24\]
+ core.ndc.col_out\[25\] core.ndc.col_out\[26\] core.ndc.col_out\[27\] core.ndc.col_out\[28\]
+ core.ndc.col_out\[29\] core.ndc.col_out\[30\] core.ndc.col_out\[31\] VDD VSS ctop_nmatrix_analog
+ adc_array_matrix_12bit
X_2327_ VSS VDD core.osr.next_result_w\[11\] _0349_ VDD VSS sky130_fd_sc_hd__clkbuf_1
X_2258_ VSS VDD _0285_ _0271_ _0287_ _0286_ VDD VSS sky130_fd_sc_hd__nand3_1
XFILLER_84_123 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_84_145 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
X_2189_ VDD VSS _0226_ core.cnb.average_sum_r\[2\] VDD VSS sky130_fd_sc_hd__inv_2
XANTENNA__1500__A VSS VDD _1057_ VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1976__A0 VSS VDD _1197_ VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_4_105 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XFILLER_108_63 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XANTENNA_input17_A VSS VDD config_1_in[9] VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_84_99 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
XFILLER_90_137 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XANTENNA__2506__A VSS VDD _0208_ VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__3107__CLK VSS VDD clknet_2_3__leaf_clk_dig_dummy VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_83_9 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XANTENNA__1719__B1 VSS VDD _1075_ VDD VSS sky130_fd_sc_hd__diode_2
X_1560_ VDD VSS _1114_ _1044_ VDD VSS sky130_fd_sc_hd__buf_2
Xclkbuf_2_2__f_clk_dig_dummy VSS VDD clknet_0_clk_dig_dummy clknet_2_2__leaf_clk_dig_dummy
+ VDD VSS sky130_fd_sc_hd__clkbuf_16
X_1491_ VSS VDD _1050_ _1051_ VDD VSS sky130_fd_sc_hd__clkbuf_2
X_3161_ VSS VDD net62 core.osr.next_result_w\[1\] net74 core.osr.result_r\[1\] VDD
+ VSS sky130_fd_sc_hd__dfrtp_1
X_2112_ VSS VDD _0165_ _0164_ _0163_ _0162_ VDD VSS sky130_fd_sc_hd__and3_1
X_3092_ VSS VDD _0976_ _0977_ _0689_ VDD VSS sky130_fd_sc_hd__nand2_1
XFILLER_54_329 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
X_2043_ VSS VDD _1403_ _0124_ _1163_ VDD VSS sky130_fd_sc_hd__nand2_1
XFILLER_50_513 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
X_2945_ VSS VDD _0831_ _0837_ _0836_ VDD VSS sky130_fd_sc_hd__nand2_1
XANTENNA__1958__B1 VSS VDD _1047_ VDD VSS sky130_fd_sc_hd__diode_2
X_2876_ VSS VDD _0769_ _0768_ _0764_ _0770_ VDD VSS sky130_fd_sc_hd__nor3_1
X_1827_ VSS VDD _1317_ _1318_ core.cnb.data_register_r\[10\] VDD VSS sky130_fd_sc_hd__nand2_1
X_1758_ VDD VSS _1273_ _1125_ _1217_ _1121_ _1193_ core.ndc.col_out\[22\] VDD VSS
+ sky130_fd_sc_hd__a221o_2
X_1689_ VSS VDD _1206_ _1103_ _1225_ _1199_ VDD VSS sky130_fd_sc_hd__a21oi_2
XANTENNA_nmat_col[8] VSS VDD core.ndc.col_out\[8\] VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA_input9_A VSS VDD config_1_in[1] VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_57_123 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XANTENNA__2045__B VSS VDD _0125_ VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_119_62 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XANTENNA__2996__A VSS VDD _1113_ VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_91_435 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
Xgenblk1\[26\].buf_p_coln VSS VDD pmatrix_col_core_n_buffered\[26\] core.pdc.col_out_n\[26\]
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
X_2730_ VSS VDD _0530_ _0626_ _0627_ VDD VSS sky130_fd_sc_hd__nor2_1
X_2661_ VSS VDD core.osr.next_result_w\[6\] _0540_ _0565_ _0528_ VDD VSS sky130_fd_sc_hd__o21ai_1
X_1612_ VDD VSS _1154_ core.ndc.col_out\[6\] _1152_ _1159_ _1155_ _1157_ VDD VSS sky130_fd_sc_hd__a221o_4
XFILLER_5_30 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
X_2592_ VDD VSS _0507_ core.cnb.data_register_r\[9\] VDD VSS sky130_fd_sc_hd__inv_2
X_1543_ VSS VDD _1099_ _1067_ _1054_ _1098_ VDD VSS sky130_fd_sc_hd__mux2_1
XFILLER_5_96 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
X_1474_ VDD VSS _1034_ _1033_ VDD VSS sky130_fd_sc_hd__buf_2
XFILLER_39_145 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
X_3144_ VSS VDD net56 _0034_ net68 net38 VDD VSS sky130_fd_sc_hd__dfrtp_1
X_3075_ VDD VSS _0833_ _0831_ _0918_ _0961_ VDD VSS sky130_fd_sc_hd__a21oi_1
XFILLER_54_137 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
X_2026_ VSS VDD _1064_ _0111_ _0110_ _1224_ core.pdc.col_out_n\[11\] _0112_ VDD VSS
+ sky130_fd_sc_hd__o221a_1
XFILLER_90_490 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XANTENNA__1985__A VSS VDD _0081_ VDD VSS sky130_fd_sc_hd__diode_2
X_2928_ VSS VDD _0819_ _0809_ _0806_ _0820_ VDD VSS sky130_fd_sc_hd__nor3_1
XANTENNA_genblk1\[9\].buf_n_coln_A VSS VDD core.ndc.col_out_n\[9\] VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_40_49 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
X_2859_ VSS VDD core.cnb.pswitch_out\[0\] _0753_ _0754_ VDD VSS sky130_fd_sc_hd__nor2_1
XFILLER_108_128 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_116_150 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
XFILLER_49_47 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XFILLER_105_86 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XFILLER_53_192 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XFILLER_53_181 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XANTENNA__2056__A VSS VDD _1242_ VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_2_0__f_clk_dig_dummy_A VSS VDD clknet_0_clk_dig_dummy VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_46_9 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XFILLER_122_153 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XANTENNA_genblk2\[14\].buf_p_rown_A VSS VDD core.pdc.row_out_n\[14\] VDD VSS sky130_fd_sc_hd__diode_2
Xinput9 VSS VDD net9 config_1_in[1] VDD VSS sky130_fd_sc_hd__clkbuf_1
XFILLER_49_487 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
X_2713_ VSS VDD _0610_ _0540_ _0612_ _0611_ VDD VSS sky130_fd_sc_hd__nand3_1
X_2644_ VSS VDD core.osr.next_result_w\[8\] _0550_ _1002_ VDD VSS sky130_fd_sc_hd__nand2_1
XFILLER_65_1 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
X_2575_ VSS VDD _0495_ core.cnb.result_out\[4\] _0480_ _0494_ VDD VSS sky130_fd_sc_hd__mux2_1
X_1526_ VDD VSS _1084_ _1083_ VDD VSS sky130_fd_sc_hd__inv_2
XANTENNA__2889__B2 VSS VDD _0758_ VDD VSS sky130_fd_sc_hd__diode_2
X_1457_ VDD VSS _1021_ _1020_ VDD VSS sky130_fd_sc_hd__inv_2
X_3127_ VSS VDD clknet_2_3__leaf_clk_dig_dummy core.cnb.next_average_sum_w\[0\] net90
+ core.cnb.average_sum_r\[0\] VDD VSS sky130_fd_sc_hd__dfrtp_1
XFILLER_27_137 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
Xgenblk1\[23\].buf_n_coln VSS VDD nmatrix_col_core_n_buffered\[23\] core.ndc.col_out_n\[23\]
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
XFILLER_55_479 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
X_3058_ VSS VDD _0945_ _0799_ _0693_ _0472_ VDD VSS sky130_fd_sc_hd__mux2_1
X_2009_ VDD VSS _0099_ _0100_ VDD VSS sky130_fd_sc_hd__clkinv_2
XFILLER_136_7 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_4_5 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_116_41 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XANTENNA__1552__A1 VSS VDD _1091_ VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1552__B2 VSS VDD _1102_ VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_116_85 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
XFILLER_18_137 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XFILLER_46_479 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
X_2360_ VDD VSS _0378_ core.osr.result_r\[16\] _0377_ VDD VSS sky130_fd_sc_hd__or2_1
XANTENNA__1543__A1 VSS VDD _1067_ VDD VSS sky130_fd_sc_hd__diode_2
X_2291_ VDD VSS _0316_ _0315_ VDD VSS sky130_fd_sc_hd__inv_2
XANTENNA__2099__A2 VSS VDD _1173_ VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_2_97 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
X_2627_ VSS VDD _1002_ _0535_ VDD VSS sky130_fd_sc_hd__clkbuf_2
X_2558_ VSS VDD _0481_ core.cnb.result_out\[1\] _0480_ _0479_ VDD VSS sky130_fd_sc_hd__mux2_1
X_2489_ VSS VDD net64 _0435_ core.osr.data_valid_r VDD VSS sky130_fd_sc_hd__nand2_1
X_1509_ VSS VDD _1067_ _1046_ _1066_ VDD VSS sky130_fd_sc_hd__nor2_4
XANTENNA__2318__B VSS VDD core.cnb.result_out\[11\] VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__3140__CLK VSS VDD clknet_2_0__leaf_clk_dig_dummy VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__2988__B VSS VDD _1113_ VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1525__A1 VSS VDD _1076_ VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_93_349 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
X_1860_ VDD VSS core.cnb.data_register_r\[8\] _1304_ core.cnb.data_register_r\[11\]
+ net14 _1345_ VDD VSS sky130_fd_sc_hd__or4_1
Xinput12 VSS VDD net12 config_1_in[4] VDD VSS sky130_fd_sc_hd__clkbuf_1
X_1791_ VSS VDD _1272_ _1175_ _1295_ VDD VSS sky130_fd_sc_hd__nor2_1
Xinput23 VDD VSS net23 config_2_in[14] VDD VSS sky130_fd_sc_hd__dlymetal6s2s_1
Xinput34 VSS VDD net34 rst_n VDD VSS sky130_fd_sc_hd__clkbuf_1
X_2412_ VSS VDD _1013_ _0417_ _0419_ VDD VSS sky130_fd_sc_hd__nor2_1
X_2343_ VDD VSS core.osr.next_result_w\[13\] _0363_ VDD VSS sky130_fd_sc_hd__inv_2
XANTENNA__3103__RESET_B VSS VDD net85 VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_96_132 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
X_2274_ VDD VSS _0290_ _0294_ _0300_ _0301_ VDD VSS sky130_fd_sc_hd__a21oi_1
XFILLER_78_891 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
X_1989_ VSS VDD _0086_ _0085_ _0082_ _0080_ VDD VSS sky130_fd_sc_hd__and3_1
XFILLER_57_25 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XFILLER_69_891 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XFILLER_87_165 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XFILLER_87_176 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XFILLER_113_64 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XFILLER_73_24 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XANTENNA__1691__B1 VSS VDD _1035_ VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__2064__A VSS VDD _0125_ VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_132_1 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XANTENNA__1994__A1 VSS VDD _1242_ VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_7_136 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XANTENNA_genblk2\[1\].buf_p_rowonn_A VSS VDD core.pdc.rowon_out_n\[1\] VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_98_65 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XFILLER_93_113 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XANTENNA_genblk2\[2\].buf_n_rowonn_A VSS VDD core.ndc.rowon_out_n\[2\] VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__3186__CLK VSS VDD clknet_2_1__leaf_clk_dig_dummy VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_75_883 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XANTENNA__1682__B1 VSS VDD _1137_ VDD VSS sky130_fd_sc_hd__diode_2
X_2961_ VDD VSS _0853_ _0742_ VDD VSS sky130_fd_sc_hd__inv_2
X_1912_ VSS VDD _1024_ core.ndc.rowon_out_n\[15\] _1331_ VDD VSS sky130_fd_sc_hd__nand2_1
XFILLER_8_41 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
X_2892_ VSS VDD _0666_ _0785_ _0702_ VDD VSS sky130_fd_sc_hd__nand2_1
X_1843_ VDD VSS _1324_ _1331_ VDD VSS sky130_fd_sc_hd__clkinv_2
X_1774_ VDD VSS _1284_ _1095_ VDD VSS sky130_fd_sc_hd__buf_2
Xgenblk2\[11\].buf_n_rowonn VSS VDD nmatrix_rowon_core_n_buffered\[11\] core.ndc.rowon_out_n\[11\]
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
X_2326_ VDD VSS _0349_ _0347_ _0348_ VDD VSS sky130_fd_sc_hd__and2_1
X_2257_ VSS VDD _0284_ _0286_ _0283_ VDD VSS sky130_fd_sc_hd__nand2_1
XFILLER_84_135 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XFILLER_66_883 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
X_2188_ VSS VDD core.cnb.next_average_sum_w\[1\] _0225_ VDD VSS sky130_fd_sc_hd__clkbuf_1
XFILLER_92_190 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
XANTENNA__1976__A1 VSS VDD _1208_ VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA_genblk2\[7\].buf_n_rown_A VSS VDD core.ndc.row_out_n\[7\] VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA_pmat_rowoff_n[0] VSS VDD core.pdc.rowoff_out_n\[0\] VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_68_35 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_48_305 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XFILLER_75_113 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_124_85 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XANTENNA__1664__B1 VSS VDD _1035_ VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_56_393 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XANTENNA__1719__A1 VSS VDD _1064_ VDD VSS sky130_fd_sc_hd__diode_2
X_1490_ VDD VSS core.cnb.data_register_r\[7\] _1050_ VDD VSS sky130_fd_sc_hd__clkinv_2
X_3160_ VSS VDD net63 core.osr.next_result_w\[0\] net81 core.osr.result_r\[0\] VDD
+ VSS sky130_fd_sc_hd__dfrtp_1
X_3091_ VSS VDD _0975_ _0976_ _0691_ VDD VSS sky130_fd_sc_hd__nand2_1
X_2111_ VSS VDD _1413_ _0164_ _1101_ VDD VSS sky130_fd_sc_hd__nand2_1
X_2042_ VSS VDD _0089_ _0123_ _1279_ VDD VSS sky130_fd_sc_hd__nand2_1
Xgenblk1\[28\].buf_n_coln VDD VSS core.ndc.col_out_n\[28\] nmatrix_col_core_n_buffered\[28\]
+ VDD VSS sky130_fd_sc_hd__buf_6
XFILLER_50_525 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
Xobstruction1 VSS VDD scboundary
X_2944_ VSS VDD _0834_ _0836_ _0835_ VDD VSS sky130_fd_sc_hd__nand2_1
XANTENNA__1958__A1 VSS VDD _1057_ VDD VSS sky130_fd_sc_hd__diode_2
X_2875_ VSS VDD _0685_ _0695_ _0769_ _0693_ VDD VSS sky130_fd_sc_hd__nand3_1
X_1826_ VSS VDD core.cnb.data_register_r\[9\] _1071_ _1317_ VDD VSS sky130_fd_sc_hd__nor2_1
X_1757_ VSS VDD _1272_ _1225_ _1273_ VDD VSS sky130_fd_sc_hd__nor2_1
X_1688_ VSS VDD _1074_ _1224_ VDD VSS sky130_fd_sc_hd__clkbuf_2
XANTENNA_nmat_col[7] VSS VDD core.ndc.col_out\[7\] VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_89_249 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
XFILLER_38_38 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
X_2309_ VSS VDD _0326_ _0333_ _0332_ VDD VSS sky130_fd_sc_hd__nand2_1
XFILLER_85_422 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XANTENNA__2438__A2 VSS VDD _1340_ VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1511__A VSS VDD _1037_ VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__2610__A2 VSS VDD core.osr.next_result_w\[3\] VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_119_41 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
Xgenblk1\[30\].buf_n_coln VSS VDD nmatrix_col_core_n_buffered\[30\] core.ndc.col_out_n\[30\]
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
XANTENNA__2061__B VSS VDD _1093_ VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_119_96 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_135_40 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_48_102 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_48_135 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XFILLER_95_44 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_95_77 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XFILLER_91_414 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XFILLER_56_190 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
XANTENNA__2062__B1 VSS VDD _1075_ VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__2252__A VSS VDD core.cnb.result_out\[5\] VDD VSS sky130_fd_sc_hd__diode_2
X_2660_ VSS VDD _0561_ _0041_ _0564_ VDD VSS sky130_fd_sc_hd__nand2_1
X_1611_ VDD VSS _1159_ _1158_ VDD VSS sky130_fd_sc_hd__inv_2
X_2591_ VSS VDD _0030_ _0506_ VDD VSS sky130_fd_sc_hd__clkbuf_1
X_1542_ VDD VSS _1098_ _1097_ VDD VSS sky130_fd_sc_hd__inv_2
X_1473_ VDD VSS _1032_ _1033_ VDD VSS sky130_fd_sc_hd__clkinv_2
XFILLER_10_1 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
X_3143_ VSS VDD clknet_2_0__leaf_clk_dig_dummy _0033_ net79 core.cnb.result_out\[11\]
+ VDD VSS sky130_fd_sc_hd__dfrtp_2
X_3074_ VSS VDD _0960_ _0959_ _0958_ _0918_ _1312_ VDD VSS sky130_fd_sc_hd__a211o_1
X_2025_ VSS VDD _0101_ _0112_ _1093_ VDD VSS sky130_fd_sc_hd__nand2_1
X_2927_ VSS VDD _0815_ _0726_ _0819_ _0818_ VDD VSS sky130_fd_sc_hd__nand3_1
XANTENNA__1985__B VSS VDD _1275_ VDD VSS sky130_fd_sc_hd__diode_2
Xgenblk2\[8\].buf_n_rowonn VSS VDD nmatrix_rowon_core_n_buffered\[8\] core.ndc.rowon_out_n\[8\]
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
X_2858_ VSS VDD _0727_ _0752_ _0753_ VDD VSS sky130_fd_sc_hd__nor2_1
Xgenblk2\[1\].buf_p_rown VSS VDD pmatrix_row_core_n_buffered\[1\] core.pdc.row_out_n\[1\]
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
X_1809_ VSS VDD net14 _1301_ _1302_ VDD VSS sky130_fd_sc_hd__nor2_1
X_2789_ VDD VSS _0685_ _0684_ VDD VSS sky130_fd_sc_hd__inv_2
XANTENNA__1506__A VSS VDD _1034_ VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1619__A0 VSS VDD _1161_ VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1416__A VSS VDD core.cnb.data_register_r\[1\] VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_49_477 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
X_2712_ VDD VSS _0348_ _0347_ _0528_ _0611_ VDD VSS sky130_fd_sc_hd__a21o_1
X_2643_ VSS VDD _0039_ _0548_ _0540_ _0547_ _0549_ VDD VSS sky130_fd_sc_hd__a31o_1
X_2574_ VSS VDD _0492_ _0494_ _0493_ VDD VSS sky130_fd_sc_hd__nand2_1
X_1525_ VSS VDD _1083_ _1076_ _1078_ _1080_ _1082_ VDD VSS sky130_fd_sc_hd__o211a_1
X_1456_ VSS VDD _1019_ _1020_ _0983_ VDD VSS sky130_fd_sc_hd__nor2_2
X_3126_ VSS VDD clknet_2_2__leaf_clk_dig_dummy core.cnb.next_average_counter_w\[4\]
+ net89 core.cnb.average_counter_r\[4\] VDD VSS sky130_fd_sc_hd__dfrtp_1
XFILLER_27_149 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
X_3057_ VSS VDD _0942_ _0944_ _0902_ VDD VSS sky130_fd_sc_hd__nand2_1
X_2008_ VSS VDD _1131_ _0098_ _0099_ VDD VSS sky130_fd_sc_hd__nor2_1
XFILLER_50_141 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XANTENNA__2026__B1 VSS VDD _1064_ VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1552__A2 VSS VDD _1096_ VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_76_46 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_132_85 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XANTENNA__2017__A0 VSS VDD _1137_ VDD VSS sky130_fd_sc_hd__diode_2
X_2290_ VSS VDD core.osr.result_r\[9\] _0315_ core.cnb.result_out\[9\] VDD VSS sky130_fd_sc_hd__nand2_1
XFILLER_110_146 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XFILLER_32_141 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
XANTENNA__2143__C VSS VDD core.cnb.sampled_avg_control_r\[2\] VDD VSS sky130_fd_sc_hd__diode_2
X_2626_ VSS VDD core.osr.next_result_w\[8\] _0534_ _0533_ VDD VSS sky130_fd_sc_hd__nand2_1
XANTENNA__2440__A VSS VDD _1342_ VDD VSS sky130_fd_sc_hd__diode_2
X_2557_ VSS VDD _0438_ _0480_ VDD VSS sky130_fd_sc_hd__clkbuf_2
X_2488_ VDD VSS core.cnb.next_conv_finished_w _0434_ VDD VSS sky130_fd_sc_hd__inv_2
X_1508_ VDD VSS _1066_ _1065_ VDD VSS sky130_fd_sc_hd__inv_2
X_1439_ VDD VSS _1003_ _1002_ VDD VSS sky130_fd_sc_hd__inv_2
XFILLER_87_347 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
X_3109_ VSS VDD clknet_2_3__leaf_clk_dig_dummy _0009_ net90 core.cnb.shift_register_r\[7\]
+ VDD VSS sky130_fd_sc_hd__dfrtp_1
XFILLER_15_108 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XFILLER_62_59 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_51_461 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_51_483 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XANTENNA__2334__B VSS VDD _0241_ VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_127_41 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XANTENNA__1525__A2 VSS VDD _1078_ VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_14_141 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
Xinput13 VSS VDD net13 config_1_in[5] VDD VSS sky130_fd_sc_hd__clkbuf_1
X_1790_ VDD VSS _1294_ _1109_ VDD VSS sky130_fd_sc_hd__inv_2
Xinput24 VSS VDD config_2_in[15] net24 VDD VSS sky130_fd_sc_hd__clkbuf_2
Xinput35 VSS VDD net35 start_conversion_in VDD VSS sky130_fd_sc_hd__clkbuf_1
X_2411_ VDD VSS _0418_ core.osr.next_sample_count_w\[6\] VDD VSS sky130_fd_sc_hd__clkinv_2
X_2342_ VSS VDD _0360_ _0363_ _0362_ VDD VSS sky130_fd_sc_hd__nand2_1
XFILLER_96_144 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
X_2273_ VDD VSS _0300_ _0299_ VDD VSS sky130_fd_sc_hd__inv_2
XANTENNA__1604__A VSS VDD _1092_ VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_52_269 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
X_1988_ VSS VDD _0084_ _0085_ _1235_ VDD VSS sky130_fd_sc_hd__nand2_1
XANTENNA__2170__A VSS VDD _0210_ VDD VSS sky130_fd_sc_hd__diode_2
X_2609_ VSS VDD _1009_ _1018_ _0520_ VDD VSS sky130_fd_sc_hd__nor2_1
XANTENNA_nmat_col[29] VSS VDD core.ndc.col_out\[29\] VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1514__A VSS VDD net15 VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_113_43 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XANTENNA__1691__A1 VSS VDD _1224_ VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_113_98 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XFILLER_11_100 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XANTENNA__1424__A VSS VDD _0983_ VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1682__A1 VSS VDD _1078_ VDD VSS sky130_fd_sc_hd__diode_2
X_2960_ VSS VDD _0850_ _0852_ _0851_ VDD VSS sky130_fd_sc_hd__nand2_1
X_1911_ VSS VDD _1378_ _1379_ _1369_ VDD VSS sky130_fd_sc_hd__nand2_1
X_2891_ VSS VDD _0784_ _0783_ _0470_ VDD VSS sky130_fd_sc_hd__nand2_2
X_1842_ VSS VDD _1325_ _1328_ _1330_ core.pdc.row_out_n\[4\] VDD VSS sky130_fd_sc_hd__o21a_1
XANTENNA__3086__A VSS VDD _1342_ VDD VSS sky130_fd_sc_hd__diode_2
X_1773_ VDD VSS core.ndc.col_out_n\[24\] core.ndc.col_out\[24\] VDD VSS sky130_fd_sc_hd__clkinv_2
Xgenblk2\[6\].buf_p_rown VSS VDD pmatrix_row_core_n_buffered\[6\] core.pdc.row_out_n\[6\]
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
XFILLER_69_122 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
X_2325_ VDD VSS _0348_ core.cnb.result_out\[11\] _0255_ VDD VSS sky130_fd_sc_hd__or2_1
XANTENNA__3130__CLK VSS VDD clknet_2_3__leaf_clk_dig_dummy VDD VSS sky130_fd_sc_hd__diode_2
X_2256_ VDD VSS _0285_ _0283_ _0284_ VDD VSS sky130_fd_sc_hd__or2_1
XFILLER_27_29 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
X_2187_ VSS VDD _0225_ _0224_ _0223_ _0209_ VDD VSS sky130_fd_sc_hd__and3_1
XFILLER_53_501 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XANTENNA__1988__B VSS VDD _1235_ VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__2165__A VSS VDD _0208_ VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_43_39 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XFILLER_68_25 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XFILLER_124_64 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
XANTENNA_nmat_sample VSS VDD sample_nmatrix_cgen VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_75_125 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XANTENNA__1664__A1 VSS VDD _1075_ VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_129_105 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
Xgenblk1\[1\].buf_p_coln VSS VDD pmatrix_col_core_n_buffered\[1\] core.pdc.col_out_n\[1\]
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
X_3090_ VSS VDD _0972_ _0975_ _0974_ VDD VSS sky130_fd_sc_hd__nand2_1
X_2110_ VSS VDD _1411_ _0163_ _1177_ VDD VSS sky130_fd_sc_hd__nand2_1
XFILLER_12_5 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
X_2041_ VDD VSS core.pdc.col_out_n\[13\] core.pdc.col_out\[13\] VDD VSS sky130_fd_sc_hd__clkinv_2
X_2943_ VDD VSS _0835_ _0829_ VDD VSS sky130_fd_sc_hd__inv_2
Xobstruction2 VSS VDD scboundary
X_2874_ VSS VDD _0662_ _0664_ _0768_ _0767_ VDD VSS sky130_fd_sc_hd__o21ai_1
XFILLER_88_1 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
X_1825_ VDD VSS core.pdc.rowoff_out_n\[8\] _1316_ VDD VSS sky130_fd_sc_hd__buf_2
X_1756_ VSS VDD _1110_ _1272_ VDD VSS sky130_fd_sc_hd__clkbuf_2
X_1687_ VDD VSS core.ndc.col_out_n\[11\] core.ndc.col_out\[11\] VDD VSS sky130_fd_sc_hd__clkinv_2
XANTENNA__1591__B1 VSS VDD _1088_ VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA_nmat_col[6] VSS VDD core.ndc.col_out\[6\] VDD VSS sky130_fd_sc_hd__diode_2
X_2308_ VDD VSS _0332_ _0330_ VDD VSS sky130_fd_sc_hd__inv_2
X_2239_ VDD VSS _0251_ core.cnb.result_out\[3\] _0269_ _0270_ VDD VSS sky130_fd_sc_hd__a21o_1
XFILLER_53_342 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XFILLER_54_16 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XANTENNA__2623__A VSS VDD _0394_ VDD VSS sky130_fd_sc_hd__diode_2
Xgenblk2\[3\].buf_n_rown VSS VDD nmatrix_row_core_n_buffered\[3\] core.ndc.row_out_n\[3\]
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
XFILLER_134_141 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_119_75 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_79_35 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_102_3 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_79_57 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_135_52 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XFILLER_48_114 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XANTENNA_input22_A VSS VDD config_2_in[13] VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_91_404 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
XFILLER_91_426 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
XFILLER_28_94 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_56_180 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
XANTENNA__2062__A1 VSS VDD _1064_ VDD VSS sky130_fd_sc_hd__diode_2
X_1610_ VDD VSS _1158_ _1073_ _1119_ VDD VSS sky130_fd_sc_hd__or2_1
X_2590_ VSS VDD _0506_ core.cnb.result_out\[8\] _0480_ _0505_ VDD VSS sky130_fd_sc_hd__mux2_1
X_1541_ VSS VDD _1047_ _1097_ _1057_ VDD VSS sky130_fd_sc_hd__nand2_1
X_1472_ VSS VDD core.cnb.data_register_r\[8\] _1032_ net15 VDD VSS sky130_fd_sc_hd__nor2_2
X_3142_ VSS VDD clknet_2_1__leaf_clk_dig_dummy _0032_ net81 core.cnb.result_out\[10\]
+ VDD VSS sky130_fd_sc_hd__dfrtp_1
X_3073_ VDD VSS _0958_ _0831_ _0856_ _0959_ VDD VSS sky130_fd_sc_hd__a21oi_1
XANTENNA__2427__B VSS VDD core.pdc.rowoff_out_n\[0\] VDD VSS sky130_fd_sc_hd__diode_2
X_2024_ VDD VSS _0083_ _1409_ _1208_ _0111_ VDD VSS sky130_fd_sc_hd__a21oi_1
XFILLER_50_389 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
X_2926_ VSS VDD _0649_ _0817_ _0818_ _0724_ VDD VSS sky130_fd_sc_hd__nand3_2
X_2857_ VSS VDD _0743_ _0745_ _0752_ _0751_ VDD VSS sky130_fd_sc_hd__nand3_1
X_1808_ VDD VSS _1301_ core.cnb.data_register_r\[11\] VDD VSS sky130_fd_sc_hd__inv_2
X_2788_ VSS VDD _0680_ _0683_ _0684_ VDD VSS sky130_fd_sc_hd__nor2_1
X_1739_ VDD VSS core.ndc.col_out\[18\] core.ndc.col_out_n\[18\] VDD VSS sky130_fd_sc_hd__inv_2
XFILLER_49_27 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XANTENNA__1522__A VSS VDD _1079_ VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_65_59 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_121_76 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XFILLER_14_63 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XFILLER_14_41 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XANTENNA__2044__A1 VSS VDD _1161_ VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__2072__B VSS VDD _1275_ VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1555__B1 VSS VDD _1088_ VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_36_106 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_55_81 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
X_2711_ VSS VDD _0607_ _0610_ _0609_ VDD VSS sky130_fd_sc_hd__nand2_1
X_2642_ VDD VSS _0393_ _0542_ core.osr.next_result_w\[1\] _0549_ net49 VDD VSS sky130_fd_sc_hd__a22o_1
X_2573_ VSS VDD _0489_ _0493_ _1200_ VDD VSS sky130_fd_sc_hd__nand2_1
XANTENNA__1607__A VSS VDD _1101_ VDD VSS sky130_fd_sc_hd__diode_2
X_1524_ VDD VSS _1081_ _1082_ VDD VSS sky130_fd_sc_hd__clkinv_2
X_1455_ VDD VSS _1019_ _1018_ VDD VSS sky130_fd_sc_hd__inv_2
X_3125_ VSS VDD clknet_2_3__leaf_clk_dig_dummy core.cnb.next_average_counter_w\[3\]
+ net89 core.cnb.average_counter_r\[3\] VDD VSS sky130_fd_sc_hd__dfrtp_1
X_3056_ VSS VDD _0689_ _0943_ _0058_ _1312_ VDD VSS sky130_fd_sc_hd__o21ai_1
XFILLER_35_18 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
X_2007_ VSS VDD _1389_ _1229_ _1161_ _0098_ VDD VSS sky130_fd_sc_hd__mux2_2
XANTENNA__2026__A1 VSS VDD _1224_ VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_50_186 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
X_2909_ VSS VDD _0798_ _0801_ _0800_ VDD VSS sky130_fd_sc_hd__nand2_1
XANTENNA__1517__A VSS VDD _1074_ VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1537__B1 VSS VDD _1075_ VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_104_111 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XANTENNA_fanout72_A VSS VDD net73 VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_46_404 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
XFILLER_26_150 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
XFILLER_92_68 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XFILLER_41_142 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XANTENNA__2017__A1 VSS VDD _1133_ VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_110_114 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_24_109 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XANTENNA_genblk2\[10\].buf_p_rown_A VSS VDD core.pdc.row_out_n\[10\] VDD VSS sky130_fd_sc_hd__diode_2
X_2625_ VSS VDD _1000_ _0533_ VDD VSS sky130_fd_sc_hd__clkbuf_2
X_2556_ VSS VDD _0477_ _0479_ _0478_ VDD VSS sky130_fd_sc_hd__nand2_1
X_2487_ VSS VDD _0220_ _0434_ core.cnb.is_holding_result_w VDD VSS sky130_fd_sc_hd__nand2_1
X_1507_ VSS VDD core.cnb.data_register_r\[4\] _1065_ _1044_ VDD VSS sky130_fd_sc_hd__nor2_2
X_1438_ VSS VDD _1000_ _1002_ _0989_ VDD VSS sky130_fd_sc_hd__nor2_2
XANTENNA__2168__A VSS VDD _0210_ VDD VSS sky130_fd_sc_hd__diode_2
X_3108_ VSS VDD clknet_2_3__leaf_clk_dig_dummy _0008_ net90 core.cnb.shift_register_r\[6\]
+ VDD VSS sky130_fd_sc_hd__dfrtp_1
X_3039_ VSS VDD _0856_ _0927_ _0924_ VDD VSS sky130_fd_sc_hd__nand2_1
XFILLER_51_473 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XFILLER_102_89 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XFILLER_127_53 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XFILLER_87_57 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
Xgenblk1\[6\].buf_p_coln VSS VDD pmatrix_col_core_n_buffered\[6\] core.pdc.col_out_n\[6\]
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
XANTENNA__2078__A VSS VDD _0065_ VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_36_61 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
XANTENNA__1710__A VSS VDD _1117_ VDD VSS sky130_fd_sc_hd__diode_2
Xinput14 VDD VSS net14 config_1_in[6] VDD VSS sky130_fd_sc_hd__buf_2
Xinput25 VSS VDD net25 config_2_in[1] VDD VSS sky130_fd_sc_hd__clkbuf_1
X_2410_ VSS VDD _1021_ _0417_ _0416_ _0418_ VDD VSS sky130_fd_sc_hd__or3b_1
X_2341_ VSS VDD _0355_ _0362_ _0361_ VDD VSS sky130_fd_sc_hd__nand2_1
X_2272_ VSS VDD _0297_ _0299_ _0298_ VDD VSS sky130_fd_sc_hd__and2b_1
XANTENNA__3091__B VSS VDD _0691_ VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__3183__RESET_B VSS VDD net86 VDD VSS sky130_fd_sc_hd__diode_2
X_1987_ VSS VDD _0084_ _1036_ _1053_ _1390_ _0083_ VDD VSS sky130_fd_sc_hd__a31o_1
Xgenblk2\[8\].buf_n_rown VSS VDD nmatrix_row_core_n_buffered\[8\] core.ndc.row_out_n\[8\]
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
X_2608_ VSS VDD _0518_ _0519_ VDD VSS sky130_fd_sc_hd__clkbuf_2
X_2539_ VSS VDD _0188_ _0463_ _0235_ VDD VSS sky130_fd_sc_hd__nand2_1
XANTENNA_nmat_col[28] VSS VDD core.ndc.col_out\[28\] VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_57_49 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
XANTENNA__2626__A VSS VDD core.osr.next_result_w\[8\] VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_83_384 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XFILLER_113_77 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_7_127 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XFILLER_138_41 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_138_85 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_98_23 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XANTENNA__1705__A VSS VDD core.ndc.col_out_n\[13\] VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__2536__A VSS VDD _0438_ VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1682__A2 VSS VDD _1135_ VDD VSS sky130_fd_sc_hd__diode_2
X_1910_ VSS VDD _1355_ _1378_ _1342_ VDD VSS sky130_fd_sc_hd__nand2_1
XFILLER_63_81 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
X_2890_ VSS VDD _0759_ _0783_ _0770_ VDD VSS sky130_fd_sc_hd__nand2_1
X_1841_ VSS VDD _1329_ _1330_ _1302_ VDD VSS sky130_fd_sc_hd__nand2_1
XANTENNA__2271__A VSS VDD core.cnb.result_out\[7\] VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__3086__B VSS VDD _0799_ VDD VSS sky130_fd_sc_hd__diode_2
X_1772_ VSS VDD core.ndc.col_out_n\[24\] _1283_ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xgenblk1\[3\].buf_n_coln VDD VSS core.ndc.col_out_n\[3\] nmatrix_col_core_n_buffered\[3\]
+ VDD VSS sky130_fd_sc_hd__buf_6
X_2324_ VSS VDD _0345_ _0271_ _0347_ _0346_ VDD VSS sky130_fd_sc_hd__nand3_1
XFILLER_69_134 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
X_2255_ VSS VDD _0277_ _0284_ _0273_ VDD VSS sky130_fd_sc_hd__nand2_1
Xpmat_sample_buf_n VSS VDD pmat_sample_switch_n_buffered core.cnb.enable_loop_out
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
X_2186_ VDD VSS core.cnb.average_sum_r\[0\] core.cnb.comparator_in core.cnb.average_sum_r\[1\]
+ _0224_ VDD VSS sky130_fd_sc_hd__a21o_1
XANTENNA__2622__A1 VSS VDD _0254_ VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_4_119 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XFILLER_88_410 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XFILLER_108_55 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XFILLER_88_454 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XANTENNA__3162__D VSS VDD core.osr.next_result_w\[2\] VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_75_137 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XFILLER_56_351 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_17_74 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XANTENNA__2613__B2 VSS VDD core.osr.next_result_w\[2\] VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_33_40 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XANTENNA__2129__B1 VSS VDD _1121_ VDD VSS sky130_fd_sc_hd__diode_2
X_2040_ VSS VDD core.pdc.col_out_n\[13\] _0122_ VDD VSS sky130_fd_sc_hd__clkbuf_1
XFILLER_47_373 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
X_2942_ VSS VDD _0753_ _0832_ _0834_ _0833_ VDD VSS sky130_fd_sc_hd__nand3_1
X_2873_ VDD VSS _0767_ _0708_ _0766_ VDD VSS sky130_fd_sc_hd__and2_1
XFILLER_90_90 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
X_1824_ VDD VSS _1316_ _1302_ VDD VSS sky130_fd_sc_hd__inv_2
X_1755_ VDD VSS core.ndc.col_out\[21\] core.ndc.col_out_n\[21\] VDD VSS sky130_fd_sc_hd__inv_2
XANTENNA__1591__A1 VSS VDD _1105_ VDD VSS sky130_fd_sc_hd__diode_2
X_1686_ VSS VDD _1223_ core.ndc.col_out_n\[11\] VDD VSS sky130_fd_sc_hd__clkbuf_2
XANTENNA_nmat_col[5] VSS VDD core.ndc.col_out\[5\] VDD VSS sky130_fd_sc_hd__diode_2
X_2307_ VSS VDD _0326_ _0331_ _0330_ VDD VSS sky130_fd_sc_hd__or2b_1
X_2238_ VSS VDD _0269_ _0268_ _0267_ _0988_ VDD VSS sky130_fd_sc_hd__and3_1
X_2169_ VSS VDD core.cnb.next_average_counter_w\[1\] _0211_ VDD VSS sky130_fd_sc_hd__clkbuf_1
XFILLER_72_129 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XFILLER_110_34 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XFILLER_119_150 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
XFILLER_119_87 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XFILLER_134_153 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XFILLER_79_47 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XANTENNA__1582__A1 VSS VDD _1079_ VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_95_24 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XFILLER_95_57 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XANTENNA_input15_A VSS VDD config_1_in[7] VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1702__B VSS VDD _1235_ VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_91_449 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XFILLER_44_61 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XANTENNA__2598__B1 VSS VDD _1022_ VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__3120__CLK VSS VDD clknet_2_0__leaf_clk_dig_dummy VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__3011__A1 VSS VDD _1053_ VDD VSS sky130_fd_sc_hd__diode_2
X_1540_ VDD VSS _1096_ _1095_ VDD VSS sky130_fd_sc_hd__buf_2
X_1471_ VSS VDD core.ndc.rowoff_out_n\[0\] core.ndc.row_out_n\[0\] core.ndc.rowon_out_n\[0\]
+ VDD VSS sky130_fd_sc_hd__nand2_1
X_3141_ VSS VDD clknet_2_0__leaf_clk_dig_dummy _0031_ net77 core.cnb.result_out\[9\]
+ VDD VSS sky130_fd_sc_hd__dfrtp_1
XFILLER_54_107 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XANTENNA_nmat_col_n[29] VSS VDD nmatrix_col_core_n_buffered\[29\] VDD VSS sky130_fd_sc_hd__diode_2
X_3072_ VSS VDD _0958_ _0833_ _0726_ _0910_ VDD VSS sky130_fd_sc_hd__and3_1
XFILLER_54_129 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
X_2023_ VDD VSS _0110_ _0108_ VDD VSS sky130_fd_sc_hd__inv_2
XFILLER_50_302 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
X_2925_ VSS VDD _0659_ _0816_ _0699_ _0817_ VDD VSS sky130_fd_sc_hd__nor3_1
X_2856_ VDD VSS _0751_ _0750_ VDD VSS sky130_fd_sc_hd__inv_2
X_1807_ VSS VDD core.cnb.data_register_r\[8\] _1300_ VDD VSS sky130_fd_sc_hd__clkbuf_2
X_2787_ VSS VDD _0640_ _0683_ _0682_ VDD VSS sky130_fd_sc_hd__nand2_1
X_1738_ VSS VDD _1035_ _1231_ _1260_ _1259_ core.ndc.col_out_n\[18\] _1261_ VDD VSS
+ sky130_fd_sc_hd__o221a_2
X_1669_ VSS VDD _1209_ _1197_ _1054_ _1208_ VDD VSS sky130_fd_sc_hd__mux2_1
XANTENNA_input7_A VSS VDD config_1_in[14] VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1803__A VSS VDD core.ndc.col_out\[31\] VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1867__A2 VSS VDD _1325_ VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_121_11 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XFILLER_121_33 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XANTENNA__2634__A VSS VDD _0983_ VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__3143__CLK VSS VDD clknet_2_0__leaf_clk_dig_dummy VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_14_53 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XFILLER_14_75 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XFILLER_30_74 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XANTENNA__1555__A1 VSS VDD _1037_ VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_30_85 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XFILLER_122_134 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
XANTENNA__1432__B VSS VDD _0995_ VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_36_118 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_55_93 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
X_2710_ VDD VSS _0609_ _0608_ VDD VSS sky130_fd_sc_hd__inv_2
X_2641_ VDD VSS _0548_ _0537_ core.osr.next_result_w\[3\] VDD VSS sky130_fd_sc_hd__or2_1
X_2572_ VDD VSS _0492_ _1200_ _0489_ VDD VSS sky130_fd_sc_hd__or2_1
X_1523_ VSS VDD core.cnb.data_register_r\[7\] _1081_ _1058_ VDD VSS sky130_fd_sc_hd__nand2_1
X_1454_ VSS VDD _1018_ _1006_ _1017_ VDD VSS sky130_fd_sc_hd__nand2_2
XANTENNA__1623__A VSS VDD _1128_ VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA_pmat_sample_buf_A VSS VDD net55 VDD VSS sky130_fd_sc_hd__diode_2
X_3124_ VSS VDD clknet_2_2__leaf_clk_dig_dummy core.cnb.next_average_counter_w\[2\]
+ net89 core.cnb.average_counter_r\[2\] VDD VSS sky130_fd_sc_hd__dfrtp_1
X_3055_ VSS VDD _0905_ _0943_ _0942_ _0781_ _0936_ VDD VSS sky130_fd_sc_hd__o211ai_1
X_2006_ VDD VSS core.pdc.col_out_n\[8\] core.pdc.col_out\[8\] VDD VSS sky130_fd_sc_hd__clkinv_2
XFILLER_50_110 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
X_2908_ VSS VDD _0799_ _0800_ _0796_ VDD VSS sky130_fd_sc_hd__nand2_1
XANTENNA__2982__B1 VSS VDD _1114_ VDD VSS sky130_fd_sc_hd__diode_2
X_2839_ VSS VDD _0733_ _0730_ _0734_ _0731_ VDD VSS sky130_fd_sc_hd__nand3_1
XANTENNA__1537__A1 VSS VDD _1064_ VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_104_123 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_116_55 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XANTENNA_fanout65_A VSS VDD net66 VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_18_129 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
Xgenblk2\[4\].buf_n_rowonn VSS VDD nmatrix_rowon_core_n_buffered\[4\] core.ndc.rowon_out_n\[4\]
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
XFILLER_92_25 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XANTENNA_nmat_rowon_n[1] VSS VDD nmatrix_rowon_core_n_buffered\[1\] VDD VSS sky130_fd_sc_hd__diode_2
Xgenblk1\[8\].buf_n_coln VDD VSS core.ndc.col_out_n\[8\] nmatrix_col_core_n_buffered\[8\]
+ VDD VSS sky130_fd_sc_hd__buf_6
XFILLER_110_104 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
XFILLER_110_126 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XANTENNA__3189__CLK VSS VDD clknet_2_1__leaf_clk_dig_dummy VDD VSS sky130_fd_sc_hd__diode_2
X_2624_ VSS VDD _0037_ _0531_ _0529_ _0532_ VDD VSS sky130_fd_sc_hd__a21bo_1
XANTENNA__1618__A VSS VDD _1163_ VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_63_1 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
X_2555_ VSS VDD _0474_ _0478_ core.cnb.pswitch_out\[1\] VDD VSS sky130_fd_sc_hd__nand2_1
X_2486_ VDD VSS _0001_ sample_nmatrix_cgen VDD VSS sky130_fd_sc_hd__inv_2
X_1506_ VDD VSS _1064_ _1034_ VDD VSS sky130_fd_sc_hd__buf_2
X_1437_ VSS VDD _1000_ _1001_ core.osr.osr_mode_r\[0\] VDD VSS sky130_fd_sc_hd__nor2_2
X_3107_ VSS VDD clknet_2_3__leaf_clk_dig_dummy _0007_ net88 core.cnb.shift_register_r\[5\]
+ VDD VSS sky130_fd_sc_hd__dfrtp_1
XFILLER_55_235 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
X_3038_ VSS VDD _0925_ _0926_ _0475_ VDD VSS sky130_fd_sc_hd__nand2_1
XANTENNA__2184__A VSS VDD core.cnb.comparator_in VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1758__A1 VSS VDD _1121_ VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1758__B2 VSS VDD _1125_ VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_11_21 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XANTENNA__1528__A VSS VDD _1079_ VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_87_25 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XFILLER_87_69 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XANTENNA__1710__B VSS VDD _1060_ VDD VSS sky130_fd_sc_hd__diode_2
Xinput15 VDD VSS net15 config_1_in[7] VDD VSS sky130_fd_sc_hd__buf_2
Xinput26 VSS VDD net26 config_2_in[2] VDD VSS sky130_fd_sc_hd__clkbuf_1
X_2340_ VDD VSS _0361_ core.osr.result_r\[13\] VDD VSS sky130_fd_sc_hd__inv_2
XFILLER_96_102 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
X_2271_ VSS VDD core.cnb.result_out\[7\] _0298_ core.osr.result_r\[7\] VDD VSS sky130_fd_sc_hd__nand2_1
XFILLER_78_883 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XFILLER_20_135 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
X_1986_ VDD VSS _0083_ _1206_ VDD VSS sky130_fd_sc_hd__inv_2
X_2607_ VDD VSS _0518_ _1001_ VDD VSS sky130_fd_sc_hd__inv_2
X_2538_ VSS VDD _0178_ _0222_ _0462_ _0187_ VDD VSS sky130_fd_sc_hd__nand3_1
XFILLER_87_113 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
X_2469_ VDD VSS core.ndc.rowoff_out_n\[15\] _0432_ VDD VSS sky130_fd_sc_hd__inv_2
XFILLER_69_883 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XFILLER_113_23 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_113_89 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XANTENNA__1530__B VSS VDD _1085_ VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_11_113 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_7_106 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
XFILLER_22_53 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_138_53 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_138_97 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
X_1840_ VSS VDD _1326_ _1023_ _1329_ VDD VSS sky130_fd_sc_hd__nor2_1
XFILLER_8_77 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
X_1771_ VSS VDD _1283_ _1282_ _1281_ _1280_ VDD VSS sky130_fd_sc_hd__and3_1
X_2323_ VSS VDD _0338_ _0328_ _0346_ _0343_ VDD VSS sky130_fd_sc_hd__nand3_1
X_2254_ VDD VSS _0283_ _0281_ _0282_ VDD VSS sky130_fd_sc_hd__and2_1
X_2185_ VSS VDD _0218_ core.cnb.average_sum_r\[1\] _0222_ _0223_ VDD VSS sky130_fd_sc_hd__or3b_1
XANTENNA__1631__A VSS VDD _1072_ VDD VSS sky130_fd_sc_hd__diode_2
X_1969_ VDD VSS _0070_ _0069_ VDD VSS sky130_fd_sc_hd__inv_2
XANTENNA__1806__A VSS VDD core.pdc.rowon_out_n\[0\] VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_108_78 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
XFILLER_88_433 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_88_477 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XANTENNA__1649__B1 VSS VDD _1082_ VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1541__A VSS VDD _1047_ VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_84_59 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XFILLER_56_385 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
XANTENNA__2091__B VSS VDD _1101_ VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__2129__A1 VSS VDD _1126_ VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_47_385 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
XFILLER_74_81 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
X_2941_ VDD VSS _0833_ _0806_ VDD VSS sky130_fd_sc_hd__inv_2
X_2872_ VSS VDD _0765_ _0766_ _0635_ VDD VSS sky130_fd_sc_hd__nand2_1
X_1823_ VSS VDD _1315_ core.pdc.row_out_n\[1\] _1307_ VDD VSS sky130_fd_sc_hd__nor2_2
X_1754_ VSS VDD _1271_ core.ndc.col_out_n\[21\] VDD VSS sky130_fd_sc_hd__clkbuf_2
XANTENNA__1591__A2 VSS VDD _1104_ VDD VSS sky130_fd_sc_hd__diode_2
X_1685_ VSS VDD _1223_ _1222_ _1219_ _1218_ VDD VSS sky130_fd_sc_hd__and3_1
XANTENNA_nmat_col[4] VSS VDD core.ndc.col_out\[4\] VDD VSS sky130_fd_sc_hd__diode_2
X_2306_ VSS VDD _0327_ _0329_ _0330_ VDD VSS sky130_fd_sc_hd__nor2_1
X_2237_ VDD VSS _0268_ _0266_ _0263_ VDD VSS sky130_fd_sc_hd__or2_1
XANTENNA__2457__A VSS VDD core.ndc.row_out_n\[2\] VDD VSS sky130_fd_sc_hd__diode_2
X_2168_ VSS VDD _0211_ _0191_ _0182_ _0210_ VDD VSS sky130_fd_sc_hd__and3_1
XFILLER_53_333 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
X_2099_ VDD VSS _0081_ _1173_ core.pdc.col_out\[25\] _0079_ _1096_ _0157_ VDD VSS
+ sky130_fd_sc_hd__a221o_1
XFILLER_134_121 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XANTENNA__1536__A VSS VDD _1091_ VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1582__A2 VSS VDD _1113_ VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_95_69 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XFILLER_63_108 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XFILLER_84_491 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_44_95 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XFILLER_44_73 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XANTENNA__2598__A1 VSS VDD _1328_ VDD VSS sky130_fd_sc_hd__diode_2
Xgenblk2\[12\].buf_p_rowonn VSS VDD pmatrix_rowon_core_n_buffered\[12\] core.pdc.rowon_out_n\[12\]
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
XFILLER_125_121 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_60_94 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
X_1470_ VSS VDD _1031_ core.ndc.rowon_out_n\[0\] _1030_ VDD VSS sky130_fd_sc_hd__nand2_4
X_3140_ VSS VDD clknet_2_0__leaf_clk_dig_dummy _0030_ net81 core.cnb.result_out\[8\]
+ VDD VSS sky130_fd_sc_hd__dfrtp_1
XANTENNA_nmat_col_n[28] VSS VDD nmatrix_col_core_n_buffered\[28\] VDD VSS sky130_fd_sc_hd__diode_2
X_3071_ VSS VDD _0936_ _0957_ _0956_ VDD VSS sky130_fd_sc_hd__nand2_1
X_2022_ VDD VSS core.pdc.col_out_n\[10\] core.pdc.col_out\[10\] VDD VSS sky130_fd_sc_hd__clkinv_2
XFILLER_62_130 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XANTENNA_genblk2\[8\].buf_p_rown_A VSS VDD core.pdc.row_out_n\[8\] VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_93_1 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
X_2924_ VDD VSS _0816_ _0645_ VDD VSS sky130_fd_sc_hd__inv_2
X_2855_ VSS VDD _0454_ _0749_ _0750_ VDD VSS sky130_fd_sc_hd__nor2_1
X_1806_ VSS VDD core.pdc.rowon_out_n\[0\] core.pdc.row_out_n\[0\] core.pdc.rowoff_out_n\[0\]
+ VDD VSS sky130_fd_sc_hd__nand2_1
X_2786_ VSS VDD _0681_ _0659_ _0682_ VDD VSS sky130_fd_sc_hd__nor2_1
XANTENNA_genblk2\[13\].buf_p_rowonn_A VSS VDD core.pdc.rowon_out_n\[13\] VDD VSS sky130_fd_sc_hd__diode_2
X_1737_ VDD VSS _1261_ _1074_ _1204_ VDD VSS sky130_fd_sc_hd__or2_1
XFILLER_131_113 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
X_1668_ VSS VDD _1206_ _1207_ _1208_ VDD VSS sky130_fd_sc_hd__nor2_1
X_1599_ VDD VSS _1149_ _1148_ VDD VSS sky130_fd_sc_hd__inv_2
XFILLER_105_35 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_105_57 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XANTENNA__3168__D VSS VDD core.osr.next_result_w\[8\] VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_91_225 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
X_2640_ VSS VDD _0544_ _0545_ _0547_ _0546_ VDD VSS sky130_fd_sc_hd__nand3_1
XANTENNA__2560__A VSS VDD core.cnb.data_register_r\[2\] VDD VSS sky130_fd_sc_hd__diode_2
X_2571_ VSS VDD _0025_ _0439_ _0489_ _0490_ _0491_ VDD VSS sky130_fd_sc_hd__o31a_1
X_1522_ VDD VSS _1080_ _1079_ VDD VSS sky130_fd_sc_hd__inv_2
X_1453_ VDD VSS _1017_ _1016_ VDD VSS sky130_fd_sc_hd__inv_2
XFILLER_87_509 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_113_124 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
X_3123_ VSS VDD clknet_2_2__leaf_clk_dig_dummy core.cnb.next_average_counter_w\[1\]
+ net88 core.cnb.average_counter_r\[1\] VDD VSS sky130_fd_sc_hd__dfrtp_1
XFILLER_27_108 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
X_3054_ VSS VDD _0941_ _0942_ _0905_ VDD VSS sky130_fd_sc_hd__nand2_1
X_2005_ VSS VDD _1035_ _0072_ _0094_ _1126_ core.pdc.col_out_n\[8\] _0097_ VDD VSS
+ sky130_fd_sc_hd__o221a_1
XFILLER_50_122 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
X_2907_ VDD VSS _0784_ _0799_ VDD VSS sky130_fd_sc_hd__buf_6
XANTENNA__2470__A VSS VDD core.pdc.row_out_n\[1\] VDD VSS sky130_fd_sc_hd__diode_2
X_2838_ VSS VDD _0638_ _0658_ _0733_ VDD VSS sky130_fd_sc_hd__nor2_1
X_2769_ VSS VDD _0662_ _0664_ _0665_ _0658_ VDD VSS sky130_fd_sc_hd__o21ai_1
XANTENNA__2734__A1 VSS VDD core.cnb.result_out\[11\] VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_104_135 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XFILLER_116_67 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XANTENNA__3110__CLK VSS VDD clknet_2_3__leaf_clk_dig_dummy VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_132_66 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XANTENNA_fanout58_A VSS VDD net67 VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_26_141 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XFILLER_92_37 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_54_494 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XFILLER_41_85 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XANTENNA_nmat_rowon_n[0] VSS VDD nmatrix_rowon_core_n_buffered\[0\] VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_2_13 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_49_266 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_92_501 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
Xgenblk2\[9\].buf_p_rowonn VSS VDD pmatrix_rowon_core_n_buffered\[9\] core.pdc.rowon_out_n\[9\]
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
XFILLER_32_111 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_82_81 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
X_2623_ VSS VDD _0394_ _0532_ net47 VDD VSS sky130_fd_sc_hd__nand2_1
X_2554_ VDD VSS _0477_ core.cnb.pswitch_out\[1\] _0474_ VDD VSS sky130_fd_sc_hd__or2_1
X_1505_ VDD VSS core.ndc.col_out\[0\] core.ndc.col_out_n\[0\] VDD VSS sky130_fd_sc_hd__inv_2
XFILLER_99_133 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XANTENNA__1634__A VSS VDD _1179_ VDD VSS sky130_fd_sc_hd__diode_2
X_2485_ VSS VDD sample_pmatrix_cgen _0000_ VDD VSS sky130_fd_sc_hd__inv_1
X_1436_ VDD VSS _1000_ _0994_ VDD VSS sky130_fd_sc_hd__inv_2
XANTENNA__3133__CLK VSS VDD clknet_2_0__leaf_clk_dig_dummy VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_101_116 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
X_3106_ VSS VDD clknet_2_2__leaf_clk_dig_dummy _0006_ net88 core.cnb.shift_register_r\[4\]
+ VDD VSS sky130_fd_sc_hd__dfrtp_1
XFILLER_83_501 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
X_3037_ VSS VDD _0831_ _0925_ _0924_ VDD VSS sky130_fd_sc_hd__nand2_1
XFILLER_62_29 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XANTENNA__1809__A VSS VDD net14 VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1758__A2 VSS VDD _1193_ VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_127_7 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XANTENNA__1528__B VSS VDD _1085_ VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_11_88 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_93_309 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_36_85 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
Xinput16 VSS VDD net16 config_1_in[8] VDD VSS sky130_fd_sc_hd__clkbuf_1
Xinput27 VSS VDD net27 config_2_in[3] VDD VSS sky130_fd_sc_hd__clkbuf_1
XANTENNA_genblk1\[1\].buf_n_coln_A VSS VDD core.ndc.col_out_n\[1\] VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_42_7 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_35_6 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
X_2270_ VSS VDD core.cnb.result_out\[7\] core.osr.result_r\[7\] _0297_ VDD VSS sky130_fd_sc_hd__nor2_1
XFILLER_20_125 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
X_1985_ VSS VDD _0081_ _0082_ _1275_ VDD VSS sky130_fd_sc_hd__nand2_1
X_2606_ VSS VDD _1003_ _0517_ VDD VSS sky130_fd_sc_hd__clkbuf_2
XANTENNA__3121__RESET_B VSS VDD net86 VDD VSS sky130_fd_sc_hd__diode_2
X_2537_ VSS VDD _0460_ _0461_ VDD VSS sky130_fd_sc_hd__clkbuf_2
X_2468_ VDD VSS _0432_ core.ndc.row_out_n\[15\] core.ndc.rowon_out_n\[15\] VDD VSS
+ sky130_fd_sc_hd__and2_1
XFILLER_87_125 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
X_1419_ VDD VSS _0982_ _0983_ VDD VSS sky130_fd_sc_hd__clkinv_2
X_2399_ VSS VDD core.osr.sample_count_r\[4\] _0405_ _0409_ VDD VSS sky130_fd_sc_hd__nor2_1
XFILLER_56_501 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XFILLER_113_57 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XFILLER_51_272 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XFILLER_11_125 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XANTENNA__1539__A VSS VDD _1072_ VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__3179__CLK VSS VDD net58 VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_22_65 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_138_65 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_47_501 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XANTENNA__2864__B1 VSS VDD core.cnb.data_register_r\[1\] VDD VSS sky130_fd_sc_hd__diode_2
X_1770_ VSS VDD _1172_ _1282_ _1095_ VDD VSS sky130_fd_sc_hd__nand2_1
X_2322_ VSS VDD _0339_ _0345_ _0344_ VDD VSS sky130_fd_sc_hd__nand2_1
X_2253_ VSS VDD core.cnb.result_out\[5\] _0282_ core.osr.result_r\[5\] VDD VSS sky130_fd_sc_hd__nand2_1
XANTENNA_cgen_sample_n_in VSS VDD net54 VDD VSS sky130_fd_sc_hd__diode_2
X_2184_ VDD VSS _0222_ core.cnb.comparator_in VDD VSS sky130_fd_sc_hd__inv_2
XANTENNA__2727__B VSS VDD _1002_ VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_53_515 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XANTENNA__2462__B VSS VDD core.ndc.rowon_out_n\[9\] VDD VSS sky130_fd_sc_hd__diode_2
X_1968_ VSS VDD _0069_ _1105_ _1104_ _1403_ _1088_ VDD VSS sky130_fd_sc_hd__a31o_1
X_1899_ VDD VSS core.pdc.rowon_out_n\[3\] _1371_ VDD VSS sky130_fd_sc_hd__inv_2
XANTENNA__1806__B VSS VDD core.pdc.rowoff_out_n\[0\] VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_88_445 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
XFILLER_48_309 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XFILLER_75_106 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
XANTENNA__1649__A1 VSS VDD _1128_ VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1541__B VSS VDD _1057_ VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_123_1 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
XFILLER_47_397 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
X_2940_ VSS VDD _0809_ _0819_ _0832_ VDD VSS sky130_fd_sc_hd__nor2_1
X_2871_ VSS VDD core.cnb.shift_register_r\[4\] _0705_ _0765_ VDD VSS sky130_fd_sc_hd__nor2_1
X_1822_ VSS VDD _1311_ _1314_ _1315_ VDD VSS sky130_fd_sc_hd__nor2_1
XFILLER_90_81 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XFILLER_128_141 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
X_1753_ VSS VDD _1271_ _1209_ _1034_ _1139_ VDD VSS sky130_fd_sc_hd__mux2_1
X_1684_ VSS VDD _1221_ _1222_ _1177_ VDD VSS sky130_fd_sc_hd__nand2_1
XANTENNA_nmat_col[3] VSS VDD core.ndc.col_out\[3\] VDD VSS sky130_fd_sc_hd__diode_2
X_2305_ VDD VSS _0329_ _0328_ VDD VSS sky130_fd_sc_hd__inv_2
XANTENNA__1642__A VSS VDD _1117_ VDD VSS sky130_fd_sc_hd__diode_2
X_2236_ VSS VDD _0263_ _0267_ _0266_ VDD VSS sky130_fd_sc_hd__nand2_1
XANTENNA__2457__B VSS VDD core.ndc.rowon_out_n\[2\] VDD VSS sky130_fd_sc_hd__diode_2
X_2167_ VSS VDD _0210_ core.cnb.next_average_counter_w\[0\] core.cnb.average_counter_r\[0\]
+ VDD VSS sky130_fd_sc_hd__nand2_1
X_2098_ VSS VDD _0065_ _0115_ _0157_ VDD VSS sky130_fd_sc_hd__nor2_1
XANTENNA__2473__A VSS VDD core.pdc.row_out_n\[4\] VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1567__B1 VSS VDD _1075_ VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_134_133 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
XANTENNA__1536__B VSS VDD _1093_ VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_0_113 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XFILLER_71_120 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_125_133 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XFILLER_5_68 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
X_3070_ VSS VDD _0904_ _0948_ _0956_ VDD VSS sky130_fd_sc_hd__nor2_1
X_2021_ VSS VDD _1064_ _0076_ _0106_ _1224_ core.pdc.col_out_n\[10\] _0109_ VDD VSS
+ sky130_fd_sc_hd__o221a_1
XFILLER_47_194 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
X_2923_ VSS VDD _0750_ _0814_ _0815_ VDD VSS sky130_fd_sc_hd__nor2_1
X_2854_ VSS VDD _0748_ _0749_ _0649_ VDD VSS sky130_fd_sc_hd__nand2_1
X_1805_ VSS VDD _1030_ core.pdc.rowoff_out_n\[0\] _1027_ VDD VSS sky130_fd_sc_hd__nand2_1
X_2785_ VSS VDD _0644_ _0681_ _0642_ VDD VSS sky130_fd_sc_hd__nand2_1
XFILLER_116_100 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
X_1736_ VDD VSS _1260_ _1124_ VDD VSS sky130_fd_sc_hd__inv_2
X_1667_ VSS VDD _1113_ _1057_ _1207_ VDD VSS sky130_fd_sc_hd__nor2_1
XFILLER_131_125 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
X_1598_ VSS VDD _1148_ _1147_ _1077_ _1146_ VDD VSS sky130_fd_sc_hd__mux2_1
XFILLER_105_47 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XFILLER_45_109 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
X_2219_ VSS VDD _0251_ _0252_ VDD VSS sky130_fd_sc_hd__clkbuf_2
XANTENNA__2277__A1 VSS VDD core.cnb.result_out\[7\] VDD VSS sky130_fd_sc_hd__diode_2
X_3199_ VSS VDD net64 core.osr.next_sample_count_w\[7\] net77 core.osr.sample_count_r\[7\]
+ VDD VSS sky130_fd_sc_hd__dfrtp_1
XFILLER_121_68 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XFILLER_121_57 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XFILLER_81_39 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XANTENNA__1547__A VSS VDD _1078_ VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_39_41 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XANTENNA_input20_A VSS VDD config_2_in[11] VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_91_237 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_44_153 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
X_2570_ VDD VSS _0491_ core.cnb.result_out\[3\] _0461_ VDD VSS sky130_fd_sc_hd__or2_1
X_1521_ VSS VDD _1079_ _1044_ _1055_ VDD VSS sky130_fd_sc_hd__nand2_2
X_1452_ VDD VSS _1003_ _1007_ _1016_ _1010_ _1012_ _1015_ VDD VSS sky130_fd_sc_hd__a221o_1
XFILLER_113_136 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
X_3122_ VDD VSS core.cnb.average_counter_r\[0\] net88 core.cnb.next_average_counter_w\[0\]
+ clknet_2_2__leaf_clk_dig_dummy VDD VSS sky130_fd_sc_hd__dfstp_1
X_3053_ VSS VDD _0937_ _0941_ _0940_ VDD VSS sky130_fd_sc_hd__nand2_1
X_2004_ VSS VDD _0096_ _0097_ _1284_ VDD VSS sky130_fd_sc_hd__nand2_1
XANTENNA__2431__B2 VSS VDD core.ndc.row_bottotop_n\[10\] VDD VSS sky130_fd_sc_hd__diode_2
X_2906_ VSS VDD _0795_ _0798_ _0797_ VDD VSS sky130_fd_sc_hd__nand2_1
XANTENNA__2470__B VSS VDD core.pdc.rowon_out_n\[1\] VDD VSS sky130_fd_sc_hd__diode_2
X_2837_ VSS VDD _0729_ _0730_ _0732_ _0731_ VDD VSS sky130_fd_sc_hd__nand3_1
X_2768_ VSS VDD _0640_ _0647_ _0664_ _0663_ VDD VSS sky130_fd_sc_hd__nand3_1
X_2699_ VSS VDD _0596_ _0597_ _0599_ _0598_ VDD VSS sky130_fd_sc_hd__nand3_1
X_1719_ VSS VDD _1075_ _1246_ _1183_ _1064_ core.ndc.col_out_n\[15\] _1248_ VDD VSS
+ sky130_fd_sc_hd__o221a_2
XANTENNA__1942__A0 VSS VDD _1067_ VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_116_79 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XFILLER_132_34 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XANTENNA_cgen_start_conv_in VSS VDD net35 VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_132_78 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
XFILLER_54_473 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XFILLER_92_49 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XFILLER_41_134 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XFILLER_41_97 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XANTENNA__1724__B VSS VDD _1213_ VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_2_25 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
Xgenblk1\[10\].buf_p_coln VSS VDD pmatrix_col_core_n_buffered\[10\] core.pdc.col_out_n\[10\]
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
XFILLER_2_69 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_92_513 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XANTENNA__2555__B VSS VDD core.cnb.pswitch_out\[1\] VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_32_123 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
X_2622_ VDD VSS _0530_ _0254_ _1018_ _0531_ VDD VSS sky130_fd_sc_hd__a21oi_1
X_2553_ VSS VDD _0476_ _0461_ core.cnb.result_out\[0\] _0474_ _0022_ VDD VSS sky130_fd_sc_hd__o22a_1
X_1504_ VSS VDD core.ndc.col_out_n\[0\] _1063_ _1049_ _1035_ VDD VSS sky130_fd_sc_hd__o21a_2
X_2484_ VDD VSS core.cnb.enable_loop_out net55 VDD VSS sky130_fd_sc_hd__inv_2
X_1435_ VDD VSS _0999_ core.osr.sample_count_r\[4\] VDD VSS sky130_fd_sc_hd__inv_2
X_3105_ VSS VDD clknet_2_2__leaf_clk_dig_dummy _0005_ net88 core.cnb.shift_register_r\[3\]
+ VDD VSS sky130_fd_sc_hd__dfrtp_1
X_3036_ VDD VSS _0924_ _0923_ VDD VSS sky130_fd_sc_hd__inv_2
XANTENNA__1650__A VSS VDD _1077_ VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__2465__B VSS VDD _1325_ VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_102_15 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
XFILLER_102_59 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XANTENNA__2481__A VSS VDD core.pdc.row_out_n\[14\] VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA_fanout70_A VSS VDD net83 VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA_genblk1\[16\].buf_n_coln_A VSS VDD core.ndc.col_out_n\[16\] VDD VSS sky130_fd_sc_hd__diode_2
Xinput17 VSS VDD net17 config_1_in[9] VDD VSS sky130_fd_sc_hd__clkbuf_1
Xinput28 VDD VSS net28 config_2_in[4] VDD VSS sky130_fd_sc_hd__dlymetal6s2s_1
Xgenblk2\[0\].buf_n_rowonn VSS VDD nmatrix_rowon_core_n_buffered\[0\] core.ndc.rowon_out_n\[0\]
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
Xgenblk2\[14\].buf_p_rown VSS VDD pmatrix_row_core_n_buffered\[14\] core.pdc.row_out_n\[14\]
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
XANTENNA__2566__A VSS VDD core.cnb.data_register_r\[1\] VDD VSS sky130_fd_sc_hd__diode_2
X_1984_ VSS VDD _0081_ _1112_ _1409_ _1118_ VDD VSS sky130_fd_sc_hd__mux2_1
X_2605_ VDD VSS _0395_ _0516_ _0995_ _0034_ net38 VDD VSS sky130_fd_sc_hd__a22o_1
XANTENNA_nmat_col[25] VSS VDD core.ndc.col_out\[25\] VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1645__A VSS VDD _1187_ VDD VSS sky130_fd_sc_hd__diode_2
X_2536_ VDD VSS _0460_ _0438_ VDD VSS sky130_fd_sc_hd__inv_2
X_2467_ VSS VDD core.ndc.row_out_n\[14\] core.ndc.rowoff_out_n\[14\] core.ndc.rowon_out_n\[14\]
+ VDD VSS sky130_fd_sc_hd__nand2_1
XANTENNA_genblk1\[6\].buf_p_coln_A VSS VDD core.pdc.col_out_n\[6\] VDD VSS sky130_fd_sc_hd__diode_2
X_1418_ VDD VSS net11 net13 net12 _0982_ VDD VSS sky130_fd_sc_hd__or3_1
XFILLER_87_137 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
X_2398_ VDD VSS core.osr.next_sample_count_w\[3\] _0408_ VDD VSS sky130_fd_sc_hd__inv_2
XFILLER_83_365 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
X_3019_ VSS VDD _0804_ _0870_ _0907_ VDD VSS sky130_fd_sc_hd__nor2_1
XFILLER_51_251 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XFILLER_11_137 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_138_77 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
XANTENNA__2864__B2 VSS VDD _0758_ VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_63_40 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XANTENNA__2833__B VSS VDD _0637_ VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_8_13 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XANTENNA__3123__CLK VSS VDD clknet_2_2__leaf_clk_dig_dummy VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_40_5 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
X_2321_ VDD VSS _0344_ _0343_ VDD VSS sky130_fd_sc_hd__inv_2
XANTENNA__2552__B1 VSS VDD core.cnb.pswitch_out\[0\] VDD VSS sky130_fd_sc_hd__diode_2
X_2252_ VDD VSS _0281_ core.cnb.result_out\[5\] core.osr.result_r\[5\] VDD VSS sky130_fd_sc_hd__or2_1
X_2183_ VDD VSS core.cnb.comparator_in core.cnb.next_average_sum_w\[0\] _0221_ VDD
+ VSS sky130_fd_sc_hd__xor2_1
XFILLER_138_109 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
X_1967_ VDD VSS _0068_ _1407_ VDD VSS sky130_fd_sc_hd__inv_2
X_1898_ VSS VDD _1370_ _1309_ _1371_ _1305_ VDD VSS sky130_fd_sc_hd__o21ai_2
XFILLER_108_25 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XFILLER_108_47 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
Xgenblk2\[11\].buf_n_rown VSS VDD nmatrix_row_core_n_buffered\[11\] core.ndc.row_out_n\[11\]
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
XFILLER_68_29 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
X_2519_ VSS VDD _0451_ core.cnb.shift_register_r\[13\] _0219_ core.cnb.shift_register_r\[12\]
+ VDD VSS sky130_fd_sc_hd__mux2_1
XFILLER_56_321 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_56_365 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_33_87 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XANTENNA__2534__A0 VSS VDD core.cnb.sampled_avg_control_r\[2\] VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_58_40 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
X_2870_ VSS VDD _0702_ _0764_ _0763_ VDD VSS sky130_fd_sc_hd__nand2_1
XFILLER_71_891 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
X_1821_ VDD VSS _1314_ _1313_ VDD VSS sky130_fd_sc_hd__inv_2
X_1752_ VDD VSS core.ndc.col_out_n\[20\] core.ndc.col_out\[20\] VDD VSS sky130_fd_sc_hd__clkinv_2
X_1683_ VDD VSS _1221_ _1220_ VDD VSS sky130_fd_sc_hd__inv_2
XANTENNA_nmat_col[2] VSS VDD core.ndc.col_out\[2\] VDD VSS sky130_fd_sc_hd__diode_2
X_2304_ VSS VDD core.osr.result_r\[10\] _0328_ core.cnb.result_out\[10\] VDD VSS sky130_fd_sc_hd__nand2_1
X_2235_ VDD VSS _0266_ _0264_ _0265_ VDD VSS sky130_fd_sc_hd__and2_1
X_2166_ VSS VDD _0209_ _0210_ VDD VSS sky130_fd_sc_hd__clkbuf_2
XANTENNA__3169__CLK VSS VDD net66 VDD VSS sky130_fd_sc_hd__diode_2
X_2097_ VDD VSS core.pdc.col_out_n\[24\] core.pdc.col_out\[24\] VDD VSS sky130_fd_sc_hd__inv_2
XFILLER_62_891 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
X_2999_ VSS VDD _0763_ _0888_ _0695_ VDD VSS sky130_fd_sc_hd__nand2_1
XANTENNA__1567__A1 VSS VDD _1064_ VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_88_298 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
Xgenblk1\[15\].buf_p_coln VSS VDD pmatrix_col_core_n_buffered\[15\] core.pdc.col_out_n\[15\]
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
XFILLER_71_132 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XFILLER_60_41 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_69_50 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
XANTENNA__1743__A VSS VDD _1227_ VDD VSS sky130_fd_sc_hd__diode_2
X_2020_ VSS VDD _0108_ _0109_ _1093_ VDD VSS sky130_fd_sc_hd__nand2_1
XFILLER_90_441 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XFILLER_90_463 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
X_2922_ VSS VDD _0737_ _0811_ _0814_ _0813_ VDD VSS sky130_fd_sc_hd__nand3_1
XANTENNA__1918__A VSS VDD _1381_ VDD VSS sky130_fd_sc_hd__diode_2
X_2853_ VSS VDD _0646_ _0673_ _0747_ _0748_ VDD VSS sky130_fd_sc_hd__nor3_1
X_1804_ VSS VDD core.pdc.rowon_out_n\[0\] _1025_ _1031_ VDD VSS sky130_fd_sc_hd__nand2_2
X_2784_ VDD VSS _0680_ _0679_ VDD VSS sky130_fd_sc_hd__inv_2
X_1735_ VSS VDD _1110_ _1259_ VDD VSS sky130_fd_sc_hd__clkbuf_2
XANTENNA__1637__B VSS VDD _1096_ VDD VSS sky130_fd_sc_hd__diode_2
X_1666_ VSS VDD _1206_ _1059_ _1052_ VDD VSS sky130_fd_sc_hd__nand2_2
XFILLER_131_137 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
X_1597_ VSS VDD _1123_ _1147_ _1068_ VDD VSS sky130_fd_sc_hd__nand2_1
X_2218_ VDD VSS _0251_ _0988_ VDD VSS sky130_fd_sc_hd__inv_2
X_3198_ VSS VDD net64 core.osr.next_sample_count_w\[6\] net77 core.osr.sample_count_r\[6\]
+ VDD VSS sky130_fd_sc_hd__dfrtp_1
X_2149_ VDD VSS _0193_ _0190_ _0192_ VDD VSS sky130_fd_sc_hd__or2_1
XFILLER_53_121 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XANTENNA__2484__A VSS VDD net55 VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_107_145 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
XFILLER_30_99 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XANTENNA__2268__A2 VSS VDD _0255_ VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_91_205 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_55_30 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XANTENNA_input13_A VSS VDD config_1_in[5] VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_91_249 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
X_1520_ VDD VSS _1078_ _1077_ VDD VSS sky130_fd_sc_hd__buf_2
X_1451_ VDD VSS core.osr.sample_count_r\[8\] _0992_ _1014_ _1015_ VDD VSS sky130_fd_sc_hd__a21o_1
XANTENNA__2569__A VSS VDD _1395_ VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1473__A VSS VDD _1032_ VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_113_148 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
Xgenblk1\[12\].buf_n_coln VDD VSS core.ndc.col_out_n\[12\] nmatrix_col_core_n_buffered\[12\]
+ VDD VSS sky130_fd_sc_hd__buf_6
X_3121_ VSS VDD clknet_2_2__leaf_clk_dig_dummy _0021_ net86 core.cnb.sampled_avg_control_r\[2\]
+ VDD VSS sky130_fd_sc_hd__dfrtp_2
XANTENNA__2259__A2 VSS VDD _0240_ VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_48_460 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
X_3052_ VDD VSS _0940_ _0939_ VDD VSS sky130_fd_sc_hd__inv_2
XFILLER_48_482 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
X_2003_ VDD VSS _0096_ _0095_ VDD VSS sky130_fd_sc_hd__inv_2
XANTENNA__3186__RESET_B VSS VDD net85 VDD VSS sky130_fd_sc_hd__diode_2
X_2905_ VDD VSS _0797_ _0796_ VDD VSS sky130_fd_sc_hd__inv_2
XANTENNA__1648__A VSS VDD core.ndc.col_out_n\[8\] VDD VSS sky130_fd_sc_hd__diode_2
X_2836_ VDD VSS _0731_ _0724_ VDD VSS sky130_fd_sc_hd__dlymetal6s2s_1
X_2767_ VSS VDD core.cnb.shift_register_r\[9\] _0633_ _0663_ VDD VSS sky130_fd_sc_hd__nor2_1
X_2698_ VSS VDD core.osr.next_result_w\[14\] _0598_ _0535_ VDD VSS sky130_fd_sc_hd__nand2_1
X_1718_ VSS VDD _1247_ _1248_ _1093_ VDD VSS sky130_fd_sc_hd__nand2_1
XFILLER_104_104 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XANTENNA__2479__A VSS VDD core.pdc.rowon_out_n\[12\] VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_116_14 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XANTENNA_nmat_rowon_n[12] VSS VDD nmatrix_rowon_core_n_buffered\[12\] VDD VSS sky130_fd_sc_hd__diode_2
X_1649_ VDD VSS core.cnb.data_register_r\[7\] _1128_ _1082_ _1191_ VDD VSS sky130_fd_sc_hd__a21o_1
XANTENNA_genblk2\[4\].buf_p_rown_A VSS VDD core.pdc.row_out_n\[4\] VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA_input5_A VSS VDD config_1_in[12] VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_132_13 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_132_46 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XFILLER_41_113 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_41_32 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XANTENNA__2186__A1 VSS VDD core.cnb.comparator_in VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_89_393 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_92_525 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XANTENNA__1740__B VSS VDD _1152_ VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_82_61 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
X_2621_ VSS VDD _1009_ _0530_ VDD VSS sky130_fd_sc_hd__clkbuf_2
X_2552_ VDD VSS _0475_ _0461_ core.cnb.pswitch_out\[0\] _0476_ VDD VSS sky130_fd_sc_hd__a21oi_1
XANTENNA__1915__B VSS VDD core.ndc.rowon_bottotop_n\[5\] VDD VSS sky130_fd_sc_hd__diode_2
X_1503_ VDD VSS _1063_ _1062_ VDD VSS sky130_fd_sc_hd__inv_2
XFILLER_99_124 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
X_2483_ VDD VSS _0433_ core.pdc.rowoff_out_n\[15\] VDD VSS sky130_fd_sc_hd__clkinv_2
X_1434_ VSS VDD _0996_ _0998_ core.osr.sample_count_r\[0\] VDD VSS sky130_fd_sc_hd__nand2_1
X_3104_ VSS VDD clknet_2_2__leaf_clk_dig_dummy _0004_ net88 core.cnb.shift_register_r\[2\]
+ VDD VSS sky130_fd_sc_hd__dfrtp_2
XFILLER_83_525 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
X_3035_ VSS VDD _0853_ _0923_ _0827_ VDD VSS sky130_fd_sc_hd__nand2_1
XFILLER_23_113 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_23_135 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XANTENNA__2481__B VSS VDD core.pdc.rowon_out_n\[14\] VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_51_499 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XANTENNA__1612__B1 VSS VDD _1155_ VDD VSS sky130_fd_sc_hd__diode_2
X_2819_ VSS VDD _0692_ _0714_ _0713_ VDD VSS sky130_fd_sc_hd__nand2_1
XFILLER_11_35 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
XFILLER_11_57 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_127_57 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_127_79 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_87_17 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XFILLER_87_39 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_86_330 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_36_21 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
XANTENNA_fanout63_A VSS VDD net66 VDD VSS sky130_fd_sc_hd__diode_2
Xinput18 VSS VDD net18 config_2_in[0] VDD VSS sky130_fd_sc_hd__clkbuf_1
Xinput29 VDD VSS net29 config_2_in[5] VDD VSS sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__2566__B VSS VDD core.cnb.data_register_r\[0\] VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_92_322 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
X_1983_ VSS VDD _0079_ _0080_ _1279_ VDD VSS sky130_fd_sc_hd__nand2_1
X_2604_ VSS VDD _0279_ _1018_ _0516_ VDD VSS sky130_fd_sc_hd__nor2_1
XANTENNA__1645__B VSS VDD _1188_ VDD VSS sky130_fd_sc_hd__diode_2
X_2535_ VSS VDD _0021_ _0459_ VDD VSS sky130_fd_sc_hd__clkbuf_1
X_2466_ VSS VDD core.ndc.row_out_n\[13\] core.ndc.rowoff_out_n\[13\] core.ndc.rowon_out_n\[13\]
+ VDD VSS sky130_fd_sc_hd__nand2_1
Xgenblk2\[5\].buf_p_rowonn VSS VDD pmatrix_rowon_core_n_buffered\[5\] core.pdc.rowon_bottotop_n\[5\]
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
XFILLER_87_149 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
X_1417_ VDD VSS core.cnb.pswitch_out\[0\] core.cnb.data_register_r\[0\] VDD VSS sky130_fd_sc_hd__inv_2
X_2397_ VDD VSS _0404_ _0403_ _0407_ _0408_ VDD VSS sky130_fd_sc_hd__a21o_1
XANTENNA__2476__B VSS VDD core.pdc.rowon_out_n\[9\] VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_56_525 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XFILLER_83_333 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
X_3018_ VSS VDD _0895_ _0879_ _0906_ VDD VSS sky130_fd_sc_hd__nor2_1
XFILLER_11_149 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
XFILLER_78_127 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XFILLER_47_525 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XFILLER_86_171 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XANTENNA__2616__A2 VSS VDD _0395_ VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_63_96 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XANTENNA__1746__A VSS VDD core.ndc.col_out_n\[19\] VDD VSS sky130_fd_sc_hd__diode_2
Xgenblk1\[22\].buf_p_coln VSS VDD pmatrix_col_core_n_buffered\[22\] core.pdc.col_out_n\[22\]
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
XANTENNA__2001__B1 VSS VDD _1053_ VDD VSS sky130_fd_sc_hd__diode_2
X_2320_ VSS VDD _0340_ _0342_ _0343_ VDD VSS sky130_fd_sc_hd__nor2_1
X_2251_ VDD VSS _0280_ core.cnb.result_out\[5\] VDD VSS sky130_fd_sc_hd__inv_2
XANTENNA__1481__A VSS VDD core.ndc.rowon_out_n\[0\] VDD VSS sky130_fd_sc_hd__diode_2
X_2182_ VSS VDD _0218_ _0220_ _0221_ VDD VSS sky130_fd_sc_hd__nor2_1
XFILLER_92_141 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
X_1966_ VDD VSS core.pdc.col_out\[3\] core.pdc.col_out_n\[3\] VDD VSS sky130_fd_sc_hd__clkinv_2
X_1897_ VSS VDD _1338_ _1370_ _1369_ VDD VSS sky130_fd_sc_hd__nand2_1
XFILLER_108_37 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
X_2518_ VSS VDD _0013_ _0450_ VDD VSS sky130_fd_sc_hd__clkbuf_1
XFILLER_88_425 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XANTENNA__2487__A VSS VDD _0220_ VDD VSS sky130_fd_sc_hd__diode_2
X_2449_ VDD VSS core.pdc.rowoff_out_n\[5\] _1369_ _1384_ core.ndc.rowon_out_n\[10\]
+ VDD VSS sky130_fd_sc_hd__a21o_1
XFILLER_84_29 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
XFILLER_56_333 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XFILLER_83_141 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XFILLER_56_377 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XFILLER_17_89 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XFILLER_33_77 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XFILLER_33_99 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XANTENNA__2534__A1 VSS VDD net10 VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_58_52 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
Xclkbuf_2_0__f_clk_dig_dummy VSS VDD clknet_0_clk_dig_dummy clknet_2_0__leaf_clk_dig_dummy
+ VDD VSS sky130_fd_sc_hd__clkbuf_16
Xgenblk1\[17\].buf_n_coln VDD VSS core.ndc.col_out_n\[17\] nmatrix_col_core_n_buffered\[17\]
+ VDD VSS sky130_fd_sc_hd__buf_6
XFILLER_47_300 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_47_355 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_74_130 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
X_1820_ VSS VDD _1313_ core.cnb.data_register_r\[9\] _1022_ _1312_ VDD VSS sky130_fd_sc_hd__and3_1
X_1751_ VSS VDD core.ndc.col_out_n\[20\] _1270_ VDD VSS sky130_fd_sc_hd__clkbuf_1
X_1682_ VSS VDD _1135_ _1078_ _1220_ _1137_ VDD VSS sky130_fd_sc_hd__a21oi_2
XANTENNA_nmat_col[1] VSS VDD core.ndc.col_out\[1\] VDD VSS sky130_fd_sc_hd__diode_2
X_2303_ VSS VDD core.osr.result_r\[10\] core.cnb.result_out\[10\] _0327_ VDD VSS sky130_fd_sc_hd__nor2_1
XANTENNA__1923__B VSS VDD core.ndc.rowoff_out_n\[5\] VDD VSS sky130_fd_sc_hd__diode_2
X_2234_ VSS VDD core.cnb.result_out\[3\] _0265_ core.osr.result_r\[3\] VDD VSS sky130_fd_sc_hd__nand2_1
X_2165_ VDD VSS _0209_ _0208_ VDD VSS sky130_fd_sc_hd__inv_2
XFILLER_93_461 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
X_2096_ VDD VSS _0092_ _1275_ core.pdc.col_out\[24\] _0087_ _1102_ _0156_ VDD VSS
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_81 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
X_2998_ VSS VDD _0884_ _0887_ _0877_ VDD VSS sky130_fd_sc_hd__nand2_1
X_1949_ VDD VSS _1403_ _1389_ VDD VSS sky130_fd_sc_hd__inv_2
XFILLER_135_57 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XANTENNA__3113__CLK VSS VDD clknet_2_3__leaf_clk_dig_dummy VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_88_288 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
XFILLER_28_33 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_28_77 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XFILLER_56_163 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XFILLER_84_450 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XFILLER_71_100 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XFILLER_44_21 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
XFILLER_100_71 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_60_53 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XFILLER_125_102 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
XANTENNA_nmat_col_n[25] VSS VDD nmatrix_col_core_n_buffered\[25\] VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_85_50 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
XFILLER_85_72 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
X_2921_ VSS VDD _0812_ _0730_ _0813_ _0724_ VDD VSS sky130_fd_sc_hd__nand3_1
X_2852_ VSS VDD _0633_ _0747_ _0746_ VDD VSS sky130_fd_sc_hd__nand2_1
X_1803_ VDD VSS core.ndc.col_out_n\[31\] core.ndc.col_out\[31\] VDD VSS sky130_fd_sc_hd__inv_2
X_2783_ VSS VDD core.cnb.shift_register_r\[15\] _0678_ _0679_ VDD VSS sky130_fd_sc_hd__nor2_1
X_1734_ VDD VSS core.ndc.col_out\[17\] core.ndc.col_out_n\[17\] VDD VSS sky130_fd_sc_hd__inv_2
X_1665_ VDD VSS core.ndc.col_out\[9\] core.ndc.col_out_n\[9\] VDD VSS sky130_fd_sc_hd__inv_2
XANTENNA__3136__CLK VSS VDD clknet_2_0__leaf_clk_dig_dummy VDD VSS sky130_fd_sc_hd__diode_2
X_1596_ VDD VSS _1146_ _1145_ VDD VSS sky130_fd_sc_hd__inv_2
XFILLER_131_149 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
XANTENNA__1653__B VSS VDD _1104_ VDD VSS sky130_fd_sc_hd__diode_2
X_2217_ VSS VDD _0239_ _0248_ _0250_ _0243_ VDD VSS sky130_fd_sc_hd__o21ai_1
XFILLER_38_141 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
X_3197_ VSS VDD net64 core.osr.next_sample_count_w\[5\] net80 core.osr.sample_count_r\[5\]
+ VDD VSS sky130_fd_sc_hd__dfrtp_1
X_2148_ VDD VSS _0192_ _0184_ _0191_ VDD VSS sky130_fd_sc_hd__or2_1
XFILLER_121_48 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XFILLER_53_133 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
X_2079_ VDD VSS _1102_ _0108_ core.pdc.col_out\[20\] _1125_ _0146_ _0147_ VDD VSS
+ sky130_fd_sc_hd__a221o_1
XANTENNA__2434__B1 VSS VDD _1328_ VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_107_113 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XANTENNA_fanout93_A VSS VDD net94 VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_91_217 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
XFILLER_55_53 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
X_1450_ VSS VDD _0986_ _1014_ _1013_ VDD VSS sky130_fd_sc_hd__nand2_1
X_3120_ VSS VDD clknet_2_0__leaf_clk_dig_dummy _0020_ net85 core.cnb.sampled_avg_control_r\[1\]
+ VDD VSS sky130_fd_sc_hd__dfrtp_1
X_3051_ VSS VDD _0938_ _0939_ _0893_ VDD VSS sky130_fd_sc_hd__nand2_1
XFILLER_48_494 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
X_2002_ VSS VDD _1082_ _1403_ _1191_ _0095_ VDD VSS sky130_fd_sc_hd__o21a_1
XFILLER_50_136 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XFILLER_91_1 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
X_2904_ VSS VDD _0648_ _0796_ _0763_ VDD VSS sky130_fd_sc_hd__nand2_1
X_2835_ VSS VDD _0660_ _0730_ VDD VSS sky130_fd_sc_hd__clkbuf_2
X_2766_ VSS VDD _0660_ _0662_ _0661_ VDD VSS sky130_fd_sc_hd__nand2_1
X_2697_ VSS VDD core.osr.next_result_w\[16\] _0597_ _0533_ VDD VSS sky130_fd_sc_hd__nand2_1
X_1717_ VDD VSS _1247_ _1070_ VDD VSS sky130_fd_sc_hd__inv_2
XANTENNA__2479__B VSS VDD core.pdc.row_out_n\[12\] VDD VSS sky130_fd_sc_hd__diode_2
X_1648_ VDD VSS core.ndc.col_out\[8\] core.ndc.col_out_n\[8\] VDD VSS sky130_fd_sc_hd__inv_2
X_1579_ VDD VSS _1130_ _1125_ _1106_ _1121_ _1124_ core.ndc.col_out\[4\] VDD VSS sky130_fd_sc_hd__a221o_2
XANTENNA__2495__A VSS VDD _0208_ VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_92_29 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
Xgenblk1\[27\].buf_p_coln VSS VDD pmatrix_col_core_n_buffered\[27\] core.pdc.col_out_n\[27\]
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
XFILLER_89_361 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_66_41 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
XFILLER_66_85 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XFILLER_82_51 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
X_2620_ VSS VDD _0527_ _0529_ _0528_ VDD VSS sky130_fd_sc_hd__nand2_1
X_2551_ VSS VDD _0472_ _0475_ VDD VSS sky130_fd_sc_hd__clkbuf_2
X_2482_ VDD VSS _0433_ core.pdc.row_out_n\[15\] core.pdc.rowon_out_n\[15\] VDD VSS
+ sky130_fd_sc_hd__and2_1
X_1502_ VSS VDD _1053_ _1061_ _1062_ VDD VSS sky130_fd_sc_hd__nor2_1
X_1433_ VDD VSS _0997_ core.osr.sample_count_r\[0\] _0996_ VDD VSS sky130_fd_sc_hd__or2_1
XFILLER_101_108 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XFILLER_55_206 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
X_3103_ VSS VDD clknet_2_0__leaf_clk_dig_dummy _0003_ net85 core.cnb.is_holding_result_w
+ VDD VSS sky130_fd_sc_hd__dfrtp_1
X_3034_ VSS VDD _0915_ _0921_ _0922_ VDD VSS sky130_fd_sc_hd__nor2_1
XFILLER_23_103 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XFILLER_51_445 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XANTENNA__1612__A1 VSS VDD _1152_ VDD VSS sky130_fd_sc_hd__diode_2
X_2818_ VSS VDD _0697_ _0704_ _0713_ _0712_ VDD VSS sky130_fd_sc_hd__nand3_1
X_2749_ VSS VDD core.cnb.shift_register_r\[14\] _0645_ core.cnb.shift_register_r\[15\]
+ VDD VSS sky130_fd_sc_hd__nor2_2
XFILLER_11_69 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XFILLER_127_69 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
XFILLER_100_141 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XFILLER_86_342 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XANTENNA__1569__A VSS VDD _1101_ VDD VSS sky130_fd_sc_hd__diode_2
Xinput19 VDD VSS net19 config_2_in[10] VDD VSS sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__2566__C VSS VDD _1076_ VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_92_345 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
XFILLER_52_209 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XFILLER_92_378 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XANTENNA__1842__A1 VSS VDD _1325_ VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1479__A VSS VDD net15 VDD VSS sky130_fd_sc_hd__diode_2
X_1982_ VDD VSS _0079_ _0066_ VDD VSS sky130_fd_sc_hd__inv_2
Xgenblk1\[24\].buf_n_coln VSS VDD nmatrix_col_core_n_buffered\[24\] core.ndc.col_out_n\[24\]
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
X_2603_ VSS VDD _0033_ _0515_ VDD VSS sky130_fd_sc_hd__clkbuf_1
XFILLER_54_1 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
X_2534_ VSS VDD _0459_ net10 net54 core.cnb.sampled_avg_control_r\[2\] VDD VSS sky130_fd_sc_hd__mux2_1
X_2465_ VSS VDD _1338_ core.ndc.rowoff_out_n\[12\] _1325_ VDD VSS sky130_fd_sc_hd__nand2_1
X_2396_ VSS VDD _0394_ _0407_ _0406_ VDD VSS sky130_fd_sc_hd__nand2_1
X_1416_ VDD VSS core.cnb.pswitch_out\[1\] core.cnb.data_register_r\[1\] VDD VSS sky130_fd_sc_hd__inv_2
XANTENNA__1661__B VSS VDD _1202_ VDD VSS sky130_fd_sc_hd__diode_2
X_3017_ VDD VSS _0905_ _0904_ VDD VSS sky130_fd_sc_hd__inv_2
XANTENNA__2086__A1 VSS VDD _0101_ VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__2086__B2 VSS VDD _1096_ VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1833__A1 VSS VDD core.pdc.rowoff_out_n\[8\] VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__3170__RESET_B VSS VDD net73 VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_51_286 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_22_13 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XFILLER_93_109 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XFILLER_63_20 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XANTENNA__3026__B1 VSS VDD _1117_ VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA_genblk2\[0\].buf_n_rowonn_A VSS VDD core.ndc.rowon_out_n\[0\] VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1588__A0 VSS VDD _1133_ VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_6_132 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XANTENNA_genblk1\[12\].buf_n_coln_A VSS VDD core.ndc.col_out_n\[12\] VDD VSS sky130_fd_sc_hd__diode_2
X_2250_ VDD VSS core.osr.next_result_w\[4\] _0279_ VDD VSS sky130_fd_sc_hd__inv_2
XANTENNA__1762__A VSS VDD _1187_ VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_26_5 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XANTENNA__1481__B VSS VDD _1040_ VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__2577__B VSS VDD _1114_ VDD VSS sky130_fd_sc_hd__diode_2
X_2181_ VDD VSS _0220_ _0219_ VDD VSS sky130_fd_sc_hd__buf_2
XANTENNA__1512__A0 VSS VDD _1067_ VDD VSS sky130_fd_sc_hd__diode_2
X_1965_ VDD VSS _1121_ _1411_ core.pdc.col_out\[3\] _1125_ _1413_ _0067_ VDD VSS sky130_fd_sc_hd__a221o_1
XANTENNA__1579__B1 VSS VDD _1106_ VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__2532__S VSS VDD net54 VDD VSS sky130_fd_sc_hd__diode_2
X_1896_ VDD VSS _1369_ _1362_ VDD VSS sky130_fd_sc_hd__dlymetal6s2s_1
X_2517_ VSS VDD _0450_ core.cnb.shift_register_r\[12\] _0444_ core.cnb.shift_register_r\[11\]
+ VDD VSS sky130_fd_sc_hd__mux2_1
X_2448_ VSS VDD _1336_ _1385_ core.ndc.rowon_out_n\[9\] core.pdc.rowon_bottotop_n\[5\]
+ VDD VSS sky130_fd_sc_hd__a21oi_2
X_2379_ VSS VDD _1020_ _0393_ VDD VSS sky130_fd_sc_hd__clkbuf_2
XFILLER_83_164 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XFILLER_17_57 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XANTENNA__2008__A VSS VDD _1131_ VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_3_113 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_58_64 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XFILLER_66_109 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
XFILLER_47_312 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XFILLER_114_70 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
XFILLER_47_323 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_74_85 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_130_80 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XFILLER_90_73 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XANTENNA__1757__A VSS VDD _1272_ VDD VSS sky130_fd_sc_hd__diode_2
X_1750_ VSS VDD _1270_ _1269_ _1268_ _1267_ VDD VSS sky130_fd_sc_hd__and3_1
X_1681_ VSS VDD _1212_ _1219_ _1173_ VDD VSS sky130_fd_sc_hd__nand2_1
XANTENNA_nmat_col[0] VSS VDD core.ndc.col_out\[0\] VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA_nmat_analog_in VSS VDD ANTENNA_nmat_analog_in/DIODE VDD VSS sky130_fd_sc_hd__diode_2
X_2302_ VSS VDD _0323_ _0326_ _0325_ VDD VSS sky130_fd_sc_hd__nand2_1
X_2233_ VDD VSS _0264_ core.cnb.result_out\[3\] core.osr.result_r\[3\] VDD VSS sky130_fd_sc_hd__or2_1
X_2164_ VSS VDD _0207_ _0208_ _0204_ VDD VSS sky130_fd_sc_hd__nand2_4
XFILLER_93_473 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
X_2095_ VSS VDD _0065_ _0135_ _0156_ VDD VSS sky130_fd_sc_hd__nor2_1
XANTENNA__1667__A VSS VDD _1113_ VDD VSS sky130_fd_sc_hd__diode_2
X_2997_ VSS VDD _0056_ _0885_ _0781_ _0884_ _0886_ VDD VSS sky130_fd_sc_hd__a31o_1
X_1948_ VDD VSS core.pdc.col_out_n\[1\] core.pdc.col_out\[1\] VDD VSS sky130_fd_sc_hd__clkinv_2
X_1879_ VSS VDD _1348_ _1357_ core.pdc.row_out_n\[13\] _1336_ VDD VSS sky130_fd_sc_hd__a21oi_4
XFILLER_135_69 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_28_45 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_100_61 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
XFILLER_60_76 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XFILLER_47_153 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_85_84 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XFILLER_90_421 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
X_2920_ VSS VDD _0638_ _0708_ _0812_ VDD VSS sky130_fd_sc_hd__nor2_1
Xgenblk2\[14\].buf_n_rowonn VSS VDD nmatrix_rowon_core_n_buffered\[14\] core.ndc.rowon_out_n\[14\]
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
XFILLER_90_498 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
X_2851_ VDD VSS _0746_ core.cnb.shift_register_r\[9\] VDD VSS sky130_fd_sc_hd__inv_2
X_1802_ VDD VSS _1062_ core.ndc.col_out\[31\] _1126_ _1299_ _1251_ _1296_ VDD VSS
+ sky130_fd_sc_hd__a221o_4
X_2782_ VDD VSS _0678_ core.cnb.shift_register_r\[14\] VDD VSS sky130_fd_sc_hd__inv_2
X_1733_ VDD VSS core.ndc.col_out_n\[17\] _1258_ VDD VSS sky130_fd_sc_hd__buf_2
X_1664_ VSS VDD _1035_ _1198_ _1194_ _1075_ core.ndc.col_out_n\[9\] _1205_ VDD VSS
+ sky130_fd_sc_hd__o221a_2
XANTENNA__1934__B VSS VDD _1069_ VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_131_106 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
X_1595_ VSS VDD _1045_ _1145_ _1079_ VDD VSS sky130_fd_sc_hd__nand2_1
XANTENNA__2111__A VSS VDD _1413_ VDD VSS sky130_fd_sc_hd__diode_2
X_2216_ VDD VSS _0239_ _0248_ _0243_ _0249_ VDD VSS sky130_fd_sc_hd__or3_1
X_3196_ VSS VDD net63 core.osr.next_sample_count_w\[4\] net77 core.osr.sample_count_r\[4\]
+ VDD VSS sky130_fd_sc_hd__dfrtp_1
X_2147_ VSS VDD core.cnb.average_counter_r\[1\] _0191_ core.cnb.average_counter_r\[0\]
+ VDD VSS sky130_fd_sc_hd__nand2_1
XFILLER_93_281 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
X_2078_ VSS VDD _0065_ _0095_ _0147_ VDD VSS sky130_fd_sc_hd__nor2_1
XANTENNA__2434__A1 VSS VDD core.pdc.rowoff_out_n\[8\] VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__2434__B2 VSS VDD _1325_ VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1945__A0 VSS VDD _1069_ VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_107_125 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XANTENNA_fanout86_A VSS VDD net87 VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1860__A VSS VDD net14 VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_44_134 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
XFILLER_44_145 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XANTENNA_genblk2\[5\].buf_n_rowonn_A VSS VDD core.ndc.rowon_bottotop_n\[5\] VDD VSS
+ sky130_fd_sc_hd__diode_2
XFILLER_111_82 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
Xgenblk1\[29\].buf_n_coln VDD VSS core.ndc.col_out_n\[29\] nmatrix_col_core_n_buffered\[29\]
+ VDD VSS sky130_fd_sc_hd__buf_6
XANTENNA_clkbuf_0_clk_dig_dummy_A VSS VDD cgen/clk_dig_out VDD VSS sky130_fd_sc_hd__diode_2
X_3050_ VSS VDD _0877_ _0894_ _0938_ VDD VSS sky130_fd_sc_hd__nand2b_1
XFILLER_96_94 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XANTENNA__2585__B VSS VDD _1067_ VDD VSS sky130_fd_sc_hd__diode_2
X_2001_ VSS VDD _1162_ _1409_ _0094_ _1053_ VDD VSS sky130_fd_sc_hd__a21oi_2
XFILLER_90_273 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XFILLER_90_284 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
X_2903_ VDD VSS _0795_ _0784_ VDD VSS sky130_fd_sc_hd__inv_2
X_2834_ VSS VDD _0636_ _0728_ _0729_ VDD VSS sky130_fd_sc_hd__nor2_1
XANTENNA__3103__CLK VSS VDD clknet_2_0__leaf_clk_dig_dummy VDD VSS sky130_fd_sc_hd__diode_2
X_2765_ VSS VDD core.cnb.shift_register_r\[16\] _0638_ _0661_ VDD VSS sky130_fd_sc_hd__nor2_1
X_2696_ VSS VDD _0519_ _0356_ _0528_ _0596_ VDD VSS sky130_fd_sc_hd__o21a_1
X_1716_ VSS VDD _1164_ _1127_ _1246_ VDD VSS sky130_fd_sc_hd__nor2_1
X_1647_ VSS VDD _1190_ core.ndc.col_out_n\[8\] VDD VSS sky130_fd_sc_hd__clkbuf_2
XFILLER_116_49 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
X_1578_ VSS VDD _1126_ _1129_ _1130_ VDD VSS sky130_fd_sc_hd__nor2_1
Xgenblk1\[31\].buf_n_coln VDD VSS core.ndc.col_out_n\[31\] nmatrix_col_core_n_buffered\[31\]
+ VDD VSS sky130_fd_sc_hd__buf_6
X_3179_ VSS VDD net58 core.osr.next_result_w\[19\] net70 core.osr.result_r\[19\] VDD
+ VSS sky130_fd_sc_hd__dfrtp_1
XFILLER_54_421 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XFILLER_25_13 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_25_57 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XANTENNA__2016__A VSS VDD core.pdc.col_out_n\[9\] VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_89_373 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_49_215 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XFILLER_49_248 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
XANTENNA__1590__A VSS VDD _1131_ VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_66_97 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_122_81 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XANTENNA__3126__CLK VSS VDD clknet_2_2__leaf_clk_dig_dummy VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_32_137 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XANTENNA__1749__B VSS VDD _1177_ VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_82_85 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
X_2550_ VSS VDD core.cnb.data_register_r\[0\] _0473_ _0474_ VDD VSS sky130_fd_sc_hd__nor2_1
X_2481_ VSS VDD core.pdc.row_out_n\[14\] core.pdc.rowoff_out_n\[14\] core.pdc.rowon_out_n\[14\]
+ VDD VSS sky130_fd_sc_hd__nand2_1
X_1501_ VSS VDD _1054_ _1061_ _1060_ VDD VSS sky130_fd_sc_hd__nand2_1
X_1432_ VSS VDD _0992_ _0996_ _0995_ VDD VSS sky130_fd_sc_hd__nand2_1
X_3102_ VDD VSS core.cnb.is_sampling_w net84 _0002_ clknet_2_0__leaf_clk_dig_dummy
+ VDD VSS sky130_fd_sc_hd__dfstp_1
Xgenblk2\[2\].buf_p_rown VSS VDD pmatrix_row_core_n_buffered\[2\] core.pdc.row_out_n\[2\]
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
XFILLER_83_505 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
X_3033_ VSS VDD _0895_ _0920_ _0921_ VDD VSS sky130_fd_sc_hd__nor2_1
XFILLER_51_413 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_102_29 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XANTENNA__1675__A VSS VDD _1138_ VDD VSS sky130_fd_sc_hd__diode_2
X_2817_ VDD VSS _0712_ _0711_ VDD VSS sky130_fd_sc_hd__inv_2
X_2748_ VSS VDD core.cnb.shift_register_r\[13\] _0644_ core.cnb.shift_register_r\[12\]
+ VDD VSS sky130_fd_sc_hd__nor2_2
X_2679_ VDD VSS _1008_ _0367_ _0524_ _0581_ VDD VSS sky130_fd_sc_hd__a21oi_1
XFILLER_86_321 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
XFILLER_86_387 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XFILLER_77_52 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XANTENNA__2566__D VSS VDD _0482_ VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1842__A2 VSS VDD _1328_ VDD VSS sky130_fd_sc_hd__diode_2
X_1981_ VDD VSS core.pdc.col_out_n\[5\] core.pdc.col_out\[5\] VDD VSS sky130_fd_sc_hd__clkinv_2
XFILLER_61_3 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
X_2602_ VSS VDD _0515_ core.cnb.result_out\[11\] _0438_ _0514_ VDD VSS sky130_fd_sc_hd__mux2_1
X_2533_ VSS VDD _0020_ _0458_ VDD VSS sky130_fd_sc_hd__clkbuf_1
XFILLER_47_1 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
X_2464_ VSS VDD core.ndc.row_out_n\[11\] core.ndc.rowoff_out_n\[11\] core.ndc.rowon_out_n\[11\]
+ VDD VSS sky130_fd_sc_hd__nand2_1
X_2395_ VDD VSS _0406_ _0405_ VDD VSS sky130_fd_sc_hd__inv_2
XFILLER_3_60 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XFILLER_56_505 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
X_3016_ VSS VDD _0902_ _0904_ _0903_ VDD VSS sky130_fd_sc_hd__nand2_1
XANTENNA__2086__A2 VSS VDD _1173_ VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA_genblk2\[9\].buf_p_rowonn_A VSS VDD core.pdc.rowon_out_n\[9\] VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_51_298 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_22_25 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XFILLER_98_29 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
XANTENNA__2010__A2 VSS VDD _1395_ VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__2013__B VSS VDD _1101_ VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_47_505 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_47_88 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XFILLER_63_32 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XANTENNA__1588__A1 VSS VDD _1137_ VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_6_100 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XANTENNA__1762__B VSS VDD _1275_ VDD VSS sky130_fd_sc_hd__diode_2
X_2180_ VSS VDD _0208_ _0219_ VDD VSS sky130_fd_sc_hd__clkbuf_2
XANTENNA__1512__A1 VSS VDD _1069_ VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_74_891 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XANTENNA__1579__A1 VSS VDD _1121_ VDD VSS sky130_fd_sc_hd__diode_2
X_1964_ VSS VDD _0065_ _0066_ _0067_ VDD VSS sky130_fd_sc_hd__nor2_1
XANTENNA__1579__B2 VSS VDD _1125_ VDD VSS sky130_fd_sc_hd__diode_2
X_1895_ VSS VDD _1305_ core.ndc.rowon_bottotop_n\[5\] _1308_ VDD VSS sky130_fd_sc_hd__nor2_2
X_2516_ VSS VDD _0012_ _0449_ VDD VSS sky130_fd_sc_hd__clkbuf_1
X_2447_ VSS VDD _1374_ core.ndc.rowon_out_n\[8\] core.pdc.rowon_out_n\[15\] VDD VSS
+ sky130_fd_sc_hd__nand2_1
XFILLER_124_38 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
X_2378_ VSS VDD core.osr.next_result_w\[19\] _0392_ VDD VSS sky130_fd_sc_hd__clkbuf_1
XFILLER_17_25 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_83_154 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XFILLER_65_891 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XANTENNA__2008__B VSS VDD _0098_ VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_33_57 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_33_46 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
Xgenblk2\[1\].buf_p_rowonn VSS VDD pmatrix_rowon_core_n_buffered\[1\] core.pdc.rowon_out_n\[1\]
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
XFILLER_3_125 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XFILLER_109_3 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XANTENNA__1863__A VSS VDD _1347_ VDD VSS sky130_fd_sc_hd__diode_2
Xcgen VDD comp/clk cgen/clk_dig_out net18 net25 net26 net27 net28 net29 net30 net31
+ net32 net33 net19 net20 net21 net22 net23 net3 net4 net5 net6 net7 net8 core.cnb.enable_loop_out
+ net24 decision_finish_comp_n net54 sample_nmatrix_cgen net55 sample_pmatrix_cgen
+ net35 VSS adc_clkgen_with_edgedetect
XFILLER_87_471 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XANTENNA_input29_A VSS VDD config_2_in[5] VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_74_97 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_71_883 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XFILLER_128_134 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
XFILLER_128_123 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
X_1680_ VSS VDD _1217_ _1218_ _1152_ VDD VSS sky130_fd_sc_hd__nand2_1
X_2301_ VDD VSS _0325_ _0324_ VDD VSS sky130_fd_sc_hd__inv_2
X_2232_ VSS VDD _0261_ _0263_ _0257_ VDD VSS sky130_fd_sc_hd__nand2_1
X_2163_ VSS VDD _0205_ _0207_ _0206_ VDD VSS sky130_fd_sc_hd__nand2_1
XFILLER_80_113 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
X_2094_ VDD VSS core.pdc.col_out_n\[23\] core.pdc.col_out\[23\] VDD VSS sky130_fd_sc_hd__clkinv_2
XFILLER_62_883 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XFILLER_9_81 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XANTENNA__1667__B VSS VDD _1057_ VDD VSS sky130_fd_sc_hd__diode_2
X_2996_ VSS VDD _1113_ _0689_ _0886_ VDD VSS sky130_fd_sc_hd__nor2_1
X_1947_ VSS VDD _1259_ _1399_ _1397_ _1224_ core.pdc.col_out_n\[1\] _1402_ VDD VSS
+ sky130_fd_sc_hd__o221a_1
X_1878_ VSS VDD core.ndc.rowoff_out_n\[8\] _1314_ _1357_ VDD VSS sky130_fd_sc_hd__nor2_1
XANTENNA__1683__A VSS VDD _1220_ VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_88_246 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XFILLER_28_57 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_71_113 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XFILLER_125_148 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XFILLER_47_165 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XANTENNA__3032__B VSS VDD _1104_ VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_90_411 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
Xgenblk2\[7\].buf_p_rown VSS VDD pmatrix_row_core_n_buffered\[7\] core.pdc.row_out_n\[7\]
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
XFILLER_90_433 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XFILLER_90_455 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XFILLER_90_477 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
X_2850_ VSS VDD _0744_ _0731_ _0745_ _0725_ VDD VSS sky130_fd_sc_hd__nand3_1
X_1801_ VSS VDD _1272_ _1084_ _1299_ VDD VSS sky130_fd_sc_hd__nor2_1
X_2781_ VSS VDD _0666_ _0677_ _0676_ VDD VSS sky130_fd_sc_hd__nand2_1
X_1732_ VSS VDD _1258_ _1257_ _1256_ _1255_ VDD VSS sky130_fd_sc_hd__and3_1
XFILLER_116_126 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
X_1663_ VDD VSS _1205_ _1110_ _1204_ VDD VSS sky130_fd_sc_hd__or2_1
X_1594_ VSS VDD _1074_ _1143_ _1144_ VDD VSS sky130_fd_sc_hd__nor2_1
XANTENNA__2111__B VSS VDD _1101_ VDD VSS sky130_fd_sc_hd__diode_2
X_2215_ VSS VDD _0246_ _0248_ _0247_ VDD VSS sky130_fd_sc_hd__nand2_1
XFILLER_85_249 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
X_3195_ VSS VDD net63 core.osr.next_sample_count_w\[3\] net77 core.osr.sample_count_r\[3\]
+ VDD VSS sky130_fd_sc_hd__dfrtp_1
X_2146_ VDD VSS _0190_ core.cnb.average_counter_r\[3\] VDD VSS sky130_fd_sc_hd__inv_2
XANTENNA__2682__A2 VSS VDD core.osr.next_result_w\[8\] VDD VSS sky130_fd_sc_hd__diode_2
X_2077_ VDD VSS _0146_ _0111_ VDD VSS sky130_fd_sc_hd__inv_2
XANTENNA__3182__CLK VSS VDD clknet_2_1__leaf_clk_dig_dummy VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1678__A VSS VDD core.ndc.col_out_n\[10\] VDD VSS sky130_fd_sc_hd__diode_2
X_2979_ VSS VDD _0868_ _0870_ _0869_ VDD VSS sky130_fd_sc_hd__nand2_1
XFILLER_30_25 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XANTENNA__1945__A1 VSS VDD _1067_ VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1860__B VSS VDD core.cnb.data_register_r\[8\] VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_55_22 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
Xgenblk1\[2\].buf_p_coln VSS VDD pmatrix_col_core_n_buffered\[2\] core.pdc.col_out_n\[2\]
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
XANTENNA__1770__B VSS VDD _1095_ VDD VSS sky130_fd_sc_hd__diode_2
X_2000_ VDD VSS core.pdc.col_out_n\[7\] core.pdc.col_out\[7\] VDD VSS sky130_fd_sc_hd__clkinv_2
X_2902_ VSS VDD _0053_ _0794_ _0781_ _0793_ _1076_ _0688_ VDD VSS sky130_fd_sc_hd__a32o_1
X_2833_ VSS VDD _0668_ _0728_ _0637_ VDD VSS sky130_fd_sc_hd__nand2_1
XFILLER_77_1 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
X_2764_ VSS VDD _0646_ _0660_ _0659_ VDD VSS sky130_fd_sc_hd__nor2_2
X_1715_ VDD VSS core.ndc.col_out\[14\] core.ndc.col_out_n\[14\] VDD VSS sky130_fd_sc_hd__inv_2
X_2695_ VSS VDD _0593_ _0594_ _0045_ _0595_ VDD VSS sky130_fd_sc_hd__nand3_1
X_1646_ VSS VDD _1190_ _1189_ _1185_ _1181_ VDD VSS sky130_fd_sc_hd__and3_1
XANTENNA__2122__A VSS VDD _1396_ VDD VSS sky130_fd_sc_hd__diode_2
X_1577_ VSS VDD _1128_ _1127_ _1129_ _1082_ VDD VSS sky130_fd_sc_hd__a21oi_2
Xgenblk2\[4\].buf_n_rown VSS VDD nmatrix_row_core_n_buffered\[4\] core.ndc.row_out_n\[4\]
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
XANTENNA__1680__B VSS VDD _1152_ VDD VSS sky130_fd_sc_hd__diode_2
X_3178_ VSS VDD net58 core.osr.next_result_w\[18\] net69 core.osr.result_r\[18\] VDD
+ VSS sky130_fd_sc_hd__dfrtp_1
X_2129_ VDD VSS _1126_ _1393_ core.pdc.col_out\[31\] _1121_ _1391_ _0175_ VDD VSS
+ sky130_fd_sc_hd__a221o_1
XFILLER_25_25 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
XFILLER_25_69 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XANTENNA__3099__S VSS VDD _0241_ VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_41_57 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XANTENNA_input11_A VSS VDD config_1_in[3] VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_122_60 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XANTENNA__2207__A VSS VDD _0240_ VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__2582__A1 VSS VDD core.cnb.result_out\[6\] VDD VSS sky130_fd_sc_hd__diode_2
X_2480_ VSS VDD core.pdc.rowon_out_n\[13\] core.pdc.rowoff_out_n\[13\] core.pdc.row_out_n\[13\]
+ VDD VSS sky130_fd_sc_hd__nand2_1
XFILLER_56_6 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XANTENNA__2582__B2 VSS VDD _1104_ VDD VSS sky130_fd_sc_hd__diode_2
X_1500_ VSS VDD _1059_ _1060_ _1057_ VDD VSS sky130_fd_sc_hd__nor2_2
X_1431_ VSS VDD _0993_ _0994_ _0995_ VDD VSS sky130_fd_sc_hd__nor2_1
X_3101_ VSS VDD clknet_2_0__leaf_clk_dig_dummy core.cnb.next_conv_finished_w net84
+ net37 VDD VSS sky130_fd_sc_hd__dfrtp_1
XFILLER_55_219 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
X_3032_ VSS VDD _0917_ _1104_ _0920_ _0919_ VDD VSS sky130_fd_sc_hd__nand3_1
XFILLER_83_517 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XFILLER_51_425 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
X_2816_ VSS VDD _0710_ _0711_ _0664_ VDD VSS sky130_fd_sc_hd__nand2_1
XANTENNA__1956__A VSS VDD core.pdc.col_out\[2\] VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1675__B VSS VDD _1177_ VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_127_16 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
X_2747_ VSS VDD _0641_ _0643_ _0642_ VDD VSS sky130_fd_sc_hd__nand2_1
X_2678_ VSS VDD _0578_ _0579_ _0043_ _0580_ VDD VSS sky130_fd_sc_hd__nand3_1
X_1629_ VSS VDD _1085_ _1043_ _1118_ _1175_ VDD VSS sky130_fd_sc_hd__o21a_1
XANTENNA_input3_A VSS VDD config_1_in[10] VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_86_300 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XFILLER_46_219 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XFILLER_117_71 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XANTENNA_cgen_ena_in VSS VDD core.cnb.enable_loop_out VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_92_358 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
XFILLER_93_85 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
X_1980_ VSS VDD _1259_ _0076_ _0074_ _1224_ core.pdc.col_out_n\[5\] _0078_ VDD VSS
+ sky130_fd_sc_hd__o221a_1
XANTENNA__1776__A VSS VDD _1033_ VDD VSS sky130_fd_sc_hd__diode_2
X_2601_ VDD VSS _1309_ _0514_ _0513_ VDD VSS sky130_fd_sc_hd__xor2_1
X_2532_ VSS VDD _0458_ net9 net54 core.cnb.sampled_avg_control_r\[1\] VDD VSS sky130_fd_sc_hd__mux2_1
X_2463_ VSS VDD core.ndc.row_out_n\[10\] core.ndc.rowoff_out_n\[10\] core.ndc.rowon_out_n\[10\]
+ VDD VSS sky130_fd_sc_hd__nand2_1
X_2394_ VSS VDD _0403_ _0404_ _0405_ VDD VSS sky130_fd_sc_hd__nor2_1
XFILLER_56_517 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
X_3015_ VSS VDD _0901_ _0903_ _1312_ VDD VSS sky130_fd_sc_hd__nand2_1
XFILLER_83_325 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XFILLER_91_380 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_138_15 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XANTENNA_genblk1\[8\].buf_n_coln_A VSS VDD core.ndc.col_out_n\[8\] VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__2010__A3 VSS VDD _1085_ VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__3116__CLK VSS VDD clknet_2_2__leaf_clk_dig_dummy VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_47_517 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XANTENNA_fanout61_A VSS VDD net67 VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_6_112 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_88_85 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XANTENNA_genblk2\[13\].buf_p_rown_A VSS VDD core.pdc.row_out_n\[13\] VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_92_155 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
X_1963_ VSS VDD _0066_ _1170_ _1400_ _1145_ VDD VSS sky130_fd_sc_hd__mux2_1
X_1894_ VSS VDD core.pdc.rowon_out_n\[2\] _1366_ _1368_ VDD VSS sky130_fd_sc_hd__nand2_2
XANTENNA__1579__A2 VSS VDD _1124_ VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__2528__A1 VSS VDD net54 VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__3139__CLK VSS VDD clknet_2_0__leaf_clk_dig_dummy VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_108_29 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
X_2515_ VSS VDD _0449_ core.cnb.shift_register_r\[11\] _0444_ core.cnb.shift_register_r\[10\]
+ VDD VSS sky130_fd_sc_hd__mux2_1
X_2446_ VSS VDD core.ndc.rowon_out_n\[7\] _0429_ VDD VSS sky130_fd_sc_hd__clkbuf_1
XANTENNA__2130__A VSS VDD core.pdc.col_out\[31\] VDD VSS sky130_fd_sc_hd__diode_2
X_2377_ VSS VDD _0392_ _0391_ _0240_ _0390_ VDD VSS sky130_fd_sc_hd__and3_1
XFILLER_68_141 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
Xgenblk1\[7\].buf_p_coln VSS VDD pmatrix_col_core_n_buffered\[7\] core.pdc.col_out_n\[7\]
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
XFILLER_137_113 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_33_69 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XFILLER_58_77 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XANTENNA__2694__B VSS VDD core.cnb.result_out\[7\] VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__2455__B1 VSS VDD core.pdc.rowon_out_n\[0\] VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_23_91 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_99_95 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
X_2300_ VDD VSS _0315_ _0306_ _0314_ _0324_ VDD VSS sky130_fd_sc_hd__a21oi_1
X_2231_ VDD VSS _0252_ core.cnb.result_out\[2\] _0262_ core.osr.next_result_w\[2\]
+ VDD VSS sky130_fd_sc_hd__a21o_1
X_2162_ VSS VDD core.cnb.shift_register_r\[4\] core.cnb.shift_register_r\[5\] _0206_
+ VDD VSS sky130_fd_sc_hd__nor2_1
Xgenblk2\[9\].buf_n_rown VSS VDD nmatrix_row_core_n_buffered\[9\] core.ndc.row_out_n\[9\]
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
X_2093_ VSS VDD core.pdc.col_out_n\[23\] _0155_ VDD VSS sky130_fd_sc_hd__clkbuf_1
XFILLER_0_95 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_80_125 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
XANTENNA__3189__RESET_B VSS VDD net81 VDD VSS sky130_fd_sc_hd__diode_2
X_2995_ VSS VDD _0883_ _0885_ _0879_ VDD VSS sky130_fd_sc_hd__nand2_1
XFILLER_119_135 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
XFILLER_9_93 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XANTENNA__3118__RESET_B VSS VDD net86 VDD VSS sky130_fd_sc_hd__diode_2
X_1946_ VSS VDD _1401_ _1402_ _1155_ VDD VSS sky130_fd_sc_hd__nand2_1
X_1877_ VSS VDD _1356_ core.pdc.row_out_n\[12\] _1354_ VDD VSS sky130_fd_sc_hd__nor2_2
XANTENNA__1964__A VSS VDD _0065_ VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_0_107 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XFILLER_0_118 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XFILLER_88_214 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
X_2429_ VSS VDD _1342_ _1314_ _0426_ VDD VSS sky130_fd_sc_hd__nor2_1
XFILLER_28_69 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XANTENNA__2019__B VSS VDD _1135_ VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1858__B VSS VDD core.ndc.rowoff_out_n\[0\] VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_100_85 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_69_32 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
Xgenblk1\[4\].buf_n_coln VDD VSS core.ndc.col_out_n\[4\] nmatrix_col_core_n_buffered\[4\]
+ VDD VSS sky130_fd_sc_hd__buf_6
XFILLER_62_114 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
XFILLER_85_97 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
XFILLER_50_309 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XANTENNA__1768__B VSS VDD _1279_ VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1651__A1 VSS VDD _1077_ VDD VSS sky130_fd_sc_hd__diode_2
X_1800_ VDD VSS core.ndc.col_out\[30\] core.ndc.col_out_n\[30\] VDD VSS sky130_fd_sc_hd__clkinv_2
XFILLER_86_6 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
X_2780_ VDD VSS _0676_ _0675_ VDD VSS sky130_fd_sc_hd__inv_2
X_1731_ VSS VDD _1165_ _1257_ _1188_ VDD VSS sky130_fd_sc_hd__nand2_1
X_1662_ VSS VDD _1043_ _1203_ _1204_ _1199_ VDD VSS sky130_fd_sc_hd__o21ai_1
X_1593_ VSS VDD _1142_ _1103_ _1143_ _1141_ VDD VSS sky130_fd_sc_hd__o21ai_2
XFILLER_85_206 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
X_3194_ VSS VDD net62 core.osr.next_sample_count_w\[2\] net75 core.osr.sample_count_r\[2\]
+ VDD VSS sky130_fd_sc_hd__dfrtp_1
XFILLER_22_1 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
X_2214_ VSS VDD core.cnb.result_out\[1\] _0247_ core.osr.result_r\[1\] VDD VSS sky130_fd_sc_hd__nand2_1
X_2145_ VDD VSS _0179_ _0188_ _0189_ _0185_ VDD VSS sky130_fd_sc_hd__o21bai_1
XFILLER_53_103 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XFILLER_53_147 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
X_2076_ VDD VSS core.pdc.col_out_n\[19\] core.pdc.col_out\[19\] VDD VSS sky130_fd_sc_hd__clkinv_2
XFILLER_53_169 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
X_2978_ VSS VDD _0865_ _0866_ _0869_ _1114_ VDD VSS sky130_fd_sc_hd__nand3_1
X_1929_ VSS VDD _1387_ core.pdc.rowon_out_n\[15\] VDD VSS sky130_fd_sc_hd__clkbuf_2
XANTENNA__1694__A VSS VDD _1105_ VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_39_13 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_130_141 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XANTENNA__1869__A VSS VDD net14 VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_71_88 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XANTENNA__1936__A2 VSS VDD _1284_ VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_121_130 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XANTENNA__2649__B1 VSS VDD _0394_ VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_90_220 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XANTENNA__1779__A VSS VDD core.ndc.col_out\[25\] VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__3074__B1 VSS VDD _1312_ VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_90_253 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
X_2901_ VSS VDD _0792_ _0794_ _0791_ VDD VSS sky130_fd_sc_hd__nand2_1
X_2832_ VDD VSS _0727_ _0726_ VDD VSS sky130_fd_sc_hd__inv_2
X_2763_ VSS VDD _0659_ _0650_ _0641_ VDD VSS sky130_fd_sc_hd__nand2_2
X_1714_ VDD VSS core.ndc.col_out_n\[14\] _1245_ VDD VSS sky130_fd_sc_hd__buf_2
X_2694_ VSS VDD _0542_ _0595_ core.cnb.result_out\[7\] VDD VSS sky130_fd_sc_hd__nand2_1
X_1645_ VSS VDD _1187_ _1189_ _1188_ VDD VSS sky130_fd_sc_hd__nand2_1
XANTENNA__2122__B VSS VDD _1188_ VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_116_29 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
X_1576_ VSS VDD _1057_ _1128_ _1087_ VDD VSS sky130_fd_sc_hd__nor2_2
Xgenblk2\[10\].buf_n_rowonn VSS VDD nmatrix_rowon_core_n_buffered\[10\] core.ndc.rowon_out_n\[10\]
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
XANTENNA__1961__B VSS VDD _1088_ VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_112_141 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
X_3177_ VSS VDD net57 core.osr.next_result_w\[17\] net69 core.osr.result_r\[17\] VDD
+ VSS sky130_fd_sc_hd__dfrtp_1
XANTENNA__2792__B VSS VDD _0208_ VDD VSS sky130_fd_sc_hd__diode_2
X_2128_ VDD VSS _0175_ _1401_ _1092_ VDD VSS sky130_fd_sc_hd__and2_1
X_2059_ VSS VDD core.pdc.col_out_n\[15\] _0137_ VDD VSS sky130_fd_sc_hd__clkbuf_1
XFILLER_41_69 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XANTENNA__2967__B VSS VDD _1076_ VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_106_95 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_122_50 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
XFILLER_122_72 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
XANTENNA__1599__A VSS VDD _1148_ VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_15_81 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XANTENNA__2582__A2 VSS VDD _0439_ VDD VSS sky130_fd_sc_hd__diode_2
X_1430_ VSS VDD core.osr.osr_mode_r\[2\] _0990_ _0994_ VDD VSS sky130_fd_sc_hd__nor2_1
XANTENNA__3172__CLK VSS VDD net58 VDD VSS sky130_fd_sc_hd__diode_2
X_3100_ VSS VDD _0064_ _0981_ VDD VSS sky130_fd_sc_hd__clkbuf_1
X_3031_ VSS VDD _0918_ _0919_ _0916_ VDD VSS sky130_fd_sc_hd__nand2_1
XFILLER_51_437 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XANTENNA__2117__B VSS VDD _1235_ VDD VSS sky130_fd_sc_hd__diode_2
X_2815_ VSS VDD _0709_ _0660_ _0710_ _0661_ VDD VSS sky130_fd_sc_hd__nand3_1
XANTENNA__2133__A VSS VDD core.cnb.sampled_avg_control_r\[2\] VDD VSS sky130_fd_sc_hd__diode_2
X_2746_ VDD VSS _0642_ core.cnb.shift_register_r\[16\] VDD VSS sky130_fd_sc_hd__inv_2
X_2677_ VSS VDD core.osr.next_result_w\[5\] _0580_ _0542_ VDD VSS sky130_fd_sc_hd__nand2_1
XANTENNA__1972__A VSS VDD _0065_ VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1781__B1 VSS VDD _1035_ VDD VSS sky130_fd_sc_hd__diode_2
X_1628_ VSS VDD _1172_ _1174_ _1173_ VDD VSS sky130_fd_sc_hd__nand2_1
X_1559_ VDD VSS _1113_ core.cnb.data_register_r\[6\] VDD VSS sky130_fd_sc_hd__inv_2
XFILLER_86_367 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_14_128 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_77_21 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_93_97 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
X_2600_ VSS VDD _1328_ _0501_ _0513_ VDD VSS sky130_fd_sc_hd__nor2_1
X_2531_ VSS VDD _0019_ _0457_ VDD VSS sky130_fd_sc_hd__clkbuf_1
X_2462_ VSS VDD core.ndc.row_out_n\[9\] core.ndc.rowoff_out_n\[9\] core.ndc.rowon_out_n\[9\]
+ VDD VSS sky130_fd_sc_hd__nand2_1
X_2393_ VDD VSS _0404_ _0401_ VDD VSS sky130_fd_sc_hd__inv_2
XFILLER_3_95 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
X_3014_ VDD VSS _0902_ _1312_ _0901_ VDD VSS sky130_fd_sc_hd__or2_1
XFILLER_83_337 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_83_359 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
X_2729_ VSS VDD _0624_ _0626_ _0625_ VDD VSS sky130_fd_sc_hd__nand2_1
Xgenblk2\[7\].buf_n_rowonn VSS VDD nmatrix_rowon_core_n_buffered\[7\] core.ndc.rowon_out_n\[7\]
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
XANTENNA__2310__B VSS VDD _0255_ VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_47_46 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XFILLER_86_197 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XANTENNA_fanout54_A VSS VDD net55 VDD VSS sky130_fd_sc_hd__diode_2
Xgenblk1\[9\].buf_n_coln VDD VSS core.ndc.col_out_n\[9\] nmatrix_col_core_n_buffered\[9\]
+ VDD VSS sky130_fd_sc_hd__buf_6
XFILLER_137_1 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_6_124 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XFILLER_12_71 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_88_75 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XFILLER_88_97 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_92_167 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
X_1962_ VSS VDD _1110_ _0065_ VDD VSS sky130_fd_sc_hd__clkbuf_2
X_1893_ VDD VSS _1368_ _1367_ VDD VSS sky130_fd_sc_hd__inv_2
XANTENNA__1984__A0 VSS VDD _1118_ VDD VSS sky130_fd_sc_hd__diode_2
X_2514_ VSS VDD _0011_ _0448_ VDD VSS sky130_fd_sc_hd__clkbuf_1
X_2445_ VDD VSS _0429_ _1351_ _1364_ VDD VSS sky130_fd_sc_hd__or2_1
X_2376_ VSS VDD _0391_ core.osr.result_r\[18\] core.osr.result_r\[19\] _0384_ VDD
+ VSS sky130_fd_sc_hd__nand3b_1
XFILLER_56_337 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XFILLER_137_125 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_58_12 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XFILLER_47_337 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_114_95 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_139_81 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
X_2230_ VSS VDD _0262_ _0261_ _0260_ _0255_ VDD VSS sky130_fd_sc_hd__and3_1
X_2161_ VSS VDD core.cnb.shift_register_r\[2\] core.cnb.shift_register_r\[3\] _0205_
+ VDD VSS sky130_fd_sc_hd__nor2_1
XFILLER_93_421 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_65_134 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
X_2092_ VSS VDD _0155_ _0154_ _0153_ _0152_ VDD VSS sky130_fd_sc_hd__and3_1
XFILLER_0_41 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
X_2994_ VDD VSS _0884_ _0879_ _0883_ VDD VSS sky130_fd_sc_hd__or2_1
XANTENNA__3106__CLK VSS VDD clknet_2_2__leaf_clk_dig_dummy VDD VSS sky130_fd_sc_hd__diode_2
X_1945_ VSS VDD _1401_ _1067_ _1400_ _1069_ VDD VSS sky130_fd_sc_hd__mux2_1
XFILLER_119_29 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
X_1876_ VSS VDD _1311_ _1355_ _1356_ VDD VSS sky130_fd_sc_hd__nor2_1
X_2428_ VSS VDD _1334_ _1315_ core.ndc.row_out_n\[9\] VDD VSS sky130_fd_sc_hd__nor2_1
X_2359_ VDD VSS _0373_ _0377_ VDD VSS sky130_fd_sc_hd__buf_6
XFILLER_56_123 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XFILLER_52_351 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XFILLER_60_13 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_100_97 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_60_57 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XANTENNA__2051__A VSS VDD _1396_ VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA_input34_A VSS VDD rst_n VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_87_281 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_47_178 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XANTENNA__3129__CLK VSS VDD clknet_2_3__leaf_clk_dig_dummy VDD VSS sky130_fd_sc_hd__diode_2
X_1730_ VSS VDD _1100_ _1256_ _1213_ VDD VSS sky130_fd_sc_hd__nand2_1
X_1661_ VSS VDD _1043_ _1203_ _1202_ VDD VSS sky130_fd_sc_hd__nand2_1
X_1592_ VSS VDD _1103_ _1142_ _1112_ VDD VSS sky130_fd_sc_hd__nand2_1
X_3193_ VSS VDD net62 core.osr.next_sample_count_w\[1\] net75 core.osr.sample_count_r\[1\]
+ VDD VSS sky130_fd_sc_hd__dfrtp_1
X_2213_ VSS VDD _0244_ _0246_ _0245_ VDD VSS sky130_fd_sc_hd__nand2_1
X_2144_ VDD VSS _0188_ _0187_ VDD VSS sky130_fd_sc_hd__inv_2
X_2075_ VSS VDD core.pdc.col_out_n\[19\] _0145_ VDD VSS sky130_fd_sc_hd__clkbuf_1
XFILLER_53_159 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XANTENNA__2136__A VSS VDD core.cnb.sampled_avg_control_r\[2\] VDD VSS sky130_fd_sc_hd__diode_2
X_2977_ VSS VDD _0867_ _0868_ _1087_ VDD VSS sky130_fd_sc_hd__nand2_1
X_1928_ VDD VSS _1387_ _1038_ _1030_ VDD VSS sky130_fd_sc_hd__or2_1
XFILLER_30_38 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
X_1859_ VSS VDD _1325_ _1318_ _1344_ VDD VSS sky130_fd_sc_hd__nor2_1
XFILLER_122_109 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XFILLER_115_150 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XFILLER_130_153 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XANTENNA__2658__A1 VSS VDD core.osr.next_result_w\[3\] VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_44_126 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XFILLER_55_57 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XANTENNA__3083__A1 VSS VDD _0758_ VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_121_142 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XANTENNA__2649__A1 VSS VDD core.osr.next_result_w\[2\] VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_96_75 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XFILLER_35_137 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_90_232 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_90_265 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
X_2900_ VDD VSS _0793_ _0791_ _0792_ VDD VSS sky130_fd_sc_hd__or2_1
XANTENNA__1795__A VSS VDD _1272_ VDD VSS sky130_fd_sc_hd__diode_2
X_2831_ VSS VDD _0725_ _0723_ _0726_ _0724_ VDD VSS sky130_fd_sc_hd__nand3_2
X_2762_ VSS VDD _0206_ _0657_ _0658_ core.cnb.shift_register_r\[7\] VDD VSS sky130_fd_sc_hd__nand3_1
X_1713_ VSS VDD _1245_ _1244_ _1241_ _1239_ VDD VSS sky130_fd_sc_hd__and3_1
X_2693_ VSS VDD _0395_ _0594_ net40 VDD VSS sky130_fd_sc_hd__nand2_1
X_1644_ VDD VSS _1188_ _1032_ VDD VSS sky130_fd_sc_hd__buf_2
X_1575_ VSS VDD _1053_ _1042_ _1127_ VDD VSS sky130_fd_sc_hd__nor2_1
XFILLER_112_120 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
X_3176_ VSS VDD net56 core.osr.next_result_w\[16\] net68 core.osr.result_r\[16\] VDD
+ VSS sky130_fd_sc_hd__dfrtp_1
XFILLER_26_115 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
X_2127_ VDD VSS core.pdc.col_out_n\[30\] core.pdc.col_out\[30\] VDD VSS sky130_fd_sc_hd__clkinv_2
X_2058_ VSS VDD _0137_ _0136_ _0132_ _0130_ VDD VSS sky130_fd_sc_hd__and3_1
XANTENNA__3173__RESET_B VSS VDD net73 VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA_fanout84_A VSS VDD net85 VDD VSS sky130_fd_sc_hd__diode_2
Xgenblk2\[15\].buf_p_rowonn VSS VDD pmatrix_rowon_core_n_buffered\[15\] core.pdc.rowon_out_n\[15\]
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
XFILLER_106_85 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XANTENNA__1854__A2 VSS VDD _1340_ VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__3056__A1 VSS VDD _1312_ VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_82_99 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_31_92 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
X_3030_ VDD VSS _0918_ _0847_ VDD VSS sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_51_449 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_31_140 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
X_2814_ VSS VDD _0706_ _0709_ _0708_ VDD VSS sky130_fd_sc_hd__nand2_1
XFILLER_82_1 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
X_2745_ VSS VDD core.cnb.shift_register_r\[10\] core.cnb.shift_register_r\[11\] _0641_
+ VDD VSS sky130_fd_sc_hd__nor2_1
X_2676_ VSS VDD _0395_ _0579_ net53 VDD VSS sky130_fd_sc_hd__nand2_1
XANTENNA__1781__A1 VSS VDD _1259_ VDD VSS sky130_fd_sc_hd__diode_2
X_1627_ VSS VDD _1032_ _1173_ VDD VSS sky130_fd_sc_hd__clkbuf_2
XANTENNA__1972__B VSS VDD _0072_ VDD VSS sky130_fd_sc_hd__diode_2
X_1558_ VDD VSS _1112_ _1111_ VDD VSS sky130_fd_sc_hd__inv_2
X_1489_ VSS VDD _1037_ _1048_ _1049_ VDD VSS sky130_fd_sc_hd__nor2_1
XFILLER_86_379 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
X_3159_ VSS VDD net62 _0049_ net74 net44 VDD VSS sky130_fd_sc_hd__dfrtp_1
XANTENNA__2043__B VSS VDD _1163_ VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_117_51 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XFILLER_77_33 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XFILLER_93_65 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
X_2530_ VSS VDD _0457_ net2 net54 core.cnb.sampled_avg_control_r\[0\] VDD VSS sky130_fd_sc_hd__mux2_1
X_2461_ VSS VDD core.ndc.row_out_n\[7\] core.ndc.rowoff_out_n\[7\] core.ndc.rowon_out_n\[7\]
+ VDD VSS sky130_fd_sc_hd__nand2_1
X_2392_ VDD VSS _0403_ core.osr.sample_count_r\[3\] VDD VSS sky130_fd_sc_hd__inv_2
X_3013_ VSS VDD _0697_ _0900_ _0901_ _0847_ VDD VSS sky130_fd_sc_hd__o21ai_1
XFILLER_83_349 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XFILLER_77_891 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XANTENNA__2128__B VSS VDD _1092_ VDD VSS sky130_fd_sc_hd__diode_2
X_2728_ VSS VDD core.osr.next_result_w\[15\] _0625_ _0568_ VDD VSS sky130_fd_sc_hd__nand2_1
X_2659_ VDD VSS _0564_ _0563_ VDD VSS sky130_fd_sc_hd__inv_2
XANTENNA__2703__B1 VSS VDD core.osr.next_result_w\[8\] VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_86_154 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_68_891 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XANTENNA__2038__B VSS VDD _1095_ VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_128_61 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XFILLER_74_883 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
X_1961_ VSS VDD _1413_ _1412_ _1088_ VDD VSS sky130_fd_sc_hd__nand2_2
X_1892_ VSS VDD _1362_ _1029_ _1367_ VDD VSS sky130_fd_sc_hd__nor2_1
XANTENNA__1984__A1 VSS VDD _1112_ VDD VSS sky130_fd_sc_hd__diode_2
X_2513_ VSS VDD _0448_ core.cnb.shift_register_r\[10\] _0444_ core.cnb.shift_register_r\[9\]
+ VDD VSS sky130_fd_sc_hd__mux2_1
X_2444_ VDD VSS core.ndc.rowon_out_n\[6\] _0428_ VDD VSS sky130_fd_sc_hd__inv_2
XFILLER_124_19 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
X_2375_ VSS VDD _0390_ _0383_ core.osr.result_r\[18\] _0377_ core.osr.result_r\[19\]
+ VDD VSS sky130_fd_sc_hd__a31o_1
XFILLER_56_305 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XFILLER_17_17 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
XFILLER_52_500 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_65_883 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XANTENNA__3185__CLK VSS VDD clknet_2_1__leaf_clk_dig_dummy VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1672__B1 VSS VDD _1206_ VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_137_137 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XANTENNA__1975__A1 VSS VDD _1141_ VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_114_85 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
XFILLER_90_55 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_128_104 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XFILLER_23_71 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XFILLER_99_53 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XFILLER_99_86 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
Xclkbuf_0_clk_dig_dummy VSS VDD cgen/clk_dig_out clknet_0_clk_dig_dummy VDD VSS sky130_fd_sc_hd__clkbuf_16
X_2160_ VDD VSS _0204_ _0203_ VDD VSS sky130_fd_sc_hd__inv_2
XFILLER_17_5 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_48_90 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
X_2091_ VSS VDD _0096_ _0154_ _1101_ VDD VSS sky130_fd_sc_hd__nand2_1
XFILLER_93_433 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_0_53 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XFILLER_93_477 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_46_382 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XANTENNA__1798__A VSS VDD _1272_ VDD VSS sky130_fd_sc_hd__diode_2
X_2993_ VSS VDD _0882_ _0883_ _0868_ VDD VSS sky130_fd_sc_hd__nand2_1
XFILLER_9_40 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
X_1944_ VSS VDD _1388_ _1400_ VDD VSS sky130_fd_sc_hd__clkbuf_2
X_1875_ VDD VSS _1355_ _1024_ VDD VSS sky130_fd_sc_hd__inv_2
X_2427_ VSS VDD _1337_ core.ndc.row_out_n\[8\] core.pdc.rowoff_out_n\[0\] VDD VSS
+ sky130_fd_sc_hd__nand2_1
XFILLER_88_238 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
X_2358_ VDD VSS core.osr.next_result_w\[15\] _0376_ VDD VSS sky130_fd_sc_hd__inv_2
XFILLER_56_113 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
X_2289_ VSS VDD core.osr.result_r\[9\] core.cnb.result_out\[9\] _0314_ VDD VSS sky130_fd_sc_hd__nor2_1
XFILLER_60_25 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XANTENNA__2051__B VSS VDD _1152_ VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_107_3 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_109_85 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XFILLER_125_40 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XANTENNA_input27_A VSS VDD config_2_in[3] VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_87_293 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
XANTENNA__2242__A VSS VDD core.cnb.result_out\[4\] VDD VSS sky130_fd_sc_hd__diode_2
X_1660_ VDD VSS _1202_ _1201_ VDD VSS sky130_fd_sc_hd__inv_2
X_1591_ VDD VSS _1104_ _1105_ _1088_ _1141_ VDD VSS sky130_fd_sc_hd__a21o_1
XFILLER_124_151 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XANTENNA__2896__B VSS VDD _1076_ VDD VSS sky130_fd_sc_hd__diode_2
X_3192_ VDD VSS core.osr.sample_count_r\[0\] net74 core.osr.next_sample_count_w\[0\]
+ net62 VDD VSS sky130_fd_sc_hd__dfstp_1
X_2212_ VDD VSS _0245_ core.osr.result_r\[1\] VDD VSS sky130_fd_sc_hd__inv_2
X_2143_ VSS VDD _0176_ _0186_ _0187_ core.cnb.sampled_avg_control_r\[2\] VDD VSS sky130_fd_sc_hd__nand3_1
XFILLER_93_230 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XFILLER_93_241 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
X_2074_ VSS VDD _0145_ _0144_ _0143_ _0142_ VDD VSS sky130_fd_sc_hd__and3_1
XFILLER_14_29 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
X_2976_ VSS VDD _0865_ _0867_ _0866_ VDD VSS sky130_fd_sc_hd__nand2_1
X_1927_ VSS VDD core.pdc.rowon_out_n\[14\] core.ndc.rowon_out_n\[0\] _1386_ VDD VSS
+ sky130_fd_sc_hd__nand2_2
XFILLER_30_17 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
X_1858_ VSS VDD _1343_ core.pdc.row_out_n\[8\] core.ndc.rowoff_out_n\[0\] VDD VSS
+ sky130_fd_sc_hd__nand2_1
X_1789_ VDD VSS core.ndc.col_out_n\[27\] core.ndc.col_out\[27\] VDD VSS sky130_fd_sc_hd__clkinv_2
XANTENNA__1991__A VSS VDD core.pdc.col_out_n\[6\] VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_130_110 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_89_525 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XFILLER_55_36 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XFILLER_55_69 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XANTENNA__1885__B VSS VDD core.ndc.rowon_out_n\[0\] VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_29_81 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XFILLER_35_149 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XFILLER_90_244 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
Xgenblk2\[10\].buf_p_rown VSS VDD pmatrix_row_core_n_buffered\[10\] core.pdc.row_out_n\[10\]
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
X_2830_ VDD VSS _0725_ _0649_ VDD VSS sky130_fd_sc_hd__buf_2
X_2761_ VDD VSS _0657_ core.cnb.shift_register_r\[6\] VDD VSS sky130_fd_sc_hd__inv_2
X_2692_ VDD VSS _0588_ _0592_ _0593_ _0591_ VDD VSS sky130_fd_sc_hd__o21bai_1
X_1712_ VDD VSS _1244_ _1034_ _1243_ VDD VSS sky130_fd_sc_hd__or2_1
XFILLER_6_41 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
X_1643_ VSS VDD _1186_ _1113_ _1187_ _1043_ VDD VSS sky130_fd_sc_hd__o21ai_2
X_1574_ VDD VSS _1126_ _1110_ VDD VSS sky130_fd_sc_hd__buf_2
XFILLER_86_506 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_112_110 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
X_3175_ VSS VDD net58 core.osr.next_result_w\[15\] net70 core.osr.result_r\[15\] VDD
+ VSS sky130_fd_sc_hd__dfrtp_1
XFILLER_26_127 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
X_2126_ VSS VDD core.pdc.col_out_n\[30\] _0174_ VDD VSS sky130_fd_sc_hd__clkbuf_1
XFILLER_54_447 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
X_2057_ VDD VSS _0136_ _1034_ _0135_ VDD VSS sky130_fd_sc_hd__or2_1
XANTENNA__1986__A VSS VDD _1206_ VDD VSS sky130_fd_sc_hd__diode_2
X_2959_ VSS VDD _0776_ _0791_ _0851_ VDD VSS sky130_fd_sc_hd__nor2_1
XANTENNA__3142__RESET_B VSS VDD net81 VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__3119__CLK VSS VDD clknet_2_0__leaf_clk_dig_dummy VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_106_53 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XFILLER_106_64 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XFILLER_66_57 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XFILLER_17_149 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XANTENNA__2057__A VSS VDD _1034_ VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_122_85 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_40_141 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XFILLER_31_152 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
X_2813_ VSS VDD _0707_ _0708_ _0206_ VDD VSS sky130_fd_sc_hd__nand2_1
XANTENNA__2007__A0 VSS VDD _1161_ VDD VSS sky130_fd_sc_hd__diode_2
X_2744_ VDD VSS _0639_ _0640_ VDD VSS sky130_fd_sc_hd__buf_6
X_2675_ VDD VSS _0573_ _0577_ _0578_ _0576_ VDD VSS sky130_fd_sc_hd__o21bai_1
XANTENNA__1781__A2 VSS VDD _1220_ VDD VSS sky130_fd_sc_hd__diode_2
X_1626_ VDD VSS _1172_ _1171_ VDD VSS sky130_fd_sc_hd__inv_2
X_1557_ VSS VDD _1085_ _1065_ _1111_ VDD VSS sky130_fd_sc_hd__nor2_1
XFILLER_98_141 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
X_1488_ VSS VDD _1043_ _1048_ _1047_ VDD VSS sky130_fd_sc_hd__nand2_1
X_3158_ VSS VDD net60 _0048_ net74 net43 VDD VSS sky130_fd_sc_hd__dfrtp_1
XFILLER_36_49 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
X_2109_ VDD VSS _0161_ _0162_ VDD VSS sky130_fd_sc_hd__clkinv_2
X_3089_ VSS VDD _0966_ _0973_ _0974_ _0969_ VDD VSS sky130_fd_sc_hd__nand3_1
XFILLER_22_130 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XANTENNA__2978__C VSS VDD _1114_ VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_93_77 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
XANTENNA_genblk2\[2\].buf_n_rown_A VSS VDD core.ndc.row_out_n\[2\] VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1565__S VSS VDD _1077_ VDD VSS sky130_fd_sc_hd__diode_2
X_2460_ VSS VDD core.ndc.row_out_n\[6\] core.ndc.rowoff_out_n\[6\] core.ndc.rowon_out_n\[6\]
+ VDD VSS sky130_fd_sc_hd__nand2_1
X_2391_ VDD VSS core.osr.next_sample_count_w\[2\] _0402_ VDD VSS sky130_fd_sc_hd__inv_2
XFILLER_3_53 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XANTENNA_nmat_en_bit_n[2] VSS VDD core.cnb.pswitch_out\[2\] VDD VSS sky130_fd_sc_hd__diode_2
X_3012_ VSS VDD _0799_ _0900_ _0697_ VDD VSS sky130_fd_sc_hd__nand2_1
XFILLER_51_214 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XFILLER_51_225 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_22_29 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_138_29 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
X_2727_ VSS VDD core.osr.next_result_w\[17\] _0624_ _1002_ VDD VSS sky130_fd_sc_hd__nand2_1
XANTENNA__1983__B VSS VDD _1279_ VDD VSS sky130_fd_sc_hd__diode_2
X_2658_ VDD VSS _0393_ core.osr.next_result_w\[3\] _0562_ _0563_ net51 VDD VSS sky130_fd_sc_hd__a22o_1
X_1609_ VSS VDD _1076_ _1156_ _1145_ _1157_ VDD VSS sky130_fd_sc_hd__o21a_1
X_2589_ VSS VDD _0503_ _0505_ _0504_ VDD VSS sky130_fd_sc_hd__nand2_1
XFILLER_47_26 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_86_133 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
XANTENNA_input1_A VSS VDD clk_vcm VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_103_43 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
Xgenblk1\[11\].buf_p_coln VSS VDD pmatrix_col_core_n_buffered\[11\] core.pdc.col_out_n\[11\]
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
XFILLER_5_1 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XFILLER_88_44 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_37_81 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
X_1960_ VSS VDD _1409_ _1412_ _1036_ VDD VSS sky130_fd_sc_hd__nand2_1
XFILLER_53_91 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
X_1891_ VDD VSS _1366_ _1365_ VDD VSS sky130_fd_sc_hd__inv_2
X_2512_ VSS VDD _0010_ _0447_ VDD VSS sky130_fd_sc_hd__clkbuf_1
XFILLER_52_3 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
X_2443_ VSS VDD _1379_ _0428_ _1368_ VDD VSS sky130_fd_sc_hd__nand2_1
X_2374_ VSS VDD core.osr.next_result_w\[18\] _0389_ VDD VSS sky130_fd_sc_hd__clkbuf_1
XFILLER_83_169 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XFILLER_52_512 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_137_105 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
XFILLER_137_149 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
XANTENNA_genblk1\[19\].buf_n_coln_A VSS VDD core.ndc.col_out_n\[19\] VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_87_497 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XFILLER_55_361 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XFILLER_74_57 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
Xgenblk2\[3\].buf_n_rowonn VSS VDD nmatrix_rowon_core_n_buffered\[3\] core.ndc.rowon_out_n\[3\]
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
XANTENNA__2065__A VSS VDD _0065_ VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_130_85 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
Xgenblk2\[15\].buf_p_rown VSS VDD pmatrix_row_core_n_buffered\[15\] core.pdc.row_out_n\[15\]
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
XFILLER_90_67 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XFILLER_23_83 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
X_2090_ VSS VDD _0139_ _0153_ _1235_ VDD VSS sky130_fd_sc_hd__nand2_1
XFILLER_93_445 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XFILLER_46_350 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
XFILLER_46_361 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XFILLER_93_489 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
X_2992_ VSS VDD _0863_ _0882_ _0881_ VDD VSS sky130_fd_sc_hd__nand2_1
XFILLER_9_52 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XANTENNA_genblk1\[9\].buf_p_coln_A VSS VDD core.pdc.col_out_n\[9\] VDD VSS sky130_fd_sc_hd__diode_2
X_1943_ VDD VSS _1399_ _1398_ VDD VSS sky130_fd_sc_hd__inv_2
X_1874_ VSS VDD core.ndc.rowoff_out_n\[8\] _1349_ _1354_ VDD VSS sky130_fd_sc_hd__nor2_1
XANTENNA__1753__S VSS VDD _1034_ VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_88_206 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
X_2426_ VSS VDD _1343_ core.ndc.row_out_n\[7\] _1361_ VDD VSS sky130_fd_sc_hd__nand2_1
XFILLER_88_228 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
X_2357_ VSS VDD _0369_ _0376_ _0375_ VDD VSS sky130_fd_sc_hd__nand2_1
X_2288_ VDD VSS _0313_ core.osr.next_result_w\[8\] _0252_ _0312_ VDD VSS sky130_fd_sc_hd__o21ai_4
XFILLER_84_445 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XANTENNA__3167__RESET_B VSS VDD net73 VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_56_169 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
XFILLER_44_49 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XANTENNA__1501__B VSS VDD _1060_ VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_100_33 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XFILLER_109_97 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_125_52 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XANTENNA__1899__A VSS VDD _1371_ VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_90_404 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XANTENNA__3175__CLK VSS VDD net58 VDD VSS sky130_fd_sc_hd__diode_2
X_1590_ VSS VDD _1131_ _1139_ _1140_ VDD VSS sky130_fd_sc_hd__nor2_1
X_2211_ VDD VSS _0244_ core.cnb.result_out\[1\] VDD VSS sky130_fd_sc_hd__inv_2
X_3191_ VDD VSS core.cnb.data_register_r\[11\] net82 _0061_ clknet_2_1__leaf_clk_dig_dummy
+ VDD VSS sky130_fd_sc_hd__dfstp_2
X_2142_ VDD VSS _0186_ core.cnb.sampled_avg_control_r\[0\] VDD VSS sky130_fd_sc_hd__inv_2
XFILLER_38_114 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_93_253 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
X_2073_ VDD VSS _0144_ _1033_ _0113_ VDD VSS sky130_fd_sc_hd__or2_1
Xgenblk2\[12\].buf_n_rown VSS VDD nmatrix_row_core_n_buffered\[12\] core.ndc.row_out_n\[12\]
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
XFILLER_46_191 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
X_2975_ VSS VDD _0795_ _0866_ _0864_ VDD VSS sky130_fd_sc_hd__nand2_1
X_1926_ VSS VDD _1385_ _1386_ _1027_ VDD VSS sky130_fd_sc_hd__nand2_1
XFILLER_30_29 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
X_1857_ VDD VSS _1342_ _1024_ _1336_ _1343_ VDD VSS sky130_fd_sc_hd__a21o_1
X_1788_ VSS VDD core.ndc.col_out_n\[27\] _1293_ VDD VSS sky130_fd_sc_hd__clkbuf_1
XFILLER_130_122 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_39_49 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
X_2409_ VSS VDD _0414_ _0417_ core.osr.sample_count_r\[6\] VDD VSS sky130_fd_sc_hd__nand2_1
XFILLER_44_106 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_71_14 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_106_152 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XFILLER_48_401 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XFILLER_48_434 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XFILLER_48_445 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XFILLER_29_93 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XANTENNA__1609__A1 VSS VDD _1076_ VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_84_6 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XANTENNA__2253__A VSS VDD core.cnb.result_out\[5\] VDD VSS sky130_fd_sc_hd__diode_2
X_2760_ VSS VDD _0648_ _0656_ _0655_ VDD VSS sky130_fd_sc_hd__nand2_1
X_2691_ VSS VDD core.osr.next_result_w\[9\] _1019_ _0592_ _0537_ VDD VSS sky130_fd_sc_hd__o21ai_1
X_1711_ VSS VDD _1243_ _1202_ _1054_ _1242_ VDD VSS sky130_fd_sc_hd__mux2_1
XANTENNA__3068__B VSS VDD _0799_ VDD VSS sky130_fd_sc_hd__diode_2
X_1642_ VSS VDD _1116_ _1186_ _1117_ VDD VSS sky130_fd_sc_hd__nor2_2
XFILLER_6_53 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
X_1573_ VSS VDD _1095_ _1125_ VDD VSS sky130_fd_sc_hd__clkbuf_2
XANTENNA__3084__A VSS VDD _1022_ VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_86_518 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
X_3174_ VSS VDD net58 core.osr.next_result_w\[14\] net70 core.osr.result_r\[14\] VDD
+ VSS sky130_fd_sc_hd__dfrtp_1
X_2125_ VSS VDD _0174_ _0173_ _0171_ _0170_ VDD VSS sky130_fd_sc_hd__and3_1
X_2056_ VSS VDD _1242_ _0134_ _0135_ VDD VSS sky130_fd_sc_hd__nor2_1
XFILLER_41_109 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
X_2958_ VSS VDD _0849_ _0850_ _0755_ VDD VSS sky130_fd_sc_hd__nand2_1
Xgenblk1\[16\].buf_p_coln VSS VDD pmatrix_col_core_n_buffered\[16\] core.pdc.col_out_n\[16\]
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
X_1909_ VSS VDD _1340_ core.pdc.rowon_out_n\[7\] core.pdc.rowoff_out_n\[8\] VDD VSS
+ sky130_fd_sc_hd__nand2_1
X_2889_ VSS VDD _0052_ _0782_ _0781_ _0780_ _0482_ _0758_ VDD VSS sky130_fd_sc_hd__a32o_1
XFILLER_103_122 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XANTENNA__3182__RESET_B VSS VDD net86 VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_106_76 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XFILLER_122_97 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_15_40 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XANTENNA__2073__A VSS VDD _1033_ VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1417__A VSS VDD core.cnb.data_register_r\[0\] VDD VSS sky130_fd_sc_hd__diode_2
Xoutput50 VDD VSS result_out[6] net50 VDD VSS sky130_fd_sc_hd__buf_2
XFILLER_48_286 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
X_2812_ VSS VDD core.cnb.shift_register_r\[7\] _0657_ _0707_ VDD VSS sky130_fd_sc_hd__nor2_1
XFILLER_72_90 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XANTENNA__2007__A1 VSS VDD _1229_ VDD VSS sky130_fd_sc_hd__diode_2
X_2743_ VSS VDD _0636_ _0638_ _0639_ VDD VSS sky130_fd_sc_hd__nor2_1
XFILLER_68_1 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
X_2674_ VSS VDD core.osr.next_result_w\[7\] _1019_ _0577_ _0537_ VDD VSS sky130_fd_sc_hd__o21ai_1
X_1625_ VSS VDD _1156_ _1171_ _1170_ VDD VSS sky130_fd_sc_hd__nand2_1
X_1556_ VDD VSS _1110_ _1039_ VDD VSS sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_100_125 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
X_1487_ VSS VDD _1046_ _1047_ _1044_ VDD VSS sky130_fd_sc_hd__nor2_2
X_3157_ VSS VDD net59 _0047_ net72 net42 VDD VSS sky130_fd_sc_hd__dfrtp_1
X_2108_ VSS VDD _1131_ _0091_ _0161_ VDD VSS sky130_fd_sc_hd__nor2_1
X_3088_ VDD VSS _0973_ _0971_ VDD VSS sky130_fd_sc_hd__inv_2
XANTENNA__1997__A VSS VDD _0091_ VDD VSS sky130_fd_sc_hd__diode_2
X_2039_ VSS VDD _0122_ _0121_ _0119_ _0117_ VDD VSS sky130_fd_sc_hd__and3_1
XFILLER_52_16 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_50_462 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_89_120 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
XFILLER_77_57 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XFILLER_92_329 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XANTENNA__1700__A VSS VDD _1034_ VDD VSS sky130_fd_sc_hd__diode_2
Xgenblk1\[13\].buf_n_coln VDD VSS core.ndc.col_out_n\[13\] nmatrix_col_core_n_buffered\[13\]
+ VDD VSS sky130_fd_sc_hd__buf_6
XFILLER_9_113 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XANTENNA__1996__B1 VSS VDD _1045_ VDD VSS sky130_fd_sc_hd__diode_2
Xgenblk2\[11\].buf_p_rowonn VSS VDD pmatrix_rowon_core_n_buffered\[11\] core.pdc.rowon_out_n\[11\]
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
XFILLER_3_21 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
X_2390_ VDD VSS _0401_ core.osr.is_last_sample _0400_ _0402_ VDD VSS sky130_fd_sc_hd__or3_1
XANTENNA_nmat_en_bit_n[1] VSS VDD core.cnb.pswitch_out\[1\] VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_3_87 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XANTENNA__3081__B VSS VDD _0691_ VDD VSS sky130_fd_sc_hd__diode_2
X_3011_ VSS VDD _0689_ _0899_ _0057_ _1053_ VDD VSS sky130_fd_sc_hd__o21ai_1
XFILLER_91_351 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XANTENNA__3109__CLK VSS VDD clknet_2_3__leaf_clk_dig_dummy VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA_genblk2\[7\].buf_p_rown_A VSS VDD core.pdc.row_out_n\[7\] VDD VSS sky130_fd_sc_hd__diode_2
X_2726_ VSS VDD core.osr.next_result_w\[19\] _0623_ _0533_ VDD VSS sky130_fd_sc_hd__nand2_1
XANTENNA__2441__A VSS VDD core.pdc.rowon_bottotop_n\[5\] VDD VSS sky130_fd_sc_hd__diode_2
X_2657_ VSS VDD _0983_ _0562_ VDD VSS sky130_fd_sc_hd__clkbuf_2
X_1608_ VSS VDD _1043_ _1156_ _1045_ VDD VSS sky130_fd_sc_hd__nand2_1
X_2588_ VSS VDD _0501_ _0504_ _1300_ VDD VSS sky130_fd_sc_hd__nand2_1
X_1539_ VSS VDD _1072_ _1095_ VDD VSS sky130_fd_sc_hd__clkbuf_2
XFILLER_103_11 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_103_66 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XANTENNA__1520__A VSS VDD _1077_ VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_10_134 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
XFILLER_128_85 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_88_34 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
XFILLER_88_56 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XFILLER_37_93 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
X_1890_ VSS VDD _1338_ _1028_ _1365_ VDD VSS sky130_fd_sc_hd__nor2_1
XANTENNA__2261__A VSS VDD core.cnb.result_out\[6\] VDD VSS sky130_fd_sc_hd__diode_2
X_2511_ VSS VDD _0447_ core.cnb.shift_register_r\[9\] _0444_ core.cnb.shift_register_r\[8\]
+ VDD VSS sky130_fd_sc_hd__mux2_1
X_2442_ VSS VDD core.ndc.rowoff_out_n\[5\] core.ndc.rowon_out_n\[4\] _1311_ VDD VSS
+ sky130_fd_sc_hd__nand2_1
X_2373_ VSS VDD _0389_ _0240_ _0388_ _0387_ VDD VSS sky130_fd_sc_hd__and3_1
XFILLER_83_137 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XFILLER_52_524 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XFILLER_91_181 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
X_2709_ VSS VDD _0363_ _1011_ _0608_ _0518_ VDD VSS sky130_fd_sc_hd__o21ai_1
XANTENNA__1515__A VSS VDD _1072_ VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_74_115 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XFILLER_74_69 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_90_13 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XFILLER_135_1 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
XFILLER_46_395 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
X_2991_ VDD VSS _0881_ _0880_ VDD VSS sky130_fd_sc_hd__inv_2
X_1942_ VSS VDD _1398_ _1098_ _1394_ _1067_ VDD VSS sky130_fd_sc_hd__mux2_1
X_1873_ VDD VSS core.pdc.row_out_n\[11\] _1353_ VDD VSS sky130_fd_sc_hd__inv_2
Xgenblk2\[8\].buf_p_rowonn VSS VDD pmatrix_rowon_core_n_buffered\[8\] core.pdc.rowon_out_n\[8\]
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
XFILLER_134_109 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
X_2425_ VDD VSS core.ndc.row_out_n\[6\] _0425_ VDD VSS sky130_fd_sc_hd__inv_2
X_2356_ VDD VSS _0375_ _0374_ VDD VSS sky130_fd_sc_hd__inv_2
X_2287_ VSS VDD _0252_ _0313_ core.cnb.result_out\[8\] VDD VSS sky130_fd_sc_hd__nand2_1
XFILLER_71_107 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XFILLER_109_32 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_47_104 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XANTENNA__2530__A0 VSS VDD core.cnb.sampled_avg_control_r\[0\] VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_87_262 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
Xgenblk1\[23\].buf_p_coln VSS VDD pmatrix_col_core_n_buffered\[23\] core.pdc.col_out_n\[23\]
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
XFILLER_18_95 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XFILLER_109_150 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XANTENNA_genblk1\[0\].buf_n_coln_A VSS VDD core.ndc.col_out_n\[0\] VDD VSS sky130_fd_sc_hd__diode_2
X_2210_ VDD VSS _0243_ core.osr.result_r\[0\] VDD VSS sky130_fd_sc_hd__inv_2
X_3190_ VSS VDD clknet_2_1__leaf_clk_dig_dummy _0060_ net81 core.cnb.data_register_r\[10\]
+ VDD VSS sky130_fd_sc_hd__dfrtp_2
X_2141_ VDD VSS _0184_ _0183_ _0177_ _0185_ VDD VSS sky130_fd_sc_hd__a21oi_1
XFILLER_38_126 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_93_265 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
X_2072_ VSS VDD _0084_ _0143_ _1275_ VDD VSS sky130_fd_sc_hd__nand2_1
X_2974_ VDD VSS _0472_ _0783_ _0864_ _0865_ VDD VSS sky130_fd_sc_hd__a21o_1
X_1925_ VSS VDD _1029_ _1385_ _1023_ VDD VSS sky130_fd_sc_hd__nand2_1
X_1856_ VDD VSS _1342_ _1301_ VDD VSS sky130_fd_sc_hd__buf_2
X_1787_ VSS VDD _1293_ _1292_ _1291_ _1290_ VDD VSS sky130_fd_sc_hd__and3_1
XFILLER_115_142 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XFILLER_89_505 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_130_134 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
XFILLER_39_28 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
X_2408_ VSS VDD core.osr.sample_count_r\[6\] _0414_ _0416_ VDD VSS sky130_fd_sc_hd__nor2_1
X_2339_ VDD VSS _0360_ _0359_ _0271_ VDD VSS sky130_fd_sc_hd__and2_1
XFILLER_29_137 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_44_118 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XFILLER_111_11 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XFILLER_71_26 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XANTENNA__2579__B1 VSS VDD core.cnb.result_out\[5\] VDD VSS sky130_fd_sc_hd__diode_2
Xgenblk1\[18\].buf_n_coln VDD VSS core.ndc.col_out_n\[18\] nmatrix_col_core_n_buffered\[18\]
+ VDD VSS sky130_fd_sc_hd__buf_6
XFILLER_20_41 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XFILLER_106_131 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
XFILLER_136_41 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_20_85 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
XFILLER_136_85 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XANTENNA__1857__A2 VSS VDD _1342_ VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA_input32_A VSS VDD config_2_in[8] VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__3142__CLK VSS VDD clknet_2_1__leaf_clk_dig_dummy VDD VSS sky130_fd_sc_hd__diode_2
X_2690_ VSS VDD _0589_ _0591_ _0590_ VDD VSS sky130_fd_sc_hd__nand2_1
XFILLER_61_81 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
X_1710_ VSS VDD _1060_ _1242_ _1117_ VDD VSS sky130_fd_sc_hd__nor2_2
X_1641_ VDD VSS _1184_ _1185_ VDD VSS sky130_fd_sc_hd__clkinv_2
XFILLER_6_65 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
X_1572_ VSS VDD _1124_ _1068_ _1078_ _1123_ VDD VSS sky130_fd_sc_hd__o21a_2
XFILLER_112_134 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
Xgenblk1\[20\].buf_n_coln VSS VDD nmatrix_col_core_n_buffered\[20\] core.ndc.col_out_n\[20\]
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
X_3173_ VSS VDD net61 core.osr.next_result_w\[13\] net73 core.osr.result_r\[13\] VDD
+ VSS sky130_fd_sc_hd__dfrtp_1
XANTENNA__1613__A VSS VDD core.ndc.col_out\[6\] VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_13_1 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
X_2124_ VDD VSS _0172_ _0173_ VDD VSS sky130_fd_sc_hd__clkinv_2
X_2055_ VDD VSS _0134_ _0133_ VDD VSS sky130_fd_sc_hd__inv_2
XANTENNA__2444__A VSS VDD _0428_ VDD VSS sky130_fd_sc_hd__diode_2
X_2957_ VSS VDD _0846_ core.cnb.data_register_r\[1\] _0849_ _0848_ VDD VSS sky130_fd_sc_hd__nand3_1
X_2888_ VSS VDD _0779_ _0782_ _0777_ VDD VSS sky130_fd_sc_hd__nand2_1
X_1908_ VSS VDD core.pdc.rowon_out_n\[6\] _1377_ VDD VSS sky130_fd_sc_hd__clkbuf_1
X_1839_ VDD VSS _1327_ _1328_ VDD VSS sky130_fd_sc_hd__clkinv_2
XFILLER_103_101 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XFILLER_103_134 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
Xclkbuf_2_3__f_clk_dig_dummy VSS VDD clknet_0_clk_dig_dummy clknet_2_3__leaf_clk_dig_dummy
+ VDD VSS sky130_fd_sc_hd__clkbuf_16
XFILLER_66_15 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_17_129 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XFILLER_15_52 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XANTENNA__2073__B VSS VDD _0113_ VDD VSS sky130_fd_sc_hd__diode_2
Xoutput51 VDD VSS result_out[7] net51 VDD VSS sky130_fd_sc_hd__buf_2
Xoutput40 VDD VSS result_out[11] net40 VDD VSS sky130_fd_sc_hd__buf_2
X_2811_ VSS VDD _0635_ core.cnb.shift_register_r\[4\] _0706_ _0705_ VDD VSS sky130_fd_sc_hd__nand3_1
X_2742_ VSS VDD _0638_ _0205_ _0637_ VDD VSS sky130_fd_sc_hd__nand2_2
X_2673_ VSS VDD _0574_ _0576_ _0575_ VDD VSS sky130_fd_sc_hd__nand2_1
X_1624_ VSS VDD _1169_ _1170_ _1045_ VDD VSS sky130_fd_sc_hd__nand2_1
X_1555_ VSS VDD _1088_ _1037_ _1109_ _1103_ VDD VSS sky130_fd_sc_hd__o21ai_2
X_1486_ VDD VSS _1046_ _1045_ VDD VSS sky130_fd_sc_hd__inv_2
XFILLER_100_137 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
X_3156_ VSS VDD net59 _0046_ net71 net41 VDD VSS sky130_fd_sc_hd__dfrtp_1
XANTENNA__3188__CLK VSS VDD clknet_2_1__leaf_clk_dig_dummy VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_54_235 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
X_3087_ VSS VDD _0970_ _0972_ _0971_ VDD VSS sky130_fd_sc_hd__nand2_1
X_2107_ VDD VSS core.pdc.col_out\[27\] core.pdc.col_out_n\[27\] VDD VSS sky130_fd_sc_hd__clkinv_2
X_2038_ VSS VDD _0120_ _0121_ _1095_ VDD VSS sky130_fd_sc_hd__nand2_1
XANTENNA_fanout82_A VSS VDD net83 VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_77_69 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XFILLER_133_31 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XANTENNA__2068__B VSS VDD _1155_ VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__2084__A VSS VDD _1039_ VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_9_125 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_3_33 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XANTENNA_nmat_en_bit_n[0] VSS VDD core.cnb.pswitch_out\[0\] VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_95_102 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
X_3010_ VSS VDD _0897_ _0781_ _0899_ _0898_ VDD VSS sky130_fd_sc_hd__nand3_1
XFILLER_77_883 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XFILLER_91_363 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
X_2725_ VSS VDD _0616_ _0048_ _0622_ VDD VSS sky130_fd_sc_hd__nand2_1
X_2656_ VSS VDD _0559_ _0540_ _0561_ _0560_ VDD VSS sky130_fd_sc_hd__nand3_1
X_1607_ VDD VSS _1155_ _1101_ VDD VSS sky130_fd_sc_hd__buf_2
X_2587_ VDD VSS _0503_ _0502_ VDD VSS sky130_fd_sc_hd__inv_2
X_1538_ VDD VSS core.ndc.col_out\[1\] core.ndc.col_out_n\[1\] VDD VSS sky130_fd_sc_hd__inv_2
XFILLER_86_102 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
X_1469_ VDD VSS _1031_ net14 VDD VSS sky130_fd_sc_hd__inv_2
XFILLER_68_883 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XFILLER_86_179 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
X_3139_ VSS VDD clknet_2_0__leaf_clk_dig_dummy _0029_ net79 core.cnb.result_out\[7\]
+ VDD VSS sky130_fd_sc_hd__dfrtp_2
XFILLER_103_23 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XANTENNA__1801__A VSS VDD _1272_ VDD VSS sky130_fd_sc_hd__diode_2
Xgenblk1\[28\].buf_p_coln VSS VDD pmatrix_col_core_n_buffered\[28\] core.pdc.col_out_n\[28\]
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
XFILLER_103_78 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XFILLER_103_89 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_12_42 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XFILLER_128_97 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
Xgenblk1\[30\].buf_p_coln VSS VDD pmatrix_col_core_n_buffered\[30\] core.pdc.col_out_n\[30\]
+ VDD VSS sky130_fd_sc_hd__clkbuf_1
X_2510_ VSS VDD _0009_ _0446_ VDD VSS sky130_fd_sc_hd__clkbuf_1
X_2441_ VSS VDD _1382_ core.ndc.rowon_out_n\[3\] core.pdc.rowon_bottotop_n\[5\] VDD
+ VSS sky130_fd_sc_hd__nor2_2
X_2372_ VDD VSS _0383_ _0377_ core.osr.result_r\[18\] _0388_ VDD VSS sky130_fd_sc_hd__a21o_1
XANTENNA__2449__A2 VSS VDD core.pdc.rowoff_out_n\[5\] VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_83_116 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XANTENNA__1621__A VSS VDD _1131_ VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_91_193 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
X_2708_ VSS VDD _0606_ _0607_ _0519_ VDD VSS sky130_fd_sc_hd__nand2_1
X_2639_ VSS VDD _0518_ _0288_ _0537_ _0546_ VDD VSS sky130_fd_sc_hd__o21a_1
XFILLER_59_113 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_87_477 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XANTENNA__2627__A VSS VDD _1002_ VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1531__A VSS VDD _1088_ VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__2612__A2 VSS VDD _0395_ VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_128_118 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XFILLER_139_41 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XANTENNA__2081__B VSS VDD _1284_ VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_139_85 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XANTENNA__1706__A VSS VDD _1227_ VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA_nmat_rowoff_n[5] VSS VDD core.ndc.rowoff_out_n\[5\] VDD VSS sky130_fd_sc_hd__diode_2
Xgenblk1\[25\].buf_n_coln VDD VSS core.ndc.col_out_n\[25\] nmatrix_col_core_n_buffered\[25\]
+ VDD VSS sky130_fd_sc_hd__buf_6
XFILLER_48_60 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_0_12 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
X_2990_ VSS VDD _0802_ _0880_ _0869_ VDD VSS sky130_fd_sc_hd__nand2_1
X_1941_ VDD VSS _1397_ _1396_ VDD VSS sky130_fd_sc_hd__inv_2
X_1872_ VDD VSS _1353_ _1350_ _1352_ VDD VSS sky130_fd_sc_hd__or2_2
XFILLER_43_1 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
X_2424_ VDD VSS _0425_ _1360_ _1346_ VDD VSS sky130_fd_sc_hd__or2_1
X_2355_ VDD VSS _0374_ _0251_ _0373_ VDD VSS sky130_fd_sc_hd__or2_1
X_2286_ VSS VDD _0310_ _0312_ _0311_ VDD VSS sky130_fd_sc_hd__nand2_1
XFILLER_44_29 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XFILLER_109_11 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_109_44 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_109_77 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XANTENNA__3163__D VSS VDD core.osr.next_result_w\[3\] VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_85_25 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XFILLER_55_171 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XANTENNA_genblk1\[15\].buf_n_coln_A VSS VDD core.ndc.col_out_n\[15\] VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_34_40 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XFILLER_70_141 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XANTENNA__1572__A2 VSS VDD _1078_ VDD VSS sky130_fd_sc_hd__diode_2
X_2140_ VDD VSS _0184_ core.cnb.average_counter_r\[2\] VDD VSS sky130_fd_sc_hd__inv_2
XFILLER_38_149 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
X_2071_ VSS VDD _0081_ _0142_ _1213_ VDD VSS sky130_fd_sc_hd__nand2_1
XFILLER_93_277 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XFILLER_46_182 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
XFILLER_93_299 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
X_2973_ VSS VDD _0864_ _0697_ _0655_ _0764_ VDD VSS sky130_fd_sc_hd__nand3b_1
X_1924_ VSS VDD _1384_ core.pdc.rowon_out_n\[13\] _1364_ VDD VSS sky130_fd_sc_hd__nor2_2
X_1855_ VSS VDD core.pdc.row_out_n\[7\] _1337_ _1341_ VDD VSS sky130_fd_sc_hd__nand2_2
X_1786_ VSS VDD _1106_ _1292_ _1188_ VDD VSS sky130_fd_sc_hd__nand2_1
XFILLER_89_517 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XANTENNA_genblk2\[2\].buf_p_rowonn_A VSS VDD core.pdc.rowon_out_n\[2\] VDD VSS sky130_fd_sc_hd__diode_2
X_2407_ VDD VSS _0415_ core.osr.next_sample_count_w\[5\] VDD VSS sky130_fd_sc_hd__clkinv_2
X_2338_ VSS VDD _0353_ _0359_ _0358_ VDD VSS sky130_fd_sc_hd__nand2_1
XANTENNA__2177__A VSS VDD _0210_ VDD VSS sky130_fd_sc_hd__diode_2
X_2269_ VSS VDD _0296_ core.osr.next_result_w\[6\] VDD VSS sky130_fd_sc_hd__clkbuf_2
XANTENNA__2276__B1 VSS VDD _0255_ VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA_nmat_col_n[9] VSS VDD nmatrix_col_core_n_buffered\[9\] VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_71_38 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XANTENNA_genblk2\[3\].buf_n_rowonn_A VSS VDD core.ndc.rowon_out_n\[3\] VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_136_53 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_20_64 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_96_35 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
XFILLER_136_97 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XANTENNA_input25_A VSS VDD config_2_in[1] VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_45_50 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
X_1640_ VSS VDD _1039_ _1183_ _1184_ VDD VSS sky130_fd_sc_hd__nor2_1
XANTENNA__2550__A VSS VDD core.cnb.data_register_r\[0\] VDD VSS sky130_fd_sc_hd__diode_2
X_1571_ VSS VDD _1122_ _1123_ _1051_ VDD VSS sky130_fd_sc_hd__nand2_1
X_3172_ VSS VDD net58 core.osr.next_result_w\[12\] net70 core.osr.result_r\[12\] VDD
+ VSS sky130_fd_sc_hd__dfrtp_1
X_2123_ VSS VDD _1039_ _1410_ _0172_ VDD VSS sky130_fd_sc_hd__nor2_1
X_2054_ VSS VDD _1400_ _0133_ _1052_ VDD VSS sky130_fd_sc_hd__nand2_1
XFILLER_34_141 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
X_2956_ VSS VDD _0820_ _0848_ _0847_ VDD VSS sky130_fd_sc_hd__nand2_1
X_1907_ VDD VSS _1377_ _1374_ _1376_ VDD VSS sky130_fd_sc_hd__and2_1
X_2887_ VSS VDD _0757_ _0781_ VDD VSS sky130_fd_sc_hd__clkbuf_2
X_1838_ VSS VDD _1326_ _1319_ _1327_ VDD VSS sky130_fd_sc_hd__nor2_1
X_1769_ VSS VDD _1249_ _1281_ _1213_ VDD VSS sky130_fd_sc_hd__nand2_1
XFILLER_103_113 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XFILLER_103_146 VDD VSS VDD VSS sky130_fd_sc_hd__decap_8
XANTENNA__2497__B1 VSS VDD _0439_ VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__3120__RESET_B VSS VDD net85 VDD VSS sky130_fd_sc_hd__diode_2
Xoutput52 VDD VSS result_out[8] net52 VDD VSS sky130_fd_sc_hd__buf_2
Xoutput41 VDD VSS result_out[12] net41 VDD VSS sky130_fd_sc_hd__buf_2
XFILLER_48_200 VDD VSS VDD VSS sky130_fd_sc_hd__decap_6
XFILLER_48_222 VSS VDD VDD VSS sky130_fd_sc_hd__decap_4
XFILLER_91_501 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
XFILLER_56_93 VDD VSS VDD VSS sky130_fd_sc_hd__decap_3
X_2810_ VDD VSS _0705_ core.cnb.shift_register_r\[5\] VDD VSS sky130_fd_sc_hd__inv_2
X_2741_ VSS VDD net54 _0637_ core.cnb.is_holding_result_w VDD VSS sky130_fd_sc_hd__nor2_2
X_2672_ VSS VDD core.osr.next_result_w\[9\] _0575_ _0568_ VDD VSS sky130_fd_sc_hd__nand2_1
XANTENNA__1608__B VSS VDD _1045_ VDD VSS sky130_fd_sc_hd__diode_2
X_1623_ VDD VSS _1169_ _1128_ VDD VSS sky130_fd_sc_hd__inv_2
X_1554_ VSS VDD _1048_ _1108_ _1097_ VDD VSS sky130_fd_sc_hd__nand2_1
X_1485_ VSS VDD _1045_ core.cnb.data_register_r\[6\] core.cnb.data_register_r\[7\]
+ VDD VSS sky130_fd_sc_hd__nor2_4
.ends


