magic
tech sky130A
magscale 1 2
timestamp 1515178157
<< checkpaint >>
rect -1260 -1260 5600 2840
<< nwell >>
rect 200 1210 4128 1356
rect 180 370 4150 1210
rect 200 224 4128 370
<< pwell >>
rect 624 1384 1136 1526
rect 3204 1384 3716 1526
rect 624 54 1136 196
rect 3204 54 3716 196
<< varactor >>
rect 330 400 4010 1180
<< psubdiff >>
rect 650 1472 1110 1500
rect 650 1438 693 1472
rect 727 1438 761 1472
rect 795 1438 829 1472
rect 863 1438 897 1472
rect 931 1438 965 1472
rect 999 1438 1033 1472
rect 1067 1438 1110 1472
rect 650 1410 1110 1438
rect 3230 1472 3690 1500
rect 3230 1438 3273 1472
rect 3307 1438 3341 1472
rect 3375 1438 3409 1472
rect 3443 1438 3477 1472
rect 3511 1438 3545 1472
rect 3579 1438 3613 1472
rect 3647 1438 3690 1472
rect 3230 1410 3690 1438
rect 650 142 1110 170
rect 650 108 693 142
rect 727 108 761 142
rect 795 108 829 142
rect 863 108 897 142
rect 931 108 965 142
rect 999 108 1033 142
rect 1067 108 1110 142
rect 650 80 1110 108
rect 3230 142 3690 170
rect 3230 108 3273 142
rect 3307 108 3341 142
rect 3375 108 3409 142
rect 3443 108 3477 142
rect 3511 108 3545 142
rect 3579 108 3613 142
rect 3647 108 3690 142
rect 3230 80 3690 108
<< nsubdiff >>
rect 330 1282 4010 1320
rect 330 1248 521 1282
rect 555 1248 589 1282
rect 623 1248 657 1282
rect 691 1248 725 1282
rect 759 1248 793 1282
rect 827 1248 861 1282
rect 895 1248 929 1282
rect 963 1248 997 1282
rect 1031 1248 1065 1282
rect 1099 1248 1133 1282
rect 1167 1248 1201 1282
rect 1235 1248 1269 1282
rect 1303 1248 1337 1282
rect 1371 1248 1405 1282
rect 1439 1248 1473 1282
rect 1507 1248 1541 1282
rect 1575 1248 1609 1282
rect 1643 1248 1677 1282
rect 1711 1248 1745 1282
rect 1779 1248 1813 1282
rect 1847 1248 1881 1282
rect 1915 1248 1949 1282
rect 1983 1248 2017 1282
rect 2051 1248 2085 1282
rect 2119 1248 2153 1282
rect 2187 1248 2221 1282
rect 2255 1248 2289 1282
rect 2323 1248 2357 1282
rect 2391 1248 2425 1282
rect 2459 1248 2493 1282
rect 2527 1248 2561 1282
rect 2595 1248 2629 1282
rect 2663 1248 2697 1282
rect 2731 1248 2765 1282
rect 2799 1248 2833 1282
rect 2867 1248 2901 1282
rect 2935 1248 2969 1282
rect 3003 1248 3037 1282
rect 3071 1248 3105 1282
rect 3139 1248 3173 1282
rect 3207 1248 3241 1282
rect 3275 1248 3309 1282
rect 3343 1248 3377 1282
rect 3411 1248 3445 1282
rect 3479 1248 3513 1282
rect 3547 1248 3581 1282
rect 3615 1248 3649 1282
rect 3683 1248 3717 1282
rect 3751 1248 3785 1282
rect 3819 1248 4010 1282
rect 330 1180 4010 1248
rect 330 332 4010 400
rect 330 298 521 332
rect 555 298 589 332
rect 623 298 657 332
rect 691 298 725 332
rect 759 298 793 332
rect 827 298 861 332
rect 895 298 929 332
rect 963 298 997 332
rect 1031 298 1065 332
rect 1099 298 1133 332
rect 1167 298 1201 332
rect 1235 298 1269 332
rect 1303 298 1337 332
rect 1371 298 1405 332
rect 1439 298 1473 332
rect 1507 298 1541 332
rect 1575 298 1609 332
rect 1643 298 1677 332
rect 1711 298 1745 332
rect 1779 298 1813 332
rect 1847 298 1881 332
rect 1915 298 1949 332
rect 1983 298 2017 332
rect 2051 298 2085 332
rect 2119 298 2153 332
rect 2187 298 2221 332
rect 2255 298 2289 332
rect 2323 298 2357 332
rect 2391 298 2425 332
rect 2459 298 2493 332
rect 2527 298 2561 332
rect 2595 298 2629 332
rect 2663 298 2697 332
rect 2731 298 2765 332
rect 2799 298 2833 332
rect 2867 298 2901 332
rect 2935 298 2969 332
rect 3003 298 3037 332
rect 3071 298 3105 332
rect 3139 298 3173 332
rect 3207 298 3241 332
rect 3275 298 3309 332
rect 3343 298 3377 332
rect 3411 298 3445 332
rect 3479 298 3513 332
rect 3547 298 3581 332
rect 3615 298 3649 332
rect 3683 298 3717 332
rect 3751 298 3785 332
rect 3819 298 4010 332
rect 330 260 4010 298
<< psubdiffcont >>
rect 693 1438 727 1472
rect 761 1438 795 1472
rect 829 1438 863 1472
rect 897 1438 931 1472
rect 965 1438 999 1472
rect 1033 1438 1067 1472
rect 3273 1438 3307 1472
rect 3341 1438 3375 1472
rect 3409 1438 3443 1472
rect 3477 1438 3511 1472
rect 3545 1438 3579 1472
rect 3613 1438 3647 1472
rect 693 108 727 142
rect 761 108 795 142
rect 829 108 863 142
rect 897 108 931 142
rect 965 108 999 142
rect 1033 108 1067 142
rect 3273 108 3307 142
rect 3341 108 3375 142
rect 3409 108 3443 142
rect 3477 108 3511 142
rect 3545 108 3579 142
rect 3613 108 3647 142
<< nsubdiffcont >>
rect 521 1248 555 1282
rect 589 1248 623 1282
rect 657 1248 691 1282
rect 725 1248 759 1282
rect 793 1248 827 1282
rect 861 1248 895 1282
rect 929 1248 963 1282
rect 997 1248 1031 1282
rect 1065 1248 1099 1282
rect 1133 1248 1167 1282
rect 1201 1248 1235 1282
rect 1269 1248 1303 1282
rect 1337 1248 1371 1282
rect 1405 1248 1439 1282
rect 1473 1248 1507 1282
rect 1541 1248 1575 1282
rect 1609 1248 1643 1282
rect 1677 1248 1711 1282
rect 1745 1248 1779 1282
rect 1813 1248 1847 1282
rect 1881 1248 1915 1282
rect 1949 1248 1983 1282
rect 2017 1248 2051 1282
rect 2085 1248 2119 1282
rect 2153 1248 2187 1282
rect 2221 1248 2255 1282
rect 2289 1248 2323 1282
rect 2357 1248 2391 1282
rect 2425 1248 2459 1282
rect 2493 1248 2527 1282
rect 2561 1248 2595 1282
rect 2629 1248 2663 1282
rect 2697 1248 2731 1282
rect 2765 1248 2799 1282
rect 2833 1248 2867 1282
rect 2901 1248 2935 1282
rect 2969 1248 3003 1282
rect 3037 1248 3071 1282
rect 3105 1248 3139 1282
rect 3173 1248 3207 1282
rect 3241 1248 3275 1282
rect 3309 1248 3343 1282
rect 3377 1248 3411 1282
rect 3445 1248 3479 1282
rect 3513 1248 3547 1282
rect 3581 1248 3615 1282
rect 3649 1248 3683 1282
rect 3717 1248 3751 1282
rect 3785 1248 3819 1282
rect 521 298 555 332
rect 589 298 623 332
rect 657 298 691 332
rect 725 298 759 332
rect 793 298 827 332
rect 861 298 895 332
rect 929 298 963 332
rect 997 298 1031 332
rect 1065 298 1099 332
rect 1133 298 1167 332
rect 1201 298 1235 332
rect 1269 298 1303 332
rect 1337 298 1371 332
rect 1405 298 1439 332
rect 1473 298 1507 332
rect 1541 298 1575 332
rect 1609 298 1643 332
rect 1677 298 1711 332
rect 1745 298 1779 332
rect 1813 298 1847 332
rect 1881 298 1915 332
rect 1949 298 1983 332
rect 2017 298 2051 332
rect 2085 298 2119 332
rect 2153 298 2187 332
rect 2221 298 2255 332
rect 2289 298 2323 332
rect 2357 298 2391 332
rect 2425 298 2459 332
rect 2493 298 2527 332
rect 2561 298 2595 332
rect 2629 298 2663 332
rect 2697 298 2731 332
rect 2765 298 2799 332
rect 2833 298 2867 332
rect 2901 298 2935 332
rect 2969 298 3003 332
rect 3037 298 3071 332
rect 3105 298 3139 332
rect 3173 298 3207 332
rect 3241 298 3275 332
rect 3309 298 3343 332
rect 3377 298 3411 332
rect 3445 298 3479 332
rect 3513 298 3547 332
rect 3581 298 3615 332
rect 3649 298 3683 332
rect 3717 298 3751 332
rect 3785 298 3819 332
<< poly >>
rect 210 1042 330 1180
rect 210 1008 248 1042
rect 282 1008 330 1042
rect 210 952 330 1008
rect 210 918 248 952
rect 282 918 330 952
rect 210 862 330 918
rect 210 828 248 862
rect 282 828 330 862
rect 210 762 330 828
rect 210 728 248 762
rect 282 728 330 762
rect 210 672 330 728
rect 210 638 248 672
rect 282 638 330 672
rect 210 582 330 638
rect 210 548 248 582
rect 282 548 330 582
rect 210 400 330 548
rect 4010 1032 4120 1180
rect 4010 998 4058 1032
rect 4092 998 4120 1032
rect 4010 942 4120 998
rect 4010 908 4058 942
rect 4092 908 4120 942
rect 4010 852 4120 908
rect 4010 818 4058 852
rect 4092 818 4120 852
rect 4010 752 4120 818
rect 4010 718 4058 752
rect 4092 718 4120 752
rect 4010 662 4120 718
rect 4010 628 4058 662
rect 4092 628 4120 662
rect 4010 572 4120 628
rect 4010 538 4058 572
rect 4092 538 4120 572
rect 4010 400 4120 538
<< polycont >>
rect 248 1008 282 1042
rect 248 918 282 952
rect 248 828 282 862
rect 248 728 282 762
rect 248 638 282 672
rect 248 548 282 582
rect 4058 998 4092 1032
rect 4058 908 4092 942
rect 4058 818 4092 852
rect 4058 718 4092 752
rect 4058 628 4092 662
rect 4058 538 4092 572
<< locali >>
rect 650 1500 1110 1580
rect 3230 1500 3690 1580
rect 80 1472 4260 1500
rect 80 1438 693 1472
rect 727 1438 761 1472
rect 795 1438 829 1472
rect 863 1438 897 1472
rect 931 1438 965 1472
rect 999 1438 1033 1472
rect 1067 1438 3273 1472
rect 3307 1438 3341 1472
rect 3375 1438 3409 1472
rect 3443 1438 3477 1472
rect 3511 1438 3545 1472
rect 3579 1438 3613 1472
rect 3647 1438 4260 1472
rect 80 1420 4260 1438
rect 80 160 160 1420
rect 650 1410 1110 1420
rect 3230 1410 3690 1420
rect 320 1282 4020 1300
rect 320 1267 521 1282
rect 555 1267 589 1282
rect 320 1233 347 1267
rect 381 1233 419 1267
rect 453 1233 507 1267
rect 555 1248 579 1267
rect 623 1248 657 1282
rect 691 1267 725 1282
rect 759 1267 793 1282
rect 701 1248 725 1267
rect 773 1248 793 1267
rect 827 1267 861 1282
rect 541 1233 579 1248
rect 613 1233 667 1248
rect 701 1233 739 1248
rect 773 1233 827 1248
rect 895 1267 929 1282
rect 895 1248 899 1267
rect 963 1248 997 1282
rect 1031 1248 1065 1282
rect 1099 1248 1133 1282
rect 1167 1248 1201 1282
rect 1235 1248 1269 1282
rect 1303 1248 1337 1282
rect 1371 1248 1405 1282
rect 1439 1248 1473 1282
rect 1507 1248 1541 1282
rect 1575 1248 1609 1282
rect 1643 1248 1677 1282
rect 1711 1248 1745 1282
rect 1779 1248 1813 1282
rect 1847 1248 1881 1282
rect 1915 1248 1949 1282
rect 1983 1248 2017 1282
rect 2051 1248 2085 1282
rect 2119 1248 2153 1282
rect 2187 1248 2221 1282
rect 2255 1248 2289 1282
rect 2323 1248 2357 1282
rect 2391 1248 2425 1282
rect 2459 1248 2493 1282
rect 2527 1248 2561 1282
rect 2595 1248 2629 1282
rect 2663 1248 2697 1282
rect 2731 1248 2765 1282
rect 2799 1248 2833 1282
rect 2867 1248 2901 1282
rect 2935 1248 2969 1282
rect 3003 1248 3037 1282
rect 3071 1248 3105 1282
rect 3139 1248 3173 1282
rect 3207 1248 3241 1282
rect 3275 1248 3309 1282
rect 3343 1248 3377 1282
rect 3411 1267 3445 1282
rect 3441 1248 3445 1267
rect 3479 1267 3513 1282
rect 861 1233 899 1248
rect 933 1233 3407 1248
rect 3441 1233 3479 1248
rect 3547 1267 3581 1282
rect 3615 1267 3649 1282
rect 3547 1248 3567 1267
rect 3615 1248 3639 1267
rect 3683 1248 3717 1282
rect 3751 1267 3785 1282
rect 3819 1267 4020 1282
rect 3761 1248 3785 1267
rect 3513 1233 3567 1248
rect 3601 1233 3639 1248
rect 3673 1233 3727 1248
rect 3761 1233 3799 1248
rect 3833 1233 3887 1267
rect 3921 1233 3959 1267
rect 3993 1233 4020 1267
rect 320 1180 4020 1233
rect 240 1100 800 1140
rect 240 1042 350 1100
rect 840 1060 910 1180
rect 240 1008 248 1042
rect 282 1008 350 1042
rect 390 1020 910 1060
rect 240 980 350 1008
rect 240 952 800 980
rect 240 918 248 952
rect 302 940 800 952
rect 302 918 350 940
rect 240 862 350 918
rect 840 900 910 1020
rect 240 828 248 862
rect 302 828 350 862
rect 390 860 910 900
rect 240 820 350 828
rect 950 830 990 1140
rect 1030 880 1070 1180
rect 1110 830 1150 1140
rect 1190 880 1230 1180
rect 1270 830 1310 1140
rect 1350 880 1390 1180
rect 1430 830 1470 1140
rect 1510 880 1550 1180
rect 1590 830 1630 1140
rect 1670 880 1710 1180
rect 1750 830 1790 1140
rect 1830 880 1870 1180
rect 1910 830 1950 1140
rect 1990 880 2030 1180
rect 2070 830 2110 1140
rect 2150 880 2190 1180
rect 2230 830 2270 1140
rect 2310 880 2350 1180
rect 2390 830 2430 1140
rect 2470 880 2510 1180
rect 2550 830 2590 1140
rect 2630 880 2670 1180
rect 2710 830 2750 1140
rect 2790 880 2830 1180
rect 2870 830 2910 1140
rect 2950 880 2990 1180
rect 3030 830 3070 1140
rect 3110 880 3150 1180
rect 3190 830 3230 1140
rect 3270 880 3310 1180
rect 3350 830 3390 1140
rect 3430 1060 3500 1180
rect 3540 1100 4100 1140
rect 3430 1020 3950 1060
rect 3990 1032 4100 1100
rect 3430 900 3500 1020
rect 3990 998 4058 1032
rect 4092 998 4100 1032
rect 3990 980 4100 998
rect 3540 942 4100 980
rect 3540 940 4038 942
rect 3990 908 4038 940
rect 4092 908 4100 942
rect 3430 860 3940 900
rect 950 820 3390 830
rect 3990 852 4100 908
rect 3990 820 4038 852
rect 240 818 4038 820
rect 4092 818 4100 852
rect 240 762 4100 818
rect 240 728 248 762
rect 302 760 4100 762
rect 302 728 350 760
rect 240 672 350 728
rect 950 750 3390 760
rect 390 680 910 720
rect 240 638 248 672
rect 302 640 350 672
rect 302 638 800 640
rect 240 600 800 638
rect 240 582 350 600
rect 240 548 248 582
rect 282 548 350 582
rect 840 560 910 680
rect 240 480 350 548
rect 390 520 910 560
rect 240 440 800 480
rect 840 400 910 520
rect 950 440 990 750
rect 1030 400 1070 700
rect 1110 440 1150 750
rect 1190 400 1230 700
rect 1270 440 1310 750
rect 1350 400 1390 700
rect 1430 440 1470 750
rect 1510 400 1550 700
rect 1590 440 1630 750
rect 1670 400 1710 700
rect 1750 440 1790 750
rect 1830 400 1870 700
rect 1910 440 1950 750
rect 1990 400 2030 700
rect 2070 450 2110 750
rect 2150 400 2190 700
rect 2230 450 2270 750
rect 2310 400 2350 700
rect 2390 440 2430 750
rect 2470 400 2510 700
rect 2550 440 2590 750
rect 2630 400 2670 700
rect 2710 440 2750 750
rect 2790 400 2830 700
rect 2870 440 2910 750
rect 2950 400 2990 700
rect 3030 440 3070 750
rect 3110 400 3150 700
rect 3190 440 3230 750
rect 3270 400 3310 700
rect 3350 440 3390 750
rect 3990 752 4100 760
rect 3430 680 3940 720
rect 3990 718 4038 752
rect 4092 718 4100 752
rect 3430 560 3500 680
rect 3990 662 4100 718
rect 3990 640 4038 662
rect 3540 628 4038 640
rect 4092 628 4100 662
rect 3540 600 4100 628
rect 3990 572 4100 600
rect 3430 520 3950 560
rect 3990 538 4058 572
rect 4092 538 4100 572
rect 3430 400 3500 520
rect 3990 480 4100 538
rect 3540 440 4100 480
rect 320 347 4020 400
rect 320 313 347 347
rect 381 313 419 347
rect 453 313 507 347
rect 541 332 579 347
rect 613 332 667 347
rect 701 332 739 347
rect 773 332 827 347
rect 555 313 579 332
rect 320 298 521 313
rect 555 298 589 313
rect 623 298 657 332
rect 701 313 725 332
rect 773 313 793 332
rect 691 298 725 313
rect 759 298 793 313
rect 861 332 899 347
rect 933 332 3407 347
rect 3441 332 3479 347
rect 827 298 861 313
rect 895 313 899 332
rect 895 298 929 313
rect 963 298 997 332
rect 1031 298 1065 332
rect 1099 298 1133 332
rect 1167 298 1201 332
rect 1235 298 1269 332
rect 1303 298 1337 332
rect 1371 298 1405 332
rect 1439 298 1473 332
rect 1507 298 1541 332
rect 1575 298 1609 332
rect 1643 298 1677 332
rect 1711 298 1745 332
rect 1779 298 1813 332
rect 1847 298 1881 332
rect 1915 298 1949 332
rect 1983 298 2017 332
rect 2051 298 2085 332
rect 2119 298 2153 332
rect 2187 298 2221 332
rect 2255 298 2289 332
rect 2323 298 2357 332
rect 2391 298 2425 332
rect 2459 298 2493 332
rect 2527 298 2561 332
rect 2595 298 2629 332
rect 2663 298 2697 332
rect 2731 298 2765 332
rect 2799 298 2833 332
rect 2867 298 2901 332
rect 2935 298 2969 332
rect 3003 298 3037 332
rect 3071 298 3105 332
rect 3139 298 3173 332
rect 3207 298 3241 332
rect 3275 298 3309 332
rect 3343 298 3377 332
rect 3441 313 3445 332
rect 3411 298 3445 313
rect 3513 332 3567 347
rect 3601 332 3639 347
rect 3673 332 3727 347
rect 3761 332 3799 347
rect 3479 298 3513 313
rect 3547 313 3567 332
rect 3615 313 3639 332
rect 3547 298 3581 313
rect 3615 298 3649 313
rect 3683 298 3717 332
rect 3761 313 3785 332
rect 3833 313 3887 347
rect 3921 313 3959 347
rect 3993 313 4020 347
rect 3751 298 3785 313
rect 3819 298 4020 313
rect 320 280 4020 298
rect 650 160 1110 170
rect 3230 160 3690 170
rect 4180 160 4260 1420
rect 80 142 4260 160
rect 80 108 693 142
rect 727 108 761 142
rect 795 108 829 142
rect 863 108 897 142
rect 931 108 965 142
rect 999 108 1033 142
rect 1067 108 3273 142
rect 3307 108 3341 142
rect 3375 108 3409 142
rect 3443 108 3477 142
rect 3511 108 3545 142
rect 3579 108 3613 142
rect 3647 108 4260 142
rect 80 80 4260 108
rect 650 0 1110 80
rect 3230 0 3690 80
<< viali >>
rect 347 1233 381 1267
rect 419 1233 453 1267
rect 507 1248 521 1267
rect 521 1248 541 1267
rect 579 1248 589 1267
rect 589 1248 613 1267
rect 667 1248 691 1267
rect 691 1248 701 1267
rect 739 1248 759 1267
rect 759 1248 773 1267
rect 507 1233 541 1248
rect 579 1233 613 1248
rect 667 1233 701 1248
rect 739 1233 773 1248
rect 827 1233 861 1267
rect 899 1248 929 1267
rect 929 1248 933 1267
rect 3407 1248 3411 1267
rect 3411 1248 3441 1267
rect 899 1233 933 1248
rect 3407 1233 3441 1248
rect 3479 1233 3513 1267
rect 3567 1248 3581 1267
rect 3581 1248 3601 1267
rect 3639 1248 3649 1267
rect 3649 1248 3673 1267
rect 3727 1248 3751 1267
rect 3751 1248 3761 1267
rect 3799 1248 3819 1267
rect 3819 1248 3833 1267
rect 3567 1233 3601 1248
rect 3639 1233 3673 1248
rect 3727 1233 3761 1248
rect 3799 1233 3833 1248
rect 3887 1233 3921 1267
rect 3959 1233 3993 1267
rect 268 918 282 952
rect 282 918 302 952
rect 268 828 282 862
rect 282 828 302 862
rect 4038 908 4058 942
rect 4058 908 4072 942
rect 4038 818 4058 852
rect 4058 818 4072 852
rect 268 728 282 762
rect 282 728 302 762
rect 268 638 282 672
rect 282 638 302 672
rect 4038 718 4058 752
rect 4058 718 4072 752
rect 4038 628 4058 662
rect 4058 628 4072 662
rect 347 313 381 347
rect 419 313 453 347
rect 507 332 541 347
rect 579 332 613 347
rect 667 332 701 347
rect 739 332 773 347
rect 507 313 521 332
rect 521 313 541 332
rect 579 313 589 332
rect 589 313 613 332
rect 667 313 691 332
rect 691 313 701 332
rect 739 313 759 332
rect 759 313 773 332
rect 827 313 861 347
rect 899 332 933 347
rect 3407 332 3441 347
rect 899 313 929 332
rect 929 313 933 332
rect 3407 313 3411 332
rect 3411 313 3441 332
rect 3479 313 3513 347
rect 3567 332 3601 347
rect 3639 332 3673 347
rect 3727 332 3761 347
rect 3799 332 3833 347
rect 3567 313 3581 332
rect 3581 313 3601 332
rect 3639 313 3649 332
rect 3649 313 3673 332
rect 3727 313 3751 332
rect 3751 313 3761 332
rect 3799 313 3819 332
rect 3819 313 3833 332
rect 3887 313 3921 347
rect 3959 313 3993 347
<< metal1 >>
rect 0 1550 640 1580
rect 0 1370 30 1550
rect 210 1370 430 1550
rect 610 1370 640 1550
rect 0 1340 640 1370
rect 1120 1550 3220 1580
rect 1120 1370 1150 1550
rect 1330 1370 1370 1550
rect 1550 1370 2080 1550
rect 2260 1370 2790 1550
rect 2970 1370 3010 1550
rect 3190 1370 3220 1550
rect 1120 1340 3220 1370
rect 3700 1550 4340 1580
rect 3700 1370 3730 1550
rect 3910 1370 4130 1550
rect 4310 1370 4340 1550
rect 3700 1340 4340 1370
rect 0 1310 460 1340
rect 0 1280 2080 1310
rect 0 1267 960 1280
rect 0 1233 347 1267
rect 381 1233 419 1267
rect 453 1233 507 1267
rect 541 1233 579 1267
rect 613 1233 667 1267
rect 701 1233 739 1267
rect 773 1233 827 1267
rect 861 1233 899 1267
rect 933 1233 960 1267
rect 2110 1250 2230 1340
rect 3880 1310 4340 1340
rect 2260 1280 4340 1310
rect 3380 1267 4340 1280
rect 0 1230 960 1233
rect 0 1050 30 1230
rect 210 1190 960 1230
rect 990 1220 3350 1250
rect 3380 1233 3407 1267
rect 3441 1233 3479 1267
rect 3513 1233 3567 1267
rect 3601 1233 3639 1267
rect 3673 1233 3727 1267
rect 3761 1233 3799 1267
rect 3833 1233 3887 1267
rect 3921 1233 3959 1267
rect 3993 1233 4340 1267
rect 3380 1230 4340 1233
rect 210 1050 240 1190
rect 330 1180 2080 1190
rect 0 1010 240 1050
rect 0 952 330 980
rect 0 921 268 952
rect 0 869 30 921
rect 82 869 94 921
rect 146 869 158 921
rect 210 918 268 921
rect 302 918 330 952
rect 210 869 330 918
rect 360 910 390 1180
rect 0 862 330 869
rect 0 828 268 862
rect 302 850 330 862
rect 420 850 450 1150
rect 480 910 510 1180
rect 540 850 570 1150
rect 600 910 630 1180
rect 660 850 690 1150
rect 720 910 750 1180
rect 840 1160 2080 1180
rect 780 850 810 1150
rect 840 1070 960 1160
rect 2110 1130 2230 1220
rect 3380 1190 4130 1230
rect 2260 1180 4010 1190
rect 2260 1160 3500 1180
rect 990 1100 3350 1130
rect 840 1040 2080 1070
rect 840 950 960 1040
rect 2110 1010 2230 1100
rect 3380 1070 3500 1160
rect 2260 1040 3500 1070
rect 990 980 3350 1010
rect 840 920 2080 950
rect 840 880 960 920
rect 2110 890 2230 980
rect 3380 950 3500 1040
rect 2260 920 3500 950
rect 990 860 3350 890
rect 3380 880 3500 920
rect 302 830 810 850
rect 2110 830 2230 860
rect 3530 850 3560 1150
rect 3590 910 3620 1180
rect 3650 850 3680 1150
rect 3710 910 3740 1180
rect 3770 850 3800 1150
rect 3830 910 3860 1180
rect 3890 850 3920 1150
rect 3950 910 3980 1180
rect 4100 1050 4130 1190
rect 4310 1050 4340 1230
rect 4100 1010 4340 1050
rect 4010 942 4340 970
rect 4010 908 4038 942
rect 4072 921 4340 942
rect 4072 908 4130 921
rect 4010 869 4130 908
rect 4182 869 4194 921
rect 4246 869 4258 921
rect 4310 869 4340 921
rect 4010 852 4340 869
rect 4010 850 4038 852
rect 3530 830 4038 850
rect 302 828 4038 830
rect 0 818 4038 828
rect 4072 818 4340 852
rect 0 762 4340 818
rect 0 728 268 762
rect 302 752 4340 762
rect 302 728 4038 752
rect 0 718 4038 728
rect 4072 718 4340 752
rect 0 711 4340 718
rect 0 659 30 711
rect 82 659 94 711
rect 146 659 158 711
rect 210 690 4130 711
rect 210 672 330 690
rect 210 659 268 672
rect 0 638 268 659
rect 302 638 330 672
rect 0 610 330 638
rect 0 530 240 570
rect 0 350 30 530
rect 210 390 240 530
rect 360 400 390 660
rect 420 430 450 690
rect 480 400 510 660
rect 540 430 570 690
rect 600 400 630 660
rect 660 430 690 690
rect 720 400 750 660
rect 780 430 810 690
rect 840 630 2080 660
rect 840 540 960 630
rect 2110 600 2230 690
rect 2260 630 3500 660
rect 990 570 3350 600
rect 840 510 2080 540
rect 840 420 960 510
rect 2110 480 2230 570
rect 3380 540 3500 630
rect 2260 510 3500 540
rect 990 450 3350 480
rect 840 400 2080 420
rect 330 390 2080 400
rect 210 350 960 390
rect 2110 360 2230 450
rect 3380 420 3500 510
rect 3530 430 3560 690
rect 2260 400 3500 420
rect 3590 400 3620 660
rect 3650 430 3680 690
rect 3710 400 3740 660
rect 3770 430 3800 690
rect 3830 400 3860 660
rect 3890 430 3920 690
rect 4010 662 4130 690
rect 3950 400 3980 660
rect 4010 628 4038 662
rect 4072 659 4130 662
rect 4182 659 4194 711
rect 4246 659 4258 711
rect 4310 659 4340 711
rect 4072 628 4340 659
rect 4010 600 4340 628
rect 4100 530 4340 570
rect 2260 390 4010 400
rect 4100 390 4130 530
rect 0 347 960 350
rect 0 313 347 347
rect 381 313 419 347
rect 453 313 507 347
rect 541 313 579 347
rect 613 313 667 347
rect 701 313 739 347
rect 773 313 827 347
rect 861 313 899 347
rect 933 313 960 347
rect 990 330 3350 360
rect 3380 350 4130 390
rect 4310 350 4340 530
rect 3380 347 4340 350
rect 0 300 960 313
rect 0 270 2080 300
rect 0 240 460 270
rect 2110 240 2230 330
rect 3380 313 3407 347
rect 3441 313 3479 347
rect 3513 313 3567 347
rect 3601 313 3639 347
rect 3673 313 3727 347
rect 3761 313 3799 347
rect 3833 313 3887 347
rect 3921 313 3959 347
rect 3993 313 4340 347
rect 3380 300 4340 313
rect 2260 270 4340 300
rect 3880 240 4340 270
rect 0 210 640 240
rect 0 30 30 210
rect 210 30 430 210
rect 610 30 640 210
rect 0 0 640 30
rect 1120 210 3220 240
rect 1120 30 1150 210
rect 1330 30 1370 210
rect 1550 30 2080 210
rect 2260 30 2790 210
rect 2970 30 3010 210
rect 3190 30 3220 210
rect 1120 0 3220 30
rect 3700 210 4340 240
rect 3700 30 3730 210
rect 3910 30 4130 210
rect 4310 30 4340 210
rect 3700 0 4340 30
<< via1 >>
rect 30 1370 210 1550
rect 430 1370 610 1550
rect 1150 1370 1330 1550
rect 1370 1370 1550 1550
rect 2080 1370 2260 1550
rect 2790 1370 2970 1550
rect 3010 1370 3190 1550
rect 3730 1370 3910 1550
rect 4130 1370 4310 1550
rect 30 1050 210 1230
rect 30 869 82 921
rect 94 869 146 921
rect 158 869 210 921
rect 4130 1050 4310 1230
rect 4130 869 4182 921
rect 4194 869 4246 921
rect 4258 869 4310 921
rect 30 659 82 711
rect 94 659 146 711
rect 158 659 210 711
rect 30 350 210 530
rect 4130 659 4182 711
rect 4194 659 4246 711
rect 4258 659 4310 711
rect 4130 350 4310 530
rect 30 30 210 210
rect 430 30 610 210
rect 1150 30 1330 210
rect 1370 30 1550 210
rect 2080 30 2260 210
rect 2790 30 2970 210
rect 3010 30 3190 210
rect 3730 30 3910 210
rect 4130 30 4310 210
<< metal2 >>
rect 0 1550 640 1580
rect 0 1370 30 1550
rect 210 1370 430 1550
rect 610 1370 640 1550
rect 0 1340 640 1370
rect 1120 1550 3220 1580
rect 1120 1370 1150 1550
rect 1330 1370 1370 1550
rect 1550 1370 2080 1550
rect 2260 1370 2790 1550
rect 2970 1370 3010 1550
rect 3190 1370 3220 1550
rect 0 1230 390 1340
rect 1120 1300 3220 1370
rect 3700 1550 4340 1580
rect 3700 1370 3730 1550
rect 3910 1370 4130 1550
rect 4310 1370 4340 1550
rect 3700 1340 4340 1370
rect 0 1050 30 1230
rect 210 1150 390 1230
rect 420 1180 3920 1300
rect 3950 1230 4340 1340
rect 210 1120 790 1150
rect 210 1050 390 1120
rect 820 1090 880 1180
rect 420 1060 880 1090
rect 0 1030 390 1050
rect 0 1010 790 1030
rect 280 1000 790 1010
rect 0 921 240 970
rect 0 869 30 921
rect 82 869 94 921
rect 146 869 158 921
rect 210 869 240 921
rect 0 711 240 869
rect 0 659 30 711
rect 82 659 94 711
rect 146 659 158 711
rect 210 659 240 711
rect 0 610 240 659
rect 280 880 390 1000
rect 820 970 880 1060
rect 420 940 880 970
rect 280 820 790 880
rect 820 850 880 940
rect 910 820 940 1150
rect 970 850 1000 1180
rect 1030 820 1060 1150
rect 1090 850 1120 1180
rect 1150 820 1180 1150
rect 1210 850 1240 1180
rect 1270 820 1300 1150
rect 1330 850 1360 1180
rect 1390 820 1420 1150
rect 1450 850 1480 1180
rect 1510 820 1540 1150
rect 1570 850 1600 1180
rect 1630 820 1660 1150
rect 1690 850 1720 1180
rect 1750 820 1780 1150
rect 1810 850 1840 1180
rect 1870 820 1900 1150
rect 1930 850 1960 1180
rect 1990 820 2020 1150
rect 2050 850 2080 1180
rect 2110 820 2230 1150
rect 2260 850 2290 1180
rect 2320 820 2350 1150
rect 2380 850 2410 1180
rect 2440 820 2470 1150
rect 2500 850 2530 1180
rect 2560 820 2590 1150
rect 2620 850 2650 1180
rect 2680 820 2710 1150
rect 2740 850 2770 1180
rect 2800 820 2830 1150
rect 2860 850 2890 1180
rect 2920 820 2950 1150
rect 2980 850 3010 1180
rect 3040 820 3070 1150
rect 3100 850 3130 1180
rect 3160 820 3190 1150
rect 3220 850 3250 1180
rect 3280 820 3310 1150
rect 3340 850 3370 1180
rect 3400 820 3430 1150
rect 3460 1090 3520 1180
rect 3950 1150 4130 1230
rect 3550 1120 4130 1150
rect 3460 1060 3920 1090
rect 3460 970 3520 1060
rect 3950 1050 4130 1120
rect 4310 1050 4340 1230
rect 3950 1030 4340 1050
rect 3550 1010 4340 1030
rect 3550 1000 4060 1010
rect 3460 940 3920 970
rect 3460 850 3520 940
rect 3950 880 4060 1000
rect 3550 820 4060 880
rect 280 760 4060 820
rect 280 670 790 760
rect 280 580 390 670
rect 820 640 880 730
rect 420 610 880 640
rect 280 570 790 580
rect 0 550 790 570
rect 0 530 390 550
rect 0 350 30 530
rect 210 460 390 530
rect 820 520 880 610
rect 420 490 880 520
rect 210 430 790 460
rect 210 350 390 430
rect 820 400 880 490
rect 910 430 940 760
rect 970 400 1000 730
rect 1030 430 1060 760
rect 1090 400 1120 730
rect 1150 430 1180 760
rect 1210 400 1240 730
rect 1270 430 1300 760
rect 1330 400 1360 730
rect 1390 430 1420 760
rect 1450 400 1480 730
rect 1510 430 1540 760
rect 1570 400 1600 730
rect 1630 430 1660 760
rect 1690 400 1720 730
rect 1750 430 1780 760
rect 1810 400 1840 730
rect 1870 430 1900 760
rect 1930 400 1960 730
rect 1990 430 2020 760
rect 2050 400 2080 730
rect 2110 430 2230 760
rect 2260 400 2290 730
rect 2320 430 2350 760
rect 2380 400 2410 730
rect 2440 430 2470 760
rect 2500 400 2530 730
rect 2560 430 2590 760
rect 2620 400 2650 730
rect 2680 430 2710 760
rect 2740 400 2770 730
rect 2800 430 2830 760
rect 2860 400 2890 730
rect 2920 430 2950 760
rect 2980 400 3010 730
rect 3040 430 3070 760
rect 3100 400 3130 730
rect 3160 430 3190 760
rect 3220 400 3250 730
rect 3280 430 3310 760
rect 3340 400 3370 730
rect 3400 430 3430 760
rect 3460 640 3520 730
rect 3550 670 4060 760
rect 3460 610 3920 640
rect 3460 520 3520 610
rect 3950 580 4060 670
rect 4100 921 4340 970
rect 4100 869 4130 921
rect 4182 869 4194 921
rect 4246 869 4258 921
rect 4310 869 4340 921
rect 4100 711 4340 869
rect 4100 659 4130 711
rect 4182 659 4194 711
rect 4246 659 4258 711
rect 4310 659 4340 711
rect 4100 610 4340 659
rect 3550 570 4060 580
rect 3550 550 4340 570
rect 3950 530 4340 550
rect 3460 490 3920 520
rect 3460 400 3520 490
rect 3950 460 4130 530
rect 3550 430 4130 460
rect 0 240 390 350
rect 420 280 3920 400
rect 3950 350 4130 430
rect 4310 350 4340 530
rect 0 210 640 240
rect 0 30 30 210
rect 210 30 430 210
rect 610 30 640 210
rect 0 0 640 30
rect 1120 210 3220 280
rect 3950 240 4340 350
rect 1120 30 1150 210
rect 1330 30 1370 210
rect 1550 30 2080 210
rect 2260 30 2790 210
rect 2970 30 3010 210
rect 3190 30 3220 210
rect 1120 0 3220 30
rect 3700 210 4340 240
rect 3700 30 3730 210
rect 3910 30 4130 210
rect 4310 30 4340 210
rect 3700 0 4340 30
<< metal3 >>
rect 0 1547 640 1580
rect 0 1403 33 1547
rect 177 1403 453 1547
rect 597 1403 640 1547
rect 1120 1527 3220 1580
rect 1120 1463 1173 1527
rect 1237 1463 1333 1527
rect 1397 1463 2943 1527
rect 3007 1463 3103 1527
rect 3167 1463 3220 1527
rect 1120 1410 3220 1463
rect 3700 1547 4340 1580
rect 0 1330 640 1403
rect 3700 1403 3743 1547
rect 3887 1403 4163 1547
rect 4307 1403 4340 1547
rect 3700 1330 4340 1403
rect 0 1287 4340 1330
rect 0 1143 33 1287
rect 177 1143 4163 1287
rect 4307 1143 4340 1287
rect 0 1100 4340 1143
rect 0 982 170 1030
rect 0 918 53 982
rect 117 918 170 982
rect 0 902 170 918
rect 0 838 53 902
rect 117 838 170 902
rect 0 742 170 838
rect 0 678 53 742
rect 117 678 170 742
rect 0 662 170 678
rect 0 598 53 662
rect 117 598 170 662
rect 0 550 170 598
rect 250 480 4090 1100
rect 4170 982 4340 1030
rect 4170 918 4223 982
rect 4287 918 4340 982
rect 4170 902 4340 918
rect 4170 838 4223 902
rect 4287 838 4340 902
rect 4170 742 4340 838
rect 4170 678 4223 742
rect 4287 678 4340 742
rect 4170 662 4340 678
rect 4170 598 4223 662
rect 4287 598 4340 662
rect 4170 550 4340 598
rect 0 437 4340 480
rect 0 293 33 437
rect 177 293 4163 437
rect 4307 293 4340 437
rect 0 250 4340 293
rect 0 177 640 250
rect 0 33 33 177
rect 177 33 453 177
rect 597 33 640 177
rect 3700 177 4340 250
rect 0 0 640 33
rect 1120 117 3220 170
rect 1120 53 1173 117
rect 1237 53 1333 117
rect 1397 53 2943 117
rect 3007 53 3103 117
rect 3167 53 3220 117
rect 1120 0 3220 53
rect 3700 33 3743 177
rect 3887 33 4163 177
rect 4307 33 4340 177
rect 3700 0 4340 33
<< via3 >>
rect 33 1403 177 1547
rect 453 1403 597 1547
rect 1173 1463 1237 1527
rect 1333 1463 1397 1527
rect 2943 1463 3007 1527
rect 3103 1463 3167 1527
rect 3743 1403 3887 1547
rect 4163 1403 4307 1547
rect 33 1143 177 1287
rect 4163 1143 4307 1287
rect 53 918 117 982
rect 53 838 117 902
rect 53 678 117 742
rect 53 598 117 662
rect 4223 918 4287 982
rect 4223 838 4287 902
rect 4223 678 4287 742
rect 4223 598 4287 662
rect 33 293 177 437
rect 4163 293 4307 437
rect 33 33 177 177
rect 453 33 597 177
rect 1173 53 1237 117
rect 1333 53 1397 117
rect 2943 53 3007 117
rect 3103 53 3167 117
rect 3743 33 3887 177
rect 4163 33 4307 177
<< mimcap >>
rect 280 1262 4060 1300
rect 280 318 338 1262
rect 4002 318 4060 1262
rect 280 280 4060 318
<< mimcapcontact >>
rect 338 318 4002 1262
<< metal4 >>
rect 0 1547 630 1580
rect 0 1403 33 1547
rect 177 1403 453 1547
rect 597 1403 630 1547
rect 0 1370 630 1403
rect 1120 1527 3220 1580
rect 1120 1463 1173 1527
rect 1237 1463 1333 1527
rect 1397 1463 2943 1527
rect 3007 1463 3103 1527
rect 3167 1463 3220 1527
rect 0 1287 210 1370
rect 1120 1290 3220 1463
rect 3710 1547 4340 1580
rect 3710 1403 3743 1547
rect 3887 1403 4163 1547
rect 4307 1403 4340 1547
rect 3710 1370 4340 1403
rect 0 1143 33 1287
rect 177 1143 210 1287
rect 0 1110 210 1143
rect 290 1262 4050 1290
rect 290 1030 338 1262
rect 0 982 338 1030
rect 0 918 53 982
rect 117 918 338 982
rect 0 902 338 918
rect 0 838 53 902
rect 117 838 338 902
rect 0 742 338 838
rect 0 678 53 742
rect 117 678 338 742
rect 0 662 338 678
rect 0 598 53 662
rect 117 598 338 662
rect 0 550 338 598
rect 0 437 210 470
rect 0 293 33 437
rect 177 293 210 437
rect 0 210 210 293
rect 290 318 338 550
rect 4002 1030 4050 1262
rect 4130 1287 4340 1370
rect 4130 1143 4163 1287
rect 4307 1143 4340 1287
rect 4130 1110 4340 1143
rect 4002 982 4340 1030
rect 4002 918 4223 982
rect 4287 918 4340 982
rect 4002 902 4340 918
rect 4002 838 4223 902
rect 4287 838 4340 902
rect 4002 742 4340 838
rect 4002 678 4223 742
rect 4287 678 4340 742
rect 4002 662 4340 678
rect 4002 598 4223 662
rect 4287 598 4340 662
rect 4002 550 4340 598
rect 4002 318 4050 550
rect 290 290 4050 318
rect 4130 437 4340 470
rect 4130 293 4163 437
rect 4307 293 4340 437
rect 0 177 630 210
rect 0 33 33 177
rect 177 33 453 177
rect 597 33 630 177
rect 0 0 630 33
rect 1120 117 3220 290
rect 4130 210 4340 293
rect 1120 53 1173 117
rect 1237 53 1333 117
rect 1397 53 2943 117
rect 3007 53 3103 117
rect 3167 53 3220 117
rect 1120 0 3220 53
rect 3710 177 4340 210
rect 3710 33 3743 177
rect 3887 33 4163 177
rect 4307 33 4340 177
rect 3710 0 4340 33
<< labels >>
flabel metal1 s 4100 1010 4340 1580 3 FreeSans 200 90 0 0 nmoscap_bot
port 1 nsew
flabel metal1 s 4100 0 4340 570 3 FreeSans 200 90 0 0 nmoscap_bot
port 1 nsew
flabel metal1 s 0 0 240 570 7 FreeSans 200 90 0 0 nmoscap_bot
port 1 nsew
flabel metal1 s 0 1010 240 1580 7 FreeSans 200 90 0 0 nmoscap_bot
port 1 nsew
flabel metal1 s 3700 1340 4340 1580 1 FreeSans 400 0 0 0 nmoscap_bot
port 1 nsew
flabel metal1 s 3700 0 4340 240 5 FreeSans 400 0 0 0 nmoscap_bot
port 1 nsew
flabel metal1 s 0 1340 640 1580 1 FreeSans 400 0 0 0 nmoscap_bot
port 1 nsew
flabel metal1 s 0 0 640 240 5 FreeSans 400 0 0 0 nmoscap_bot
port 1 nsew
flabel metal1 s 4100 600 4340 970 3 FreeSans 400 90 0 0 nmoscap_top
port 2 nsew
flabel metal1 s 0 610 240 980 7 FreeSans 400 90 0 0 nmoscap_top
port 2 nsew
flabel metal1 s 1120 1340 3220 1580 1 FreeSans 400 0 0 0 nmoscap_top
port 2 nsew
flabel metal1 s 1120 0 3220 240 5 FreeSans 400 0 0 0 nmoscap_top
port 2 nsew
flabel locali s 3230 1500 3690 1580 1 FreeSans 400 0 0 0 pwell
port 3 nsew
flabel locali s 650 1500 1110 1580 1 FreeSans 400 0 0 0 pwell
port 3 nsew
flabel locali s 3230 0 3690 80 5 FreeSans 400 0 0 0 pwell
port 3 nsew
flabel locali s 650 0 1110 80 5 FreeSans 400 0 0 0 pwell
port 3 nsew
flabel metal3 s 4090 1100 4340 1580 3 FreeSans 400 90 0 0 mimcap_bot
port 4 nsew
flabel metal3 s 4090 0 4340 480 3 FreeSans 400 90 0 0 mimcap_bot
port 4 nsew
flabel metal3 s 0 0 250 480 7 FreeSans 400 90 0 0 mimcap_bot
port 4 nsew
flabel metal3 s 0 1100 250 1580 7 FreeSans 400 90 0 0 mimcap_bot
port 4 nsew
flabel metal3 s 3700 1340 4340 1580 1 FreeSans 400 0 0 0 mimcap_bot
port 4 nsew
flabel metal3 s 0 1340 640 1580 1 FreeSans 400 0 0 0 mimcap_bot
port 4 nsew
flabel metal3 s 3700 0 4340 240 5 FreeSans 400 0 0 0 mimcap_bot
port 4 nsew
flabel metal3 s 0 0 640 240 5 FreeSans 400 0 0 0 mimcap_bot
port 4 nsew
flabel metal3 s 0 550 170 1030 7 FreeSans 400 90 0 0 mimcap_top
port 5 nsew
flabel metal3 s 4170 550 4340 1030 3 FreeSans 400 90 0 0 mimcap_top
port 5 nsew
flabel metal3 s 1120 1410 3220 1580 1 FreeSans 400 0 0 0 mimcap_top
port 5 nsew
flabel metal3 s 1120 0 3220 170 5 FreeSans 400 0 0 0 mimcap_top
port 5 nsew
<< properties >>
string FIXED_BBOX 0 0 4340 1580
string GDS_END 99242
string GDS_FILE adc_top.gds.gz
string GDS_START 5926
<< end >>
