magic
tech sky130A
magscale 1 2
timestamp 1695298289
<< error_p >>
rect -29 181 29 187
rect -29 147 -17 181
rect -29 141 29 147
rect -127 -147 -69 -141
rect 69 -147 127 -141
rect -127 -181 -115 -147
rect 69 -181 81 -147
rect -127 -187 -69 -181
rect 69 -187 127 -181
<< nwell >>
rect -314 -319 314 319
<< pmos >>
rect -118 -100 -78 100
rect -20 -100 20 100
rect 78 -100 118 100
<< pdiff >>
rect -176 88 -118 100
rect -176 -88 -164 88
rect -130 -88 -118 88
rect -176 -100 -118 -88
rect -78 88 -20 100
rect -78 -88 -66 88
rect -32 -88 -20 88
rect -78 -100 -20 -88
rect 20 88 78 100
rect 20 -88 32 88
rect 66 -88 78 88
rect 20 -100 78 -88
rect 118 88 176 100
rect 118 -88 130 88
rect 164 -88 176 88
rect 118 -100 176 -88
<< pdiffc >>
rect -164 -88 -130 88
rect -66 -88 -32 88
rect 32 -88 66 88
rect 130 -88 164 88
<< nsubdiff >>
rect -278 249 -182 283
rect 182 249 278 283
rect -278 187 -244 249
rect 244 187 278 249
rect -278 -249 -244 -187
rect 244 -249 278 -187
rect -278 -283 -182 -249
rect 182 -283 278 -249
<< nsubdiffcont >>
rect -182 249 182 283
rect -278 -187 -244 187
rect 244 -187 278 187
rect -182 -283 182 -249
<< poly >>
rect -33 181 33 197
rect -33 147 -17 181
rect 17 147 33 181
rect -33 131 33 147
rect -118 100 -78 126
rect -20 100 20 131
rect 78 100 118 126
rect -118 -131 -78 -100
rect -20 -126 20 -100
rect 78 -131 118 -100
rect -131 -147 -65 -131
rect -131 -181 -115 -147
rect -81 -181 -65 -147
rect -131 -197 -65 -181
rect 65 -147 131 -131
rect 65 -181 81 -147
rect 115 -181 131 -147
rect 65 -197 131 -181
<< polycont >>
rect -17 147 17 181
rect -115 -181 -81 -147
rect 81 -181 115 -147
<< locali >>
rect -278 249 -182 283
rect 182 249 278 283
rect -278 187 -244 249
rect 244 187 278 249
rect -33 147 -17 181
rect 17 147 33 181
rect -164 88 -130 104
rect -164 -104 -130 -88
rect -66 88 -32 104
rect -66 -104 -32 -88
rect 32 88 66 104
rect 32 -104 66 -88
rect 130 88 164 104
rect 130 -104 164 -88
rect -131 -181 -115 -147
rect -81 -181 -65 -147
rect 65 -181 81 -147
rect 115 -181 131 -147
rect -278 -249 -244 -187
rect 244 -249 278 -187
rect -278 -283 -182 -249
rect 182 -283 278 -249
<< viali >>
rect -17 147 17 181
rect -164 -88 -130 88
rect -66 -88 -32 88
rect 32 -88 66 88
rect 130 -88 164 88
rect -115 -181 -81 -147
rect 81 -181 115 -147
<< metal1 >>
rect -29 181 29 187
rect -29 147 -17 181
rect 17 147 29 181
rect -29 141 29 147
rect -170 88 -124 100
rect -170 -88 -164 88
rect -130 -88 -124 88
rect -170 -100 -124 -88
rect -72 88 -26 100
rect -72 -88 -66 88
rect -32 -88 -26 88
rect -72 -100 -26 -88
rect 26 88 72 100
rect 26 -88 32 88
rect 66 -88 72 88
rect 26 -100 72 -88
rect 124 88 170 100
rect 124 -88 130 88
rect 164 -88 170 88
rect 124 -100 170 -88
rect -127 -147 -69 -141
rect -127 -181 -115 -147
rect -81 -181 -69 -147
rect -127 -187 -69 -181
rect 69 -147 127 -141
rect 69 -181 81 -147
rect 115 -181 127 -147
rect 69 -187 127 -181
<< properties >>
string FIXED_BBOX -261 -266 261 266
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 1 l 0.2 m 1 nf 3 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
