magic
tech sky130A
magscale 1 2
timestamp 1696841769
<< metal4 >>
rect -549 6239 549 6280
rect -549 5761 293 6239
rect 529 5761 549 6239
rect -549 5720 549 5761
rect -549 5439 549 5480
rect -549 4961 293 5439
rect 529 4961 549 5439
rect -549 4920 549 4961
rect -549 4639 549 4680
rect -549 4161 293 4639
rect 529 4161 549 4639
rect -549 4120 549 4161
rect -549 3839 549 3880
rect -549 3361 293 3839
rect 529 3361 549 3839
rect -549 3320 549 3361
rect -549 3039 549 3080
rect -549 2561 293 3039
rect 529 2561 549 3039
rect -549 2520 549 2561
rect -549 2239 549 2280
rect -549 1761 293 2239
rect 529 1761 549 2239
rect -549 1720 549 1761
rect -549 1439 549 1480
rect -549 961 293 1439
rect 529 961 549 1439
rect -549 920 549 961
rect -549 639 549 680
rect -549 161 293 639
rect 529 161 549 639
rect -549 120 549 161
rect -549 -161 549 -120
rect -549 -639 293 -161
rect 529 -639 549 -161
rect -549 -680 549 -639
rect -549 -961 549 -920
rect -549 -1439 293 -961
rect 529 -1439 549 -961
rect -549 -1480 549 -1439
rect -549 -1761 549 -1720
rect -549 -2239 293 -1761
rect 529 -2239 549 -1761
rect -549 -2280 549 -2239
rect -549 -2561 549 -2520
rect -549 -3039 293 -2561
rect 529 -3039 549 -2561
rect -549 -3080 549 -3039
rect -549 -3361 549 -3320
rect -549 -3839 293 -3361
rect 529 -3839 549 -3361
rect -549 -3880 549 -3839
rect -549 -4161 549 -4120
rect -549 -4639 293 -4161
rect 529 -4639 549 -4161
rect -549 -4680 549 -4639
rect -549 -4961 549 -4920
rect -549 -5439 293 -4961
rect 529 -5439 549 -4961
rect -549 -5480 549 -5439
rect -549 -5761 549 -5720
rect -549 -6239 293 -5761
rect 529 -6239 549 -5761
rect -549 -6280 549 -6239
<< via4 >>
rect 293 5761 529 6239
rect 293 4961 529 5439
rect 293 4161 529 4639
rect 293 3361 529 3839
rect 293 2561 529 3039
rect 293 1761 529 2239
rect 293 961 529 1439
rect 293 161 529 639
rect 293 -639 529 -161
rect 293 -1439 529 -961
rect 293 -2239 529 -1761
rect 293 -3039 529 -2561
rect 293 -3839 529 -3361
rect 293 -4639 529 -4161
rect 293 -5439 529 -4961
rect 293 -6239 529 -5761
<< mimcap2 >>
rect -469 6160 -69 6200
rect -469 5840 -429 6160
rect -109 5840 -69 6160
rect -469 5800 -69 5840
rect -469 5360 -69 5400
rect -469 5040 -429 5360
rect -109 5040 -69 5360
rect -469 5000 -69 5040
rect -469 4560 -69 4600
rect -469 4240 -429 4560
rect -109 4240 -69 4560
rect -469 4200 -69 4240
rect -469 3760 -69 3800
rect -469 3440 -429 3760
rect -109 3440 -69 3760
rect -469 3400 -69 3440
rect -469 2960 -69 3000
rect -469 2640 -429 2960
rect -109 2640 -69 2960
rect -469 2600 -69 2640
rect -469 2160 -69 2200
rect -469 1840 -429 2160
rect -109 1840 -69 2160
rect -469 1800 -69 1840
rect -469 1360 -69 1400
rect -469 1040 -429 1360
rect -109 1040 -69 1360
rect -469 1000 -69 1040
rect -469 560 -69 600
rect -469 240 -429 560
rect -109 240 -69 560
rect -469 200 -69 240
rect -469 -240 -69 -200
rect -469 -560 -429 -240
rect -109 -560 -69 -240
rect -469 -600 -69 -560
rect -469 -1040 -69 -1000
rect -469 -1360 -429 -1040
rect -109 -1360 -69 -1040
rect -469 -1400 -69 -1360
rect -469 -1840 -69 -1800
rect -469 -2160 -429 -1840
rect -109 -2160 -69 -1840
rect -469 -2200 -69 -2160
rect -469 -2640 -69 -2600
rect -469 -2960 -429 -2640
rect -109 -2960 -69 -2640
rect -469 -3000 -69 -2960
rect -469 -3440 -69 -3400
rect -469 -3760 -429 -3440
rect -109 -3760 -69 -3440
rect -469 -3800 -69 -3760
rect -469 -4240 -69 -4200
rect -469 -4560 -429 -4240
rect -109 -4560 -69 -4240
rect -469 -4600 -69 -4560
rect -469 -5040 -69 -5000
rect -469 -5360 -429 -5040
rect -109 -5360 -69 -5040
rect -469 -5400 -69 -5360
rect -469 -5840 -69 -5800
rect -469 -6160 -429 -5840
rect -109 -6160 -69 -5840
rect -469 -6200 -69 -6160
<< mimcap2contact >>
rect -429 5840 -109 6160
rect -429 5040 -109 5360
rect -429 4240 -109 4560
rect -429 3440 -109 3760
rect -429 2640 -109 2960
rect -429 1840 -109 2160
rect -429 1040 -109 1360
rect -429 240 -109 560
rect -429 -560 -109 -240
rect -429 -1360 -109 -1040
rect -429 -2160 -109 -1840
rect -429 -2960 -109 -2640
rect -429 -3760 -109 -3440
rect -429 -4560 -109 -4240
rect -429 -5360 -109 -5040
rect -429 -6160 -109 -5840
<< metal5 >>
rect -429 6184 -109 6400
rect 251 6239 571 6400
rect -453 6160 -85 6184
rect -453 5840 -429 6160
rect -109 5840 -85 6160
rect -453 5816 -85 5840
rect -429 5384 -109 5816
rect 251 5761 293 6239
rect 529 5761 571 6239
rect 251 5439 571 5761
rect -453 5360 -85 5384
rect -453 5040 -429 5360
rect -109 5040 -85 5360
rect -453 5016 -85 5040
rect -429 4584 -109 5016
rect 251 4961 293 5439
rect 529 4961 571 5439
rect 251 4639 571 4961
rect -453 4560 -85 4584
rect -453 4240 -429 4560
rect -109 4240 -85 4560
rect -453 4216 -85 4240
rect -429 3784 -109 4216
rect 251 4161 293 4639
rect 529 4161 571 4639
rect 251 3839 571 4161
rect -453 3760 -85 3784
rect -453 3440 -429 3760
rect -109 3440 -85 3760
rect -453 3416 -85 3440
rect -429 2984 -109 3416
rect 251 3361 293 3839
rect 529 3361 571 3839
rect 251 3039 571 3361
rect -453 2960 -85 2984
rect -453 2640 -429 2960
rect -109 2640 -85 2960
rect -453 2616 -85 2640
rect -429 2184 -109 2616
rect 251 2561 293 3039
rect 529 2561 571 3039
rect 251 2239 571 2561
rect -453 2160 -85 2184
rect -453 1840 -429 2160
rect -109 1840 -85 2160
rect -453 1816 -85 1840
rect -429 1384 -109 1816
rect 251 1761 293 2239
rect 529 1761 571 2239
rect 251 1439 571 1761
rect -453 1360 -85 1384
rect -453 1040 -429 1360
rect -109 1040 -85 1360
rect -453 1016 -85 1040
rect -429 584 -109 1016
rect 251 961 293 1439
rect 529 961 571 1439
rect 251 639 571 961
rect -453 560 -85 584
rect -453 240 -429 560
rect -109 240 -85 560
rect -453 216 -85 240
rect -429 -216 -109 216
rect 251 161 293 639
rect 529 161 571 639
rect 251 -161 571 161
rect -453 -240 -85 -216
rect -453 -560 -429 -240
rect -109 -560 -85 -240
rect -453 -584 -85 -560
rect -429 -1016 -109 -584
rect 251 -639 293 -161
rect 529 -639 571 -161
rect 251 -961 571 -639
rect -453 -1040 -85 -1016
rect -453 -1360 -429 -1040
rect -109 -1360 -85 -1040
rect -453 -1384 -85 -1360
rect -429 -1816 -109 -1384
rect 251 -1439 293 -961
rect 529 -1439 571 -961
rect 251 -1761 571 -1439
rect -453 -1840 -85 -1816
rect -453 -2160 -429 -1840
rect -109 -2160 -85 -1840
rect -453 -2184 -85 -2160
rect -429 -2616 -109 -2184
rect 251 -2239 293 -1761
rect 529 -2239 571 -1761
rect 251 -2561 571 -2239
rect -453 -2640 -85 -2616
rect -453 -2960 -429 -2640
rect -109 -2960 -85 -2640
rect -453 -2984 -85 -2960
rect -429 -3416 -109 -2984
rect 251 -3039 293 -2561
rect 529 -3039 571 -2561
rect 251 -3361 571 -3039
rect -453 -3440 -85 -3416
rect -453 -3760 -429 -3440
rect -109 -3760 -85 -3440
rect -453 -3784 -85 -3760
rect -429 -4216 -109 -3784
rect 251 -3839 293 -3361
rect 529 -3839 571 -3361
rect 251 -4161 571 -3839
rect -453 -4240 -85 -4216
rect -453 -4560 -429 -4240
rect -109 -4560 -85 -4240
rect -453 -4584 -85 -4560
rect -429 -5016 -109 -4584
rect 251 -4639 293 -4161
rect 529 -4639 571 -4161
rect 251 -4961 571 -4639
rect -453 -5040 -85 -5016
rect -453 -5360 -429 -5040
rect -109 -5360 -85 -5040
rect -453 -5384 -85 -5360
rect -429 -5816 -109 -5384
rect 251 -5439 293 -4961
rect 529 -5439 571 -4961
rect 251 -5761 571 -5439
rect -453 -5840 -85 -5816
rect -453 -6160 -429 -5840
rect -109 -6160 -85 -5840
rect -453 -6184 -85 -6160
rect -429 -6400 -109 -6184
rect 251 -6239 293 -5761
rect 529 -6239 571 -5761
rect 251 -6400 571 -6239
<< properties >>
string FIXED_BBOX -549 5720 11 6280
string gencell sky130_fd_pr__cap_mim_m3_2
string library sky130
string parameters w 2.0 l 2.0 val 9.52 carea 2.00 cperi 0.19 nx 1 ny 16 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
