magic
tech sky130A
magscale 1 2
timestamp 1695375165
<< pwell >>
rect -363 -310 363 310
<< nmos >>
rect -167 -100 -127 100
rect -69 -100 -29 100
rect 29 -100 69 100
rect 127 -100 167 100
<< ndiff >>
rect -225 88 -167 100
rect -225 -88 -213 88
rect -179 -88 -167 88
rect -225 -100 -167 -88
rect -127 88 -69 100
rect -127 -88 -115 88
rect -81 -88 -69 88
rect -127 -100 -69 -88
rect -29 88 29 100
rect -29 -88 -17 88
rect 17 -88 29 88
rect -29 -100 29 -88
rect 69 88 127 100
rect 69 -88 81 88
rect 115 -88 127 88
rect 69 -100 127 -88
rect 167 88 225 100
rect 167 -88 179 88
rect 213 -88 225 88
rect 167 -100 225 -88
<< ndiffc >>
rect -213 -88 -179 88
rect -115 -88 -81 88
rect -17 -88 17 88
rect 81 -88 115 88
rect 179 -88 213 88
<< psubdiff >>
rect -327 240 -231 274
rect 231 240 327 274
rect -327 178 -293 240
rect 293 178 327 240
rect -327 -240 -293 -178
rect 293 -240 327 -178
rect -327 -274 -231 -240
rect 231 -274 327 -240
<< psubdiffcont >>
rect -231 240 231 274
rect -327 -178 -293 178
rect 293 -178 327 178
rect -231 -274 231 -240
<< poly >>
rect -87 192 -21 208
rect -87 158 -71 192
rect -37 158 -21 192
rect -87 142 -21 158
rect 21 192 87 208
rect 21 158 37 192
rect 71 158 87 192
rect 21 142 87 158
rect -167 100 -127 126
rect -69 100 -29 142
rect 29 100 69 142
rect 127 100 167 126
rect -167 -122 -127 -100
rect -193 -138 -127 -122
rect -69 -126 -29 -100
rect 29 -126 69 -100
rect 127 -122 167 -100
rect -193 -172 -177 -138
rect -143 -172 -127 -138
rect -193 -188 -127 -172
rect 127 -138 193 -122
rect 127 -172 143 -138
rect 177 -172 193 -138
rect 127 -188 193 -172
<< polycont >>
rect -71 158 -37 192
rect 37 158 71 192
rect -177 -172 -143 -138
rect 143 -172 177 -138
<< locali >>
rect -327 240 -231 274
rect 231 240 327 274
rect -327 178 -293 240
rect -87 158 -71 192
rect -37 158 -21 192
rect 21 158 37 192
rect 71 158 87 192
rect 293 178 327 240
rect -213 88 -179 104
rect -213 -104 -179 -88
rect -115 88 -81 104
rect -115 -104 -81 -88
rect -17 88 17 104
rect -17 -104 17 -88
rect 81 88 115 104
rect 81 -104 115 -88
rect 179 88 213 104
rect 179 -104 213 -88
rect -193 -172 -177 -138
rect -143 -172 -127 -138
rect 127 -172 143 -138
rect 177 -172 293 -138
rect -327 -240 -293 -178
rect 127 -178 293 -172
rect 127 -180 327 -178
rect 293 -240 327 -180
rect -327 -274 -231 -240
rect 231 -274 327 -240
<< viali >>
rect -213 -88 -179 88
rect -115 -88 -81 88
rect -17 -88 17 88
rect 81 -88 115 88
rect 179 -88 213 88
<< metal1 >>
rect -219 88 -173 100
rect -219 -88 -213 88
rect -179 -88 -173 88
rect -219 -100 -173 -88
rect -121 88 -75 100
rect -121 -88 -115 88
rect -81 -88 -75 88
rect -121 -100 -75 -88
rect -23 88 23 100
rect -23 -88 -17 88
rect 17 -88 23 88
rect -23 -100 23 -88
rect 75 88 121 100
rect 75 -88 81 88
rect 115 -88 121 88
rect 75 -100 121 -88
rect 173 88 219 100
rect 173 -88 179 88
rect 213 -88 219 88
rect 173 -100 219 -88
<< properties >>
string FIXED_BBOX -310 -257 310 257
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 1 l 0.2 m 1 nf 4 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
