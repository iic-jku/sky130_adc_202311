magic
tech sky130A
magscale 1 2
timestamp 1698999411
<< nwell >>
rect -10 48 408 452
<< pwell >>
rect 0 -244 398 -90
rect -68 -332 408 -244
<< nmos >>
rect 88 -216 118 -116
rect 184 -216 214 -116
rect 280 -216 310 -116
<< pmos >>
rect 88 110 118 310
rect 184 110 214 310
rect 280 110 310 310
<< ndiff >>
rect 26 -152 88 -116
rect 26 -186 38 -152
rect 72 -186 88 -152
rect 26 -216 88 -186
rect 118 -149 184 -116
rect 118 -183 134 -149
rect 168 -183 184 -149
rect 118 -216 184 -183
rect 214 -149 280 -116
rect 214 -183 230 -149
rect 264 -183 280 -149
rect 214 -216 280 -183
rect 310 -149 372 -116
rect 310 -183 326 -149
rect 360 -183 372 -149
rect 310 -216 372 -183
<< pdiff >>
rect 26 295 88 310
rect 26 261 38 295
rect 72 261 88 295
rect 26 227 88 261
rect 26 193 38 227
rect 72 193 88 227
rect 26 159 88 193
rect 26 125 38 159
rect 72 125 88 159
rect 26 110 88 125
rect 118 295 184 310
rect 118 261 134 295
rect 168 261 184 295
rect 118 227 184 261
rect 118 193 134 227
rect 168 193 184 227
rect 118 159 184 193
rect 118 125 134 159
rect 168 125 184 159
rect 118 110 184 125
rect 214 295 280 310
rect 214 261 230 295
rect 264 261 280 295
rect 214 227 280 261
rect 214 193 230 227
rect 264 193 280 227
rect 214 159 280 193
rect 214 125 230 159
rect 264 125 280 159
rect 214 110 280 125
rect 310 295 372 310
rect 310 261 326 295
rect 360 261 372 295
rect 310 227 372 261
rect 310 193 326 227
rect 360 193 372 227
rect 310 159 372 193
rect 310 125 326 159
rect 360 125 372 159
rect 310 110 372 125
<< ndiffc >>
rect 38 -186 72 -152
rect 134 -183 168 -149
rect 230 -183 264 -149
rect 326 -183 360 -149
<< pdiffc >>
rect 38 261 72 295
rect 38 193 72 227
rect 38 125 72 159
rect 134 261 168 295
rect 134 193 168 227
rect 134 125 168 159
rect 230 261 264 295
rect 230 193 264 227
rect 230 125 264 159
rect 326 261 360 295
rect 326 193 360 227
rect 326 125 360 159
<< psubdiff >>
rect -42 -304 -16 -270
rect 18 -304 52 -270
rect 86 -304 120 -270
rect 154 -304 188 -270
rect 222 -304 256 -270
rect 290 -304 324 -270
rect 358 -304 382 -270
rect -42 -306 382 -304
<< nsubdiff >>
rect 26 414 372 416
rect 26 380 52 414
rect 86 380 128 414
rect 162 380 204 414
rect 238 380 280 414
rect 314 380 372 414
rect 26 378 372 380
<< psubdiffcont >>
rect -16 -304 18 -270
rect 52 -304 86 -270
rect 120 -304 154 -270
rect 188 -304 222 -270
rect 256 -304 290 -270
rect 324 -304 358 -270
<< nsubdiffcont >>
rect 52 380 86 414
rect 128 380 162 414
rect 204 380 238 414
rect 280 380 314 414
<< poly >>
rect 88 310 118 336
rect 184 310 214 336
rect 280 310 310 336
rect 88 28 118 110
rect 184 84 214 110
rect 280 84 310 110
rect 184 48 310 84
rect 68 11 128 28
rect 68 -23 78 11
rect 112 -23 128 11
rect 68 -40 128 -23
rect 216 11 274 48
rect 216 -23 226 11
rect 260 -23 274 11
rect 88 -116 118 -40
rect 216 -70 274 -23
rect 184 -100 310 -70
rect 184 -116 214 -100
rect 280 -116 310 -100
rect 88 -242 118 -216
rect 184 -242 214 -216
rect 280 -242 310 -216
<< polycont >>
rect 78 -23 112 11
rect 226 -23 260 11
<< locali >>
rect -42 414 408 416
rect -42 380 52 414
rect 86 380 128 414
rect 162 380 204 414
rect 238 380 280 414
rect 314 380 408 414
rect -42 378 408 380
rect 38 295 72 314
rect 38 227 72 261
rect 38 171 72 193
rect 38 106 72 125
rect 134 295 168 378
rect 134 227 168 261
rect 134 159 168 193
rect 134 106 168 125
rect 230 295 264 314
rect 230 227 264 261
rect 230 159 264 162
rect 230 106 264 125
rect 326 295 360 378
rect 326 227 360 261
rect 326 159 360 193
rect 326 106 360 125
rect 68 11 128 28
rect 68 -23 78 11
rect 112 -23 128 11
rect 68 -40 128 -23
rect 216 11 262 28
rect 216 -23 226 11
rect 260 -23 262 11
rect 216 -40 262 -23
rect 38 -143 72 -112
rect 38 -220 72 -186
rect 134 -149 168 -112
rect 134 -270 168 -183
rect 230 -149 264 -112
rect 230 -220 264 -185
rect 326 -149 360 -112
rect 326 -270 360 -183
rect -42 -304 -16 -270
rect 18 -304 52 -270
rect 86 -304 120 -270
rect 154 -304 188 -270
rect 222 -304 256 -270
rect 290 -304 324 -270
rect 358 -304 382 -270
rect -42 -306 382 -304
<< viali >>
rect 38 159 72 171
rect 38 137 72 159
rect 230 193 264 196
rect 230 162 264 193
rect 78 -23 112 11
rect 226 -23 260 11
rect 38 -152 72 -143
rect 38 -177 72 -152
rect 230 -183 264 -151
rect 230 -185 264 -183
<< metal1 >>
rect 32 171 78 198
rect 32 137 38 171
rect 72 137 78 171
rect 224 196 360 218
rect 224 162 230 196
rect 264 162 360 196
rect 224 142 360 162
rect 32 116 78 137
rect 38 84 72 116
rect 38 56 272 84
rect 68 11 128 28
rect 68 8 78 11
rect -16 -20 78 8
rect 68 -23 78 -20
rect 112 -23 128 11
rect 68 -40 128 -23
rect 214 11 272 56
rect 214 -23 226 11
rect 260 -23 272 11
rect 214 -68 272 -23
rect 38 -96 272 -68
rect 326 8 360 142
rect 326 -20 408 8
rect 38 -124 72 -96
rect 32 -143 78 -124
rect 326 -128 360 -20
rect 32 -177 38 -143
rect 72 -177 78 -143
rect 32 -198 78 -177
rect 224 -151 360 -128
rect 224 -185 230 -151
rect 264 -185 360 -151
rect 224 -204 360 -185
<< labels >>
flabel metal1 s 356 -20 408 8 0 FreeSans 200 0 0 0 out
port 1 nsew
flabel metal1 s -16 -20 34 8 0 FreeSans 200 0 0 0 in
port 2 nsew
flabel locali s -42 -306 382 -270 0 FreeSans 200 0 0 0 VSS
port 3 nsew
flabel locali s -42 378 408 416 0 FreeSans 200 0 0 0 VDD
port 4 nsew
<< end >>
