magic
tech sky130A
magscale 1 2
timestamp 1696930192
<< pwell >>
rect -455 -260 455 260
<< nmos >>
rect -255 -50 -225 50
rect -159 -50 -129 50
rect -63 -50 -33 50
rect 33 -50 63 50
rect 129 -50 159 50
rect 225 -50 255 50
<< ndiff >>
rect -317 38 -255 50
rect -317 -38 -305 38
rect -271 -38 -255 38
rect -317 -50 -255 -38
rect -225 38 -159 50
rect -225 -38 -209 38
rect -175 -38 -159 38
rect -225 -50 -159 -38
rect -129 38 -63 50
rect -129 -38 -113 38
rect -79 -38 -63 38
rect -129 -50 -63 -38
rect -33 38 33 50
rect -33 -38 -17 38
rect 17 -38 33 38
rect -33 -50 33 -38
rect 63 38 129 50
rect 63 -38 79 38
rect 113 -38 129 38
rect 63 -50 129 -38
rect 159 38 225 50
rect 159 -38 175 38
rect 209 -38 225 38
rect 159 -50 225 -38
rect 255 38 317 50
rect 255 -38 271 38
rect 305 -38 317 38
rect 255 -50 317 -38
<< ndiffc >>
rect -305 -38 -271 38
rect -209 -38 -175 38
rect -113 -38 -79 38
rect -17 -38 17 38
rect 79 -38 113 38
rect 175 -38 209 38
rect 271 -38 305 38
<< psubdiff >>
rect -419 190 -323 224
rect 323 190 419 224
rect -419 128 -385 190
rect 385 128 419 190
rect -419 -190 -385 -128
rect 385 -190 419 -128
rect -419 -224 -323 -190
rect 323 -224 419 -190
<< psubdiffcont >>
rect -323 190 323 224
rect -419 -128 -385 128
rect 385 -128 419 128
rect -323 -224 323 -190
<< poly >>
rect -255 50 -225 76
rect -159 50 -129 76
rect -63 50 -33 76
rect 33 50 63 76
rect 129 50 159 76
rect 225 50 255 76
rect -255 -72 -225 -50
rect -159 -72 -129 -50
rect -63 -72 -33 -50
rect 33 -72 63 -50
rect 129 -72 159 -50
rect 225 -72 255 -50
rect -291 -88 -225 -72
rect -291 -122 -275 -88
rect -241 -122 -225 -88
rect -291 -138 -225 -122
rect -177 -88 -111 -72
rect -177 -122 -161 -88
rect -127 -122 -111 -88
rect -177 -138 -111 -122
rect -63 -88 63 -72
rect -63 -122 -47 -88
rect 47 -122 63 -88
rect -63 -138 63 -122
rect 111 -88 177 -72
rect 111 -122 127 -88
rect 161 -122 177 -88
rect 111 -138 177 -122
rect 225 -88 291 -72
rect 225 -122 241 -88
rect 275 -122 291 -88
rect 225 -138 291 -122
<< polycont >>
rect -275 -122 -241 -88
rect -161 -122 -127 -88
rect -47 -122 47 -88
rect 127 -122 161 -88
rect 241 -122 275 -88
<< locali >>
rect -419 190 -323 224
rect 323 190 419 224
rect -419 128 -385 190
rect 385 128 419 190
rect -305 38 -271 54
rect -305 -54 -271 -38
rect -209 38 -175 54
rect -209 -54 -175 -38
rect -113 38 -79 54
rect -113 -54 -79 -38
rect -17 38 17 54
rect -17 -54 17 -38
rect 79 38 113 54
rect 79 -54 113 -38
rect 175 38 209 54
rect 175 -54 209 -38
rect 271 38 305 54
rect 271 -54 305 -38
rect -291 -122 -275 -88
rect -241 -122 -225 -88
rect -177 -122 -161 -88
rect -127 -122 -111 -88
rect -63 -122 -47 -88
rect 47 -122 63 -88
rect 111 -122 127 -88
rect 161 -122 177 -88
rect 225 -122 241 -88
rect 275 -122 291 -88
rect -419 -190 -385 -128
rect 385 -190 419 -128
rect -419 -224 -323 -190
rect 323 -224 419 -190
<< viali >>
rect -305 -38 -271 38
rect -209 -38 -175 38
rect -113 -38 -79 38
rect -17 -38 17 38
rect 79 -38 113 38
rect 175 -38 209 38
rect 271 -38 305 38
rect -161 -122 -127 -88
rect -47 -122 47 -88
rect 127 -122 161 -88
<< metal1 >>
rect -311 38 -265 50
rect -311 -38 -305 38
rect -271 -38 -265 38
rect -311 -50 -265 -38
rect -215 38 -169 50
rect -215 -38 -209 38
rect -175 -38 -169 38
rect -215 -50 -169 -38
rect -119 38 -73 50
rect -119 -38 -113 38
rect -79 -38 -73 38
rect -119 -50 -73 -38
rect -23 38 23 50
rect -23 -38 -17 38
rect 17 -38 23 38
rect -23 -50 23 -38
rect 73 38 119 50
rect 73 -38 79 38
rect 113 -38 119 38
rect 73 -50 119 -38
rect 169 38 215 50
rect 169 -38 175 38
rect 209 -38 215 38
rect 169 -50 215 -38
rect 265 38 311 50
rect 265 -38 271 38
rect 305 -38 311 38
rect 265 -50 311 -38
rect -177 -88 -111 -82
rect -177 -122 -161 -88
rect -127 -122 -111 -88
rect -177 -138 -111 -122
rect -59 -88 59 -82
rect -59 -122 -47 -88
rect 47 -122 59 -88
rect -59 -128 59 -122
rect 111 -88 177 -82
rect 111 -122 127 -88
rect 161 -122 177 -88
rect 111 -138 177 -122
<< properties >>
string FIXED_BBOX -402 -207 402 207
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 0.5 l 0.150 m 1 nf 6 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
