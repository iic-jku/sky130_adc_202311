magic
tech sky130A
magscale 1 2
timestamp 1515178157
<< checkpaint >>
rect -1298 -1308 2218 1852
<< nwell >>
rect -38 261 958 582
<< pwell >>
rect 134 157 884 203
rect 37 21 884 157
rect 37 17 59 21
rect 25 -17 59 17
<< scnmos >>
rect 115 47 145 131
rect 210 47 240 177
rect 398 47 428 131
rect 493 47 523 177
rect 681 47 711 131
rect 776 47 806 177
<< scpmoshvt >>
rect 115 413 145 497
rect 210 297 240 497
rect 398 413 428 497
rect 493 297 523 497
rect 681 413 711 497
rect 776 297 806 497
<< ndiff >>
rect 160 131 210 177
rect 63 106 115 131
rect 63 72 71 106
rect 105 72 115 106
rect 63 47 115 72
rect 145 93 210 131
rect 145 59 160 93
rect 194 59 210 93
rect 145 47 210 59
rect 240 105 292 177
rect 443 131 493 177
rect 240 71 250 105
rect 284 71 292 105
rect 240 47 292 71
rect 346 105 398 131
rect 346 71 354 105
rect 388 71 398 105
rect 346 47 398 71
rect 428 93 493 131
rect 428 59 443 93
rect 477 59 493 93
rect 428 47 493 59
rect 523 105 575 177
rect 726 131 776 177
rect 523 71 533 105
rect 567 71 575 105
rect 523 47 575 71
rect 629 105 681 131
rect 629 71 637 105
rect 671 71 681 105
rect 629 47 681 71
rect 711 93 776 131
rect 711 59 726 93
rect 760 59 776 93
rect 711 47 776 59
rect 806 105 858 177
rect 806 71 816 105
rect 850 71 858 105
rect 806 47 858 71
<< pdiff >>
rect 63 472 115 497
rect 63 438 71 472
rect 105 438 115 472
rect 63 413 115 438
rect 145 489 210 497
rect 145 455 161 489
rect 195 455 210 489
rect 145 413 210 455
rect 160 297 210 413
rect 240 477 292 497
rect 240 443 250 477
rect 284 443 292 477
rect 240 409 292 443
rect 346 472 398 497
rect 346 438 354 472
rect 388 438 398 472
rect 346 413 398 438
rect 428 489 493 497
rect 428 455 444 489
rect 478 455 493 489
rect 428 413 493 455
rect 240 375 250 409
rect 284 375 292 409
rect 240 297 292 375
rect 443 297 493 413
rect 523 477 575 497
rect 523 443 533 477
rect 567 443 575 477
rect 523 409 575 443
rect 629 472 681 497
rect 629 438 637 472
rect 671 438 681 472
rect 629 413 681 438
rect 711 489 776 497
rect 711 455 727 489
rect 761 455 776 489
rect 711 413 776 455
rect 523 375 533 409
rect 567 375 575 409
rect 523 297 575 375
rect 726 297 776 413
rect 806 477 858 497
rect 806 443 816 477
rect 850 443 858 477
rect 806 409 858 443
rect 806 375 816 409
rect 850 375 858 409
rect 806 297 858 375
<< ndiffc >>
rect 71 72 105 106
rect 160 59 194 93
rect 250 71 284 105
rect 354 71 388 105
rect 443 59 477 93
rect 533 71 567 105
rect 637 71 671 105
rect 726 59 760 93
rect 816 71 850 105
<< pdiffc >>
rect 71 438 105 472
rect 161 455 195 489
rect 250 443 284 477
rect 354 438 388 472
rect 444 455 478 489
rect 250 375 284 409
rect 533 443 567 477
rect 637 438 671 472
rect 727 455 761 489
rect 533 375 567 409
rect 816 443 850 477
rect 816 375 850 409
<< poly >>
rect 115 497 145 523
rect 210 497 240 523
rect 398 497 428 523
rect 493 497 523 523
rect 681 497 711 523
rect 776 497 806 523
rect 115 265 145 413
rect 210 265 240 297
rect 398 265 428 413
rect 493 265 523 297
rect 681 265 711 413
rect 776 265 806 297
rect 58 249 145 265
rect 58 215 68 249
rect 102 215 145 249
rect 58 199 145 215
rect 187 249 241 265
rect 187 215 197 249
rect 231 215 241 249
rect 187 199 241 215
rect 341 249 428 265
rect 341 215 351 249
rect 385 215 428 249
rect 341 199 428 215
rect 470 249 524 265
rect 470 215 480 249
rect 514 215 524 249
rect 470 199 524 215
rect 624 249 711 265
rect 624 215 634 249
rect 668 215 711 249
rect 624 199 711 215
rect 753 249 807 265
rect 753 215 763 249
rect 797 215 807 249
rect 753 199 807 215
rect 115 131 145 199
rect 210 177 240 199
rect 398 131 428 199
rect 493 177 523 199
rect 681 131 711 199
rect 776 177 806 199
rect 115 21 145 47
rect 210 21 240 47
rect 398 21 428 47
rect 493 21 523 47
rect 681 21 711 47
rect 776 21 806 47
<< polycont >>
rect 68 215 102 249
rect 197 215 231 249
rect 351 215 385 249
rect 480 215 514 249
rect 634 215 668 249
rect 763 215 797 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 920 561
rect 17 472 105 493
rect 17 438 71 472
rect 139 489 216 527
rect 139 455 161 489
rect 195 455 216 489
rect 139 442 216 455
rect 250 477 304 493
rect 284 443 304 477
rect 17 408 105 438
rect 250 409 304 443
rect 17 374 216 408
rect 17 249 115 340
rect 17 215 68 249
rect 102 215 115 249
rect 17 199 115 215
rect 149 265 216 374
rect 284 375 304 409
rect 250 335 304 375
rect 338 472 388 493
rect 338 438 354 472
rect 422 489 499 527
rect 422 455 444 489
rect 478 455 499 489
rect 422 442 499 455
rect 533 477 583 493
rect 567 443 583 477
rect 338 408 388 438
rect 533 409 583 443
rect 338 369 499 408
rect 250 299 395 335
rect 149 249 231 265
rect 149 215 197 249
rect 149 199 231 215
rect 265 249 395 299
rect 265 215 351 249
rect 385 215 395 249
rect 265 199 395 215
rect 429 265 499 369
rect 567 375 583 409
rect 533 335 583 375
rect 617 472 671 493
rect 617 438 637 472
rect 705 489 782 527
rect 705 455 727 489
rect 761 455 782 489
rect 705 442 782 455
rect 816 477 903 493
rect 850 443 903 477
rect 617 408 671 438
rect 816 409 903 443
rect 617 369 782 408
rect 533 299 678 335
rect 429 249 514 265
rect 429 215 480 249
rect 429 199 514 215
rect 548 249 678 299
rect 548 215 634 249
rect 668 215 678 249
rect 548 199 678 215
rect 712 265 782 369
rect 850 375 903 409
rect 816 299 903 375
rect 712 249 797 265
rect 712 215 763 249
rect 712 199 797 215
rect 149 165 216 199
rect 265 165 304 199
rect 429 165 499 199
rect 548 165 583 199
rect 712 165 782 199
rect 831 165 903 299
rect 17 131 216 165
rect 17 106 105 131
rect 17 72 71 106
rect 250 105 304 165
rect 17 51 105 72
rect 139 93 216 97
rect 139 59 160 93
rect 194 59 216 93
rect 139 17 216 59
rect 284 71 304 105
rect 250 51 304 71
rect 338 131 499 165
rect 338 105 388 131
rect 338 71 354 105
rect 533 105 583 165
rect 338 51 388 71
rect 422 93 499 97
rect 422 59 443 93
rect 477 59 499 93
rect 422 17 499 59
rect 567 71 583 105
rect 533 51 583 71
rect 617 131 782 165
rect 617 105 671 131
rect 617 71 637 105
rect 816 105 903 165
rect 617 51 671 71
rect 705 93 782 97
rect 705 59 726 93
rect 760 59 782 93
rect 705 17 782 59
rect 850 71 903 105
rect 816 51 903 71
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 920 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
<< metal1 >>
rect 0 561 920 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 920 561
rect 0 496 920 527
rect 0 17 920 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 920 17
rect 0 -48 920 -17
<< labels >>
flabel metal1 s 25 527 59 561 0 FreeSans 200 0 0 0 VPWR
port 1 nsew
flabel metal1 s 25 -17 59 17 0 FreeSans 200 0 0 0 VGND
port 2 nsew
flabel locali s 25 221 59 255 0 FreeSans 200 0 0 0 A
port 4 nsew
flabel locali s 861 289 895 323 0 FreeSans 200 0 0 0 X
port 3 nsew
flabel locali s 25 289 59 323 0 FreeSans 200 0 0 0 A
port 4 nsew
flabel locali s 861 357 895 391 0 FreeSans 200 0 0 0 X
port 3 nsew
flabel locali s 861 425 895 459 0 FreeSans 200 0 0 0 X
port 3 nsew
flabel locali s 861 221 895 255 0 FreeSans 200 0 0 0 X
port 3 nsew
flabel locali s 861 153 895 187 0 FreeSans 200 0 0 0 X
port 3 nsew
flabel locali s 861 85 895 119 0 FreeSans 200 0 0 0 X
port 3 nsew
rlabel comment s 0 0 0 0 4 dlymetal6s6s_1
flabel nwell s 25 527 59 561 0 FreeSans 200 0 0 0 VPB
port 6 nsew
flabel pwell s 25 -17 59 17 0 FreeSans 200 0 0 0 VNB
port 7 nsew
<< properties >>
string FIXED_BBOX 0 0 920 544
string GDS_END 205990
string GDS_FILE adc_top.gds.gz
string GDS_START 198454
string path 0.000 2.720 4.600 2.720 
<< end >>
