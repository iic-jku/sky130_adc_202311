magic
tech sky130A
magscale 1 2
timestamp 1695305941
<< error_p >>
rect -29 172 29 178
rect -29 138 -17 172
rect -29 132 29 138
rect -127 -138 -69 -132
rect 69 -138 127 -132
rect -127 -172 -115 -138
rect 69 -172 81 -138
rect -127 -178 -69 -172
rect 69 -178 127 -172
<< pwell >>
rect -314 -310 314 310
<< nmos >>
rect -118 -100 -78 100
rect -20 -100 20 100
rect 78 -100 118 100
<< ndiff >>
rect -176 88 -118 100
rect -176 -88 -164 88
rect -130 -88 -118 88
rect -176 -100 -118 -88
rect -78 88 -20 100
rect -78 -88 -66 88
rect -32 -88 -20 88
rect -78 -100 -20 -88
rect 20 88 78 100
rect 20 -88 32 88
rect 66 -88 78 88
rect 20 -100 78 -88
rect 118 88 176 100
rect 118 -88 130 88
rect 164 -88 176 88
rect 118 -100 176 -88
<< ndiffc >>
rect -164 -88 -130 88
rect -66 -88 -32 88
rect 32 -88 66 88
rect 130 -88 164 88
<< psubdiff >>
rect -278 240 278 274
rect -278 178 -244 240
rect 244 178 278 240
rect -278 -240 -244 -178
rect 244 -240 278 -178
rect -278 -274 278 -240
<< psubdiffcont >>
rect -278 -178 -244 178
rect 244 -178 278 178
<< poly >>
rect -33 172 33 188
rect -33 138 -17 172
rect 17 138 33 172
rect -118 100 -78 126
rect -33 122 33 138
rect -20 100 20 122
rect 78 100 118 126
rect -118 -122 -78 -100
rect -131 -138 -65 -122
rect -20 -126 20 -100
rect 78 -122 118 -100
rect -131 -172 -115 -138
rect -81 -172 -65 -138
rect -131 -188 -65 -172
rect 65 -138 131 -122
rect 65 -172 81 -138
rect 115 -172 131 -138
rect 65 -188 131 -172
<< polycont >>
rect -17 138 17 172
rect -115 -172 -81 -138
rect 81 -172 115 -138
<< locali >>
rect -278 240 278 274
rect -278 178 -244 240
rect 244 178 278 240
rect -33 138 -17 172
rect 17 138 33 172
rect -164 88 -130 104
rect -164 -104 -130 -88
rect -66 88 -32 104
rect -66 -104 -32 -88
rect 32 88 66 104
rect 32 -104 66 -88
rect 130 88 164 104
rect 130 -104 164 -88
rect -131 -172 -115 -138
rect -81 -172 -65 -138
rect 65 -172 81 -138
rect 115 -172 131 -138
rect -278 -240 -244 -178
rect 244 -240 278 -178
rect -278 -274 278 -240
<< viali >>
rect -17 138 17 172
rect -164 -88 -130 88
rect -66 -88 -32 88
rect 32 -88 66 88
rect 130 -88 164 88
rect -115 -172 -81 -138
rect 81 -172 115 -138
<< metal1 >>
rect -29 172 29 178
rect -29 138 -17 172
rect 17 138 29 172
rect -29 132 29 138
rect -170 88 -124 100
rect -170 -88 -164 88
rect -130 -88 -124 88
rect -170 -100 -124 -88
rect -72 88 -26 100
rect -72 -88 -66 88
rect -32 -88 -26 88
rect -72 -100 -26 -88
rect 26 88 72 100
rect 26 -88 32 88
rect 66 -88 72 88
rect 26 -100 72 -88
rect 124 88 170 100
rect 124 -88 130 88
rect 164 -88 170 88
rect 124 -100 170 -88
rect -127 -138 -69 -132
rect -127 -172 -115 -138
rect -81 -172 -69 -138
rect -127 -178 -69 -172
rect 69 -138 127 -132
rect 69 -172 81 -138
rect 115 -172 127 -138
rect 69 -178 127 -172
<< properties >>
string FIXED_BBOX -261 -257 261 257
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 1 l 0.2 m 1 nf 3 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
