magic
tech sky130A
magscale 1 2
timestamp 1697705955
<< error_p >>
rect -365 -413 -307 -407
rect 307 -413 365 -407
rect -365 -447 -353 -413
rect 307 -447 319 -413
rect -365 -453 -307 -447
rect 307 -453 365 -447
<< pwell >>
rect -647 -585 647 585
<< nmos >>
rect -447 -375 -417 375
rect -351 -375 -321 375
rect -255 -375 -225 375
rect -159 -375 -129 375
rect -63 -375 -33 375
rect 33 -375 63 375
rect 129 -375 159 375
rect 225 -375 255 375
rect 321 -375 351 375
rect 417 -375 447 375
<< ndiff >>
rect -509 363 -447 375
rect -509 -363 -497 363
rect -463 -363 -447 363
rect -509 -375 -447 -363
rect -417 363 -351 375
rect -417 -363 -401 363
rect -367 -363 -351 363
rect -417 -375 -351 -363
rect -321 363 -255 375
rect -321 -363 -305 363
rect -271 -363 -255 363
rect -321 -375 -255 -363
rect -225 363 -159 375
rect -225 -363 -209 363
rect -175 -363 -159 363
rect -225 -375 -159 -363
rect -129 363 -63 375
rect -129 -363 -113 363
rect -79 -363 -63 363
rect -129 -375 -63 -363
rect -33 363 33 375
rect -33 -363 -17 363
rect 17 -363 33 363
rect -33 -375 33 -363
rect 63 363 129 375
rect 63 -363 79 363
rect 113 -363 129 363
rect 63 -375 129 -363
rect 159 363 225 375
rect 159 -363 175 363
rect 209 -363 225 363
rect 159 -375 225 -363
rect 255 363 321 375
rect 255 -363 271 363
rect 305 -363 321 363
rect 255 -375 321 -363
rect 351 363 417 375
rect 351 -363 367 363
rect 401 -363 417 363
rect 351 -375 417 -363
rect 447 363 509 375
rect 447 -363 463 363
rect 497 -363 509 363
rect 447 -375 509 -363
<< ndiffc >>
rect -497 -363 -463 363
rect -401 -363 -367 363
rect -305 -363 -271 363
rect -209 -363 -175 363
rect -113 -363 -79 363
rect -17 -363 17 363
rect 79 -363 113 363
rect 175 -363 209 363
rect 271 -363 305 363
rect 367 -363 401 363
rect 463 -363 497 363
<< psubdiff >>
rect -611 515 -515 549
rect 515 515 611 549
rect -611 453 -577 515
rect 577 453 611 515
rect -611 -515 -577 -453
rect 577 -515 611 -453
rect -611 -549 -515 -515
rect 515 -549 611 -515
<< psubdiffcont >>
rect -515 515 515 549
rect -611 -453 -577 453
rect 577 -453 611 453
rect -515 -549 515 -515
<< poly >>
rect -447 375 -417 401
rect -351 375 -321 401
rect -255 375 -225 401
rect -159 375 -129 401
rect -63 375 -33 401
rect 33 375 63 401
rect 129 375 159 401
rect 225 375 255 401
rect 321 375 351 401
rect 417 375 447 401
rect -447 -397 -417 -375
rect -351 -397 -321 -375
rect -255 -397 -225 -375
rect -159 -397 -129 -375
rect -483 -413 -417 -397
rect -483 -447 -467 -413
rect -433 -447 -417 -413
rect -483 -463 -417 -447
rect -369 -413 -303 -397
rect -369 -447 -353 -413
rect -319 -447 -303 -413
rect -369 -463 -303 -447
rect -255 -413 -129 -397
rect -255 -447 -239 -413
rect -145 -447 -129 -413
rect -255 -463 -129 -447
rect -63 -397 -33 -375
rect 33 -397 63 -375
rect -63 -413 63 -397
rect -63 -447 -47 -413
rect 47 -447 63 -413
rect -63 -463 63 -447
rect 129 -397 159 -375
rect 225 -397 255 -375
rect 321 -397 351 -375
rect 417 -397 447 -375
rect 129 -413 255 -397
rect 129 -447 145 -413
rect 239 -447 255 -413
rect 129 -463 255 -447
rect 303 -413 369 -397
rect 303 -447 319 -413
rect 353 -447 369 -413
rect 303 -463 369 -447
rect 417 -413 483 -397
rect 417 -447 433 -413
rect 467 -447 483 -413
rect 417 -463 483 -447
<< polycont >>
rect -467 -447 -433 -413
rect -353 -447 -319 -413
rect -239 -447 -145 -413
rect -47 -447 47 -413
rect 145 -447 239 -413
rect 319 -447 353 -413
rect 433 -447 467 -413
<< locali >>
rect -611 515 -515 549
rect 515 515 611 549
rect -611 453 -577 515
rect 577 453 611 515
rect -497 363 -463 379
rect -497 -379 -463 -363
rect -401 363 -367 379
rect -401 -379 -367 -363
rect -305 363 -271 379
rect -305 -379 -271 -363
rect -209 363 -175 379
rect -209 -379 -175 -363
rect -113 363 -79 379
rect -113 -379 -79 -363
rect -17 363 17 379
rect -17 -379 17 -363
rect 79 363 113 379
rect 79 -379 113 -363
rect 175 363 209 379
rect 175 -379 209 -363
rect 271 363 305 379
rect 271 -379 305 -363
rect 367 363 401 379
rect 367 -379 401 -363
rect 463 363 497 379
rect 463 -379 497 -363
rect -483 -447 -467 -413
rect -433 -447 -417 -413
rect -369 -447 -353 -413
rect -319 -447 -303 -413
rect -255 -447 -239 -413
rect -145 -447 -129 -413
rect -63 -447 -47 -413
rect 47 -447 63 -413
rect 129 -447 145 -413
rect 239 -447 255 -413
rect 303 -447 319 -413
rect 353 -447 369 -413
rect 417 -447 433 -413
rect 467 -447 483 -413
rect -611 -515 -577 -453
rect 577 -515 611 -453
rect -611 -549 -515 -515
rect 515 -549 611 -515
<< viali >>
rect -497 -363 -463 363
rect -401 -363 -367 363
rect -305 -363 -271 363
rect -209 -363 -175 363
rect -113 -363 -79 363
rect -17 -363 17 363
rect 79 -363 113 363
rect 175 -363 209 363
rect 271 -363 305 363
rect 367 -363 401 363
rect 463 -363 497 363
rect -353 -447 -319 -413
rect -239 -447 -145 -413
rect -47 -447 47 -413
rect 145 -447 239 -413
rect 319 -447 353 -413
<< metal1 >>
rect -503 363 -457 375
rect -503 -363 -497 363
rect -463 -363 -457 363
rect -503 -375 -457 -363
rect -407 363 -361 375
rect -407 -363 -401 363
rect -367 -363 -361 363
rect -407 -375 -361 -363
rect -311 363 -265 375
rect -311 -363 -305 363
rect -271 -363 -265 363
rect -311 -375 -265 -363
rect -215 363 -169 375
rect -215 -363 -209 363
rect -175 -363 -169 363
rect -215 -375 -169 -363
rect -119 363 -73 375
rect -119 -363 -113 363
rect -79 -363 -73 363
rect -119 -375 -73 -363
rect -23 363 23 375
rect -23 -363 -17 363
rect 17 -363 23 363
rect -23 -375 23 -363
rect 73 363 119 375
rect 73 -363 79 363
rect 113 -363 119 363
rect 73 -375 119 -363
rect 169 363 215 375
rect 169 -363 175 363
rect 209 -363 215 363
rect 169 -375 215 -363
rect 265 363 311 375
rect 265 -363 271 363
rect 305 -363 311 363
rect 265 -375 311 -363
rect 361 363 407 375
rect 361 -363 367 363
rect 401 -363 407 363
rect 361 -375 407 -363
rect 457 363 503 375
rect 457 -363 463 363
rect 497 -363 503 363
rect 457 -375 503 -363
rect -365 -413 -307 -407
rect -365 -447 -353 -413
rect -319 -447 -307 -413
rect -365 -453 -307 -447
rect -251 -413 -133 -407
rect -251 -447 -239 -413
rect -145 -447 -133 -413
rect -251 -453 -133 -447
rect -59 -413 59 -407
rect -59 -447 -47 -413
rect 47 -447 59 -413
rect -59 -453 59 -447
rect 133 -413 251 -407
rect 133 -447 145 -413
rect 239 -447 251 -413
rect 133 -453 251 -447
rect 307 -413 365 -407
rect 307 -447 319 -413
rect 353 -447 365 -413
rect 307 -453 365 -447
<< properties >>
string FIXED_BBOX -594 -532 594 532
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 3.75 l 0.150 m 1 nf 10 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
