magic
tech sky130A
magscale 1 2
timestamp 1695375165
<< nwell >>
rect -363 -319 363 319
<< pmos >>
rect -167 -100 -127 100
rect -69 -100 -29 100
rect 29 -100 69 100
rect 127 -100 167 100
<< pdiff >>
rect -225 88 -167 100
rect -225 -88 -213 88
rect -179 -88 -167 88
rect -225 -100 -167 -88
rect -127 88 -69 100
rect -127 -88 -115 88
rect -81 -88 -69 88
rect -127 -100 -69 -88
rect -29 88 29 100
rect -29 -88 -17 88
rect 17 -88 29 88
rect -29 -100 29 -88
rect 69 88 127 100
rect 69 -88 81 88
rect 115 -88 127 88
rect 69 -100 127 -88
rect 167 88 225 100
rect 167 -88 179 88
rect 213 -88 225 88
rect 167 -100 225 -88
<< pdiffc >>
rect -213 -88 -179 88
rect -115 -88 -81 88
rect -17 -88 17 88
rect 81 -88 115 88
rect 179 -88 213 88
<< nsubdiff >>
rect -327 249 -231 283
rect 231 249 327 283
rect -327 187 -293 249
rect 293 187 327 249
rect -327 -249 -293 -187
rect 293 -249 327 -187
rect -327 -283 -231 -249
rect 231 -283 327 -249
<< nsubdiffcont >>
rect -231 249 231 283
rect -327 -187 -293 187
rect 293 -187 327 187
rect -231 -283 231 -249
<< poly >>
rect -69 181 69 197
rect -69 147 -53 181
rect 53 147 69 181
rect -69 131 69 147
rect -167 100 -127 126
rect -69 100 -29 131
rect 29 100 69 131
rect 127 100 167 131
rect -167 -131 -127 -100
rect -69 -131 -29 -100
rect 29 -131 69 -100
rect 127 -131 167 -100
rect -180 -147 -114 -131
rect -180 -181 -164 -147
rect -130 -181 -114 -147
rect -180 -197 -114 -181
rect 114 -147 180 -131
rect 114 -181 130 -147
rect 164 -181 180 -147
rect 114 -197 180 -181
<< polycont >>
rect -53 147 53 181
rect -164 -181 -130 -147
rect 130 -181 164 -147
<< locali >>
rect -327 249 -231 283
rect 231 249 327 283
rect -327 187 -293 249
rect 293 187 327 249
rect -69 147 -53 181
rect 53 147 69 181
rect -213 88 -179 104
rect -213 -104 -179 -88
rect -115 88 -81 104
rect -115 -104 -81 -88
rect -17 88 17 104
rect -17 -104 17 -88
rect 81 88 115 104
rect 179 99 213 104
rect 81 -104 115 -88
rect 177 88 293 99
rect 177 -88 179 88
rect 213 -88 293 88
rect 177 -101 293 -88
rect 179 -104 213 -101
rect 114 -147 293 -143
rect -180 -181 -164 -147
rect -130 -181 -114 -147
rect 114 -181 130 -147
rect 164 -181 293 -147
rect 114 -185 293 -181
rect -327 -249 -293 -187
rect 293 -249 327 -187
rect -327 -283 -231 -249
rect 231 -283 327 -249
<< viali >>
rect -53 147 53 181
rect -213 -88 -179 88
rect -115 -88 -81 88
rect -17 -88 17 88
rect 81 -88 115 88
rect 179 -88 213 88
<< metal1 >>
rect -65 181 65 187
rect -65 147 -53 181
rect 53 147 65 181
rect -65 141 65 147
rect -219 88 -173 100
rect -219 -88 -213 88
rect -179 -88 -173 88
rect -219 -100 -173 -88
rect -121 88 -75 100
rect -121 -88 -115 88
rect -81 -88 -75 88
rect -121 -100 -75 -88
rect -23 88 23 100
rect -23 -88 -17 88
rect 17 -88 23 88
rect -23 -100 23 -88
rect 75 88 121 100
rect 75 -88 81 88
rect 115 -88 121 88
rect 75 -100 121 -88
rect 173 88 219 100
rect 173 -88 179 88
rect 213 -88 219 88
rect 173 -100 219 -88
<< properties >>
string FIXED_BBOX -310 -266 310 266
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 1 l 0.2 m 1 nf 4 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
