magic
tech sky130A
magscale 1 2
timestamp 1699054381
<< metal3 >>
rect -30 60 30 117
rect -30 -117 30 -60
<< rmetal3 >>
rect -30 -60 30 60
<< properties >>
string gencell sky130_fd_pr__res_generic_m3
string library sky130
string parameters w 0.3 l 0.6 m 1 nx 1 wmin 0.30 lmin 0.30 rho 0.047 val 94.0m dummy 0 dw 0.0 term 0.0 roverlap 0
<< end >>
