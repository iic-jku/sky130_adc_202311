magic
tech sky130A
magscale 1 2
timestamp 1699972208
<< metal1 >>
rect -1624 54698 -1504 54704
rect -1624 46688 -1504 54578
rect -1252 54688 -1132 54694
rect -1630 46568 -1624 46688
rect -1504 46568 -1498 46688
rect -1252 45502 -1132 54568
rect -1258 45382 -1252 45502
rect -1132 45382 -1126 45502
rect 89942 19068 89998 19074
rect 89998 19012 95240 19068
rect 95296 19012 95302 19068
rect 89942 19006 89998 19012
rect 89942 -916 89998 -910
rect 89942 -2620 89998 -972
rect 89936 -2676 89942 -2620
rect 89998 -2676 90004 -2620
<< via1 >>
rect -1624 54578 -1504 54698
rect -1252 54568 -1132 54688
rect -1624 46568 -1504 46688
rect -1252 45382 -1132 45502
rect 89942 19012 89998 19068
rect 95240 19012 95296 19068
rect 89942 -972 89998 -916
rect 89942 -2676 89998 -2620
<< metal2 >>
rect 94070 243762 94130 243771
rect 94070 243693 94130 243702
rect 94072 154352 94128 243693
rect 95708 241404 95768 241413
rect 95708 241335 95768 241344
rect 94061 154292 94070 154352
rect 94130 154292 94139 154352
rect 94072 109933 94128 154292
rect 94852 152008 94972 152017
rect 94070 109924 94130 109933
rect 94070 109855 94130 109864
rect -1619 82306 -1509 82310
rect -1624 82301 93630 82306
rect -1624 82191 -1619 82301
rect -1509 82191 93630 82301
rect -1624 82186 93630 82191
rect 93750 82186 93759 82306
rect -1619 82182 -1509 82186
rect 94072 81862 94128 109855
rect 94425 107496 94434 107556
rect 94494 107496 94503 107556
rect -13896 81806 94128 81862
rect -13896 64 -13840 81806
rect -1266 81621 -1122 81636
rect -1266 81604 -1247 81621
rect -11806 81548 -1247 81604
rect -11806 80092 -11750 81548
rect -1266 81511 -1247 81548
rect -1137 81604 -1122 81621
rect 94436 81604 94492 107496
rect 94852 82301 94972 151888
rect 94852 82191 94857 82301
rect 94967 82191 94972 82301
rect 94852 82186 94972 82191
rect 94857 82182 94967 82186
rect -1137 81548 94492 81604
rect -1137 81511 -1122 81548
rect -1266 81498 -1122 81511
rect 88470 81103 88628 81130
rect 88470 81076 88487 81103
rect -6838 81020 88487 81076
rect -6838 80092 -6782 81020
rect 88470 80993 88487 81020
rect 88597 81076 88628 81103
rect 95710 81076 95766 241335
rect 88597 81020 95766 81076
rect 88597 80993 88628 81020
rect 88470 80974 88628 80993
rect -1624 79700 -1504 79709
rect -1624 54698 -1504 79580
rect -1252 79686 -1132 79695
rect -1630 54578 -1624 54698
rect -1504 54578 -1498 54698
rect -1252 54688 -1132 79566
rect 89940 65488 90000 65497
rect 89940 65419 90000 65428
rect -1258 54568 -1252 54688
rect -1132 54568 -1126 54688
rect -3452 53588 86 53708
rect 206 53588 215 53708
rect -4629 50324 -4519 50328
rect -3452 50324 -3332 53588
rect -3070 52092 98 52212
rect 218 52092 227 52212
rect -4634 50319 -3322 50324
rect -4634 50209 -4629 50319
rect -4519 50209 -3322 50319
rect -4634 50204 -3322 50209
rect -4629 50200 -4519 50204
rect -3973 48964 -3863 48968
rect -3070 48964 -2950 52092
rect -3978 48959 -2950 48964
rect -3978 48849 -3973 48959
rect -3863 48849 -2950 48959
rect -3978 48844 -2950 48849
rect -2740 50604 92 50724
rect 212 50604 221 50724
rect -3973 48840 -3863 48844
rect -3677 47604 -3567 47608
rect -2740 47604 -2620 50604
rect -3682 47599 -2620 47604
rect -3682 47489 -3677 47599
rect -3567 47489 -2620 47599
rect -3682 47484 -2620 47489
rect -2436 49102 92 49222
rect 212 49102 221 49222
rect -3677 47480 -3567 47484
rect -3865 46244 -3755 46248
rect -2436 46244 -2316 49102
rect -3870 46239 -2316 46244
rect -3870 46129 -3865 46239
rect -3755 46129 -2316 46239
rect -3870 46124 -2316 46129
rect -2152 47600 92 47720
rect 212 47600 221 47720
rect -3865 46120 -3755 46124
rect -3859 44884 -3749 44888
rect -2152 44884 -2032 47600
rect -1624 46688 -1504 46694
rect -1624 46227 -1504 46568
rect -1628 46117 -1619 46227
rect -1509 46117 -1500 46227
rect -1624 46112 -1504 46117
rect 88482 46060 88602 46069
rect -1252 45502 -1132 45508
rect -1252 45097 -1132 45382
rect -1256 44987 -1247 45097
rect -1137 44987 -1128 45097
rect -1252 44982 -1132 44987
rect -3864 44879 -2032 44884
rect -3864 44769 -3859 44879
rect -3749 44769 -2032 44879
rect -3864 44764 -2032 44769
rect -3859 44760 -3749 44764
rect 88482 40243 88602 45940
rect 88482 40133 88487 40243
rect 88597 40133 88602 40243
rect 88482 40128 88602 40133
rect 88487 40124 88597 40128
rect -4225 21764 -4115 21768
rect -4230 21759 -320 21764
rect -4230 21649 -4225 21759
rect -4115 21649 -320 21759
rect -4230 21644 -320 21649
rect -4225 21640 -4115 21644
rect -4225 20404 -4115 20408
rect -4230 20399 -618 20404
rect -4230 20289 -4225 20399
rect -4115 20289 -618 20399
rect -4230 20284 -618 20289
rect -4225 20280 -4115 20284
rect -4225 19044 -4115 19048
rect -4230 19039 -928 19044
rect -4230 18929 -4225 19039
rect -4115 18929 -928 19039
rect -4230 18924 -928 18929
rect -4225 18920 -4115 18924
rect -4217 17684 -4107 17688
rect -4222 17679 -1338 17684
rect -4222 17569 -4217 17679
rect -4107 17569 -1338 17679
rect -4222 17564 -1338 17569
rect -4217 17560 -4107 17564
rect -4219 16324 -4109 16328
rect -4224 16319 -1768 16324
rect -4224 16209 -4219 16319
rect -4109 16209 -1768 16319
rect -4224 16204 -1768 16209
rect -4219 16200 -4109 16204
rect -1888 11824 -1768 16204
rect -1458 13324 -1338 17564
rect -1048 14820 -928 18924
rect -738 16318 -618 20284
rect -446 17804 -326 21644
rect 89942 19068 89998 65419
rect 95228 19070 95310 19080
rect 89936 19012 89942 19068
rect 89998 19012 90004 19068
rect -446 17640 -326 17684
rect -738 16189 -618 16198
rect -1048 14630 -928 14700
rect -1458 13195 -1338 13204
rect -1888 11704 -338 11824
rect -218 11704 -209 11824
rect -13462 64 -13406 600
rect -13896 8 -13406 64
rect -13462 -2620 -13406 8
rect -11806 -2388 -11750 204
rect -10150 -2186 -10094 720
rect -8494 -1942 -8438 634
rect -6838 -1608 -6782 556
rect -5182 -1222 -5126 216
rect 89942 -916 89998 19012
rect 95228 19010 95238 19070
rect 95298 19010 95310 19070
rect 95228 19000 95310 19010
rect 89936 -972 89942 -916
rect 89998 -972 90004 -916
rect -5182 -1278 94620 -1222
rect -6838 -1664 94234 -1608
rect -8494 -1998 93822 -1942
rect -10150 -2242 93482 -2186
rect -11806 -2444 93184 -2388
rect 89942 -2620 89998 -2614
rect -13462 -2676 89942 -2620
rect 89998 -2676 92982 -2620
rect 89942 -2682 89998 -2676
rect 92926 -26148 92982 -2676
rect 92915 -26208 92924 -26148
rect 92984 -26208 92993 -26148
rect 92926 -70572 92982 -26208
rect 92915 -70632 92924 -70572
rect 92984 -70632 92993 -70572
rect 93128 -250576 93184 -2444
rect 93117 -250636 93126 -250576
rect 93186 -250636 93195 -250576
rect 93128 -295235 93184 -250636
rect 93426 -251763 93482 -2242
rect 93766 -72927 93822 -1998
rect 94178 -28495 94234 -1664
rect 94176 -28504 94236 -28495
rect 94176 -28573 94236 -28564
rect 93764 -72936 93824 -72927
rect 93764 -73005 93824 -72996
rect 93424 -251772 93484 -251763
rect 93424 -251841 93484 -251832
rect 93126 -295244 93186 -295235
rect 93126 -295313 93186 -295304
rect 94564 -296420 94620 -1278
rect 94548 -296426 94640 -296420
rect 94548 -296486 94562 -296426
rect 94622 -296486 94640 -296426
rect 94548 -296492 94640 -296486
<< via2 >>
rect 94070 243702 94130 243762
rect 95708 241344 95768 241404
rect 94070 154292 94130 154352
rect 94852 151888 94972 152008
rect 94070 109864 94130 109924
rect -1619 82191 -1509 82301
rect 93630 82186 93750 82306
rect 94434 107496 94494 107556
rect -1247 81511 -1137 81621
rect 94857 82191 94967 82301
rect 88487 80993 88597 81103
rect -1624 79580 -1504 79700
rect -1252 79566 -1132 79686
rect 89940 65428 90000 65488
rect 86 53588 206 53708
rect 98 52092 218 52212
rect -4629 50209 -4519 50319
rect -3973 48849 -3863 48959
rect 92 50604 212 50724
rect -3677 47489 -3567 47599
rect 92 49102 212 49222
rect -3865 46129 -3755 46239
rect 92 47600 212 47720
rect -1619 46117 -1509 46227
rect 88482 45940 88602 46060
rect -1247 44987 -1137 45097
rect -3859 44769 -3749 44879
rect 88487 40133 88597 40243
rect -4225 21649 -4115 21759
rect -4225 20289 -4115 20399
rect -4225 18929 -4115 19039
rect -4217 17569 -4107 17679
rect -4219 16209 -4109 16319
rect -446 17684 -326 17804
rect -738 16198 -618 16318
rect -1048 14700 -928 14820
rect -1458 13204 -1338 13324
rect -338 11704 -218 11824
rect 95238 19068 95298 19070
rect 95238 19012 95240 19068
rect 95240 19012 95296 19068
rect 95296 19012 95298 19068
rect 95238 19010 95298 19012
rect 92924 -26208 92984 -26148
rect 92924 -70632 92984 -70572
rect 93126 -250636 93186 -250576
rect 94176 -28564 94236 -28504
rect 93764 -72996 93824 -72936
rect 93424 -251832 93484 -251772
rect 93126 -295304 93186 -295244
rect 94562 -296486 94622 -296426
<< metal3 >>
rect 145344 297650 148518 297652
rect 84678 295190 84684 297650
rect 87144 295190 148518 297650
rect 84732 285130 84738 287590
rect 87198 285130 148520 287590
rect 94065 243762 94135 243767
rect 94065 243702 94070 243762
rect 94130 243702 148442 243762
rect 94065 243697 94135 243702
rect 95703 241404 95773 241409
rect 95703 241344 95708 241404
rect 95768 241344 149698 241404
rect 95703 241339 95773 241344
rect 94065 154352 94135 154357
rect 94065 154292 94070 154352
rect 94130 154292 148738 154352
rect 94065 154287 94135 154292
rect 94847 152008 94977 152013
rect 149392 152008 149698 152010
rect 94847 151888 94852 152008
rect 94972 151888 149698 152008
rect 94847 151883 94977 151888
rect 94065 109924 94135 109929
rect 94065 109864 94070 109924
rect 94130 109864 148654 109924
rect 94065 109859 94135 109864
rect 94429 107556 94499 107561
rect 94429 107496 94434 107556
rect 94494 107496 149698 107556
rect 94429 107491 94499 107496
rect 93625 82306 93755 82311
rect -1624 82301 -1504 82306
rect -1624 82191 -1619 82301
rect -1509 82191 -1504 82301
rect -1624 79705 -1504 82191
rect 93625 82186 93630 82306
rect 93750 82301 94972 82306
rect 93750 82191 94857 82301
rect 94967 82191 94972 82301
rect 93750 82186 94972 82191
rect 93625 82181 93755 82186
rect -1252 81621 -1132 81638
rect -1252 81511 -1247 81621
rect -1137 81511 -1132 81621
rect -1629 79700 -1499 79705
rect -1629 79580 -1624 79700
rect -1504 79580 -1499 79700
rect -1252 79691 -1132 81511
rect 88482 81103 88602 81130
rect 88482 80993 88487 81103
rect 88597 80993 88602 81103
rect -1629 79575 -1499 79580
rect -1257 79686 -1127 79691
rect -1257 79566 -1252 79686
rect -1132 79566 -1127 79686
rect -1257 79561 -1127 79566
rect -4292 79024 634 79144
rect -4292 73444 -4172 79024
rect -4462 73324 -4172 73444
rect -4020 77526 456 77646
rect -4020 72084 -3900 77526
rect -4572 71964 -3900 72084
rect -3840 76032 816 76152
rect -3840 70724 -3720 76032
rect -4648 70604 -3720 70724
rect -3622 74532 496 74652
rect -3622 69364 -3502 74532
rect -4488 69244 -3502 69364
rect -3424 73040 596 73160
rect -3424 68004 -3304 73040
rect -4620 67884 -3304 68004
rect -3146 71544 540 71664
rect -3146 66644 -3026 71544
rect -4506 66524 -3026 66644
rect -2894 70046 626 70166
rect -2894 65284 -2774 70046
rect -4702 65164 -2774 65284
rect -2646 68552 644 68672
rect -2646 63924 -2526 68552
rect -4428 63804 -2526 63924
rect -2400 67058 644 67178
rect -2400 62564 -2280 67058
rect -4602 62444 -2280 62564
rect -2122 65556 634 65676
rect -2122 61204 -2002 65556
rect -4500 61084 -2002 61204
rect -1892 64062 594 64182
rect -1892 59844 -1772 64062
rect -4546 59724 -1772 59844
rect -1646 62566 410 62686
rect -1646 58484 -1526 62566
rect -4534 58364 -1526 58484
rect -1396 61074 488 61194
rect -1396 57124 -1276 61074
rect -4676 57004 -1276 57124
rect -1100 59570 558 59690
rect -1100 55764 -980 59570
rect -4654 55644 -980 55764
rect -816 58078 532 58198
rect -816 54404 -696 58078
rect -4458 54284 -696 54404
rect -548 56582 576 56702
rect -548 53044 -428 56582
rect -4468 52924 -428 53044
rect -308 55088 600 55208
rect -308 51684 -188 55088
rect 81 53708 211 53713
rect 81 53588 86 53708
rect 206 53588 634 53708
rect 81 53583 211 53588
rect 93 52212 223 52217
rect 93 52092 98 52212
rect 218 52092 732 52212
rect 93 52087 223 52092
rect -4446 51564 -188 51684
rect 87 50724 217 50729
rect 87 50604 92 50724
rect 212 50604 708 50724
rect 87 50599 217 50604
rect -4634 50319 -4514 50324
rect -4634 50209 -4629 50319
rect -4519 50209 -4514 50319
rect -4634 50204 -4514 50209
rect 87 49222 217 49227
rect 87 49102 92 49222
rect 212 49102 486 49222
rect 87 49097 217 49102
rect -4526 48959 -3858 48964
rect -4526 48849 -3973 48959
rect -3863 48849 -3858 48959
rect -4526 48844 -3858 48849
rect 87 47720 217 47725
rect -4698 47599 -3562 47604
rect -4698 47489 -3677 47599
rect -3567 47489 -3562 47599
rect 87 47600 92 47720
rect 212 47600 588 47720
rect 87 47595 217 47600
rect -4698 47484 -3562 47489
rect -4458 46239 -3750 46244
rect -4458 46129 -3865 46239
rect -3755 46129 -3750 46239
rect -4458 46124 -3750 46129
rect -1624 46227 264 46232
rect -1624 46117 -1619 46227
rect -1509 46117 264 46227
rect -1624 46112 264 46117
rect 88482 46065 88602 80993
rect 89935 65488 90005 65493
rect 89935 65428 89940 65488
rect 90000 65428 147572 65488
rect 89935 65423 90005 65428
rect 93510 59508 149698 59620
rect 88477 46060 88607 46065
rect 88477 45940 88482 46060
rect 88602 45940 88607 46060
rect 88477 45935 88607 45940
rect -1252 45097 -1132 45102
rect -1252 44987 -1247 45097
rect -1137 44987 -1132 45097
rect -4538 44879 -3744 44884
rect -4538 44769 -3859 44879
rect -3749 44769 -3744 44879
rect -4538 44764 -3744 44769
rect -1252 44736 -1132 44987
rect -1252 44616 210 44736
rect 93510 44417 93622 59508
rect 84476 44297 93622 44417
rect 93510 44296 93622 44297
rect -4472 43404 -3740 43524
rect -3860 43238 -3740 43404
rect 93512 43296 93624 43298
rect -3860 43118 550 43238
rect 84414 43176 93624 43296
rect -4546 42044 -3738 42164
rect -3858 41742 -3738 42044
rect -3858 41622 486 41742
rect -4496 40684 156 40804
rect -4492 39324 -142 39444
rect -4498 37964 -418 38084
rect -4522 36604 -734 36724
rect -4434 35244 -1034 35364
rect -4628 33884 -1328 34004
rect -4498 32524 -1598 32644
rect -4428 31164 -1938 31284
rect -4492 29804 -2196 29924
rect -4480 28444 -2506 28564
rect -4498 27084 -2806 27204
rect -4458 25724 -3094 25844
rect -4516 24364 -3410 24484
rect -4516 23004 -3728 23124
rect -4678 21759 -4110 21764
rect -4678 21649 -4225 21759
rect -4115 21649 -4110 21759
rect -4678 21644 -4110 21649
rect -4542 20399 -4110 20404
rect -4542 20289 -4225 20399
rect -4115 20289 -4110 20399
rect -4542 20284 -4110 20289
rect -3848 19304 -3728 23004
rect -3530 20796 -3410 24364
rect -3214 22292 -3094 25724
rect -2926 23794 -2806 27084
rect -2626 25290 -2506 28444
rect -2316 26780 -2196 29804
rect -2058 28278 -1938 31164
rect -1718 29772 -1598 32524
rect -1448 31268 -1328 33884
rect -1154 32766 -1034 35244
rect -854 34264 -734 36604
rect -538 35758 -418 37964
rect -262 37260 -142 39324
rect 36 38752 156 40684
rect 84194 40243 88602 40248
rect 84194 40133 88487 40243
rect 88597 40133 88602 40243
rect 84194 40128 88602 40133
rect 36 38632 384 38752
rect -262 37140 550 37260
rect -538 35638 574 35758
rect -854 34144 620 34264
rect -1154 32646 468 32766
rect -1448 31148 550 31268
rect -1718 29652 504 29772
rect -2058 28158 568 28278
rect -2316 26660 438 26780
rect -2626 25170 532 25290
rect -2926 23674 568 23794
rect -3214 22172 562 22292
rect -3530 20676 562 20796
rect -3848 19184 492 19304
rect -4530 19039 -4110 19044
rect -4530 18929 -4225 19039
rect -4115 18929 -4110 19039
rect -4530 18924 -4110 18929
rect -462 17804 -302 17814
rect -462 17684 -446 17804
rect -326 17684 634 17804
rect -4464 17679 -4102 17684
rect -4464 17569 -4217 17679
rect -4107 17569 -4102 17679
rect -462 17670 -302 17684
rect -4464 17564 -4102 17569
rect -4478 16319 -4104 16324
rect -4478 16209 -4219 16319
rect -4109 16209 -4104 16319
rect -4478 16204 -4104 16209
rect -743 16318 -613 16323
rect -743 16198 -738 16318
rect -618 16198 544 16318
rect -743 16193 -613 16198
rect -4476 14844 -1628 14964
rect -4488 13484 -1868 13604
rect -4464 12124 -2230 12244
rect -4488 10764 -2526 10884
rect -4514 9404 -2858 9524
rect -4478 8044 -3142 8164
rect -4628 6684 -3486 6804
rect -3606 1348 -3486 6684
rect -3262 2854 -3142 8044
rect -2978 4336 -2858 9404
rect -2646 5836 -2526 10764
rect -2350 7340 -2230 12124
rect -1988 8834 -1868 13484
rect -1748 10324 -1628 14844
rect -1070 14820 -916 14826
rect -1070 14700 -1048 14820
rect -928 14700 562 14820
rect -1070 14690 -916 14700
rect -1463 13324 -1333 13329
rect -1463 13204 -1458 13324
rect -1338 13204 472 13324
rect -1463 13199 -1333 13204
rect 93512 13198 93624 43176
rect 95233 19070 95303 19075
rect 95233 19010 95238 19070
rect 95298 19010 147006 19070
rect 95233 19005 95303 19010
rect 93512 13086 149698 13198
rect -343 11824 -213 11829
rect -343 11704 -338 11824
rect -218 11704 474 11824
rect -343 11699 -213 11704
rect -1748 10204 588 10324
rect -1988 8714 630 8834
rect -2350 7220 660 7340
rect -2646 5716 612 5836
rect -2978 4216 518 4336
rect -3262 2734 584 2854
rect -3606 1228 658 1348
rect 92919 -26148 92989 -26143
rect 92919 -26208 92924 -26148
rect 92984 -26208 148806 -26148
rect 92919 -26213 92989 -26208
rect 94171 -28504 94241 -28499
rect 94171 -28564 94176 -28504
rect 94236 -28564 149698 -28504
rect 94171 -28569 94241 -28564
rect 92919 -70572 92989 -70567
rect 92919 -70632 92924 -70572
rect 92984 -70632 148610 -70572
rect 92919 -70637 92989 -70632
rect 93759 -72936 93829 -72931
rect 93759 -72996 93764 -72936
rect 93824 -72996 149698 -72936
rect 93759 -73001 93829 -72996
rect 84776 -153242 84782 -150782
rect 87242 -150784 147906 -150782
rect 87242 -153242 148518 -150784
rect 84776 -163144 84782 -160684
rect 87242 -163144 148518 -160684
rect 93121 -250576 93191 -250571
rect 93121 -250636 93126 -250576
rect 93186 -250636 149306 -250576
rect 93121 -250641 93191 -250636
rect 93419 -251772 93489 -251767
rect 93419 -251832 93424 -251772
rect 93484 -251832 149698 -251772
rect 93419 -251837 93489 -251832
rect 93121 -295244 93191 -295239
rect 93121 -295304 93126 -295244
rect 93186 -295304 149274 -295244
rect 93121 -295309 93191 -295304
rect 94548 -296426 94640 -296420
rect 94548 -296486 94562 -296426
rect 94622 -296486 149698 -296426
rect 94548 -296492 94640 -296486
<< via3 >>
rect 84684 295190 87144 297650
rect 84738 285130 87198 287590
rect 84782 -153242 87242 -150782
rect 84782 -163144 87242 -160684
<< metal4 >>
rect -14724 78718 -14404 86898
rect -11964 79752 -11644 86884
rect -6964 79726 -6644 86858
rect -4276 78686 -3956 86872
rect -416 79250 -96 86888
rect 3344 79850 3664 86888
rect 8144 79974 8464 86904
rect 12944 79988 13264 86904
rect 47590 85784 51542 85810
rect 17961 85721 21959 85745
rect 17961 81771 17985 85721
rect 21935 81771 21959 85721
rect 17961 79830 21959 81771
rect 47590 81834 47592 85784
rect 47590 80014 51542 81834
rect 17961 79514 18048 79830
rect 21858 79514 21959 79830
rect 17961 79415 21959 79514
rect 47586 79822 51542 80014
rect 47586 79558 47644 79822
rect 51488 79558 51542 79822
rect 47586 79452 51542 79558
rect 84644 79020 84964 86904
rect -15384 -7024 -15064 1150
rect -11304 -7010 -10984 832
rect -6304 -7024 -5984 832
rect -3616 -7036 -3296 872
rect -1076 -7032 -756 804
rect 4004 -7032 4324 678
rect 8804 -7032 9124 726
rect 13604 -7062 13924 726
rect 85304 -6874 85624 678
<< via4 >>
rect 84683 297650 87145 297651
rect 84683 295190 84684 297650
rect 84684 295190 87144 297650
rect 87144 295190 87145 297650
rect 84683 295189 87145 295190
rect 84737 287590 87199 287591
rect 84737 285130 84738 287590
rect 84738 285130 87198 287590
rect 87198 285130 87199 287590
rect 84737 285129 87199 285130
rect -14724 86898 -14404 87218
rect -11964 86884 -11644 87204
rect -6964 86858 -6644 87178
rect -4276 86872 -3956 87192
rect -416 86888 -96 87208
rect 3344 86888 3664 87208
rect 8144 86904 8464 87224
rect 12944 86904 13264 87224
rect 84644 86904 84964 87224
rect 17985 81771 21935 85721
rect 47592 81834 51542 85784
rect 18048 79514 21858 79830
rect 47644 79558 51488 79822
rect -15384 -7344 -15064 -7024
rect -11304 -7330 -10984 -7010
rect -6304 -7344 -5984 -7024
rect -3616 -7356 -3296 -7036
rect -1076 -7352 -756 -7032
rect 4004 -7352 4324 -7032
rect 8804 -7352 9124 -7032
rect 13604 -7382 13924 -7062
rect 85304 -7194 85624 -6874
rect 84781 -150782 87243 -150781
rect 84781 -153242 84782 -150782
rect 84782 -153242 87242 -150782
rect 87242 -153242 87243 -150782
rect 84781 -153243 87243 -153242
rect 84781 -160684 87243 -160683
rect 84781 -163144 84782 -160684
rect 84782 -163144 87242 -160684
rect 87242 -163144 87243 -160684
rect 84781 -163145 87243 -163144
<< metal5 >>
rect 83871 297651 87869 298237
rect 83871 295189 84683 297651
rect 87145 295189 87869 297651
rect 83871 287591 87869 295189
rect 83871 285129 84737 287591
rect 87199 285129 87869 287591
rect 83871 90739 87869 285129
rect -21565 87224 87869 90739
rect -21565 87218 8144 87224
rect -21565 86898 -14724 87218
rect -14404 87208 8144 87218
rect -14404 87204 -416 87208
rect -14404 86898 -11964 87204
rect -21565 86884 -11964 86898
rect -11644 87192 -416 87204
rect -11644 87178 -4276 87192
rect -11644 86884 -6964 87178
rect -21565 86858 -6964 86884
rect -6644 86872 -4276 87178
rect -3956 86888 -416 87192
rect -96 86888 3344 87208
rect 3664 86904 8144 87208
rect 8464 86904 12944 87224
rect 13264 86904 84644 87224
rect 84964 86904 87869 87224
rect 3664 86888 87869 86904
rect -3956 86872 87869 86888
rect -6644 86858 87869 86872
rect -21565 86741 87869 86858
rect -21565 46106 -17567 86741
rect 17961 85721 21959 86741
rect 47569 85808 51567 86741
rect 17961 81771 17985 85721
rect 21935 81771 21959 85721
rect 47568 85784 51567 85808
rect 47568 81834 47592 85784
rect 51542 81834 51567 85784
rect 47568 81810 51567 81834
rect 17961 81033 21959 81771
rect 47569 81091 51567 81810
rect 21858 79852 21918 79856
rect 18024 79830 21918 79852
rect 18024 79514 18048 79830
rect 21858 79514 21918 79830
rect 47620 79822 51512 79846
rect 47620 79558 47644 79822
rect 51488 79558 51512 79822
rect 47620 79534 51512 79558
rect 18024 79496 21918 79514
rect 18026 79482 21918 79496
rect -21565 -6715 -17567 34714
rect 17915 -6715 21913 105
rect 43279 -6715 47277 147
rect 66753 -6715 70751 183
rect -21565 -6874 87985 -6715
rect -21565 -7010 85304 -6874
rect -21565 -7024 -11304 -7010
rect -21565 -7344 -15384 -7024
rect -15064 -7330 -11304 -7024
rect -10984 -7024 85304 -7010
rect -10984 -7330 -6304 -7024
rect -15064 -7344 -6304 -7330
rect -5984 -7032 85304 -7024
rect -5984 -7036 -1076 -7032
rect -5984 -7344 -3616 -7036
rect -21565 -7356 -3616 -7344
rect -3296 -7352 -1076 -7036
rect -756 -7352 4004 -7032
rect 4324 -7352 8804 -7032
rect 9124 -7062 85304 -7032
rect 9124 -7352 13604 -7062
rect -3296 -7356 13604 -7352
rect -21565 -7382 13604 -7356
rect 13924 -7194 85304 -7062
rect 85624 -7194 87985 -6874
rect 13924 -7382 87985 -7194
rect -21565 -10713 87985 -7382
rect 83987 -150781 87985 -10713
rect 83987 -153243 84781 -150781
rect 87243 -153243 87985 -150781
rect 83987 -160683 87985 -153243
rect 83987 -163145 84781 -160683
rect 87243 -163145 87985 -160683
rect 83987 -163833 87985 -163145
use adc_bridge  adc_bridge_0
timestamp 1699972208
transform 1 0 -14308 0 1 148
box -1076 -4 11012 80000
use adc_top  adc_top_0
timestamp 1699972208
transform 1 0 0 0 1 0
box -1076 -4 85624 80516
<< labels >>
rlabel metal5 83871 87224 87869 285129 1 VDD
port 1 n
rlabel metal5 83987 -150781 87985 -7194 1 VSS
port 2 n
rlabel metal3 94494 107496 99972 107556 1 rst_n
port 3 n default input
rlabel metal3 95768 241344 99960 241404 1 clk
port 4 n default input
rlabel metal3 94972 151888 100020 152008 1 conv_start
port 5 n default input
rlabel metal3 94236 -28564 100026 -28504 1 load
port 7 n default input
rlabel metal3 93824 -72996 99996 -72936 1 dati
port 8 n default input
rlabel metal3 93484 -251832 100038 -251772 1 dato
port 9 n default output
rlabel metal3 93510 59508 99838 59620 1 inp_ana
port 12 n
rlabel metal3 93512 13086 100078 13198 1 inn_ana
port 13 n
rlabel metal3 93186 -295304 99274 -295244 1 tie0
port 10 n default output
rlabel metal3 92984 -70632 98610 -70572 1 tie1
port 11 n default output
rlabel metal3 94746 -296486 99336 -296426 1 conv_finish
port 6 n default output
<< end >>
