magic
tech sky130A
magscale 1 2
timestamp 1515178157
<< checkpaint >>
rect -1260 -1260 5260 5260
<< nwell >>
rect 180 224 3820 3776
<< pwell >>
rect 864 3804 1376 3946
rect 2624 3804 3136 3946
rect 54 2624 180 3136
rect 54 864 180 1376
rect 3820 2624 3946 3136
rect 3820 864 3946 1376
rect 864 54 1376 196
rect 2624 54 3136 196
<< varactor >>
rect 360 400 3640 3600
<< psubdiff >>
rect 890 3892 1350 3920
rect 890 3858 933 3892
rect 967 3858 1001 3892
rect 1035 3858 1069 3892
rect 1103 3858 1137 3892
rect 1171 3858 1205 3892
rect 1239 3858 1273 3892
rect 1307 3858 1350 3892
rect 890 3830 1350 3858
rect 2650 3892 3110 3920
rect 2650 3858 2693 3892
rect 2727 3858 2761 3892
rect 2795 3858 2829 3892
rect 2863 3858 2897 3892
rect 2931 3858 2965 3892
rect 2999 3858 3033 3892
rect 3067 3858 3110 3892
rect 2650 3830 3110 3858
rect 80 3067 154 3110
rect 80 3033 108 3067
rect 142 3033 154 3067
rect 80 2999 154 3033
rect 80 2965 108 2999
rect 142 2965 154 2999
rect 80 2931 154 2965
rect 80 2897 108 2931
rect 142 2897 154 2931
rect 80 2863 154 2897
rect 80 2829 108 2863
rect 142 2829 154 2863
rect 80 2795 154 2829
rect 80 2761 108 2795
rect 142 2761 154 2795
rect 80 2727 154 2761
rect 80 2693 108 2727
rect 142 2693 154 2727
rect 80 2650 154 2693
rect 80 1307 154 1350
rect 80 1273 108 1307
rect 142 1273 154 1307
rect 80 1239 154 1273
rect 80 1205 108 1239
rect 142 1205 154 1239
rect 80 1171 154 1205
rect 80 1137 108 1171
rect 142 1137 154 1171
rect 80 1103 154 1137
rect 80 1069 108 1103
rect 142 1069 154 1103
rect 80 1035 154 1069
rect 80 1001 108 1035
rect 142 1001 154 1035
rect 80 967 154 1001
rect 80 933 108 967
rect 142 933 154 967
rect 80 890 154 933
rect 3846 3067 3920 3110
rect 3846 3033 3858 3067
rect 3892 3033 3920 3067
rect 3846 2999 3920 3033
rect 3846 2965 3858 2999
rect 3892 2965 3920 2999
rect 3846 2931 3920 2965
rect 3846 2897 3858 2931
rect 3892 2897 3920 2931
rect 3846 2863 3920 2897
rect 3846 2829 3858 2863
rect 3892 2829 3920 2863
rect 3846 2795 3920 2829
rect 3846 2761 3858 2795
rect 3892 2761 3920 2795
rect 3846 2727 3920 2761
rect 3846 2693 3858 2727
rect 3892 2693 3920 2727
rect 3846 2650 3920 2693
rect 3846 1307 3920 1350
rect 3846 1273 3858 1307
rect 3892 1273 3920 1307
rect 3846 1239 3920 1273
rect 3846 1205 3858 1239
rect 3892 1205 3920 1239
rect 3846 1171 3920 1205
rect 3846 1137 3858 1171
rect 3892 1137 3920 1171
rect 3846 1103 3920 1137
rect 3846 1069 3858 1103
rect 3892 1069 3920 1103
rect 3846 1035 3920 1069
rect 3846 1001 3858 1035
rect 3892 1001 3920 1035
rect 3846 967 3920 1001
rect 3846 933 3858 967
rect 3892 933 3920 967
rect 3846 890 3920 933
rect 890 142 1350 170
rect 890 108 933 142
rect 967 108 1001 142
rect 1035 108 1069 142
rect 1103 108 1137 142
rect 1171 108 1205 142
rect 1239 108 1273 142
rect 1307 108 1350 142
rect 890 80 1350 108
rect 2650 142 3110 170
rect 2650 108 2693 142
rect 2727 108 2761 142
rect 2795 108 2829 142
rect 2863 108 2897 142
rect 2931 108 2965 142
rect 2999 108 3033 142
rect 3067 108 3110 142
rect 2650 80 3110 108
<< nsubdiff >>
rect 360 3703 3640 3740
rect 360 3669 448 3703
rect 482 3669 516 3703
rect 550 3669 584 3703
rect 618 3669 652 3703
rect 686 3669 720 3703
rect 754 3669 788 3703
rect 822 3669 856 3703
rect 890 3669 924 3703
rect 958 3669 992 3703
rect 1026 3669 1060 3703
rect 1094 3669 1128 3703
rect 1162 3669 1196 3703
rect 1230 3669 1264 3703
rect 1298 3669 1332 3703
rect 1366 3669 1400 3703
rect 1434 3669 1468 3703
rect 1502 3669 1536 3703
rect 1570 3669 1604 3703
rect 1638 3669 1672 3703
rect 1706 3669 1740 3703
rect 1774 3669 1808 3703
rect 1842 3669 1876 3703
rect 1910 3669 1944 3703
rect 1978 3669 2012 3703
rect 2046 3669 2080 3703
rect 2114 3669 2148 3703
rect 2182 3669 2216 3703
rect 2250 3669 2284 3703
rect 2318 3669 2352 3703
rect 2386 3669 2420 3703
rect 2454 3669 2488 3703
rect 2522 3669 2556 3703
rect 2590 3669 2624 3703
rect 2658 3669 2692 3703
rect 2726 3669 2760 3703
rect 2794 3669 2828 3703
rect 2862 3669 2896 3703
rect 2930 3669 2964 3703
rect 2998 3669 3032 3703
rect 3066 3669 3100 3703
rect 3134 3669 3168 3703
rect 3202 3669 3236 3703
rect 3270 3669 3304 3703
rect 3338 3669 3372 3703
rect 3406 3669 3440 3703
rect 3474 3669 3508 3703
rect 3542 3669 3640 3703
rect 360 3600 3640 3669
rect 360 330 3640 400
rect 360 296 448 330
rect 482 296 516 330
rect 550 296 584 330
rect 618 296 652 330
rect 686 296 720 330
rect 754 296 788 330
rect 822 296 856 330
rect 890 296 924 330
rect 958 296 992 330
rect 1026 296 1060 330
rect 1094 296 1128 330
rect 1162 296 1196 330
rect 1230 296 1264 330
rect 1298 296 1332 330
rect 1366 296 1400 330
rect 1434 296 1468 330
rect 1502 296 1536 330
rect 1570 296 1604 330
rect 1638 296 1672 330
rect 1706 296 1740 330
rect 1774 296 1808 330
rect 1842 296 1876 330
rect 1910 296 1944 330
rect 1978 296 2012 330
rect 2046 296 2080 330
rect 2114 296 2148 330
rect 2182 296 2216 330
rect 2250 296 2284 330
rect 2318 296 2352 330
rect 2386 296 2420 330
rect 2454 296 2488 330
rect 2522 296 2556 330
rect 2590 296 2624 330
rect 2658 296 2692 330
rect 2726 296 2760 330
rect 2794 296 2828 330
rect 2862 296 2896 330
rect 2930 296 2964 330
rect 2998 296 3032 330
rect 3066 296 3100 330
rect 3134 296 3168 330
rect 3202 296 3236 330
rect 3270 296 3304 330
rect 3338 296 3372 330
rect 3406 296 3440 330
rect 3474 296 3508 330
rect 3542 296 3640 330
rect 360 260 3640 296
<< psubdiffcont >>
rect 933 3858 967 3892
rect 1001 3858 1035 3892
rect 1069 3858 1103 3892
rect 1137 3858 1171 3892
rect 1205 3858 1239 3892
rect 1273 3858 1307 3892
rect 2693 3858 2727 3892
rect 2761 3858 2795 3892
rect 2829 3858 2863 3892
rect 2897 3858 2931 3892
rect 2965 3858 2999 3892
rect 3033 3858 3067 3892
rect 108 3033 142 3067
rect 108 2965 142 2999
rect 108 2897 142 2931
rect 108 2829 142 2863
rect 108 2761 142 2795
rect 108 2693 142 2727
rect 108 1273 142 1307
rect 108 1205 142 1239
rect 108 1137 142 1171
rect 108 1069 142 1103
rect 108 1001 142 1035
rect 108 933 142 967
rect 3858 3033 3892 3067
rect 3858 2965 3892 2999
rect 3858 2897 3892 2931
rect 3858 2829 3892 2863
rect 3858 2761 3892 2795
rect 3858 2693 3892 2727
rect 3858 1273 3892 1307
rect 3858 1205 3892 1239
rect 3858 1137 3892 1171
rect 3858 1069 3892 1103
rect 3858 1001 3892 1035
rect 3858 933 3892 967
rect 933 108 967 142
rect 1001 108 1035 142
rect 1069 108 1103 142
rect 1137 108 1171 142
rect 1205 108 1239 142
rect 1273 108 1307 142
rect 2693 108 2727 142
rect 2761 108 2795 142
rect 2829 108 2863 142
rect 2897 108 2931 142
rect 2965 108 2999 142
rect 3033 108 3067 142
<< nsubdiffcont >>
rect 448 3669 482 3703
rect 516 3669 550 3703
rect 584 3669 618 3703
rect 652 3669 686 3703
rect 720 3669 754 3703
rect 788 3669 822 3703
rect 856 3669 890 3703
rect 924 3669 958 3703
rect 992 3669 1026 3703
rect 1060 3669 1094 3703
rect 1128 3669 1162 3703
rect 1196 3669 1230 3703
rect 1264 3669 1298 3703
rect 1332 3669 1366 3703
rect 1400 3669 1434 3703
rect 1468 3669 1502 3703
rect 1536 3669 1570 3703
rect 1604 3669 1638 3703
rect 1672 3669 1706 3703
rect 1740 3669 1774 3703
rect 1808 3669 1842 3703
rect 1876 3669 1910 3703
rect 1944 3669 1978 3703
rect 2012 3669 2046 3703
rect 2080 3669 2114 3703
rect 2148 3669 2182 3703
rect 2216 3669 2250 3703
rect 2284 3669 2318 3703
rect 2352 3669 2386 3703
rect 2420 3669 2454 3703
rect 2488 3669 2522 3703
rect 2556 3669 2590 3703
rect 2624 3669 2658 3703
rect 2692 3669 2726 3703
rect 2760 3669 2794 3703
rect 2828 3669 2862 3703
rect 2896 3669 2930 3703
rect 2964 3669 2998 3703
rect 3032 3669 3066 3703
rect 3100 3669 3134 3703
rect 3168 3669 3202 3703
rect 3236 3669 3270 3703
rect 3304 3669 3338 3703
rect 3372 3669 3406 3703
rect 3440 3669 3474 3703
rect 3508 3669 3542 3703
rect 448 296 482 330
rect 516 296 550 330
rect 584 296 618 330
rect 652 296 686 330
rect 720 296 754 330
rect 788 296 822 330
rect 856 296 890 330
rect 924 296 958 330
rect 992 296 1026 330
rect 1060 296 1094 330
rect 1128 296 1162 330
rect 1196 296 1230 330
rect 1264 296 1298 330
rect 1332 296 1366 330
rect 1400 296 1434 330
rect 1468 296 1502 330
rect 1536 296 1570 330
rect 1604 296 1638 330
rect 1672 296 1706 330
rect 1740 296 1774 330
rect 1808 296 1842 330
rect 1876 296 1910 330
rect 1944 296 1978 330
rect 2012 296 2046 330
rect 2080 296 2114 330
rect 2148 296 2182 330
rect 2216 296 2250 330
rect 2284 296 2318 330
rect 2352 296 2386 330
rect 2420 296 2454 330
rect 2488 296 2522 330
rect 2556 296 2590 330
rect 2624 296 2658 330
rect 2692 296 2726 330
rect 2760 296 2794 330
rect 2828 296 2862 330
rect 2896 296 2930 330
rect 2964 296 2998 330
rect 3032 296 3066 330
rect 3100 296 3134 330
rect 3168 296 3202 330
rect 3236 296 3270 330
rect 3304 296 3338 330
rect 3372 296 3406 330
rect 3440 296 3474 330
rect 3508 296 3542 330
<< poly >>
rect 320 3150 360 3600
rect 210 2940 360 3150
rect 210 2906 259 2940
rect 293 2906 360 2940
rect 210 2872 360 2906
rect 210 2838 259 2872
rect 293 2838 360 2872
rect 210 2804 360 2838
rect 210 2770 259 2804
rect 293 2770 360 2804
rect 210 2736 360 2770
rect 210 2702 259 2736
rect 293 2702 360 2736
rect 210 2668 360 2702
rect 210 2634 259 2668
rect 293 2634 360 2668
rect 210 2600 360 2634
rect 210 2566 259 2600
rect 293 2566 360 2600
rect 210 2532 360 2566
rect 210 2498 259 2532
rect 293 2498 360 2532
rect 210 2464 360 2498
rect 210 2430 259 2464
rect 293 2430 360 2464
rect 210 2396 360 2430
rect 210 2362 259 2396
rect 293 2362 360 2396
rect 210 2328 360 2362
rect 210 2294 259 2328
rect 293 2294 360 2328
rect 210 2260 360 2294
rect 210 2226 259 2260
rect 293 2226 360 2260
rect 210 2192 360 2226
rect 210 2158 259 2192
rect 293 2158 360 2192
rect 210 2124 360 2158
rect 210 2090 259 2124
rect 293 2090 360 2124
rect 210 2056 360 2090
rect 210 2022 259 2056
rect 293 2022 360 2056
rect 210 1988 360 2022
rect 210 1954 259 1988
rect 293 1954 360 1988
rect 210 1920 360 1954
rect 210 1886 259 1920
rect 293 1886 360 1920
rect 210 1852 360 1886
rect 210 1818 259 1852
rect 293 1818 360 1852
rect 210 1784 360 1818
rect 210 1750 259 1784
rect 293 1750 360 1784
rect 210 1716 360 1750
rect 210 1682 259 1716
rect 293 1682 360 1716
rect 210 1648 360 1682
rect 210 1614 259 1648
rect 293 1614 360 1648
rect 210 1580 360 1614
rect 210 1546 259 1580
rect 293 1546 360 1580
rect 210 1512 360 1546
rect 210 1478 259 1512
rect 293 1478 360 1512
rect 210 1444 360 1478
rect 210 1410 259 1444
rect 293 1410 360 1444
rect 210 1376 360 1410
rect 210 1342 259 1376
rect 293 1342 360 1376
rect 210 1308 360 1342
rect 210 1274 259 1308
rect 293 1274 360 1308
rect 210 1240 360 1274
rect 210 1206 259 1240
rect 293 1206 360 1240
rect 210 1172 360 1206
rect 210 1138 259 1172
rect 293 1138 360 1172
rect 210 1104 360 1138
rect 210 1070 259 1104
rect 293 1070 360 1104
rect 210 840 360 1070
rect 320 400 360 840
rect 3640 3150 3680 3600
rect 3640 2940 3790 3150
rect 3640 2906 3706 2940
rect 3740 2906 3790 2940
rect 3640 2872 3790 2906
rect 3640 2838 3706 2872
rect 3740 2838 3790 2872
rect 3640 2804 3790 2838
rect 3640 2770 3706 2804
rect 3740 2770 3790 2804
rect 3640 2736 3790 2770
rect 3640 2702 3706 2736
rect 3740 2702 3790 2736
rect 3640 2668 3790 2702
rect 3640 2634 3706 2668
rect 3740 2634 3790 2668
rect 3640 2600 3790 2634
rect 3640 2566 3706 2600
rect 3740 2566 3790 2600
rect 3640 2532 3790 2566
rect 3640 2498 3706 2532
rect 3740 2498 3790 2532
rect 3640 2464 3790 2498
rect 3640 2430 3706 2464
rect 3740 2430 3790 2464
rect 3640 2396 3790 2430
rect 3640 2362 3706 2396
rect 3740 2362 3790 2396
rect 3640 2328 3790 2362
rect 3640 2294 3706 2328
rect 3740 2294 3790 2328
rect 3640 2260 3790 2294
rect 3640 2226 3706 2260
rect 3740 2226 3790 2260
rect 3640 2192 3790 2226
rect 3640 2158 3706 2192
rect 3740 2158 3790 2192
rect 3640 2124 3790 2158
rect 3640 2090 3706 2124
rect 3740 2090 3790 2124
rect 3640 2056 3790 2090
rect 3640 2022 3706 2056
rect 3740 2022 3790 2056
rect 3640 1988 3790 2022
rect 3640 1954 3706 1988
rect 3740 1954 3790 1988
rect 3640 1920 3790 1954
rect 3640 1886 3706 1920
rect 3740 1886 3790 1920
rect 3640 1852 3790 1886
rect 3640 1818 3706 1852
rect 3740 1818 3790 1852
rect 3640 1784 3790 1818
rect 3640 1750 3706 1784
rect 3740 1750 3790 1784
rect 3640 1716 3790 1750
rect 3640 1682 3706 1716
rect 3740 1682 3790 1716
rect 3640 1648 3790 1682
rect 3640 1614 3706 1648
rect 3740 1614 3790 1648
rect 3640 1580 3790 1614
rect 3640 1546 3706 1580
rect 3740 1546 3790 1580
rect 3640 1512 3790 1546
rect 3640 1478 3706 1512
rect 3740 1478 3790 1512
rect 3640 1444 3790 1478
rect 3640 1410 3706 1444
rect 3740 1410 3790 1444
rect 3640 1376 3790 1410
rect 3640 1342 3706 1376
rect 3740 1342 3790 1376
rect 3640 1308 3790 1342
rect 3640 1274 3706 1308
rect 3740 1274 3790 1308
rect 3640 1240 3790 1274
rect 3640 1206 3706 1240
rect 3740 1206 3790 1240
rect 3640 1172 3790 1206
rect 3640 1138 3706 1172
rect 3740 1138 3790 1172
rect 3640 1104 3790 1138
rect 3640 1070 3706 1104
rect 3740 1070 3790 1104
rect 3640 840 3790 1070
rect 3640 400 3680 840
<< polycont >>
rect 259 2906 293 2940
rect 259 2838 293 2872
rect 259 2770 293 2804
rect 259 2702 293 2736
rect 259 2634 293 2668
rect 259 2566 293 2600
rect 259 2498 293 2532
rect 259 2430 293 2464
rect 259 2362 293 2396
rect 259 2294 293 2328
rect 259 2226 293 2260
rect 259 2158 293 2192
rect 259 2090 293 2124
rect 259 2022 293 2056
rect 259 1954 293 1988
rect 259 1886 293 1920
rect 259 1818 293 1852
rect 259 1750 293 1784
rect 259 1682 293 1716
rect 259 1614 293 1648
rect 259 1546 293 1580
rect 259 1478 293 1512
rect 259 1410 293 1444
rect 259 1342 293 1376
rect 259 1274 293 1308
rect 259 1206 293 1240
rect 259 1138 293 1172
rect 259 1070 293 1104
rect 3706 2906 3740 2940
rect 3706 2838 3740 2872
rect 3706 2770 3740 2804
rect 3706 2702 3740 2736
rect 3706 2634 3740 2668
rect 3706 2566 3740 2600
rect 3706 2498 3740 2532
rect 3706 2430 3740 2464
rect 3706 2362 3740 2396
rect 3706 2294 3740 2328
rect 3706 2226 3740 2260
rect 3706 2158 3740 2192
rect 3706 2090 3740 2124
rect 3706 2022 3740 2056
rect 3706 1954 3740 1988
rect 3706 1886 3740 1920
rect 3706 1818 3740 1852
rect 3706 1750 3740 1784
rect 3706 1682 3740 1716
rect 3706 1614 3740 1648
rect 3706 1546 3740 1580
rect 3706 1478 3740 1512
rect 3706 1410 3740 1444
rect 3706 1342 3740 1376
rect 3706 1274 3740 1308
rect 3706 1206 3740 1240
rect 3706 1138 3740 1172
rect 3706 1070 3740 1104
<< locali >>
rect 890 3920 1350 4000
rect 2650 3920 3110 4000
rect 80 3892 3920 3920
rect 80 3858 933 3892
rect 967 3858 1001 3892
rect 1035 3858 1069 3892
rect 1103 3858 1137 3892
rect 1171 3858 1205 3892
rect 1239 3858 1273 3892
rect 1307 3858 2693 3892
rect 2727 3858 2761 3892
rect 2795 3858 2829 3892
rect 2863 3858 2897 3892
rect 2931 3858 2965 3892
rect 2999 3858 3033 3892
rect 3067 3858 3920 3892
rect 80 3840 3920 3858
rect 80 3110 160 3840
rect 890 3830 1350 3840
rect 2650 3830 3110 3840
rect 360 3703 3640 3720
rect 360 3687 448 3703
rect 482 3687 516 3703
rect 360 3653 427 3687
rect 482 3669 499 3687
rect 550 3669 584 3703
rect 618 3687 652 3703
rect 686 3687 720 3703
rect 754 3687 788 3703
rect 822 3687 856 3703
rect 621 3669 652 3687
rect 693 3669 720 3687
rect 781 3669 788 3687
rect 853 3669 856 3687
rect 890 3687 924 3703
rect 958 3687 992 3703
rect 890 3669 907 3687
rect 958 3669 979 3687
rect 1026 3669 1060 3703
rect 1094 3687 1128 3703
rect 1162 3687 1196 3703
rect 1101 3669 1128 3687
rect 1173 3669 1196 3687
rect 1230 3669 1264 3703
rect 1298 3669 1332 3703
rect 1366 3669 1400 3703
rect 1434 3669 1468 3703
rect 1502 3669 1536 3703
rect 1570 3669 1604 3703
rect 1638 3669 1672 3703
rect 1706 3669 1740 3703
rect 1774 3669 1808 3703
rect 1842 3669 1876 3703
rect 1910 3669 1944 3703
rect 1978 3669 2012 3703
rect 2046 3669 2080 3703
rect 2114 3669 2148 3703
rect 2182 3669 2216 3703
rect 2250 3669 2284 3703
rect 2318 3669 2352 3703
rect 2386 3669 2420 3703
rect 2454 3669 2488 3703
rect 2522 3669 2556 3703
rect 2590 3669 2624 3703
rect 2658 3669 2692 3703
rect 2726 3669 2760 3703
rect 2794 3687 2828 3703
rect 2794 3669 2827 3687
rect 2862 3669 2896 3703
rect 2930 3687 2964 3703
rect 2998 3687 3032 3703
rect 3066 3687 3100 3703
rect 2933 3669 2964 3687
rect 3021 3669 3032 3687
rect 3093 3669 3100 3687
rect 3134 3687 3168 3703
rect 3202 3687 3236 3703
rect 3134 3669 3147 3687
rect 3202 3669 3219 3687
rect 3270 3669 3304 3703
rect 3338 3687 3372 3703
rect 3406 3687 3440 3703
rect 3474 3687 3508 3703
rect 3542 3687 3640 3703
rect 3341 3669 3372 3687
rect 3413 3669 3440 3687
rect 3496 3669 3508 3687
rect 461 3653 499 3669
rect 533 3653 587 3669
rect 621 3653 659 3669
rect 693 3653 747 3669
rect 781 3653 819 3669
rect 853 3653 907 3669
rect 941 3653 979 3669
rect 1013 3653 1067 3669
rect 1101 3653 1139 3669
rect 1173 3653 2827 3669
rect 2861 3653 2899 3669
rect 2933 3653 2987 3669
rect 3021 3653 3059 3669
rect 3093 3653 3147 3669
rect 3181 3653 3219 3669
rect 3253 3653 3307 3669
rect 3341 3653 3379 3669
rect 3413 3653 3462 3669
rect 3496 3653 3534 3669
rect 3568 3653 3640 3687
rect 360 3600 3640 3653
rect 240 3520 1040 3560
rect 240 3400 320 3520
rect 1080 3480 1150 3600
rect 360 3440 1150 3480
rect 240 3360 1040 3400
rect 240 3240 320 3360
rect 1080 3320 1150 3440
rect 360 3280 1150 3320
rect 240 3200 1040 3240
rect 0 3067 170 3110
rect 0 3033 108 3067
rect 142 3033 170 3067
rect 0 2999 170 3033
rect 0 2965 108 2999
rect 142 2965 170 2999
rect 0 2931 170 2965
rect 0 2897 108 2931
rect 142 2897 170 2931
rect 0 2863 170 2897
rect 0 2829 108 2863
rect 142 2829 170 2863
rect 0 2795 170 2829
rect 0 2761 108 2795
rect 142 2761 170 2795
rect 0 2727 170 2761
rect 0 2693 108 2727
rect 142 2693 170 2727
rect 0 2650 170 2693
rect 240 3080 320 3200
rect 1080 3160 1150 3280
rect 360 3120 1150 3160
rect 240 3040 1040 3080
rect 240 2940 320 3040
rect 1080 3000 1150 3120
rect 360 2960 1150 3000
rect 240 2906 259 2940
rect 293 2922 320 2940
rect 297 2920 320 2922
rect 240 2888 263 2906
rect 297 2888 1040 2920
rect 240 2880 1040 2888
rect 240 2872 320 2880
rect 240 2838 259 2872
rect 293 2850 320 2872
rect 240 2816 263 2838
rect 297 2816 320 2850
rect 1080 2840 1150 2960
rect 240 2804 320 2816
rect 240 2770 259 2804
rect 293 2778 320 2804
rect 360 2800 1150 2840
rect 240 2744 263 2770
rect 297 2760 320 2778
rect 297 2744 1040 2760
rect 240 2736 1040 2744
rect 240 2702 259 2736
rect 293 2720 1040 2736
rect 293 2706 320 2720
rect 240 2672 263 2702
rect 297 2672 320 2706
rect 1080 2680 1150 2800
rect 240 2668 320 2672
rect 80 1350 160 2650
rect 240 2634 259 2668
rect 293 2634 320 2668
rect 360 2640 1150 2680
rect 240 2600 263 2634
rect 297 2600 320 2634
rect 240 2566 259 2600
rect 293 2566 1040 2600
rect 240 2562 1040 2566
rect 240 2532 263 2562
rect 297 2560 1040 2562
rect 240 2498 259 2532
rect 297 2528 320 2560
rect 293 2498 320 2528
rect 1080 2520 1150 2640
rect 240 2490 320 2498
rect 240 2464 263 2490
rect 240 2430 259 2464
rect 297 2456 320 2490
rect 360 2480 1150 2520
rect 293 2440 320 2456
rect 293 2430 1040 2440
rect 240 2418 1040 2430
rect 240 2396 263 2418
rect 297 2400 1040 2418
rect 240 2362 259 2396
rect 297 2384 320 2400
rect 293 2362 320 2384
rect 240 2346 320 2362
rect 1080 2360 1150 2480
rect 240 2328 263 2346
rect 240 2294 259 2328
rect 297 2312 320 2346
rect 360 2320 1150 2360
rect 293 2294 320 2312
rect 240 2280 320 2294
rect 240 2274 1040 2280
rect 240 2260 263 2274
rect 240 2226 259 2260
rect 297 2240 1040 2274
rect 293 2226 320 2240
rect 240 2202 320 2226
rect 240 2192 263 2202
rect 240 2158 259 2192
rect 297 2168 320 2202
rect 1080 2200 1150 2320
rect 293 2158 320 2168
rect 360 2160 1150 2200
rect 240 2130 320 2158
rect 240 2124 263 2130
rect 240 2090 259 2124
rect 297 2120 320 2130
rect 297 2096 1040 2120
rect 293 2090 1040 2096
rect 240 2080 1040 2090
rect 1080 2080 1150 2160
rect 240 2058 320 2080
rect 240 2056 263 2058
rect 240 2022 259 2056
rect 297 2040 320 2058
rect 1190 2040 1230 3560
rect 1270 2080 1310 3600
rect 1350 2040 1390 3560
rect 1430 2080 1470 3600
rect 1510 2040 1550 3560
rect 1590 2080 1630 3600
rect 1670 2040 1710 3560
rect 1750 2080 1790 3600
rect 1830 2040 1870 3560
rect 297 2024 1870 2040
rect 293 2022 1870 2024
rect 240 1988 1870 2022
rect 240 1954 259 1988
rect 293 1986 1870 1988
rect 297 1960 1870 1986
rect 240 1952 263 1954
rect 297 1952 320 1960
rect 240 1920 320 1952
rect 240 1886 259 1920
rect 293 1914 1040 1920
rect 240 1880 263 1886
rect 297 1880 1040 1914
rect 240 1852 320 1880
rect 240 1818 259 1852
rect 293 1842 320 1852
rect 240 1808 263 1818
rect 297 1808 320 1842
rect 1080 1840 1150 1920
rect 240 1784 320 1808
rect 360 1800 1150 1840
rect 240 1750 259 1784
rect 293 1770 320 1784
rect 297 1760 320 1770
rect 240 1736 263 1750
rect 297 1736 1040 1760
rect 240 1720 1040 1736
rect 240 1716 320 1720
rect 240 1682 259 1716
rect 293 1698 320 1716
rect 240 1664 263 1682
rect 297 1664 320 1698
rect 1080 1680 1150 1800
rect 240 1648 320 1664
rect 240 1614 259 1648
rect 293 1626 320 1648
rect 360 1640 1150 1680
rect 240 1592 263 1614
rect 297 1600 320 1626
rect 297 1592 1040 1600
rect 240 1580 1040 1592
rect 240 1546 259 1580
rect 293 1560 1040 1580
rect 293 1554 320 1560
rect 240 1520 263 1546
rect 297 1520 320 1554
rect 1080 1520 1150 1640
rect 240 1512 320 1520
rect 240 1478 259 1512
rect 293 1482 320 1512
rect 240 1448 263 1478
rect 297 1448 320 1482
rect 360 1480 1150 1520
rect 240 1444 320 1448
rect 240 1410 259 1444
rect 293 1440 320 1444
rect 293 1410 1040 1440
rect 240 1376 263 1410
rect 297 1400 1040 1410
rect 297 1376 320 1400
rect 0 1307 170 1350
rect 0 1273 108 1307
rect 142 1273 170 1307
rect 0 1239 170 1273
rect 0 1205 108 1239
rect 142 1205 170 1239
rect 0 1171 170 1205
rect 0 1137 108 1171
rect 142 1137 170 1171
rect 0 1103 170 1137
rect 0 1069 108 1103
rect 142 1069 170 1103
rect 0 1035 170 1069
rect 0 1001 108 1035
rect 142 1001 170 1035
rect 0 967 170 1001
rect 0 933 108 967
rect 142 933 170 967
rect 0 890 170 933
rect 240 1342 259 1376
rect 293 1342 320 1376
rect 1080 1360 1150 1480
rect 240 1338 320 1342
rect 240 1308 263 1338
rect 240 1274 259 1308
rect 297 1304 320 1338
rect 360 1320 1150 1360
rect 293 1280 320 1304
rect 293 1274 1040 1280
rect 240 1266 1040 1274
rect 240 1240 263 1266
rect 297 1240 1040 1266
rect 240 1206 259 1240
rect 297 1232 320 1240
rect 293 1206 320 1232
rect 240 1194 320 1206
rect 1080 1200 1150 1320
rect 240 1172 263 1194
rect 240 1138 259 1172
rect 297 1160 320 1194
rect 360 1160 1150 1200
rect 293 1138 320 1160
rect 240 1122 320 1138
rect 240 1104 263 1122
rect 297 1120 320 1122
rect 240 1070 259 1104
rect 297 1088 1040 1120
rect 293 1080 1040 1088
rect 293 1070 320 1080
rect 240 960 320 1070
rect 1080 1040 1150 1160
rect 360 1000 1150 1040
rect 240 920 1040 960
rect 80 160 160 890
rect 240 800 320 920
rect 1080 880 1150 1000
rect 360 840 1150 880
rect 240 760 1040 800
rect 240 640 320 760
rect 1080 720 1150 840
rect 360 680 1150 720
rect 240 600 1040 640
rect 240 480 320 600
rect 1080 560 1150 680
rect 360 520 1150 560
rect 240 440 1040 480
rect 1080 400 1150 520
rect 1190 440 1230 1960
rect 1270 400 1310 1920
rect 1350 440 1390 1960
rect 1430 400 1470 1920
rect 1510 440 1550 1960
rect 1590 400 1630 1920
rect 1670 440 1710 1960
rect 1750 400 1790 1920
rect 1830 440 1870 1960
rect 1910 400 2090 3600
rect 2130 2040 2170 3560
rect 2210 2080 2250 3600
rect 2290 2040 2330 3560
rect 2370 2080 2410 3600
rect 2450 2040 2490 3560
rect 2530 2080 2570 3600
rect 2610 2040 2650 3560
rect 2690 2080 2730 3600
rect 2770 2040 2810 3560
rect 2850 3480 2920 3600
rect 2960 3520 3760 3560
rect 2850 3440 3640 3480
rect 2850 3320 2920 3440
rect 3680 3400 3760 3520
rect 2960 3360 3760 3400
rect 2850 3280 3640 3320
rect 2850 3160 2920 3280
rect 3680 3240 3760 3360
rect 2960 3200 3760 3240
rect 2850 3120 3640 3160
rect 2850 3000 2920 3120
rect 3680 3080 3760 3200
rect 3840 3110 3920 3840
rect 2960 3040 3760 3080
rect 2850 2960 3640 3000
rect 2850 2840 2920 2960
rect 3680 2940 3760 3040
rect 3680 2922 3706 2940
rect 3680 2920 3703 2922
rect 2960 2888 3703 2920
rect 3740 2906 3760 2940
rect 3737 2888 3760 2906
rect 2960 2880 3760 2888
rect 3680 2872 3760 2880
rect 3680 2850 3706 2872
rect 2850 2800 3640 2840
rect 3680 2816 3703 2850
rect 3740 2838 3760 2872
rect 3737 2816 3760 2838
rect 3680 2804 3760 2816
rect 2850 2680 2920 2800
rect 3680 2778 3706 2804
rect 3680 2760 3703 2778
rect 3740 2770 3760 2804
rect 2960 2744 3703 2760
rect 3737 2744 3760 2770
rect 2960 2736 3760 2744
rect 2960 2720 3706 2736
rect 3680 2706 3706 2720
rect 2850 2640 3640 2680
rect 3680 2672 3703 2706
rect 3740 2702 3760 2736
rect 3737 2672 3760 2702
rect 3680 2668 3760 2672
rect 2850 2520 2920 2640
rect 3680 2634 3706 2668
rect 3740 2634 3760 2668
rect 3830 3067 4000 3110
rect 3830 3033 3858 3067
rect 3892 3033 4000 3067
rect 3830 2999 4000 3033
rect 3830 2965 3858 2999
rect 3892 2965 4000 2999
rect 3830 2931 4000 2965
rect 3830 2897 3858 2931
rect 3892 2897 4000 2931
rect 3830 2863 4000 2897
rect 3830 2829 3858 2863
rect 3892 2829 4000 2863
rect 3830 2795 4000 2829
rect 3830 2761 3858 2795
rect 3892 2761 4000 2795
rect 3830 2727 4000 2761
rect 3830 2693 3858 2727
rect 3892 2693 4000 2727
rect 3830 2650 4000 2693
rect 3680 2600 3703 2634
rect 3737 2600 3760 2634
rect 2960 2566 3706 2600
rect 3740 2566 3760 2600
rect 2960 2562 3760 2566
rect 2960 2560 3703 2562
rect 3680 2528 3703 2560
rect 3737 2532 3760 2562
rect 2850 2480 3640 2520
rect 3680 2498 3706 2528
rect 3740 2498 3760 2532
rect 3680 2490 3760 2498
rect 2850 2360 2920 2480
rect 3680 2456 3703 2490
rect 3737 2464 3760 2490
rect 3680 2440 3706 2456
rect 2960 2430 3706 2440
rect 3740 2430 3760 2464
rect 2960 2418 3760 2430
rect 2960 2400 3703 2418
rect 3680 2384 3703 2400
rect 3737 2396 3760 2418
rect 3680 2362 3706 2384
rect 3740 2362 3760 2396
rect 2850 2320 3640 2360
rect 3680 2346 3760 2362
rect 2850 2200 2920 2320
rect 3680 2312 3703 2346
rect 3737 2328 3760 2346
rect 3680 2294 3706 2312
rect 3740 2294 3760 2328
rect 3680 2280 3760 2294
rect 2960 2274 3760 2280
rect 2960 2240 3703 2274
rect 3737 2260 3760 2274
rect 3680 2226 3706 2240
rect 3740 2226 3760 2260
rect 3680 2202 3760 2226
rect 2850 2160 3640 2200
rect 3680 2168 3703 2202
rect 3737 2192 3760 2202
rect 2850 2080 2920 2160
rect 3680 2158 3706 2168
rect 3740 2158 3760 2192
rect 3680 2130 3760 2158
rect 3680 2120 3703 2130
rect 3737 2124 3760 2130
rect 2960 2096 3703 2120
rect 2960 2090 3706 2096
rect 3740 2090 3760 2124
rect 2960 2080 3760 2090
rect 3680 2058 3760 2080
rect 3680 2040 3703 2058
rect 3737 2056 3760 2058
rect 2130 2024 3703 2040
rect 2130 2022 3706 2024
rect 3740 2022 3760 2056
rect 2130 1988 3760 2022
rect 2130 1986 3706 1988
rect 2130 1960 3703 1986
rect 2130 440 2170 1960
rect 2210 400 2250 1920
rect 2290 440 2330 1960
rect 2370 400 2410 1920
rect 2450 440 2490 1960
rect 2530 400 2570 1920
rect 2610 440 2650 1960
rect 2690 400 2730 1920
rect 2770 440 2810 1960
rect 3680 1952 3703 1960
rect 3740 1954 3760 1988
rect 3737 1952 3760 1954
rect 3680 1920 3760 1952
rect 2850 1840 2920 1920
rect 2960 1914 3706 1920
rect 2960 1880 3703 1914
rect 3740 1886 3760 1920
rect 3737 1880 3760 1886
rect 3680 1852 3760 1880
rect 3680 1842 3706 1852
rect 2850 1800 3640 1840
rect 3680 1808 3703 1842
rect 3740 1818 3760 1852
rect 3737 1808 3760 1818
rect 2850 1680 2920 1800
rect 3680 1784 3760 1808
rect 3680 1770 3706 1784
rect 3680 1760 3703 1770
rect 2960 1736 3703 1760
rect 3740 1750 3760 1784
rect 3737 1736 3760 1750
rect 2960 1720 3760 1736
rect 3680 1716 3760 1720
rect 3680 1698 3706 1716
rect 2850 1640 3640 1680
rect 3680 1664 3703 1698
rect 3740 1682 3760 1716
rect 3737 1664 3760 1682
rect 3680 1648 3760 1664
rect 2850 1520 2920 1640
rect 3680 1626 3706 1648
rect 3680 1600 3703 1626
rect 3740 1614 3760 1648
rect 2960 1592 3703 1600
rect 3737 1592 3760 1614
rect 2960 1580 3760 1592
rect 2960 1560 3706 1580
rect 3680 1554 3706 1560
rect 3680 1520 3703 1554
rect 3740 1546 3760 1580
rect 3737 1520 3760 1546
rect 2850 1480 3640 1520
rect 3680 1512 3760 1520
rect 3680 1482 3706 1512
rect 2850 1360 2920 1480
rect 3680 1448 3703 1482
rect 3740 1478 3760 1512
rect 3737 1448 3760 1478
rect 3680 1444 3760 1448
rect 3680 1440 3706 1444
rect 2960 1410 3706 1440
rect 3740 1410 3760 1444
rect 2960 1400 3703 1410
rect 3680 1376 3703 1400
rect 3737 1376 3760 1410
rect 2850 1320 3640 1360
rect 3680 1342 3706 1376
rect 3740 1342 3760 1376
rect 3840 1350 3920 2650
rect 3680 1338 3760 1342
rect 2850 1200 2920 1320
rect 3680 1304 3703 1338
rect 3737 1308 3760 1338
rect 3680 1280 3706 1304
rect 2960 1274 3706 1280
rect 3740 1274 3760 1308
rect 2960 1266 3760 1274
rect 2960 1240 3703 1266
rect 3737 1240 3760 1266
rect 3680 1232 3703 1240
rect 3680 1206 3706 1232
rect 3740 1206 3760 1240
rect 2850 1160 3640 1200
rect 3680 1194 3760 1206
rect 3680 1160 3703 1194
rect 3737 1172 3760 1194
rect 2850 1040 2920 1160
rect 3680 1138 3706 1160
rect 3740 1138 3760 1172
rect 3680 1122 3760 1138
rect 3680 1120 3703 1122
rect 2960 1088 3703 1120
rect 3737 1104 3760 1122
rect 2960 1080 3706 1088
rect 3680 1070 3706 1080
rect 3740 1070 3760 1104
rect 2850 1000 3640 1040
rect 2850 880 2920 1000
rect 3680 960 3760 1070
rect 2960 920 3760 960
rect 2850 840 3640 880
rect 2850 720 2920 840
rect 3680 800 3760 920
rect 3830 1307 4000 1350
rect 3830 1273 3858 1307
rect 3892 1273 4000 1307
rect 3830 1239 4000 1273
rect 3830 1205 3858 1239
rect 3892 1205 4000 1239
rect 3830 1171 4000 1205
rect 3830 1137 3858 1171
rect 3892 1137 4000 1171
rect 3830 1103 4000 1137
rect 3830 1069 3858 1103
rect 3892 1069 4000 1103
rect 3830 1035 4000 1069
rect 3830 1001 3858 1035
rect 3892 1001 4000 1035
rect 3830 967 4000 1001
rect 3830 933 3858 967
rect 3892 933 4000 967
rect 3830 890 4000 933
rect 2960 760 3760 800
rect 2850 680 3640 720
rect 2850 560 2920 680
rect 3680 640 3760 760
rect 2960 600 3760 640
rect 2850 520 3640 560
rect 2850 400 2920 520
rect 3680 480 3760 600
rect 2960 440 3760 480
rect 360 347 3640 400
rect 360 313 427 347
rect 461 330 499 347
rect 533 330 587 347
rect 621 330 659 347
rect 693 330 747 347
rect 781 330 819 347
rect 853 330 907 347
rect 941 330 979 347
rect 1013 330 1067 347
rect 1101 330 1139 347
rect 1173 330 2827 347
rect 2861 330 2899 347
rect 2933 330 2987 347
rect 3021 330 3059 347
rect 3093 330 3147 347
rect 3181 330 3219 347
rect 3253 330 3307 347
rect 3341 330 3379 347
rect 3413 330 3462 347
rect 3496 330 3534 347
rect 482 313 499 330
rect 360 296 448 313
rect 482 296 516 313
rect 550 296 584 330
rect 621 313 652 330
rect 693 313 720 330
rect 781 313 788 330
rect 853 313 856 330
rect 618 296 652 313
rect 686 296 720 313
rect 754 296 788 313
rect 822 296 856 313
rect 890 313 907 330
rect 958 313 979 330
rect 890 296 924 313
rect 958 296 992 313
rect 1026 296 1060 330
rect 1101 313 1128 330
rect 1173 313 1196 330
rect 1094 296 1128 313
rect 1162 296 1196 313
rect 1230 296 1264 330
rect 1298 296 1332 330
rect 1366 296 1400 330
rect 1434 296 1468 330
rect 1502 296 1536 330
rect 1570 296 1604 330
rect 1638 296 1672 330
rect 1706 296 1740 330
rect 1774 296 1808 330
rect 1842 296 1876 330
rect 1910 296 1944 330
rect 1978 296 2012 330
rect 2046 296 2080 330
rect 2114 296 2148 330
rect 2182 296 2216 330
rect 2250 296 2284 330
rect 2318 296 2352 330
rect 2386 296 2420 330
rect 2454 296 2488 330
rect 2522 296 2556 330
rect 2590 296 2624 330
rect 2658 296 2692 330
rect 2726 296 2760 330
rect 2794 313 2827 330
rect 2794 296 2828 313
rect 2862 296 2896 330
rect 2933 313 2964 330
rect 3021 313 3032 330
rect 3093 313 3100 330
rect 2930 296 2964 313
rect 2998 296 3032 313
rect 3066 296 3100 313
rect 3134 313 3147 330
rect 3202 313 3219 330
rect 3134 296 3168 313
rect 3202 296 3236 313
rect 3270 296 3304 330
rect 3341 313 3372 330
rect 3413 313 3440 330
rect 3496 313 3508 330
rect 3568 313 3640 347
rect 3338 296 3372 313
rect 3406 296 3440 313
rect 3474 296 3508 313
rect 3542 296 3640 313
rect 360 280 3640 296
rect 890 160 1350 170
rect 2650 160 3110 170
rect 3840 160 3920 890
rect 80 142 3920 160
rect 80 108 933 142
rect 967 108 1001 142
rect 1035 108 1069 142
rect 1103 108 1137 142
rect 1171 108 1205 142
rect 1239 108 1273 142
rect 1307 108 2693 142
rect 2727 108 2761 142
rect 2795 108 2829 142
rect 2863 108 2897 142
rect 2931 108 2965 142
rect 2999 108 3033 142
rect 3067 108 3920 142
rect 80 80 3920 108
rect 890 0 1350 80
rect 2650 0 3110 80
<< viali >>
rect 427 3669 448 3687
rect 448 3669 461 3687
rect 499 3669 516 3687
rect 516 3669 533 3687
rect 587 3669 618 3687
rect 618 3669 621 3687
rect 659 3669 686 3687
rect 686 3669 693 3687
rect 747 3669 754 3687
rect 754 3669 781 3687
rect 819 3669 822 3687
rect 822 3669 853 3687
rect 907 3669 924 3687
rect 924 3669 941 3687
rect 979 3669 992 3687
rect 992 3669 1013 3687
rect 1067 3669 1094 3687
rect 1094 3669 1101 3687
rect 1139 3669 1162 3687
rect 1162 3669 1173 3687
rect 2827 3669 2828 3687
rect 2828 3669 2861 3687
rect 2899 3669 2930 3687
rect 2930 3669 2933 3687
rect 2987 3669 2998 3687
rect 2998 3669 3021 3687
rect 3059 3669 3066 3687
rect 3066 3669 3093 3687
rect 3147 3669 3168 3687
rect 3168 3669 3181 3687
rect 3219 3669 3236 3687
rect 3236 3669 3253 3687
rect 3307 3669 3338 3687
rect 3338 3669 3341 3687
rect 3379 3669 3406 3687
rect 3406 3669 3413 3687
rect 3462 3669 3474 3687
rect 3474 3669 3496 3687
rect 3534 3669 3542 3687
rect 3542 3669 3568 3687
rect 427 3653 461 3669
rect 499 3653 533 3669
rect 587 3653 621 3669
rect 659 3653 693 3669
rect 747 3653 781 3669
rect 819 3653 853 3669
rect 907 3653 941 3669
rect 979 3653 1013 3669
rect 1067 3653 1101 3669
rect 1139 3653 1173 3669
rect 2827 3653 2861 3669
rect 2899 3653 2933 3669
rect 2987 3653 3021 3669
rect 3059 3653 3093 3669
rect 3147 3653 3181 3669
rect 3219 3653 3253 3669
rect 3307 3653 3341 3669
rect 3379 3653 3413 3669
rect 3462 3653 3496 3669
rect 3534 3653 3568 3669
rect 263 2906 293 2922
rect 293 2906 297 2922
rect 263 2888 297 2906
rect 263 2838 293 2850
rect 293 2838 297 2850
rect 263 2816 297 2838
rect 263 2770 293 2778
rect 293 2770 297 2778
rect 263 2744 297 2770
rect 263 2702 293 2706
rect 293 2702 297 2706
rect 263 2672 297 2702
rect 263 2600 297 2634
rect 263 2532 297 2562
rect 263 2528 293 2532
rect 293 2528 297 2532
rect 263 2464 297 2490
rect 263 2456 293 2464
rect 293 2456 297 2464
rect 263 2396 297 2418
rect 263 2384 293 2396
rect 293 2384 297 2396
rect 263 2328 297 2346
rect 263 2312 293 2328
rect 293 2312 297 2328
rect 263 2260 297 2274
rect 263 2240 293 2260
rect 293 2240 297 2260
rect 263 2192 297 2202
rect 263 2168 293 2192
rect 293 2168 297 2192
rect 263 2124 297 2130
rect 263 2096 293 2124
rect 293 2096 297 2124
rect 263 2056 297 2058
rect 263 2024 293 2056
rect 293 2024 297 2056
rect 263 1954 293 1986
rect 293 1954 297 1986
rect 263 1952 297 1954
rect 263 1886 293 1914
rect 293 1886 297 1914
rect 263 1880 297 1886
rect 263 1818 293 1842
rect 293 1818 297 1842
rect 263 1808 297 1818
rect 263 1750 293 1770
rect 293 1750 297 1770
rect 263 1736 297 1750
rect 263 1682 293 1698
rect 293 1682 297 1698
rect 263 1664 297 1682
rect 263 1614 293 1626
rect 293 1614 297 1626
rect 263 1592 297 1614
rect 263 1546 293 1554
rect 293 1546 297 1554
rect 263 1520 297 1546
rect 263 1478 293 1482
rect 293 1478 297 1482
rect 263 1448 297 1478
rect 263 1376 297 1410
rect 263 1308 297 1338
rect 263 1304 293 1308
rect 293 1304 297 1308
rect 263 1240 297 1266
rect 263 1232 293 1240
rect 293 1232 297 1240
rect 263 1172 297 1194
rect 263 1160 293 1172
rect 293 1160 297 1172
rect 263 1104 297 1122
rect 263 1088 293 1104
rect 293 1088 297 1104
rect 3703 2906 3706 2922
rect 3706 2906 3737 2922
rect 3703 2888 3737 2906
rect 3703 2838 3706 2850
rect 3706 2838 3737 2850
rect 3703 2816 3737 2838
rect 3703 2770 3706 2778
rect 3706 2770 3737 2778
rect 3703 2744 3737 2770
rect 3703 2702 3706 2706
rect 3706 2702 3737 2706
rect 3703 2672 3737 2702
rect 3703 2600 3737 2634
rect 3703 2532 3737 2562
rect 3703 2528 3706 2532
rect 3706 2528 3737 2532
rect 3703 2464 3737 2490
rect 3703 2456 3706 2464
rect 3706 2456 3737 2464
rect 3703 2396 3737 2418
rect 3703 2384 3706 2396
rect 3706 2384 3737 2396
rect 3703 2328 3737 2346
rect 3703 2312 3706 2328
rect 3706 2312 3737 2328
rect 3703 2260 3737 2274
rect 3703 2240 3706 2260
rect 3706 2240 3737 2260
rect 3703 2192 3737 2202
rect 3703 2168 3706 2192
rect 3706 2168 3737 2192
rect 3703 2124 3737 2130
rect 3703 2096 3706 2124
rect 3706 2096 3737 2124
rect 3703 2056 3737 2058
rect 3703 2024 3706 2056
rect 3706 2024 3737 2056
rect 3703 1954 3706 1986
rect 3706 1954 3737 1986
rect 3703 1952 3737 1954
rect 3703 1886 3706 1914
rect 3706 1886 3737 1914
rect 3703 1880 3737 1886
rect 3703 1818 3706 1842
rect 3706 1818 3737 1842
rect 3703 1808 3737 1818
rect 3703 1750 3706 1770
rect 3706 1750 3737 1770
rect 3703 1736 3737 1750
rect 3703 1682 3706 1698
rect 3706 1682 3737 1698
rect 3703 1664 3737 1682
rect 3703 1614 3706 1626
rect 3706 1614 3737 1626
rect 3703 1592 3737 1614
rect 3703 1546 3706 1554
rect 3706 1546 3737 1554
rect 3703 1520 3737 1546
rect 3703 1478 3706 1482
rect 3706 1478 3737 1482
rect 3703 1448 3737 1478
rect 3703 1376 3737 1410
rect 3703 1308 3737 1338
rect 3703 1304 3706 1308
rect 3706 1304 3737 1308
rect 3703 1240 3737 1266
rect 3703 1232 3706 1240
rect 3706 1232 3737 1240
rect 3703 1172 3737 1194
rect 3703 1160 3706 1172
rect 3706 1160 3737 1172
rect 3703 1104 3737 1122
rect 3703 1088 3706 1104
rect 3706 1088 3737 1104
rect 427 330 461 347
rect 499 330 533 347
rect 587 330 621 347
rect 659 330 693 347
rect 747 330 781 347
rect 819 330 853 347
rect 907 330 941 347
rect 979 330 1013 347
rect 1067 330 1101 347
rect 1139 330 1173 347
rect 2827 330 2861 347
rect 2899 330 2933 347
rect 2987 330 3021 347
rect 3059 330 3093 347
rect 3147 330 3181 347
rect 3219 330 3253 347
rect 3307 330 3341 347
rect 3379 330 3413 347
rect 3462 330 3496 347
rect 3534 330 3568 347
rect 427 313 448 330
rect 448 313 461 330
rect 499 313 516 330
rect 516 313 533 330
rect 587 313 618 330
rect 618 313 621 330
rect 659 313 686 330
rect 686 313 693 330
rect 747 313 754 330
rect 754 313 781 330
rect 819 313 822 330
rect 822 313 853 330
rect 907 313 924 330
rect 924 313 941 330
rect 979 313 992 330
rect 992 313 1013 330
rect 1067 313 1094 330
rect 1094 313 1101 330
rect 1139 313 1162 330
rect 1162 313 1173 330
rect 2827 313 2828 330
rect 2828 313 2861 330
rect 2899 313 2930 330
rect 2930 313 2933 330
rect 2987 313 2998 330
rect 2998 313 3021 330
rect 3059 313 3066 330
rect 3066 313 3093 330
rect 3147 313 3168 330
rect 3168 313 3181 330
rect 3219 313 3236 330
rect 3236 313 3253 330
rect 3307 313 3338 330
rect 3338 313 3341 330
rect 3379 313 3406 330
rect 3406 313 3413 330
rect 3462 313 3474 330
rect 3474 313 3496 330
rect 3534 313 3542 330
rect 3542 313 3568 330
<< metal1 >>
rect 0 3970 880 4000
rect 1360 3970 2640 4000
rect 0 3790 30 3970
rect 210 3790 350 3970
rect 530 3790 670 3970
rect 850 3790 1200 3970
rect 0 3760 880 3790
rect 0 3650 240 3760
rect 910 3730 1200 3790
rect 1360 3790 1390 3970
rect 1570 3790 1620 3970
rect 1800 3790 1846 3970
rect 2154 3790 2200 3970
rect 2380 3790 2430 3970
rect 2610 3790 2640 3970
rect 3120 3970 4000 4000
rect 3120 3960 3150 3970
rect 1360 3760 2640 3790
rect 2800 3790 3150 3960
rect 3330 3790 3470 3970
rect 3650 3790 3790 3970
rect 3970 3790 4000 3970
rect 2800 3780 4000 3790
rect 0 3470 30 3650
rect 210 3470 240 3650
rect 0 3330 240 3470
rect 0 3150 30 3330
rect 210 3150 240 3330
rect 0 3120 240 3150
rect 360 3690 1200 3730
rect 360 3687 1870 3690
rect 360 3653 427 3687
rect 461 3653 499 3687
rect 533 3653 587 3687
rect 621 3653 659 3687
rect 693 3653 747 3687
rect 781 3653 819 3687
rect 853 3653 907 3687
rect 941 3653 979 3687
rect 1013 3653 1067 3687
rect 1101 3653 1139 3687
rect 1173 3660 1870 3687
rect 1173 3653 1200 3660
rect 360 3600 1200 3653
rect 1900 3630 2100 3760
rect 2800 3730 3090 3780
rect 3120 3760 4000 3780
rect 2800 3690 3640 3730
rect 2140 3687 3640 3690
rect 2140 3660 2827 3687
rect 2800 3653 2827 3660
rect 2861 3653 2899 3687
rect 2933 3653 2987 3687
rect 3021 3653 3059 3687
rect 3093 3653 3147 3687
rect 3181 3653 3219 3687
rect 3253 3653 3307 3687
rect 3341 3653 3379 3687
rect 3413 3653 3462 3687
rect 3496 3653 3534 3687
rect 3568 3653 3640 3687
rect 1230 3600 2770 3630
rect 2800 3600 3640 3653
rect 360 3030 390 3600
rect 240 2922 390 3000
rect 240 2888 263 2922
rect 297 2888 390 2922
rect 240 2850 390 2888
rect 240 2816 263 2850
rect 297 2816 390 2850
rect 240 2778 390 2816
rect 240 2744 263 2778
rect 297 2744 390 2778
rect 240 2706 390 2744
rect 240 2672 263 2706
rect 297 2672 390 2706
rect 240 2640 390 2672
rect 0 2634 390 2640
rect 0 2608 263 2634
rect 0 2492 32 2608
rect 148 2600 263 2608
rect 297 2600 390 2634
rect 148 2562 390 2600
rect 148 2528 263 2562
rect 297 2528 390 2562
rect 148 2492 390 2528
rect 0 2490 390 2492
rect 0 2456 263 2490
rect 297 2456 390 2490
rect 0 2438 390 2456
rect 0 2322 32 2438
rect 148 2418 390 2438
rect 148 2384 263 2418
rect 297 2384 390 2418
rect 148 2346 390 2384
rect 148 2322 263 2346
rect 0 2312 263 2322
rect 297 2312 390 2346
rect 0 2274 390 2312
rect 0 2268 263 2274
rect 0 2152 32 2268
rect 148 2240 263 2268
rect 297 2240 390 2274
rect 148 2202 390 2240
rect 148 2168 263 2202
rect 297 2168 390 2202
rect 148 2152 390 2168
rect 0 2130 390 2152
rect 0 2096 263 2130
rect 297 2096 390 2130
rect 0 2090 390 2096
rect 0 1910 30 2090
rect 160 2060 390 2090
rect 420 2060 450 3570
rect 480 2090 510 3600
rect 540 2060 570 3570
rect 600 2090 630 3600
rect 660 2060 690 3570
rect 720 2090 750 3600
rect 780 2060 810 3570
rect 840 2090 870 3600
rect 900 2060 930 3570
rect 960 2090 990 3600
rect 1080 3570 1200 3600
rect 1020 2060 1050 3570
rect 1080 3540 1870 3570
rect 1080 3450 1200 3540
rect 1900 3510 2100 3600
rect 2800 3570 2920 3600
rect 2130 3540 2920 3570
rect 1230 3480 2770 3510
rect 1080 3420 1870 3450
rect 1080 3330 1200 3420
rect 1900 3390 2100 3480
rect 2800 3450 2920 3540
rect 2130 3420 2920 3450
rect 1230 3360 2770 3390
rect 1080 3300 1870 3330
rect 1080 3210 1200 3300
rect 1900 3270 2100 3360
rect 2800 3330 2920 3420
rect 2130 3300 2920 3330
rect 1230 3240 2770 3270
rect 1080 3180 1870 3210
rect 1080 3090 1200 3180
rect 1900 3150 2100 3240
rect 2800 3210 2920 3300
rect 2130 3180 2920 3210
rect 1230 3120 2770 3150
rect 1080 3060 1870 3090
rect 1080 2970 1200 3060
rect 1900 3030 2100 3120
rect 2800 3090 2920 3180
rect 2130 3060 2920 3090
rect 1230 3000 2770 3030
rect 1080 2940 1870 2970
rect 1080 2850 1200 2940
rect 1900 2910 2100 3000
rect 2800 2970 2920 3060
rect 2130 2940 2920 2970
rect 1230 2880 2770 2910
rect 1080 2820 1870 2850
rect 1080 2730 1200 2820
rect 1900 2790 2100 2880
rect 2800 2850 2920 2940
rect 2130 2820 2920 2850
rect 1230 2760 2770 2790
rect 1080 2700 1870 2730
rect 1080 2610 1200 2700
rect 1900 2670 2100 2760
rect 2800 2730 2920 2820
rect 2130 2700 2920 2730
rect 1230 2640 2770 2670
rect 1080 2580 1870 2610
rect 1080 2490 1200 2580
rect 1900 2550 2100 2640
rect 2800 2610 2920 2700
rect 2130 2580 2920 2610
rect 1230 2520 2770 2550
rect 1080 2460 1870 2490
rect 1080 2370 1200 2460
rect 1900 2430 2100 2520
rect 2800 2490 2920 2580
rect 2130 2460 2920 2490
rect 1230 2400 2770 2430
rect 1080 2340 1870 2370
rect 1080 2250 1200 2340
rect 1900 2310 2100 2400
rect 2800 2370 2920 2460
rect 2130 2340 2920 2370
rect 1230 2280 2770 2310
rect 1080 2220 1870 2250
rect 1080 2130 1200 2220
rect 1900 2190 2100 2280
rect 2800 2250 2920 2340
rect 2130 2220 2920 2250
rect 1230 2160 2770 2190
rect 1080 2090 1870 2130
rect 1900 2060 2100 2160
rect 2800 2130 2920 2220
rect 2130 2090 2920 2130
rect 2950 2060 2980 3570
rect 3010 2090 3040 3600
rect 3070 2060 3100 3570
rect 3130 2090 3160 3600
rect 3190 2060 3220 3570
rect 3250 2090 3280 3600
rect 3310 2060 3340 3570
rect 3370 2090 3400 3600
rect 3430 2060 3460 3570
rect 3490 2090 3520 3600
rect 3550 2060 3580 3570
rect 3610 3030 3640 3600
rect 3760 3650 4000 3760
rect 3760 3470 3790 3650
rect 3970 3470 4000 3650
rect 3760 3330 4000 3470
rect 3760 3150 3790 3330
rect 3970 3150 4000 3330
rect 3760 3120 4000 3150
rect 3610 2922 3760 3000
rect 3610 2888 3703 2922
rect 3737 2888 3760 2922
rect 3610 2850 3760 2888
rect 3610 2816 3703 2850
rect 3737 2816 3760 2850
rect 3610 2778 3760 2816
rect 3610 2744 3703 2778
rect 3737 2744 3760 2778
rect 3610 2706 3760 2744
rect 3610 2672 3703 2706
rect 3737 2672 3760 2706
rect 3610 2640 3760 2672
rect 3610 2634 4000 2640
rect 3610 2600 3703 2634
rect 3737 2608 4000 2634
rect 3737 2600 3852 2608
rect 3610 2562 3852 2600
rect 3610 2528 3703 2562
rect 3737 2528 3852 2562
rect 3610 2492 3852 2528
rect 3968 2492 4000 2608
rect 3610 2490 4000 2492
rect 3610 2456 3703 2490
rect 3737 2456 4000 2490
rect 3610 2438 4000 2456
rect 3610 2418 3852 2438
rect 3610 2384 3703 2418
rect 3737 2384 3852 2418
rect 3610 2346 3852 2384
rect 3610 2312 3703 2346
rect 3737 2322 3852 2346
rect 3968 2322 4000 2438
rect 3737 2312 4000 2322
rect 3610 2274 4000 2312
rect 3610 2240 3703 2274
rect 3737 2268 4000 2274
rect 3737 2240 3852 2268
rect 3610 2202 3852 2240
rect 3610 2168 3703 2202
rect 3737 2168 3852 2202
rect 3610 2152 3852 2168
rect 3968 2152 4000 2268
rect 3610 2130 4000 2152
rect 3610 2096 3703 2130
rect 3737 2096 4000 2130
rect 3610 2090 4000 2096
rect 3610 2060 3840 2090
rect 160 2058 3840 2060
rect 160 2024 263 2058
rect 297 2024 3703 2058
rect 3737 2024 3840 2058
rect 160 1986 3840 2024
rect 160 1952 263 1986
rect 297 1952 3703 1986
rect 3737 1952 3840 1986
rect 160 1940 3840 1952
rect 160 1914 390 1940
rect 160 1910 263 1914
rect 0 1880 263 1910
rect 297 1880 390 1914
rect 0 1848 390 1880
rect 0 1732 32 1848
rect 148 1842 390 1848
rect 148 1808 263 1842
rect 297 1808 390 1842
rect 148 1770 390 1808
rect 148 1736 263 1770
rect 297 1736 390 1770
rect 148 1732 390 1736
rect 0 1698 390 1732
rect 0 1678 263 1698
rect 0 1562 32 1678
rect 148 1664 263 1678
rect 297 1664 390 1698
rect 148 1626 390 1664
rect 148 1592 263 1626
rect 297 1592 390 1626
rect 148 1562 390 1592
rect 0 1554 390 1562
rect 0 1520 263 1554
rect 297 1520 390 1554
rect 0 1508 390 1520
rect 0 1392 32 1508
rect 148 1482 390 1508
rect 148 1448 263 1482
rect 297 1448 390 1482
rect 148 1410 390 1448
rect 148 1392 263 1410
rect 0 1376 263 1392
rect 297 1376 390 1410
rect 0 1360 390 1376
rect 240 1338 390 1360
rect 240 1304 263 1338
rect 297 1304 390 1338
rect 240 1266 390 1304
rect 240 1232 263 1266
rect 297 1232 390 1266
rect 240 1194 390 1232
rect 240 1160 263 1194
rect 297 1160 390 1194
rect 240 1122 390 1160
rect 240 1088 263 1122
rect 297 1088 390 1122
rect 240 1010 390 1088
rect 0 850 240 880
rect 0 670 30 850
rect 210 670 240 850
rect 0 530 240 670
rect 0 350 30 530
rect 210 350 240 530
rect 0 240 240 350
rect 360 400 390 980
rect 420 430 450 1940
rect 480 400 510 1910
rect 540 430 570 1940
rect 600 400 630 1910
rect 660 430 690 1940
rect 720 400 750 1910
rect 780 430 810 1940
rect 840 400 870 1910
rect 900 430 930 1940
rect 960 400 990 1910
rect 1020 430 1050 1940
rect 1080 1870 1870 1910
rect 1080 1780 1200 1870
rect 1900 1840 2100 1940
rect 2130 1870 2920 1910
rect 1230 1810 2770 1840
rect 1080 1750 1870 1780
rect 1080 1660 1200 1750
rect 1900 1720 2100 1810
rect 2800 1780 2920 1870
rect 2130 1750 2920 1780
rect 1230 1690 2770 1720
rect 1080 1630 1870 1660
rect 1080 1540 1200 1630
rect 1900 1600 2100 1690
rect 2800 1660 2920 1750
rect 2130 1630 2920 1660
rect 1230 1570 2770 1600
rect 1080 1510 1870 1540
rect 1080 1420 1200 1510
rect 1900 1480 2100 1570
rect 2800 1540 2920 1630
rect 2130 1510 2920 1540
rect 1230 1450 2770 1480
rect 1080 1390 1870 1420
rect 1080 1300 1200 1390
rect 1900 1360 2100 1450
rect 2800 1420 2920 1510
rect 2130 1390 2920 1420
rect 1230 1330 2770 1360
rect 1080 1270 1870 1300
rect 1080 1180 1200 1270
rect 1900 1240 2100 1330
rect 2800 1300 2920 1390
rect 2130 1270 2920 1300
rect 1230 1210 2770 1240
rect 1080 1150 1870 1180
rect 1080 1060 1200 1150
rect 1900 1120 2100 1210
rect 2800 1180 2920 1270
rect 2130 1150 2920 1180
rect 1230 1090 2770 1120
rect 1080 1030 1870 1060
rect 1080 940 1200 1030
rect 1900 1000 2100 1090
rect 2800 1060 2920 1150
rect 2130 1030 2920 1060
rect 1230 970 2770 1000
rect 1080 910 1870 940
rect 1080 820 1200 910
rect 1900 880 2100 970
rect 2800 940 2920 1030
rect 2130 910 2920 940
rect 1230 850 2770 880
rect 1080 790 1870 820
rect 1080 700 1200 790
rect 1900 760 2100 850
rect 2800 820 2920 910
rect 2130 790 2920 820
rect 1230 730 2770 760
rect 1080 670 1870 700
rect 1080 580 1200 670
rect 1900 640 2100 730
rect 2800 700 2920 790
rect 2130 670 2920 700
rect 1230 610 2770 640
rect 1080 550 1870 580
rect 1080 460 1200 550
rect 1900 520 2100 610
rect 2800 580 2920 670
rect 2130 550 2920 580
rect 1230 490 2770 520
rect 1080 430 1870 460
rect 1080 400 1200 430
rect 1900 400 2100 490
rect 2800 460 2920 550
rect 2130 430 2920 460
rect 2950 430 2980 1940
rect 2800 400 2920 430
rect 3010 400 3040 1910
rect 3070 430 3100 1940
rect 3130 400 3160 1910
rect 3190 430 3220 1940
rect 3250 400 3280 1910
rect 3310 430 3340 1940
rect 3370 400 3400 1910
rect 3430 430 3460 1940
rect 3490 400 3520 1910
rect 3550 430 3580 1940
rect 3610 1914 3840 1940
rect 3610 1880 3703 1914
rect 3737 1910 3840 1914
rect 3970 1910 4000 2090
rect 3737 1880 4000 1910
rect 3610 1848 4000 1880
rect 3610 1842 3852 1848
rect 3610 1808 3703 1842
rect 3737 1808 3852 1842
rect 3610 1770 3852 1808
rect 3610 1736 3703 1770
rect 3737 1736 3852 1770
rect 3610 1732 3852 1736
rect 3968 1732 4000 1848
rect 3610 1698 4000 1732
rect 3610 1664 3703 1698
rect 3737 1678 4000 1698
rect 3737 1664 3852 1678
rect 3610 1626 3852 1664
rect 3610 1592 3703 1626
rect 3737 1592 3852 1626
rect 3610 1562 3852 1592
rect 3968 1562 4000 1678
rect 3610 1554 4000 1562
rect 3610 1520 3703 1554
rect 3737 1520 4000 1554
rect 3610 1508 4000 1520
rect 3610 1482 3852 1508
rect 3610 1448 3703 1482
rect 3737 1448 3852 1482
rect 3610 1410 3852 1448
rect 3610 1376 3703 1410
rect 3737 1392 3852 1410
rect 3968 1392 4000 1508
rect 3737 1376 4000 1392
rect 3610 1360 4000 1376
rect 3610 1338 3760 1360
rect 3610 1304 3703 1338
rect 3737 1304 3760 1338
rect 3610 1266 3760 1304
rect 3610 1232 3703 1266
rect 3737 1232 3760 1266
rect 3610 1194 3760 1232
rect 3610 1160 3703 1194
rect 3737 1160 3760 1194
rect 3610 1122 3760 1160
rect 3610 1088 3703 1122
rect 3737 1088 3760 1122
rect 3610 1010 3760 1088
rect 3610 400 3640 980
rect 360 347 1200 400
rect 1230 370 2770 400
rect 360 313 427 347
rect 461 313 499 347
rect 533 313 587 347
rect 621 313 659 347
rect 693 313 747 347
rect 781 313 819 347
rect 853 313 907 347
rect 941 313 979 347
rect 1013 313 1067 347
rect 1101 313 1139 347
rect 1173 340 1200 347
rect 1173 313 1870 340
rect 360 310 1870 313
rect 360 270 1200 310
rect 0 210 880 240
rect 910 210 1200 270
rect 1900 240 2100 370
rect 2800 347 3640 400
rect 2800 340 2827 347
rect 2130 313 2827 340
rect 2861 313 2899 347
rect 2933 313 2987 347
rect 3021 313 3059 347
rect 3093 313 3147 347
rect 3181 313 3219 347
rect 3253 313 3307 347
rect 3341 313 3379 347
rect 3413 313 3462 347
rect 3496 313 3534 347
rect 3568 313 3640 347
rect 2130 310 3640 313
rect 2800 270 3640 310
rect 3760 850 4000 880
rect 3760 670 3790 850
rect 3970 670 4000 850
rect 3760 530 4000 670
rect 3760 350 3790 530
rect 3970 350 4000 530
rect 0 30 30 210
rect 210 30 350 210
rect 530 30 670 210
rect 850 30 1200 210
rect 1360 210 2640 240
rect 1360 30 1390 210
rect 1570 30 1610 210
rect 1790 30 1836 210
rect 2144 30 2200 210
rect 2380 30 2430 210
rect 2610 30 2640 210
rect 2800 210 3090 270
rect 3760 240 4000 350
rect 3120 210 4000 240
rect 2800 30 3150 210
rect 3330 30 3470 210
rect 3650 30 3790 210
rect 3970 30 4000 210
rect 0 0 880 30
rect 1360 0 2640 30
rect 3120 0 4000 30
<< via1 >>
rect 30 3790 210 3970
rect 350 3790 530 3970
rect 670 3790 850 3970
rect 1390 3790 1570 3970
rect 1620 3790 1800 3970
rect 1846 3790 2154 3970
rect 2200 3790 2380 3970
rect 2430 3790 2610 3970
rect 3150 3790 3330 3970
rect 3470 3790 3650 3970
rect 3790 3790 3970 3970
rect 30 3470 210 3650
rect 30 3150 210 3330
rect 32 2492 148 2608
rect 32 2322 148 2438
rect 32 2152 148 2268
rect 3790 3470 3970 3650
rect 3790 3150 3970 3330
rect 3852 2492 3968 2608
rect 3852 2322 3968 2438
rect 3852 2152 3968 2268
rect 32 1732 148 1848
rect 32 1562 148 1678
rect 32 1392 148 1508
rect 30 670 210 850
rect 30 350 210 530
rect 3852 1732 3968 1848
rect 3852 1562 3968 1678
rect 3852 1392 3968 1508
rect 3790 670 3970 850
rect 3790 350 3970 530
rect 30 30 210 210
rect 350 30 530 210
rect 670 30 850 210
rect 1390 30 1570 210
rect 1610 30 1790 210
rect 1836 30 2144 210
rect 2200 30 2380 210
rect 2430 30 2610 210
rect 3150 30 3330 210
rect 3470 30 3650 210
rect 3790 30 3970 210
<< metal2 >>
rect 0 3970 880 4000
rect 0 3790 30 3970
rect 210 3790 350 3970
rect 530 3790 670 3970
rect 850 3790 880 3970
rect 1360 3970 2640 4000
rect 1360 3820 1390 3970
rect 0 3760 880 3790
rect 980 3790 1390 3820
rect 1570 3790 1620 3970
rect 1800 3790 1846 3970
rect 2154 3790 2200 3970
rect 2380 3790 2430 3970
rect 2610 3820 2640 3970
rect 3120 3970 4000 4000
rect 2610 3790 3020 3820
rect 0 3650 242 3760
rect 980 3720 3020 3790
rect 3120 3790 3150 3970
rect 3330 3790 3470 3970
rect 3650 3790 3790 3970
rect 3970 3790 4000 3970
rect 3120 3760 4000 3790
rect 0 3470 30 3650
rect 210 3570 242 3650
rect 360 3710 3640 3720
rect 360 3600 1120 3710
rect 210 3540 1030 3570
rect 210 3470 320 3540
rect 1060 3510 1120 3600
rect 350 3480 1120 3510
rect 0 3450 320 3470
rect 0 3420 1030 3450
rect 0 3330 320 3420
rect 1060 3390 1120 3480
rect 350 3360 1120 3390
rect 0 3150 30 3330
rect 210 3300 1030 3330
rect 210 3210 320 3300
rect 1060 3270 1120 3360
rect 350 3240 1120 3270
rect 210 3180 1030 3210
rect 210 3150 320 3180
rect 1060 3150 1120 3240
rect 0 3120 320 3150
rect 350 3120 1120 3150
rect 240 3090 320 3120
rect 240 3060 1030 3090
rect 240 2970 320 3060
rect 1060 3030 1120 3120
rect 350 3000 1120 3030
rect 240 2940 1030 2970
rect 240 2850 320 2940
rect 1060 2910 1120 3000
rect 350 2880 1120 2910
rect 240 2820 1030 2850
rect 240 2730 320 2820
rect 1060 2790 1120 2880
rect 350 2760 1120 2790
rect 240 2700 1030 2730
rect 0 2608 180 2640
rect 0 2492 32 2608
rect 148 2492 180 2608
rect 0 2438 180 2492
rect 0 2322 32 2438
rect 148 2322 180 2438
rect 0 2268 180 2322
rect 0 2152 32 2268
rect 148 2152 180 2268
rect 0 1848 180 2152
rect 0 1732 32 1848
rect 148 1732 180 1848
rect 0 1678 180 1732
rect 0 1562 32 1678
rect 148 1562 180 1678
rect 0 1508 180 1562
rect 0 1392 32 1508
rect 148 1392 180 1508
rect 0 1360 180 1392
rect 240 2610 320 2700
rect 1060 2670 1120 2760
rect 350 2640 1120 2670
rect 240 2580 1030 2610
rect 240 2490 320 2580
rect 1060 2550 1120 2640
rect 350 2520 1120 2550
rect 240 2460 1030 2490
rect 240 2370 320 2460
rect 1060 2430 1120 2520
rect 350 2400 1120 2430
rect 240 2340 1030 2370
rect 240 2250 320 2340
rect 1060 2310 1120 2400
rect 350 2280 1120 2310
rect 240 2220 1030 2250
rect 240 2130 320 2220
rect 1060 2190 1120 2280
rect 350 2160 1120 2190
rect 240 2100 1030 2130
rect 240 2040 320 2100
rect 1060 2070 1120 2160
rect 1150 2040 1180 3680
rect 1210 2070 1240 3710
rect 1270 2040 1300 3680
rect 1330 2070 1360 3710
rect 1390 2040 1420 3680
rect 1450 2070 1480 3710
rect 1510 2040 1540 3680
rect 1570 2070 1600 3710
rect 1630 2040 1660 3680
rect 1690 2070 1720 3710
rect 1750 2040 1780 3680
rect 1810 2070 1840 3710
rect 1870 2040 1900 3680
rect 240 1960 1900 2040
rect 240 1900 320 1960
rect 240 1870 1030 1900
rect 240 1780 320 1870
rect 1060 1840 1120 1930
rect 350 1810 1120 1840
rect 240 1750 1030 1780
rect 240 1660 320 1750
rect 1060 1720 1120 1810
rect 350 1690 1120 1720
rect 240 1630 1030 1660
rect 240 1540 320 1630
rect 1060 1600 1120 1690
rect 350 1570 1120 1600
rect 240 1510 1030 1540
rect 240 1420 320 1510
rect 1060 1480 1120 1570
rect 350 1450 1120 1480
rect 240 1390 1030 1420
rect 240 1300 320 1390
rect 1060 1360 1120 1450
rect 350 1330 1120 1360
rect 240 1270 1030 1300
rect 240 1180 320 1270
rect 1060 1240 1120 1330
rect 350 1210 1120 1240
rect 240 1150 1030 1180
rect 240 1060 320 1150
rect 1060 1120 1120 1210
rect 350 1090 1120 1120
rect 240 1030 1030 1060
rect 240 940 320 1030
rect 1060 1000 1120 1090
rect 350 970 1120 1000
rect 240 910 1030 940
rect 240 880 320 910
rect 1060 880 1120 970
rect 0 850 320 880
rect 350 850 1120 880
rect 0 670 30 850
rect 210 820 320 850
rect 210 790 1030 820
rect 210 700 320 790
rect 1060 760 1120 850
rect 350 730 1120 760
rect 210 670 1030 700
rect 0 580 320 670
rect 1060 640 1120 730
rect 350 610 1120 640
rect 0 550 1030 580
rect 0 530 320 550
rect 0 350 30 530
rect 210 460 320 530
rect 1060 520 1120 610
rect 350 490 1120 520
rect 210 430 1030 460
rect 210 350 240 430
rect 1060 400 1120 490
rect 0 240 240 350
rect 360 290 1120 400
rect 1150 320 1180 1960
rect 1210 290 1240 1930
rect 1270 320 1300 1960
rect 1330 290 1360 1930
rect 1390 320 1420 1960
rect 1450 290 1480 1930
rect 1510 320 1540 1960
rect 1570 290 1600 1930
rect 1630 320 1660 1960
rect 1690 290 1720 1930
rect 1750 320 1780 1960
rect 1810 290 1840 1930
rect 1870 320 1900 1960
rect 1930 290 2070 3710
rect 2100 2040 2130 3680
rect 2160 2070 2190 3710
rect 2220 2040 2250 3680
rect 2280 2070 2310 3710
rect 2340 2040 2370 3680
rect 2400 2070 2430 3710
rect 2460 2040 2490 3680
rect 2520 2070 2550 3710
rect 2580 2040 2610 3680
rect 2640 2070 2670 3710
rect 2700 2040 2730 3680
rect 2760 2070 2790 3710
rect 2820 2040 2850 3680
rect 2880 3600 3640 3710
rect 3760 3650 4000 3760
rect 2880 3510 2940 3600
rect 3760 3570 3790 3650
rect 2970 3540 3790 3570
rect 2880 3480 3650 3510
rect 2880 3390 2940 3480
rect 3680 3470 3790 3540
rect 3970 3470 4000 3650
rect 3680 3450 4000 3470
rect 2970 3420 4000 3450
rect 2880 3360 3650 3390
rect 2880 3270 2940 3360
rect 3680 3330 4000 3420
rect 2970 3300 3790 3330
rect 2880 3240 3650 3270
rect 2880 3150 2940 3240
rect 3680 3210 3790 3300
rect 2970 3180 3790 3210
rect 3680 3150 3790 3180
rect 3970 3150 4000 3330
rect 2880 3120 3650 3150
rect 3680 3120 4000 3150
rect 2880 3030 2940 3120
rect 3680 3090 3760 3120
rect 2970 3060 3760 3090
rect 2880 3000 3650 3030
rect 2880 2910 2940 3000
rect 3680 2970 3760 3060
rect 2970 2940 3760 2970
rect 2880 2880 3650 2910
rect 2880 2790 2940 2880
rect 3680 2850 3760 2940
rect 2970 2820 3760 2850
rect 2880 2760 3650 2790
rect 2880 2670 2940 2760
rect 3680 2730 3760 2820
rect 2970 2700 3760 2730
rect 2880 2640 3650 2670
rect 2880 2550 2940 2640
rect 3680 2610 3760 2700
rect 2970 2580 3760 2610
rect 2880 2520 3650 2550
rect 2880 2430 2940 2520
rect 3680 2490 3760 2580
rect 2970 2460 3760 2490
rect 2880 2400 3650 2430
rect 2880 2310 2940 2400
rect 3680 2370 3760 2460
rect 2970 2340 3760 2370
rect 2880 2280 3650 2310
rect 2880 2190 2940 2280
rect 3680 2250 3760 2340
rect 2970 2220 3760 2250
rect 2880 2160 3650 2190
rect 2880 2070 2940 2160
rect 3680 2130 3760 2220
rect 2970 2100 3760 2130
rect 3680 2040 3760 2100
rect 2100 1960 3760 2040
rect 2100 320 2130 1960
rect 2160 290 2190 1930
rect 2220 320 2250 1960
rect 2280 290 2310 1930
rect 2340 320 2370 1960
rect 2400 290 2430 1930
rect 2460 320 2490 1960
rect 2520 290 2550 1930
rect 2580 320 2610 1960
rect 2640 290 2670 1930
rect 2700 320 2730 1960
rect 2760 290 2790 1930
rect 2820 320 2850 1960
rect 2880 1840 2940 1930
rect 3680 1900 3760 1960
rect 2970 1870 3760 1900
rect 2880 1810 3650 1840
rect 2880 1720 2940 1810
rect 3680 1780 3760 1870
rect 2970 1750 3760 1780
rect 2880 1690 3650 1720
rect 2880 1600 2940 1690
rect 3680 1660 3760 1750
rect 2970 1630 3760 1660
rect 2880 1570 3650 1600
rect 2880 1480 2940 1570
rect 3680 1540 3760 1630
rect 2970 1510 3760 1540
rect 2880 1450 3650 1480
rect 2880 1360 2940 1450
rect 3680 1420 3760 1510
rect 2970 1390 3760 1420
rect 2880 1330 3650 1360
rect 2880 1240 2940 1330
rect 3680 1300 3760 1390
rect 3820 2608 4000 2640
rect 3820 2492 3852 2608
rect 3968 2492 4000 2608
rect 3820 2438 4000 2492
rect 3820 2322 3852 2438
rect 3968 2322 4000 2438
rect 3820 2268 4000 2322
rect 3820 2152 3852 2268
rect 3968 2152 4000 2268
rect 3820 1848 4000 2152
rect 3820 1732 3852 1848
rect 3968 1732 4000 1848
rect 3820 1678 4000 1732
rect 3820 1562 3852 1678
rect 3968 1562 4000 1678
rect 3820 1508 4000 1562
rect 3820 1392 3852 1508
rect 3968 1392 4000 1508
rect 3820 1360 4000 1392
rect 2970 1270 3760 1300
rect 2880 1210 3650 1240
rect 2880 1120 2940 1210
rect 3680 1180 3760 1270
rect 2970 1150 3760 1180
rect 2880 1090 3650 1120
rect 2880 1000 2940 1090
rect 3680 1060 3760 1150
rect 2970 1030 3760 1060
rect 2880 970 3650 1000
rect 2880 880 2940 970
rect 3680 940 3760 1030
rect 2970 910 3760 940
rect 3680 880 3760 910
rect 2880 850 3650 880
rect 3680 850 4000 880
rect 2880 760 2940 850
rect 3680 820 3790 850
rect 2970 790 3790 820
rect 2880 730 3650 760
rect 2880 640 2940 730
rect 3680 700 3790 790
rect 2970 670 3790 700
rect 3970 670 4000 850
rect 2880 610 3650 640
rect 2880 520 2940 610
rect 3680 580 4000 670
rect 2970 550 4000 580
rect 3680 530 4000 550
rect 2880 490 3650 520
rect 2880 400 2940 490
rect 3680 460 3790 530
rect 2970 430 3790 460
rect 2880 290 3640 400
rect 360 280 3640 290
rect 3760 350 3790 430
rect 3970 350 4000 530
rect 0 210 880 240
rect 0 30 30 210
rect 210 30 350 210
rect 530 30 670 210
rect 850 30 880 210
rect 980 210 3020 280
rect 3760 240 4000 350
rect 980 180 1390 210
rect 0 0 880 30
rect 1360 30 1390 180
rect 1570 30 1610 210
rect 1790 30 1836 210
rect 2144 30 2200 210
rect 2380 30 2430 210
rect 2610 180 3020 210
rect 3120 210 4000 240
rect 2610 30 2640 180
rect 1360 0 2640 30
rect 3120 30 3150 210
rect 3330 30 3470 210
rect 3650 30 3790 210
rect 3970 30 4000 210
rect 3120 0 4000 30
<< metal3 >>
rect 0 3967 880 4000
rect 0 3823 33 3967
rect 177 3823 223 3967
rect 367 3823 513 3967
rect 657 3823 703 3967
rect 847 3823 880 3967
rect 1360 3947 2640 4000
rect 1360 3883 1413 3947
rect 1477 3883 1573 3947
rect 1637 3883 1733 3947
rect 1797 3883 2203 3947
rect 2267 3883 2363 3947
rect 2427 3883 2523 3947
rect 2587 3883 2640 3947
rect 1360 3830 2640 3883
rect 3120 3967 4000 4000
rect 0 3777 880 3823
rect 0 3633 33 3777
rect 177 3750 880 3777
rect 3120 3823 3153 3967
rect 3297 3823 3343 3967
rect 3487 3823 3633 3967
rect 3777 3823 3823 3967
rect 3967 3823 4000 3967
rect 3120 3777 4000 3823
rect 3120 3750 3823 3777
rect 177 3633 3823 3750
rect 3967 3633 4000 3777
rect 0 3487 4000 3633
rect 0 3343 33 3487
rect 177 3343 3823 3487
rect 3967 3343 4000 3487
rect 0 3297 4000 3343
rect 0 3153 33 3297
rect 177 3153 3823 3297
rect 3967 3153 4000 3297
rect 0 3120 4000 3153
rect 0 2587 170 2640
rect 0 2523 53 2587
rect 117 2523 170 2587
rect 0 2427 170 2523
rect 0 2363 53 2427
rect 117 2363 170 2427
rect 0 2267 170 2363
rect 0 2203 53 2267
rect 117 2203 170 2267
rect 0 1797 170 2203
rect 0 1733 53 1797
rect 117 1733 170 1797
rect 0 1637 170 1733
rect 0 1573 53 1637
rect 117 1573 170 1637
rect 0 1477 170 1573
rect 0 1413 53 1477
rect 117 1413 170 1477
rect 0 1360 170 1413
rect 250 880 3750 3120
rect 3830 2587 4000 2640
rect 3830 2523 3883 2587
rect 3947 2523 4000 2587
rect 3830 2427 4000 2523
rect 3830 2363 3883 2427
rect 3947 2363 4000 2427
rect 3830 2267 4000 2363
rect 3830 2203 3883 2267
rect 3947 2203 4000 2267
rect 3830 1797 4000 2203
rect 3830 1733 3883 1797
rect 3947 1733 4000 1797
rect 3830 1637 4000 1733
rect 3830 1573 3883 1637
rect 3947 1573 4000 1637
rect 3830 1477 4000 1573
rect 3830 1413 3883 1477
rect 3947 1413 4000 1477
rect 3830 1360 4000 1413
rect 0 847 4000 880
rect 0 703 33 847
rect 177 703 3823 847
rect 3967 703 4000 847
rect 0 657 4000 703
rect 0 513 33 657
rect 177 513 3823 657
rect 3967 513 4000 657
rect 0 367 4000 513
rect 0 223 33 367
rect 177 250 3823 367
rect 177 223 880 250
rect 0 177 880 223
rect 0 33 33 177
rect 177 33 223 177
rect 367 33 513 177
rect 657 33 703 177
rect 847 33 880 177
rect 3120 223 3823 250
rect 3967 223 4000 367
rect 3120 177 4000 223
rect 0 0 880 33
rect 1360 117 2640 170
rect 1360 53 1413 117
rect 1477 53 1573 117
rect 1637 53 1733 117
rect 1797 53 2203 117
rect 2267 53 2363 117
rect 2427 53 2523 117
rect 2587 53 2640 117
rect 1360 0 2640 53
rect 3120 33 3153 177
rect 3297 33 3343 177
rect 3487 33 3633 177
rect 3777 33 3823 177
rect 3967 33 4000 177
rect 3120 0 4000 33
<< via3 >>
rect 33 3823 177 3967
rect 223 3823 367 3967
rect 513 3823 657 3967
rect 703 3823 847 3967
rect 1413 3883 1477 3947
rect 1573 3883 1637 3947
rect 1733 3883 1797 3947
rect 2203 3883 2267 3947
rect 2363 3883 2427 3947
rect 2523 3883 2587 3947
rect 33 3633 177 3777
rect 3153 3823 3297 3967
rect 3343 3823 3487 3967
rect 3633 3823 3777 3967
rect 3823 3823 3967 3967
rect 3823 3633 3967 3777
rect 33 3343 177 3487
rect 3823 3343 3967 3487
rect 33 3153 177 3297
rect 3823 3153 3967 3297
rect 53 2523 117 2587
rect 53 2363 117 2427
rect 53 2203 117 2267
rect 53 1733 117 1797
rect 53 1573 117 1637
rect 53 1413 117 1477
rect 3883 2523 3947 2587
rect 3883 2363 3947 2427
rect 3883 2203 3947 2267
rect 3883 1733 3947 1797
rect 3883 1573 3947 1637
rect 3883 1413 3947 1477
rect 33 703 177 847
rect 3823 703 3967 847
rect 33 513 177 657
rect 3823 513 3967 657
rect 33 223 177 367
rect 33 33 177 177
rect 223 33 367 177
rect 513 33 657 177
rect 703 33 847 177
rect 3823 223 3967 367
rect 1413 53 1477 117
rect 1573 53 1637 117
rect 1733 53 1797 117
rect 2203 53 2267 117
rect 2363 53 2427 117
rect 2523 53 2587 117
rect 3153 33 3297 177
rect 3343 33 3487 177
rect 3633 33 3777 177
rect 3823 33 3967 177
<< mimcap >>
rect 280 3672 3720 3720
rect 280 328 328 3672
rect 3672 328 3720 3672
rect 280 280 3720 328
<< mimcapcontact >>
rect 328 328 3672 3672
<< metal4 >>
rect 0 3967 880 4000
rect 0 3823 33 3967
rect 177 3823 223 3967
rect 367 3823 513 3967
rect 657 3823 703 3967
rect 847 3823 880 3967
rect 0 3790 880 3823
rect 1360 3947 2640 4000
rect 1360 3883 1413 3947
rect 1477 3883 1573 3947
rect 1637 3883 1733 3947
rect 1797 3883 2203 3947
rect 2267 3883 2363 3947
rect 2427 3883 2523 3947
rect 2587 3883 2640 3947
rect 0 3777 210 3790
rect 0 3633 33 3777
rect 177 3633 210 3777
rect 1360 3710 2640 3883
rect 3120 3967 4000 4000
rect 3120 3823 3153 3967
rect 3297 3823 3343 3967
rect 3487 3823 3633 3967
rect 3777 3823 3823 3967
rect 3967 3823 4000 3967
rect 3120 3790 4000 3823
rect 3790 3777 4000 3790
rect 0 3487 210 3633
rect 0 3343 33 3487
rect 177 3343 210 3487
rect 0 3297 210 3343
rect 0 3153 33 3297
rect 177 3153 210 3297
rect 0 3120 210 3153
rect 290 3672 3710 3710
rect 290 2640 328 3672
rect 0 2587 328 2640
rect 0 2523 53 2587
rect 117 2523 328 2587
rect 0 2427 328 2523
rect 0 2363 53 2427
rect 117 2363 328 2427
rect 0 2267 328 2363
rect 0 2203 53 2267
rect 117 2203 328 2267
rect 0 1797 328 2203
rect 0 1733 53 1797
rect 117 1733 328 1797
rect 0 1637 328 1733
rect 0 1573 53 1637
rect 117 1573 328 1637
rect 0 1477 328 1573
rect 0 1413 53 1477
rect 117 1413 328 1477
rect 0 1360 328 1413
rect 0 847 210 880
rect 0 703 33 847
rect 177 703 210 847
rect 0 657 210 703
rect 0 513 33 657
rect 177 513 210 657
rect 0 367 210 513
rect 0 223 33 367
rect 177 223 210 367
rect 290 328 328 1360
rect 3672 2640 3710 3672
rect 3790 3633 3823 3777
rect 3967 3633 4000 3777
rect 3790 3487 4000 3633
rect 3790 3343 3823 3487
rect 3967 3343 4000 3487
rect 3790 3297 4000 3343
rect 3790 3153 3823 3297
rect 3967 3153 4000 3297
rect 3790 3120 4000 3153
rect 3672 2587 4000 2640
rect 3672 2523 3883 2587
rect 3947 2523 4000 2587
rect 3672 2427 4000 2523
rect 3672 2363 3883 2427
rect 3947 2363 4000 2427
rect 3672 2267 4000 2363
rect 3672 2203 3883 2267
rect 3947 2203 4000 2267
rect 3672 1797 4000 2203
rect 3672 1733 3883 1797
rect 3947 1733 4000 1797
rect 3672 1637 4000 1733
rect 3672 1573 3883 1637
rect 3947 1573 4000 1637
rect 3672 1477 4000 1573
rect 3672 1413 3883 1477
rect 3947 1413 4000 1477
rect 3672 1360 4000 1413
rect 3672 328 3710 1360
rect 290 290 3710 328
rect 3790 847 4000 880
rect 3790 703 3823 847
rect 3967 703 4000 847
rect 3790 657 4000 703
rect 3790 513 3823 657
rect 3967 513 4000 657
rect 3790 367 4000 513
rect 0 210 210 223
rect 0 177 880 210
rect 0 33 33 177
rect 177 33 223 177
rect 367 33 513 177
rect 657 33 703 177
rect 847 33 880 177
rect 0 0 880 33
rect 1360 117 2640 290
rect 3790 223 3823 367
rect 3967 223 4000 367
rect 3790 210 4000 223
rect 1360 53 1413 117
rect 1477 53 1573 117
rect 1637 53 1733 117
rect 1797 53 2203 117
rect 2267 53 2363 117
rect 2427 53 2523 117
rect 2587 53 2640 117
rect 1360 0 2640 53
rect 3120 177 4000 210
rect 3120 33 3153 177
rect 3297 33 3343 177
rect 3487 33 3633 177
rect 3777 33 3823 177
rect 3967 33 4000 177
rect 3120 0 4000 33
<< labels >>
flabel metal1 s 1360 0 2640 180 5 FreeSans 400 0 0 0 nmoscap_top
port 1 nsew
flabel metal1 s 1360 3820 2640 4000 1 FreeSans 400 0 0 0 nmoscap_top
port 1 nsew
flabel metal1 s 3974 1360 4000 2640 3 FreeSans 400 90 0 0 nmoscap_top
port 1 nsew
flabel metal1 s 0 1360 26 2640 7 FreeSans 400 90 0 0 nmoscap_top
port 1 nsew
flabel metal1 s 0 3120 240 4000 7 FreeSans 400 90 0 0 nmoscap_bot
port 2 nsew
flabel metal1 s 0 0 240 880 7 FreeSans 400 90 0 0 nmoscap_bot
port 2 nsew
flabel metal1 s 3760 0 4000 880 3 FreeSans 400 90 0 0 nmoscap_bot
port 2 nsew
flabel metal1 s 3760 3120 4000 4000 3 FreeSans 400 90 0 0 nmoscap_bot
port 2 nsew
flabel metal1 s 3120 3760 4000 4000 1 FreeSans 400 0 0 0 nmoscap_bot
port 2 nsew
flabel metal1 s 0 3760 880 4000 1 FreeSans 400 0 0 0 nmoscap_bot
port 2 nsew
flabel metal1 s 0 0 880 240 5 FreeSans 400 0 0 0 nmoscap_bot
port 2 nsew
flabel metal1 s 3120 0 4000 240 5 FreeSans 400 0 0 0 nmoscap_bot
port 2 nsew
flabel locali s 890 0 1350 80 5 FreeSans 400 0 0 0 pwell
port 3 nsew
flabel locali s 2650 0 3110 80 5 FreeSans 400 0 0 0 pwell
port 3 nsew
flabel locali s 2650 3920 3110 4000 1 FreeSans 400 0 0 0 pwell
port 3 nsew
flabel locali s 890 3920 1350 4000 1 FreeSans 400 0 0 0 pwell
port 3 nsew
flabel locali s 3920 2650 4000 3110 3 FreeSans 400 90 0 0 pwell
port 3 nsew
flabel locali s 3920 890 4000 1350 3 FreeSans 400 90 0 0 pwell
port 3 nsew
flabel locali s 0 890 80 1350 7 FreeSans 400 90 0 0 pwell
port 3 nsew
flabel locali s 0 2650 80 3110 7 FreeSans 400 90 0 0 pwell
port 3 nsew
flabel metal4 s 1360 3830 2640 4000 1 FreeSans 400 0 0 0 mimcap_top
port 4 nsew
flabel metal4 s 1360 0 2640 170 5 FreeSans 400 0 0 0 mimcap_top
port 4 nsew
flabel metal4 s 3830 1360 4000 2640 3 FreeSans 400 90 0 0 mimcap_top
port 4 nsew
flabel metal4 s 0 1360 170 2640 7 FreeSans 400 90 0 0 mimcap_top
port 4 nsew
flabel metal4 s 3120 0 4000 210 5 FreeSans 400 0 0 0 mimcap_bot
port 5 nsew
flabel metal4 s 0 0 880 210 5 FreeSans 400 0 0 0 mimcap_bot
port 5 nsew
flabel metal4 s 0 3790 880 4000 1 FreeSans 400 0 0 0 mimcap_bot
port 5 nsew
flabel metal4 s 3120 3790 4000 4000 1 FreeSans 400 0 0 0 mimcap_bot
port 5 nsew
flabel metal4 s 3790 3120 4000 4000 3 FreeSans 400 90 0 0 mimcap_bot
port 5 nsew
flabel metal4 s 3790 0 4000 880 3 FreeSans 400 90 0 0 mimcap_bot
port 5 nsew
flabel metal4 s 0 0 210 880 7 FreeSans 400 90 0 0 mimcap_bot
port 5 nsew
flabel metal4 s 0 3120 210 4000 7 FreeSans 400 90 0 0 mimcap_bot
port 5 nsew
<< properties >>
string FIXED_BBOX 0 0 4000 4000
string GDS_END 423956
string GDS_FILE adc_top.gds.gz
string GDS_START 206808
<< end >>
