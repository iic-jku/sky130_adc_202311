magic
tech sky130A
magscale 1 2
timestamp 1698052002
<< locali >>
rect -58 17777 1358 18777
rect -58 10919 1047 17777
rect 2410 17436 2507 17637
rect -58 9919 1418 10919
rect -58 3061 1047 9919
rect 2410 9578 2507 9779
rect -58 2061 1449 3061
rect -58 -1553 1047 2061
rect 2410 1720 2507 1921
rect -58 -2553 1415 -1553
rect -58 -4545 1047 -2553
rect 2410 -2894 2507 -2693
rect -58 -5545 1402 -4545
rect -58 -7537 1047 -5545
rect 2410 -5886 2507 -5685
rect -58 -8537 1442 -7537
rect 2410 -8878 2507 -8677
<< metal1 >>
rect 2201 17434 2299 17746
rect 2201 9576 2299 9888
rect 2201 1718 2299 2030
rect 2201 -2896 2299 -2584
rect 2201 -5888 2299 -5576
rect 2201 -8880 2299 -8568
<< metal2 >>
rect 2653 19457 3254 19467
rect 2653 19285 2689 19457
rect 3089 19285 3254 19457
rect 2653 19275 3254 19285
rect 1289 19217 1890 19227
rect 1289 19045 1459 19217
rect 1859 19045 1890 19217
rect 1289 19035 1890 19045
rect 2653 11599 3254 11609
rect 2653 11427 2689 11599
rect 3089 11427 3254 11599
rect 2653 11417 3254 11427
rect 1289 11359 1890 11369
rect 1289 11187 1459 11359
rect 1859 11187 1890 11359
rect 1289 11177 1890 11187
rect 2653 3741 3254 3751
rect 2653 3569 2689 3741
rect 3089 3569 3254 3741
rect 2653 3559 3254 3569
rect 1289 3501 1890 3511
rect 1289 3329 1459 3501
rect 1859 3329 1890 3501
rect 1289 3319 1890 3329
rect 2653 -873 3254 -863
rect 2653 -1045 2689 -873
rect 3089 -1045 3254 -873
rect 2653 -1055 3254 -1045
rect 1289 -1113 1890 -1103
rect 1289 -1285 1459 -1113
rect 1859 -1285 1890 -1113
rect 1289 -1295 1890 -1285
rect 2653 -3865 3254 -3855
rect 2653 -4037 2689 -3865
rect 3089 -4037 3254 -3865
rect 2653 -4047 3254 -4037
rect 1289 -4105 1890 -4095
rect 1289 -4277 1459 -4105
rect 1859 -4277 1890 -4105
rect 1289 -4287 1890 -4277
rect 2653 -6857 3254 -6847
rect 2653 -7029 2689 -6857
rect 3089 -7029 3254 -6857
rect 2653 -7039 3254 -7029
rect 1289 -7097 1890 -7087
rect 1289 -7269 1459 -7097
rect 1859 -7269 1890 -7097
rect 1289 -7279 1890 -7269
<< via2 >>
rect 2689 19285 3089 19457
rect 1459 19045 1859 19217
rect 2689 11427 3089 11599
rect 1459 11187 1859 11359
rect 2689 3569 3089 3741
rect 1459 3329 1859 3501
rect 2689 -1045 3089 -873
rect 1459 -1285 1859 -1113
rect 2689 -4037 3089 -3865
rect 1459 -4277 1859 -4105
rect 2689 -7029 3089 -6857
rect 1459 -7269 1859 -7097
<< metal3 >>
rect 1282 19476 1890 19482
rect 1282 19026 1288 19476
rect 1884 19026 1890 19476
rect 1282 19020 1890 19026
rect 2653 19476 3260 19482
rect 2653 19026 2659 19476
rect 3254 19026 3260 19476
rect 2653 19020 3260 19026
rect 1282 11618 1890 11624
rect 1282 11168 1288 11618
rect 1884 11168 1890 11618
rect 1282 11162 1890 11168
rect 2653 11618 3260 11624
rect 2653 11168 2659 11618
rect 3254 11168 3260 11618
rect 2653 11162 3260 11168
rect 1282 3760 1890 3766
rect 1282 3310 1288 3760
rect 1884 3310 1890 3760
rect 1282 3304 1890 3310
rect 2653 3760 3260 3766
rect 2653 3310 2659 3760
rect 3254 3310 3260 3760
rect 2653 3304 3260 3310
rect 1282 -854 1890 -848
rect 1282 -1304 1288 -854
rect 1884 -1304 1890 -854
rect 1282 -1310 1890 -1304
rect 2653 -854 3260 -848
rect 2653 -1304 2659 -854
rect 3254 -1304 3260 -854
rect 2653 -1310 3260 -1304
rect 1282 -3846 1890 -3840
rect 1282 -4296 1288 -3846
rect 1884 -4296 1890 -3846
rect 1282 -4302 1890 -4296
rect 2653 -3846 3260 -3840
rect 2653 -4296 2659 -3846
rect 3254 -4296 3260 -3846
rect 2653 -4302 3260 -4296
rect 1282 -6838 1890 -6832
rect 1282 -7288 1288 -6838
rect 1884 -7288 1890 -6838
rect 1282 -7294 1890 -7288
rect 2653 -6838 3260 -6832
rect 2653 -7288 2659 -6838
rect 3254 -7288 3260 -6838
rect 2653 -7294 3260 -7288
<< via3 >>
rect 1288 19217 1884 19476
rect 1288 19045 1459 19217
rect 1459 19045 1859 19217
rect 1859 19045 1884 19217
rect 1288 19026 1884 19045
rect 2659 19457 3254 19476
rect 2659 19285 2689 19457
rect 2689 19285 3089 19457
rect 3089 19285 3254 19457
rect 2659 19026 3254 19285
rect 1288 11359 1884 11618
rect 1288 11187 1459 11359
rect 1459 11187 1859 11359
rect 1859 11187 1884 11359
rect 1288 11168 1884 11187
rect 2659 11599 3254 11618
rect 2659 11427 2689 11599
rect 2689 11427 3089 11599
rect 3089 11427 3254 11599
rect 2659 11168 3254 11427
rect 1288 3501 1884 3760
rect 1288 3329 1459 3501
rect 1459 3329 1859 3501
rect 1859 3329 1884 3501
rect 1288 3310 1884 3329
rect 2659 3741 3254 3760
rect 2659 3569 2689 3741
rect 2689 3569 3089 3741
rect 3089 3569 3254 3741
rect 2659 3310 3254 3569
rect 1288 -1113 1884 -854
rect 1288 -1285 1459 -1113
rect 1459 -1285 1859 -1113
rect 1859 -1285 1884 -1113
rect 1288 -1304 1884 -1285
rect 2659 -873 3254 -854
rect 2659 -1045 2689 -873
rect 2689 -1045 3089 -873
rect 3089 -1045 3254 -873
rect 2659 -1304 3254 -1045
rect 1288 -4105 1884 -3846
rect 1288 -4277 1459 -4105
rect 1459 -4277 1859 -4105
rect 1859 -4277 1884 -4105
rect 1288 -4296 1884 -4277
rect 2659 -3865 3254 -3846
rect 2659 -4037 2689 -3865
rect 2689 -4037 3089 -3865
rect 3089 -4037 3254 -3865
rect 2659 -4296 3254 -4037
rect 1288 -7097 1884 -6838
rect 1288 -7269 1459 -7097
rect 1459 -7269 1859 -7097
rect 1859 -7269 1884 -7097
rect 1288 -7288 1884 -7269
rect 2659 -6857 3254 -6838
rect 2659 -7029 2689 -6857
rect 2689 -7029 3089 -6857
rect 3089 -7029 3254 -6857
rect 2659 -7288 3254 -7029
<< metal4 >>
rect -4432 19476 1943 19536
rect -4432 19026 1003 19476
rect 1884 19026 1943 19476
rect -4432 18966 1943 19026
rect 2599 19476 8974 19536
rect 2599 19026 2659 19476
rect 3540 19026 8974 19476
rect 2599 18966 8974 19026
rect -4432 17854 1943 17914
rect -4432 17404 -1397 17854
rect -516 17404 1943 17854
rect -4432 17344 1943 17404
rect 2599 17854 8974 17914
rect 2599 17404 5059 17854
rect 5940 17404 8974 17854
rect 2599 17344 8974 17404
rect -4432 16232 1943 16292
rect -4432 15782 1003 16232
rect 1884 15782 1943 16232
rect -4432 15722 1943 15782
rect 2599 16232 8974 16292
rect 2599 15782 2659 16232
rect 3540 15782 8974 16232
rect 2599 15722 8974 15782
rect -4432 14610 1943 14670
rect -4432 14160 -1397 14610
rect -516 14160 1943 14610
rect -4432 14100 1943 14160
rect 2599 14610 8974 14670
rect 2599 14160 5059 14610
rect 5940 14160 8974 14610
rect 2599 14100 8974 14160
rect -4432 12988 1943 13048
rect -4432 12538 1003 12988
rect 1884 12538 1943 12988
rect -4432 12478 1943 12538
rect 2599 12988 8974 13048
rect 2599 12538 2659 12988
rect 3540 12538 8974 12988
rect 2599 12478 8974 12538
rect -4432 11618 1943 11678
rect -4432 11168 1003 11618
rect 1884 11168 1943 11618
rect -4432 11108 1943 11168
rect 2599 11618 8974 11678
rect 2599 11168 2659 11618
rect 3540 11168 8974 11618
rect 2599 11108 8974 11168
rect -4432 9996 1943 10056
rect -4432 9546 -1397 9996
rect -516 9546 1943 9996
rect -4432 9486 1943 9546
rect 2599 9996 8974 10056
rect 2599 9546 5059 9996
rect 5940 9546 8974 9996
rect 2599 9486 8974 9546
rect -4432 8374 1943 8434
rect -4432 7924 1003 8374
rect 1884 7924 1943 8374
rect -4432 7864 1943 7924
rect 2599 8374 8974 8434
rect 2599 7924 2659 8374
rect 3540 7924 8974 8374
rect 2599 7864 8974 7924
rect -4432 6752 1943 6812
rect -4432 6302 -1397 6752
rect -516 6302 1943 6752
rect -4432 6242 1943 6302
rect 2599 6752 8974 6812
rect 2599 6302 5059 6752
rect 5940 6302 8974 6752
rect 2599 6242 8974 6302
rect -4432 5130 1943 5190
rect -4432 4680 1003 5130
rect 1884 4680 1943 5130
rect -4432 4620 1943 4680
rect 2599 5130 8974 5190
rect 2599 4680 2659 5130
rect 3540 4680 8974 5130
rect 2599 4620 8974 4680
rect -4432 3760 1943 3820
rect -4432 3310 1003 3760
rect 1884 3310 1943 3760
rect -4432 3250 1943 3310
rect 2599 3760 8974 3820
rect 2599 3310 2659 3760
rect 3540 3310 8974 3760
rect 2599 3250 8974 3310
rect -4432 2138 1943 2198
rect -4432 1688 -1397 2138
rect -516 1688 1943 2138
rect -4432 1628 1943 1688
rect 2599 2138 8974 2198
rect 2599 1688 5059 2138
rect 5940 1688 8974 2138
rect 2599 1628 8974 1688
rect -4432 516 1943 576
rect -4432 66 1003 516
rect 1884 66 1943 516
rect -4432 6 1943 66
rect 2599 516 8974 576
rect 2599 66 2659 516
rect 3540 66 8974 516
rect 2599 6 8974 66
rect -4432 -854 1943 -794
rect -4432 -1304 1003 -854
rect 1884 -1304 1943 -854
rect -4432 -1364 1943 -1304
rect 2599 -854 8974 -794
rect 2599 -1304 2659 -854
rect 3540 -1304 8974 -854
rect 2599 -1364 8974 -1304
rect -4432 -2476 1943 -2416
rect -4432 -2926 -1397 -2476
rect -516 -2926 1943 -2476
rect -4432 -2986 1943 -2926
rect 2599 -2476 8974 -2416
rect 2599 -2926 5059 -2476
rect 5940 -2926 8974 -2476
rect 2599 -2986 8974 -2926
rect -4432 -3846 1943 -3786
rect -4432 -4296 1003 -3846
rect 1884 -4296 1943 -3846
rect -4432 -4356 1943 -4296
rect 2599 -3846 8974 -3786
rect 2599 -4296 2659 -3846
rect 3540 -4296 8974 -3846
rect 2599 -4356 8974 -4296
rect -4432 -5468 1943 -5408
rect -4432 -5918 -1397 -5468
rect -516 -5918 1943 -5468
rect -4432 -5978 1943 -5918
rect 2599 -5468 8974 -5408
rect 2599 -5918 5059 -5468
rect 5940 -5918 8974 -5468
rect 2599 -5978 8974 -5918
rect -4432 -6838 1943 -6778
rect -4432 -7288 1003 -6838
rect 1884 -7288 1943 -6838
rect -4432 -7348 1943 -7288
rect 2599 -6838 8974 -6778
rect 2599 -7288 2659 -6838
rect 3540 -7288 8974 -6838
rect 2599 -7348 8974 -7288
rect -4432 -8460 1943 -8400
rect -4432 -8910 -1397 -8460
rect -516 -8910 1943 -8460
rect -4432 -8970 1943 -8910
rect 2599 -8460 8974 -8400
rect 2599 -8910 5059 -8460
rect 5940 -8910 8974 -8460
rect 2599 -8970 8974 -8910
<< via4 >>
rect 1003 19026 1288 19476
rect 1288 19026 1884 19476
rect 2659 19026 3254 19476
rect 3254 19026 3540 19476
rect -1397 17404 -516 17854
rect 5059 17404 5940 17854
rect 1003 15782 1884 16232
rect 2659 15782 3540 16232
rect -1397 14160 -516 14610
rect 5059 14160 5940 14610
rect 1003 12538 1884 12988
rect 2659 12538 3540 12988
rect 1003 11168 1288 11618
rect 1288 11168 1884 11618
rect 2659 11168 3254 11618
rect 3254 11168 3540 11618
rect -1397 9546 -516 9996
rect 5059 9546 5940 9996
rect 1003 7924 1884 8374
rect 2659 7924 3540 8374
rect -1397 6302 -516 6752
rect 5059 6302 5940 6752
rect 1003 4680 1884 5130
rect 2659 4680 3540 5130
rect 1003 3310 1288 3760
rect 1288 3310 1884 3760
rect 2659 3310 3254 3760
rect 3254 3310 3540 3760
rect -1397 1688 -516 2138
rect 5059 1688 5940 2138
rect 1003 66 1884 516
rect 2659 66 3540 516
rect 1003 -1304 1288 -854
rect 1288 -1304 1884 -854
rect 2659 -1304 3254 -854
rect 3254 -1304 3540 -854
rect -1397 -2926 -516 -2476
rect 5059 -2926 5940 -2476
rect 1003 -4296 1288 -3846
rect 1288 -4296 1884 -3846
rect 2659 -4296 3254 -3846
rect 3254 -4296 3540 -3846
rect -1397 -5918 -516 -5468
rect 5059 -5918 5940 -5468
rect 1003 -7288 1288 -6838
rect 1288 -7288 1884 -6838
rect 2659 -7288 3254 -6838
rect 3254 -7288 3540 -6838
rect -1397 -8910 -516 -8460
rect 5059 -8910 5940 -8460
<< metal5 >>
rect -1457 17854 -457 20462
rect -1457 17404 -1397 17854
rect -516 17404 -457 17854
rect -1457 14610 -457 17404
rect -1457 14160 -1397 14610
rect -516 14160 -457 14610
rect -1457 9996 -457 14160
rect 943 19476 1943 19536
rect 943 19026 1003 19476
rect 1884 19026 1943 19476
rect 943 16232 1943 19026
rect 943 15782 1003 16232
rect 1884 15782 1943 16232
rect 943 12988 1943 15782
rect 943 12538 1003 12988
rect 1884 12538 1943 12988
rect 943 12478 1943 12538
rect 2599 19476 3600 19536
rect 2599 19026 2659 19476
rect 3540 19026 3600 19476
rect 2599 16232 3600 19026
rect 2599 15782 2659 16232
rect 3540 15782 3600 16232
rect 2599 12988 3600 15782
rect 2599 12538 2659 12988
rect 3540 12538 3600 12988
rect 2599 12478 3600 12538
rect 4999 17854 5999 20462
rect 4999 17404 5059 17854
rect 5940 17404 5999 17854
rect 4999 14610 5999 17404
rect 4999 14160 5059 14610
rect 5940 14160 5999 14610
rect -1457 9546 -1397 9996
rect -516 9546 -457 9996
rect -1457 6752 -457 9546
rect -1457 6302 -1397 6752
rect -516 6302 -457 6752
rect -1457 2138 -457 6302
rect 943 11618 1943 11678
rect 943 11168 1003 11618
rect 1884 11168 1943 11618
rect 943 8374 1943 11168
rect 943 7924 1003 8374
rect 1884 7924 1943 8374
rect 943 5130 1943 7924
rect 943 4680 1003 5130
rect 1884 4680 1943 5130
rect 943 4620 1943 4680
rect 2599 11618 3600 11678
rect 2599 11168 2659 11618
rect 3540 11168 3600 11618
rect 2599 8374 3600 11168
rect 2599 7924 2659 8374
rect 3540 7924 3600 8374
rect 2599 5130 3600 7924
rect 2599 4680 2659 5130
rect 3540 4680 3600 5130
rect 2599 4620 3600 4680
rect 4999 9996 5999 14160
rect 4999 9546 5059 9996
rect 5940 9546 5999 9996
rect 4999 6752 5999 9546
rect 4999 6302 5059 6752
rect 5940 6302 5999 6752
rect -1457 1688 -1397 2138
rect -516 1688 -457 2138
rect -1457 -2476 -457 1688
rect 943 3760 1943 3820
rect 943 3310 1003 3760
rect 1884 3310 1943 3760
rect 943 516 1943 3310
rect 943 66 1003 516
rect 1884 66 1943 516
rect 943 6 1943 66
rect 2599 3760 3600 3820
rect 2599 3310 2659 3760
rect 3540 3310 3600 3760
rect 2599 516 3600 3310
rect 2599 66 2659 516
rect 3540 66 3600 516
rect 2599 6 3600 66
rect 4999 2138 5999 6302
rect 4999 1688 5059 2138
rect 5940 1688 5999 2138
rect -1457 -2926 -1397 -2476
rect -516 -2926 -457 -2476
rect -1457 -5468 -457 -2926
rect 943 -854 1943 -794
rect 943 -1304 1003 -854
rect 1884 -1304 1943 -854
rect 943 -2986 1943 -1304
rect 2599 -854 3600 -794
rect 2599 -1304 2659 -854
rect 3540 -1304 3600 -854
rect 2599 -2986 3600 -1304
rect 4999 -2476 5999 1688
rect 4999 -2926 5059 -2476
rect 5940 -2926 5999 -2476
rect -1457 -5918 -1397 -5468
rect -516 -5918 -457 -5468
rect -1457 -8460 -457 -5918
rect 943 -3846 1943 -3786
rect 943 -4296 1003 -3846
rect 1884 -4296 1943 -3846
rect 943 -5978 1943 -4296
rect 2599 -3846 3600 -3786
rect 2599 -4296 2659 -3846
rect 3540 -4296 3600 -3846
rect 2599 -5978 3600 -4296
rect 4999 -5468 5999 -2926
rect 4999 -5918 5059 -5468
rect 5940 -5918 5999 -5468
rect -1457 -8910 -1397 -8460
rect -516 -8910 -457 -8460
rect -1457 -9038 -457 -8910
rect 943 -6838 1943 -6778
rect 943 -7288 1003 -6838
rect 1884 -7288 1943 -6838
rect 943 -8970 1943 -7288
rect 2599 -6838 3600 -6778
rect 2599 -7288 2659 -6838
rect 3540 -7288 3600 -6838
rect 2599 -8970 3600 -7288
rect 4999 -8460 5999 -5918
rect 4999 -8910 5059 -8460
rect 5940 -8910 5999 -8460
rect 4999 -9038 5999 -8910
use cap_sw  cap_sw_0
timestamp 1696250317
transform 1 0 1419 0 1 17607
box -131 -40 1835 1868
use cap_sw  cap_sw_1
timestamp 1696250317
transform 1 0 1419 0 1 1891
box -131 -40 1835 1868
use cap_sw  cap_sw_2
timestamp 1696250317
transform 1 0 1419 0 1 9749
box -131 -40 1835 1868
use cap_sw  cap_sw_3
timestamp 1696250317
transform 1 0 1419 0 1 -8707
box -131 -40 1835 1868
use cap_sw  cap_sw_4
timestamp 1696250317
transform 1 0 1419 0 1 -2723
box -131 -40 1835 1868
use cap_sw  cap_sw_5
timestamp 1696250317
transform 1 0 1419 0 1 -5715
box -131 -40 1835 1868
use sky130_fd_pr__cap_mim_m3_1_H9ZJA7  sky130_fd_pr__cap_mim_m3_1_H9ZJA7_0
timestamp 1696250317
transform 0 -1 8384 -1 0 18440
box -686 -590 686 590
use sky130_fd_pr__cap_mim_m3_1_H9ZJA7  sky130_fd_pr__cap_mim_m3_1_H9ZJA7_1
timestamp 1696250317
transform 0 -1 4094 1 0 18440
box -686 -590 686 590
use sky130_fd_pr__cap_mim_m3_1_H9ZJA7  sky130_fd_pr__cap_mim_m3_1_H9ZJA7_2
timestamp 1696250317
transform 0 -1 4094 1 0 15196
box -686 -590 686 590
use sky130_fd_pr__cap_mim_m3_1_H9ZJA7  sky130_fd_pr__cap_mim_m3_1_H9ZJA7_3
timestamp 1696250317
transform 0 -1 8384 -1 0 15196
box -686 -590 686 590
use sky130_fd_pr__cap_mim_m3_1_H9ZJA7  sky130_fd_pr__cap_mim_m3_1_H9ZJA7_4
timestamp 1696250317
transform 0 -1 448 1 0 15196
box -686 -590 686 590
use sky130_fd_pr__cap_mim_m3_1_H9ZJA7  sky130_fd_pr__cap_mim_m3_1_H9ZJA7_5
timestamp 1696250317
transform 0 -1 -982 -1 0 15196
box -686 -590 686 590
use sky130_fd_pr__cap_mim_m3_1_H9ZJA7  sky130_fd_pr__cap_mim_m3_1_H9ZJA7_6
timestamp 1696250317
transform 0 -1 448 1 0 18440
box -686 -590 686 590
use sky130_fd_pr__cap_mim_m3_1_H9ZJA7  sky130_fd_pr__cap_mim_m3_1_H9ZJA7_7
timestamp 1696250317
transform 0 -1 -3842 -1 0 18440
box -686 -590 686 590
use sky130_fd_pr__cap_mim_m3_1_H9ZJA7  sky130_fd_pr__cap_mim_m3_1_H9ZJA7_8
timestamp 1696250317
transform 0 -1 4094 -1 0 16818
box -686 -590 686 590
use sky130_fd_pr__cap_mim_m3_1_H9ZJA7  sky130_fd_pr__cap_mim_m3_1_H9ZJA7_9
timestamp 1696250317
transform 0 -1 4094 -1 0 13574
box -686 -590 686 590
use sky130_fd_pr__cap_mim_m3_1_H9ZJA7  sky130_fd_pr__cap_mim_m3_1_H9ZJA7_10
timestamp 1696250317
transform 0 -1 8384 1 0 16818
box -686 -590 686 590
use sky130_fd_pr__cap_mim_m3_1_H9ZJA7  sky130_fd_pr__cap_mim_m3_1_H9ZJA7_11
timestamp 1696250317
transform 0 -1 8384 1 0 13574
box -686 -590 686 590
use sky130_fd_pr__cap_mim_m3_1_H9ZJA7  sky130_fd_pr__cap_mim_m3_1_H9ZJA7_12
timestamp 1696250317
transform 0 -1 448 -1 0 16818
box -686 -590 686 590
use sky130_fd_pr__cap_mim_m3_1_H9ZJA7  sky130_fd_pr__cap_mim_m3_1_H9ZJA7_13
timestamp 1696250317
transform 0 -1 -982 1 0 16818
box -686 -590 686 590
use sky130_fd_pr__cap_mim_m3_1_H9ZJA7  sky130_fd_pr__cap_mim_m3_1_H9ZJA7_14
timestamp 1696250317
transform 0 -1 -3842 1 0 13574
box -686 -590 686 590
use sky130_fd_pr__cap_mim_m3_1_H9ZJA7  sky130_fd_pr__cap_mim_m3_1_H9ZJA7_15
timestamp 1696250317
transform 0 -1 448 -1 0 13574
box -686 -590 686 590
use sky130_fd_pr__cap_mim_m3_1_H9ZJA7  sky130_fd_pr__cap_mim_m3_1_H9ZJA7_16
timestamp 1696250317
transform 0 -1 -982 -1 0 18440
box -686 -590 686 590
use sky130_fd_pr__cap_mim_m3_1_H9ZJA7  sky130_fd_pr__cap_mim_m3_1_H9ZJA7_17
timestamp 1696250317
transform 0 -1 -2412 1 0 18440
box -686 -590 686 590
use sky130_fd_pr__cap_mim_m3_1_H9ZJA7  sky130_fd_pr__cap_mim_m3_1_H9ZJA7_18
timestamp 1696250317
transform 0 -1 -3842 1 0 16818
box -686 -590 686 590
use sky130_fd_pr__cap_mim_m3_1_H9ZJA7  sky130_fd_pr__cap_mim_m3_1_H9ZJA7_19
timestamp 1696250317
transform 0 -1 -2412 -1 0 16818
box -686 -590 686 590
use sky130_fd_pr__cap_mim_m3_1_H9ZJA7  sky130_fd_pr__cap_mim_m3_1_H9ZJA7_20
timestamp 1696250317
transform 0 -1 -3842 -1 0 15196
box -686 -590 686 590
use sky130_fd_pr__cap_mim_m3_1_H9ZJA7  sky130_fd_pr__cap_mim_m3_1_H9ZJA7_21
timestamp 1696250317
transform 0 -1 -2412 1 0 15196
box -686 -590 686 590
use sky130_fd_pr__cap_mim_m3_1_H9ZJA7  sky130_fd_pr__cap_mim_m3_1_H9ZJA7_22
timestamp 1696250317
transform 0 -1 -982 1 0 13574
box -686 -590 686 590
use sky130_fd_pr__cap_mim_m3_1_H9ZJA7  sky130_fd_pr__cap_mim_m3_1_H9ZJA7_23
timestamp 1696250317
transform 0 -1 -2412 -1 0 13574
box -686 -590 686 590
use sky130_fd_pr__cap_mim_m3_1_H9ZJA7  sky130_fd_pr__cap_mim_m3_1_H9ZJA7_24
timestamp 1696250317
transform 0 -1 5524 -1 0 18440
box -686 -590 686 590
use sky130_fd_pr__cap_mim_m3_1_H9ZJA7  sky130_fd_pr__cap_mim_m3_1_H9ZJA7_25
timestamp 1696250317
transform 0 -1 6954 1 0 18440
box -686 -590 686 590
use sky130_fd_pr__cap_mim_m3_1_H9ZJA7  sky130_fd_pr__cap_mim_m3_1_H9ZJA7_26
timestamp 1696250317
transform 0 -1 5524 1 0 16818
box -686 -590 686 590
use sky130_fd_pr__cap_mim_m3_1_H9ZJA7  sky130_fd_pr__cap_mim_m3_1_H9ZJA7_27
timestamp 1696250317
transform 0 -1 6954 -1 0 16818
box -686 -590 686 590
use sky130_fd_pr__cap_mim_m3_1_H9ZJA7  sky130_fd_pr__cap_mim_m3_1_H9ZJA7_28
timestamp 1696250317
transform 0 -1 5524 -1 0 15196
box -686 -590 686 590
use sky130_fd_pr__cap_mim_m3_1_H9ZJA7  sky130_fd_pr__cap_mim_m3_1_H9ZJA7_29
timestamp 1696250317
transform 0 -1 6954 1 0 15196
box -686 -590 686 590
use sky130_fd_pr__cap_mim_m3_1_H9ZJA7  sky130_fd_pr__cap_mim_m3_1_H9ZJA7_30
timestamp 1696250317
transform 0 -1 5524 1 0 13574
box -686 -590 686 590
use sky130_fd_pr__cap_mim_m3_1_H9ZJA7  sky130_fd_pr__cap_mim_m3_1_H9ZJA7_31
timestamp 1696250317
transform 0 -1 6954 -1 0 13574
box -686 -590 686 590
use sky130_fd_pr__cap_mim_m3_1_H9ZJA7  sky130_fd_pr__cap_mim_m3_1_H9ZJA7_32
timestamp 1696250317
transform 0 -1 -3842 1 0 5716
box -686 -590 686 590
use sky130_fd_pr__cap_mim_m3_1_H9ZJA7  sky130_fd_pr__cap_mim_m3_1_H9ZJA7_33
timestamp 1696250317
transform 0 -1 -3842 -1 0 7338
box -686 -590 686 590
use sky130_fd_pr__cap_mim_m3_1_H9ZJA7  sky130_fd_pr__cap_mim_m3_1_H9ZJA7_34
timestamp 1696250317
transform 0 -1 -2412 -1 0 5716
box -686 -590 686 590
use sky130_fd_pr__cap_mim_m3_1_H9ZJA7  sky130_fd_pr__cap_mim_m3_1_H9ZJA7_35
timestamp 1696250317
transform 0 -1 -982 1 0 5716
box -686 -590 686 590
use sky130_fd_pr__cap_mim_m3_1_H9ZJA7  sky130_fd_pr__cap_mim_m3_1_H9ZJA7_36
timestamp 1696250317
transform 0 -1 -2412 1 0 7338
box -686 -590 686 590
use sky130_fd_pr__cap_mim_m3_1_H9ZJA7  sky130_fd_pr__cap_mim_m3_1_H9ZJA7_37
timestamp 1696250317
transform 0 -1 -982 -1 0 7338
box -686 -590 686 590
use sky130_fd_pr__cap_mim_m3_1_H9ZJA7  sky130_fd_pr__cap_mim_m3_1_H9ZJA7_38
timestamp 1696250317
transform 0 -1 448 -1 0 5716
box -686 -590 686 590
use sky130_fd_pr__cap_mim_m3_1_H9ZJA7  sky130_fd_pr__cap_mim_m3_1_H9ZJA7_39
timestamp 1696250317
transform 0 -1 448 1 0 7338
box -686 -590 686 590
use sky130_fd_pr__cap_mim_m3_1_H9ZJA7  sky130_fd_pr__cap_mim_m3_1_H9ZJA7_40
timestamp 1696250317
transform 0 -1 5524 1 0 5716
box -686 -590 686 590
use sky130_fd_pr__cap_mim_m3_1_H9ZJA7  sky130_fd_pr__cap_mim_m3_1_H9ZJA7_41
timestamp 1696250317
transform 0 -1 4094 -1 0 5716
box -686 -590 686 590
use sky130_fd_pr__cap_mim_m3_1_H9ZJA7  sky130_fd_pr__cap_mim_m3_1_H9ZJA7_42
timestamp 1696250317
transform 0 -1 5524 -1 0 7338
box -686 -590 686 590
use sky130_fd_pr__cap_mim_m3_1_H9ZJA7  sky130_fd_pr__cap_mim_m3_1_H9ZJA7_43
timestamp 1696250317
transform 0 -1 4094 1 0 7338
box -686 -590 686 590
use sky130_fd_pr__cap_mim_m3_1_H9ZJA7  sky130_fd_pr__cap_mim_m3_1_H9ZJA7_44
timestamp 1696250317
transform 0 -1 6954 -1 0 5716
box -686 -590 686 590
use sky130_fd_pr__cap_mim_m3_1_H9ZJA7  sky130_fd_pr__cap_mim_m3_1_H9ZJA7_45
timestamp 1696250317
transform 0 -1 8384 1 0 5716
box -686 -590 686 590
use sky130_fd_pr__cap_mim_m3_1_H9ZJA7  sky130_fd_pr__cap_mim_m3_1_H9ZJA7_46
timestamp 1696250317
transform 0 -1 6954 1 0 7338
box -686 -590 686 590
use sky130_fd_pr__cap_mim_m3_1_H9ZJA7  sky130_fd_pr__cap_mim_m3_1_H9ZJA7_47
timestamp 1696250317
transform 0 -1 8384 -1 0 7338
box -686 -590 686 590
use sky130_fd_pr__cap_mim_m3_1_H9ZJA7  sky130_fd_pr__cap_mim_m3_1_H9ZJA7_48
timestamp 1696250317
transform 0 -1 -3842 -1 0 2724
box -686 -590 686 590
use sky130_fd_pr__cap_mim_m3_1_H9ZJA7  sky130_fd_pr__cap_mim_m3_1_H9ZJA7_49
timestamp 1696250317
transform 0 -1 -3842 1 0 1102
box -686 -590 686 590
use sky130_fd_pr__cap_mim_m3_1_H9ZJA7  sky130_fd_pr__cap_mim_m3_1_H9ZJA7_50
timestamp 1696250317
transform 0 -1 -2412 1 0 2724
box -686 -590 686 590
use sky130_fd_pr__cap_mim_m3_1_H9ZJA7  sky130_fd_pr__cap_mim_m3_1_H9ZJA7_51
timestamp 1696250317
transform 0 -1 -2412 -1 0 1102
box -686 -590 686 590
use sky130_fd_pr__cap_mim_m3_1_H9ZJA7  sky130_fd_pr__cap_mim_m3_1_H9ZJA7_52
timestamp 1696250317
transform 0 -1 -982 -1 0 2724
box -686 -590 686 590
use sky130_fd_pr__cap_mim_m3_1_H9ZJA7  sky130_fd_pr__cap_mim_m3_1_H9ZJA7_53
timestamp 1696250317
transform 0 -1 -982 1 0 1102
box -686 -590 686 590
use sky130_fd_pr__cap_mim_m3_1_H9ZJA7  sky130_fd_pr__cap_mim_m3_1_H9ZJA7_54
timestamp 1696250317
transform 0 -1 448 1 0 2724
box -686 -590 686 590
use sky130_fd_pr__cap_mim_m3_1_H9ZJA7  sky130_fd_pr__cap_mim_m3_1_H9ZJA7_55
timestamp 1696250317
transform 0 -1 448 -1 0 1102
box -686 -590 686 590
use sky130_fd_pr__cap_mim_m3_1_H9ZJA7  sky130_fd_pr__cap_mim_m3_1_H9ZJA7_56
timestamp 1696250317
transform 0 -1 5524 -1 0 2724
box -686 -590 686 590
use sky130_fd_pr__cap_mim_m3_1_H9ZJA7  sky130_fd_pr__cap_mim_m3_1_H9ZJA7_57
timestamp 1696250317
transform 0 -1 4094 1 0 2724
box -686 -590 686 590
use sky130_fd_pr__cap_mim_m3_1_H9ZJA7  sky130_fd_pr__cap_mim_m3_1_H9ZJA7_58
timestamp 1696250317
transform 0 -1 5524 1 0 1102
box -686 -590 686 590
use sky130_fd_pr__cap_mim_m3_1_H9ZJA7  sky130_fd_pr__cap_mim_m3_1_H9ZJA7_59
timestamp 1696250317
transform 0 -1 4094 -1 0 1102
box -686 -590 686 590
use sky130_fd_pr__cap_mim_m3_1_H9ZJA7  sky130_fd_pr__cap_mim_m3_1_H9ZJA7_60
timestamp 1696250317
transform 0 -1 6954 1 0 2724
box -686 -590 686 590
use sky130_fd_pr__cap_mim_m3_1_H9ZJA7  sky130_fd_pr__cap_mim_m3_1_H9ZJA7_61
timestamp 1696250317
transform 0 -1 6954 -1 0 1102
box -686 -590 686 590
use sky130_fd_pr__cap_mim_m3_1_H9ZJA7  sky130_fd_pr__cap_mim_m3_1_H9ZJA7_62
timestamp 1696250317
transform 0 -1 8384 -1 0 2724
box -686 -590 686 590
use sky130_fd_pr__cap_mim_m3_1_H9ZJA7  sky130_fd_pr__cap_mim_m3_1_H9ZJA7_63
timestamp 1696250317
transform 0 -1 8384 1 0 1102
box -686 -590 686 590
use sky130_fd_pr__cap_mim_m3_1_H9ZJA7  sky130_fd_pr__cap_mim_m3_1_H9ZJA7_64
timestamp 1696250317
transform 0 -1 -982 -1 0 -4882
box -686 -590 686 590
use sky130_fd_pr__cap_mim_m3_1_H9ZJA7  sky130_fd_pr__cap_mim_m3_1_H9ZJA7_65
timestamp 1696250317
transform 0 -1 448 1 0 -4882
box -686 -590 686 590
use sky130_fd_pr__cap_mim_m3_1_H9ZJA7  sky130_fd_pr__cap_mim_m3_1_H9ZJA7_66
timestamp 1696250317
transform 0 -1 4094 1 0 -7874
box -686 -590 686 590
use sky130_fd_pr__cap_mim_m3_1_H9ZJA7  sky130_fd_pr__cap_mim_m3_1_H9ZJA7_68
timestamp 1696250317
transform 0 -1 448 1 0 -7874
box -686 -590 686 590
use sky130_fd_pr__cap_mim_m3_1_H9ZJA7  sky130_fd_pr__cap_mim_m3_1_H9ZJA7_70
timestamp 1696250317
transform 0 -1 5524 -1 0 -4882
box -686 -590 686 590
use sky130_fd_pr__cap_mim_m3_1_H9ZJA7  sky130_fd_pr__cap_mim_m3_1_H9ZJA7_71
timestamp 1696250317
transform 0 -1 4094 1 0 -4882
box -686 -590 686 590
use sky130_fd_pr__cap_mim_m3_1_H9ZJA7  sky130_fd_pr__cap_mim_m3_1_H9ZJA7_80
timestamp 1696250317
transform 0 -1 -3842 -1 0 -1890
box -686 -590 686 590
use sky130_fd_pr__cap_mim_m3_1_H9ZJA7  sky130_fd_pr__cap_mim_m3_1_H9ZJA7_82
timestamp 1696250317
transform 0 -1 -2412 1 0 -1890
box -686 -590 686 590
use sky130_fd_pr__cap_mim_m3_1_H9ZJA7  sky130_fd_pr__cap_mim_m3_1_H9ZJA7_84
timestamp 1696250317
transform 0 -1 -982 -1 0 -1890
box -686 -590 686 590
use sky130_fd_pr__cap_mim_m3_1_H9ZJA7  sky130_fd_pr__cap_mim_m3_1_H9ZJA7_86
timestamp 1696250317
transform 0 -1 448 1 0 -1890
box -686 -590 686 590
use sky130_fd_pr__cap_mim_m3_1_H9ZJA7  sky130_fd_pr__cap_mim_m3_1_H9ZJA7_88
timestamp 1696250317
transform 0 -1 5524 -1 0 -1890
box -686 -590 686 590
use sky130_fd_pr__cap_mim_m3_1_H9ZJA7  sky130_fd_pr__cap_mim_m3_1_H9ZJA7_89
timestamp 1696250317
transform 0 -1 4094 1 0 -1890
box -686 -590 686 590
use sky130_fd_pr__cap_mim_m3_1_H9ZJA7  sky130_fd_pr__cap_mim_m3_1_H9ZJA7_92
timestamp 1696250317
transform 0 -1 6954 1 0 -1890
box -686 -590 686 590
use sky130_fd_pr__cap_mim_m3_1_H9ZJA7  sky130_fd_pr__cap_mim_m3_1_H9ZJA7_94
timestamp 1696250317
transform 0 -1 8384 -1 0 -1890
box -686 -590 686 590
use sky130_fd_pr__cap_mim_m3_1_H9ZJA7  sky130_fd_pr__cap_mim_m3_1_H9ZJA7_96
timestamp 1696250317
transform 0 -1 -3842 -1 0 10582
box -686 -590 686 590
use sky130_fd_pr__cap_mim_m3_1_H9ZJA7  sky130_fd_pr__cap_mim_m3_1_H9ZJA7_97
timestamp 1696250317
transform 0 -1 -3842 1 0 8960
box -686 -590 686 590
use sky130_fd_pr__cap_mim_m3_1_H9ZJA7  sky130_fd_pr__cap_mim_m3_1_H9ZJA7_98
timestamp 1696250317
transform 0 -1 -2412 1 0 10582
box -686 -590 686 590
use sky130_fd_pr__cap_mim_m3_1_H9ZJA7  sky130_fd_pr__cap_mim_m3_1_H9ZJA7_99
timestamp 1696250317
transform 0 -1 -2412 -1 0 8960
box -686 -590 686 590
use sky130_fd_pr__cap_mim_m3_1_H9ZJA7  sky130_fd_pr__cap_mim_m3_1_H9ZJA7_100
timestamp 1696250317
transform 0 -1 -982 -1 0 10582
box -686 -590 686 590
use sky130_fd_pr__cap_mim_m3_1_H9ZJA7  sky130_fd_pr__cap_mim_m3_1_H9ZJA7_101
timestamp 1696250317
transform 0 -1 -982 1 0 8960
box -686 -590 686 590
use sky130_fd_pr__cap_mim_m3_1_H9ZJA7  sky130_fd_pr__cap_mim_m3_1_H9ZJA7_102
timestamp 1696250317
transform 0 -1 448 1 0 10582
box -686 -590 686 590
use sky130_fd_pr__cap_mim_m3_1_H9ZJA7  sky130_fd_pr__cap_mim_m3_1_H9ZJA7_103
timestamp 1696250317
transform 0 -1 448 -1 0 8960
box -686 -590 686 590
use sky130_fd_pr__cap_mim_m3_1_H9ZJA7  sky130_fd_pr__cap_mim_m3_1_H9ZJA7_104
timestamp 1696250317
transform 0 -1 5524 -1 0 10582
box -686 -590 686 590
use sky130_fd_pr__cap_mim_m3_1_H9ZJA7  sky130_fd_pr__cap_mim_m3_1_H9ZJA7_105
timestamp 1696250317
transform 0 -1 4094 1 0 10582
box -686 -590 686 590
use sky130_fd_pr__cap_mim_m3_1_H9ZJA7  sky130_fd_pr__cap_mim_m3_1_H9ZJA7_106
timestamp 1696250317
transform 0 -1 5524 1 0 8960
box -686 -590 686 590
use sky130_fd_pr__cap_mim_m3_1_H9ZJA7  sky130_fd_pr__cap_mim_m3_1_H9ZJA7_107
timestamp 1696250317
transform 0 -1 4094 -1 0 8960
box -686 -590 686 590
use sky130_fd_pr__cap_mim_m3_1_H9ZJA7  sky130_fd_pr__cap_mim_m3_1_H9ZJA7_108
timestamp 1696250317
transform 0 -1 6954 1 0 10582
box -686 -590 686 590
use sky130_fd_pr__cap_mim_m3_1_H9ZJA7  sky130_fd_pr__cap_mim_m3_1_H9ZJA7_109
timestamp 1696250317
transform 0 -1 6954 -1 0 8960
box -686 -590 686 590
use sky130_fd_pr__cap_mim_m3_1_H9ZJA7  sky130_fd_pr__cap_mim_m3_1_H9ZJA7_110
timestamp 1696250317
transform 0 -1 8384 -1 0 10582
box -686 -590 686 590
use sky130_fd_pr__cap_mim_m3_1_H9ZJA7  sky130_fd_pr__cap_mim_m3_1_H9ZJA7_111
timestamp 1696250317
transform 0 -1 8384 1 0 8960
box -686 -590 686 590
<< labels >>
flabel metal1 2201 17434 2299 17746 0 FreeSans 320 0 0 0 tune[5]
port 1 nsew
flabel metal5 -1457 17854 -457 20462 0 FreeSans 1600 0 0 0 vn_cap
port 8 nsew
flabel metal1 2201 9576 2299 9888 0 FreeSans 320 0 0 0 tune[4]
port 2 nsew
flabel locali 2410 9578 2507 9779 0 FreeSans 320 0 0 0 vss_cap
port 0 nsew
flabel locali 2410 17436 2507 17637 0 FreeSans 320 0 0 0 vss_cap
port 0 nsew
flabel locali 2410 1720 2507 1921 0 FreeSans 320 0 0 0 vss_cap
port 0 nsew
flabel locali 2410 -2894 2507 -2693 0 FreeSans 320 0 0 0 vss_cap
port 0 nsew
flabel metal1 2201 -2896 2299 -2584 0 FreeSans 320 0 0 0 tune[2]
port 4 nsew
flabel metal1 2201 1718 2299 2030 0 FreeSans 320 0 0 0 tune[3]
port 3 nsew
flabel locali 2410 -5886 2507 -5685 0 FreeSans 320 0 0 0 vss_cap
port 0 nsew
flabel metal1 2201 -5888 2299 -5576 0 FreeSans 320 0 0 0 tune[1]
port 5 nsew
flabel locali 2410 -8878 2507 -8677 0 FreeSans 320 0 0 0 vss_cap
port 0 nsew
flabel metal1 2201 -8880 2299 -8568 0 FreeSans 320 0 0 0 tune[0]
port 6 nsew
flabel metal5 4999 17854 5999 20462 0 FreeSans 1600 0 0 0 vp_cap
port 7 nsew
<< end >>
