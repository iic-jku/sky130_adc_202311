magic
tech sky130A
magscale 1 2
timestamp 1699972208
<< nwell >>
rect -532 261 -319 582
rect 123 395 1978 582
rect 2435 261 2650 582
<< pwell >>
rect -532 21 2648 203
<< psubdiff >>
rect -453 179 -409 203
rect -453 37 -409 61
rect 2525 179 2569 203
rect 2525 37 2569 61
<< nsubdiff >>
rect -493 384 -469 454
rect -371 384 -347 454
rect 2468 384 2492 454
rect 2590 384 2614 454
<< psubdiffcont >>
rect -453 61 -409 179
rect 2525 61 2569 179
<< nsubdiffcont >>
rect -469 384 -371 454
rect 2492 384 2590 454
<< locali >>
rect -453 454 -409 535
rect 2525 454 2569 530
rect -493 384 -469 454
rect -371 384 -347 454
rect 2468 384 2492 454
rect 2590 384 2614 454
rect -88 215 19 265
rect 2136 215 2180 265
rect -453 179 -409 203
rect -453 17 -409 61
rect 2525 179 2569 203
rect -302 17 -252 57
rect 2374 17 2424 51
rect 2525 17 2569 61
rect -409 -17 -319 17
rect 2412 -17 2525 17
<< viali >>
rect -453 535 -409 569
rect 2525 530 2569 564
rect 37 221 79 255
rect 159 216 201 250
rect 356 221 398 255
rect 499 224 541 258
rect 617 217 659 251
rect 821 215 863 249
rect 959 224 1001 258
rect 1115 224 1157 258
rect 1256 215 1293 255
rect 1456 216 1498 250
rect 1575 224 1617 258
rect 1721 215 1758 255
rect 1918 221 1960 255
rect 2034 221 2076 255
rect -453 -17 -409 17
rect 2525 -17 2569 17
<< metal1 >>
rect -532 569 2648 592
rect -532 535 -453 569
rect -409 564 2648 569
rect -409 535 2525 564
rect -532 530 2525 535
rect 2569 530 2648 564
rect -532 496 2648 530
rect 26 266 98 272
rect 26 206 32 266
rect 92 206 98 266
rect 26 199 98 206
rect 141 265 213 271
rect 141 205 147 265
rect 207 205 213 265
rect 141 199 213 205
rect 348 265 443 271
rect 348 255 377 265
rect 348 221 356 255
rect 348 205 377 221
rect 437 205 443 265
rect 601 265 673 271
rect 348 199 443 205
rect 486 258 558 264
rect 486 198 492 258
rect 552 198 558 258
rect 601 205 607 265
rect 667 205 673 265
rect 601 199 673 205
rect 809 265 903 271
rect 809 249 837 265
rect 809 215 821 249
rect 809 205 837 215
rect 897 205 903 265
rect 1213 265 1303 271
rect 809 199 903 205
rect 946 258 1018 264
rect 486 192 558 198
rect 946 198 952 258
rect 1012 198 1018 258
rect 946 192 1018 198
rect 1098 258 1170 264
rect 1098 198 1104 258
rect 1164 198 1170 258
rect 1213 205 1219 265
rect 1279 255 1303 265
rect 1293 215 1303 255
rect 1279 205 1303 215
rect 1213 199 1303 205
rect 1443 265 1515 271
rect 1443 205 1449 265
rect 1509 205 1515 265
rect 1673 265 1767 271
rect 1443 199 1515 205
rect 1558 258 1630 264
rect 1098 192 1170 198
rect 1558 198 1564 258
rect 1624 198 1630 258
rect 1673 205 1679 265
rect 1739 255 1767 265
rect 1758 215 1767 255
rect 1739 205 1767 215
rect 1673 199 1767 205
rect 1903 265 1975 271
rect 1903 205 1909 265
rect 1969 205 1975 265
rect 1903 199 1975 205
rect 2018 265 2090 271
rect 2018 205 2025 265
rect 2085 205 2090 265
rect 2018 199 2090 205
rect 1558 192 1630 198
rect -532 31 2648 48
rect -532 30 2024 31
rect -532 17 32 30
rect -532 -17 -453 17
rect -409 -17 32 17
rect -532 -30 32 -17
rect 92 -29 2024 30
rect 2084 17 2648 31
rect 2084 -17 2525 17
rect 2569 -17 2648 17
rect 2084 -29 2648 -17
rect 92 -30 2648 -29
rect -532 -48 2648 -30
<< via1 >>
rect 32 255 92 266
rect 32 221 37 255
rect 37 221 79 255
rect 79 221 92 255
rect 32 206 92 221
rect 147 250 207 265
rect 147 216 159 250
rect 159 216 201 250
rect 201 216 207 250
rect 147 205 207 216
rect 377 255 437 265
rect 377 221 398 255
rect 398 221 437 255
rect 377 205 437 221
rect 492 224 499 258
rect 499 224 541 258
rect 541 224 552 258
rect 492 198 552 224
rect 607 251 667 265
rect 607 217 617 251
rect 617 217 659 251
rect 659 217 667 251
rect 607 205 667 217
rect 837 249 897 265
rect 837 215 863 249
rect 863 215 897 249
rect 837 205 897 215
rect 952 224 959 258
rect 959 224 1001 258
rect 1001 224 1012 258
rect 952 198 1012 224
rect 1104 224 1115 258
rect 1115 224 1157 258
rect 1157 224 1164 258
rect 1104 198 1164 224
rect 1219 255 1279 265
rect 1219 215 1256 255
rect 1256 215 1279 255
rect 1219 205 1279 215
rect 1449 250 1509 265
rect 1449 216 1456 250
rect 1456 216 1498 250
rect 1498 216 1509 250
rect 1449 205 1509 216
rect 1564 224 1575 258
rect 1575 224 1617 258
rect 1617 224 1624 258
rect 1564 198 1624 224
rect 1679 255 1739 265
rect 1679 215 1721 255
rect 1721 215 1739 255
rect 1679 205 1739 215
rect 1909 255 1969 265
rect 1909 221 1918 255
rect 1918 221 1960 255
rect 1960 221 1969 255
rect 1909 205 1969 221
rect 2025 255 2085 265
rect 2025 221 2034 255
rect 2034 221 2076 255
rect 2076 221 2085 255
rect 2025 205 2085 221
rect 32 -30 92 30
rect 2024 -29 2084 31
<< metal2 >>
rect 141 922 213 1544
rect 141 838 147 922
rect 207 838 213 922
rect 26 266 98 272
rect 26 206 32 266
rect 92 206 98 266
rect 26 30 98 206
rect 141 265 213 838
rect 141 205 147 265
rect 207 205 213 265
rect 371 730 443 1544
rect 371 646 377 730
rect 437 646 443 730
rect 371 265 443 646
rect 141 199 213 205
rect 26 -30 32 30
rect 92 -30 98 30
rect 26 -847 98 -30
rect 256 -847 328 264
rect 371 205 377 265
rect 437 205 443 265
rect 601 1114 673 1544
rect 601 1030 607 1114
rect 667 1030 673 1114
rect 601 265 673 1030
rect 371 199 443 205
rect 486 258 558 264
rect 486 198 492 258
rect 552 198 558 258
rect 601 205 607 265
rect 667 205 673 265
rect 831 730 903 1544
rect 831 646 837 730
rect 897 646 903 730
rect 831 265 903 646
rect 601 199 673 205
rect 486 -102 558 198
rect 486 -186 492 -102
rect 552 -186 558 -102
rect 486 -847 558 -186
rect 716 -847 788 264
rect 831 205 837 265
rect 897 205 903 265
rect 1213 730 1285 1544
rect 1213 646 1219 730
rect 1279 646 1285 730
rect 1213 265 1285 646
rect 831 199 903 205
rect 946 258 1018 264
rect 946 198 952 258
rect 1012 198 1018 258
rect 946 -294 1018 198
rect 946 -378 952 -294
rect 1012 -378 1018 -294
rect 946 -847 1018 -378
rect 1098 258 1170 264
rect 1098 198 1104 258
rect 1164 198 1170 258
rect 1213 205 1219 265
rect 1279 205 1285 265
rect 1443 1306 1515 1544
rect 1443 1222 1449 1306
rect 1509 1222 1515 1306
rect 1443 265 1515 1222
rect 1213 199 1285 205
rect 1098 -486 1170 198
rect 1098 -570 1104 -486
rect 1164 -570 1170 -486
rect 1098 -847 1170 -570
rect 1328 -847 1400 264
rect 1443 205 1449 265
rect 1509 205 1515 265
rect 1673 730 1745 1544
rect 1673 646 1679 730
rect 1739 646 1745 730
rect 1673 265 1745 646
rect 1443 199 1515 205
rect 1558 258 1630 264
rect 1558 198 1564 258
rect 1624 198 1630 258
rect 1673 205 1679 265
rect 1739 205 1745 265
rect 1903 1498 1975 1544
rect 1903 1414 1909 1498
rect 1969 1414 1975 1498
rect 1903 265 1975 1414
rect 1673 199 1745 205
rect 1558 -678 1630 198
rect 1558 -762 1564 -678
rect 1624 -762 1630 -678
rect 1558 -847 1630 -762
rect 1788 -847 1860 264
rect 1903 205 1909 265
rect 1969 205 1975 265
rect 1903 199 1975 205
rect 2018 265 2090 271
rect 2018 205 2025 265
rect 2085 205 2090 265
rect 2018 31 2090 205
rect 2018 -29 2024 31
rect 2084 -29 2090 31
rect 2018 -847 2090 -29
<< via2 >>
rect 147 838 207 922
rect 377 646 437 730
rect 607 1030 667 1114
rect 837 646 897 730
rect 492 -186 552 -102
rect 1219 646 1279 730
rect 952 -378 1012 -294
rect 1449 1222 1509 1306
rect 1104 -570 1164 -486
rect 1679 646 1739 730
rect 1909 1414 1969 1498
rect 1564 -762 1624 -678
<< metal3 >>
rect -532 1498 2648 1504
rect -532 1414 1909 1498
rect 1969 1414 2648 1498
rect -532 1408 2648 1414
rect -532 1306 2648 1312
rect -532 1222 1449 1306
rect 1509 1222 2648 1306
rect -532 1216 2648 1222
rect -532 1114 2648 1120
rect -532 1030 607 1114
rect 667 1030 2648 1114
rect -532 1024 2648 1030
rect -532 922 2648 928
rect -532 838 147 922
rect 207 838 2648 922
rect -532 832 2648 838
rect -532 730 2648 736
rect -532 646 377 730
rect 437 646 837 730
rect 897 646 1219 730
rect 1279 646 1679 730
rect 1739 646 2648 730
rect -532 640 2648 646
rect -532 -102 2648 -96
rect -532 -186 492 -102
rect 552 -186 2648 -102
rect -532 -192 2648 -186
rect -532 -294 2648 -288
rect -532 -378 952 -294
rect 1012 -378 2648 -294
rect -532 -384 2648 -378
rect -532 -486 2648 -480
rect -532 -570 1104 -486
rect 1164 -570 2648 -486
rect -532 -576 2648 -570
rect -532 -678 2648 -672
rect -532 -762 1564 -678
rect 1624 -762 2648 -678
rect -532 -768 2648 -762
use sky130_fd_sc_hd__and2_1  sky130_fd_sc_hd__and2_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform -1 0 141 0 1 0
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  sky130_fd_sc_hd__and2_1_1
timestamp 1694700623
transform -1 0 601 0 1 0
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  sky130_fd_sc_hd__and2_1_2
timestamp 1694700623
transform 1 0 1521 0 1 0
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  sky130_fd_sc_hd__and2_1_3
timestamp 1694700623
transform -1 0 1061 0 1 0
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  sky130_fd_sc_hd__and2_1_4
timestamp 1694700623
transform 1 0 1061 0 1 0
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  sky130_fd_sc_hd__and2_1_5
timestamp 1694700623
transform 1 0 1981 0 1 0
box -38 -48 498 592
<< labels >>
flabel metal3 1975 640 2648 736 0 FreeSans 320 0 0 0 in_gc
port 2 nsew
flabel metal3 1975 832 2648 928 0 FreeSans 320 0 0 0 out_gc[0]
port 3 nsew
flabel metal3 1975 1024 2648 1120 0 FreeSans 320 0 0 0 out_gc[1]
port 4 nsew
flabel metal3 1975 1408 2648 1504 0 FreeSans 320 0 0 0 out_gc[3]
port 6 nsew
flabel metal3 1975 -192 2648 -96 0 FreeSans 320 0 0 0 en_gc[0]
port 7 nsew
flabel metal3 1975 -384 2648 -288 0 FreeSans 320 0 0 0 en_gc[1]
port 8 nsew
flabel metal3 1975 -576 2648 -480 0 FreeSans 320 0 0 0 en_gc[2]
port 9 nsew
flabel metal3 1975 -768 2648 -672 0 FreeSans 320 0 0 0 en_gc[3]
port 10 nsew
flabel metal3 1975 1216 2648 1312 0 FreeSans 320 0 0 0 out_gc[2]
port 5 nsew
flabel metal1 -532 496 2648 592 0 FreeSans 320 0 0 0 vdd_gc
port 11 nsew
flabel metal1 -532 -48 2648 48 0 FreeSans 320 0 0 0 vss_gc
port 0 nsew
<< end >>
