magic
tech sky130A
magscale 1 2
timestamp 1697705955
<< metal1 >>
rect 1721 21 1769 23
rect 2105 21 2153 23
rect 1719 15 1771 21
rect 1719 -91 1771 -85
rect 2103 15 2155 21
rect 2103 -91 2155 -85
rect 1721 -94 1769 -91
rect 2105 -94 2153 -91
rect 427 -123 475 -121
rect 811 -123 859 -121
rect 425 -129 477 -123
rect 425 -235 477 -229
rect 809 -129 861 -123
rect 809 -235 861 -229
rect 427 -238 475 -235
rect 811 -238 859 -235
<< via1 >>
rect 1719 -85 1771 15
rect 2103 -85 2155 15
rect 425 -229 477 -129
rect 809 -229 861 -129
<< metal2 >>
rect 1719 15 1771 21
rect 1717 -83 1719 13
rect 2103 15 2155 21
rect 1771 -83 1773 13
rect 2101 -83 2103 13
rect 1719 -91 1771 -85
rect 2155 -83 2157 13
rect 2103 -91 2155 -85
rect 425 -129 477 -123
rect 423 -227 425 -131
rect 809 -129 861 -123
rect 477 -227 479 -131
rect 807 -227 809 -131
rect 425 -235 477 -229
rect 861 -227 863 -131
rect 809 -235 861 -229
use osc_nfet_w15_nf4  osc_nfet_w15_nf4_0
timestamp 1697705955
transform 1 0 130 0 1 227
box -134 -465 1160 1732
use osc_nfet_w15_nf4  osc_nfet_w15_nf4_1
timestamp 1697705955
transform 1 0 1424 0 1 227
box -134 -465 1160 1732
<< end >>
