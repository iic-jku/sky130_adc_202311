magic
tech sky130A
magscale 1 2
timestamp 1699571430
<< viali >>
rect 18061 77469 18095 77503
rect 16957 77333 16991 77367
rect 17233 77333 17267 77367
rect 18245 77333 18279 77367
rect 17141 76925 17175 76959
rect 17417 76925 17451 76959
rect 17693 76925 17727 76959
rect 13921 76789 13955 76823
rect 14289 76789 14323 76823
rect 14657 76789 14691 76823
rect 15945 76789 15979 76823
rect 16221 76789 16255 76823
rect 17141 76585 17175 76619
rect 17509 76585 17543 76619
rect 17877 76585 17911 76619
rect 18245 76585 18279 76619
rect 7757 76449 7791 76483
rect 7849 76381 7883 76415
rect 8033 76381 8067 76415
rect 14933 76381 14967 76415
rect 8493 76313 8527 76347
rect 11621 76313 11655 76347
rect 15178 76313 15212 76347
rect 7205 76245 7239 76279
rect 11253 76245 11287 76279
rect 11713 76245 11747 76279
rect 16313 76245 16347 76279
rect 7573 75973 7607 76007
rect 8769 75973 8803 76007
rect 3985 75905 4019 75939
rect 4252 75905 4286 75939
rect 6929 75905 6963 75939
rect 7113 75905 7147 75939
rect 14105 75905 14139 75939
rect 14197 75905 14231 75939
rect 6837 75837 6871 75871
rect 14381 75837 14415 75871
rect 5365 75769 5399 75803
rect 8401 75701 8435 75735
rect 8861 75701 8895 75735
rect 9229 75701 9263 75735
rect 13737 75701 13771 75735
rect 15209 75429 15243 75463
rect 5733 75361 5767 75395
rect 5549 75293 5583 75327
rect 7573 75293 7607 75327
rect 15393 75293 15427 75327
rect 18061 75293 18095 75327
rect 4997 75225 5031 75259
rect 5089 75157 5123 75191
rect 5457 75157 5491 75191
rect 6193 75157 6227 75191
rect 6561 75157 6595 75191
rect 6837 75157 6871 75191
rect 7205 75157 7239 75191
rect 7757 75157 7791 75191
rect 8125 75157 8159 75191
rect 8493 75157 8527 75191
rect 9137 75157 9171 75191
rect 18245 75157 18279 75191
rect 4721 74953 4755 74987
rect 16221 74953 16255 74987
rect 5089 74885 5123 74919
rect 5181 74817 5215 74851
rect 6653 74817 6687 74851
rect 14841 74817 14875 74851
rect 15108 74817 15142 74851
rect 16865 74817 16899 74851
rect 5273 74749 5307 74783
rect 6745 74613 6779 74647
rect 17049 74613 17083 74647
rect 12081 74409 12115 74443
rect 12725 74273 12759 74307
rect 14289 74205 14323 74239
rect 12541 74137 12575 74171
rect 14534 74137 14568 74171
rect 15945 74137 15979 74171
rect 16313 74137 16347 74171
rect 12449 74069 12483 74103
rect 13645 74069 13679 74103
rect 15669 74069 15703 74103
rect 7297 73865 7331 73899
rect 7665 73729 7699 73763
rect 7757 73729 7791 73763
rect 18061 73729 18095 73763
rect 7941 73661 7975 73695
rect 18245 73525 18279 73559
rect 6653 73185 6687 73219
rect 9137 73185 9171 73219
rect 6898 73049 6932 73083
rect 8309 73049 8343 73083
rect 5549 72981 5583 73015
rect 5917 72981 5951 73015
rect 6285 72981 6319 73015
rect 8033 72981 8067 73015
rect 13185 72641 13219 72675
rect 13277 72573 13311 72607
rect 13461 72573 13495 72607
rect 12817 72437 12851 72471
rect 17049 72233 17083 72267
rect 17233 72029 17267 72063
rect 3065 71553 3099 71587
rect 3332 71553 3366 71587
rect 18061 71553 18095 71587
rect 4445 71349 4479 71383
rect 18245 71349 18279 71383
rect 10517 71077 10551 71111
rect 6009 71009 6043 71043
rect 9137 70941 9171 70975
rect 15485 70941 15519 70975
rect 6276 70873 6310 70907
rect 9382 70873 9416 70907
rect 15752 70873 15786 70907
rect 7389 70805 7423 70839
rect 16865 70805 16899 70839
rect 2053 69989 2087 70023
rect 2513 69921 2547 69955
rect 15301 69921 15335 69955
rect 3985 69853 4019 69887
rect 7113 69853 7147 69887
rect 9137 69853 9171 69887
rect 9413 69853 9447 69887
rect 15025 69853 15059 69887
rect 18061 69853 18095 69887
rect 2605 69785 2639 69819
rect 7358 69785 7392 69819
rect 2513 69717 2547 69751
rect 3065 69717 3099 69751
rect 3433 69717 3467 69751
rect 4169 69717 4203 69751
rect 4629 69717 4663 69751
rect 4997 69717 5031 69751
rect 8493 69717 8527 69751
rect 18245 69717 18279 69751
rect 9934 69445 9968 69479
rect 9689 69377 9723 69411
rect 11069 69173 11103 69207
rect 9137 68833 9171 68867
rect 14289 68765 14323 68799
rect 9404 68697 9438 68731
rect 14556 68697 14590 68731
rect 10517 68629 10551 68663
rect 15669 68629 15703 68663
rect 12449 67813 12483 67847
rect 18245 67813 18279 67847
rect 12633 67677 12667 67711
rect 18061 67677 18095 67711
rect 12081 67609 12115 67643
rect 7941 67201 7975 67235
rect 17969 67201 18003 67235
rect 17325 67133 17359 67167
rect 18061 67133 18095 67167
rect 18153 67133 18187 67167
rect 8125 66997 8159 67031
rect 17601 66997 17635 67031
rect 13820 66181 13854 66215
rect 17969 66181 18003 66215
rect 13553 66113 13587 66147
rect 17785 66113 17819 66147
rect 18061 66045 18095 66079
rect 14933 65909 14967 65943
rect 17509 65909 17543 65943
rect 4077 65637 4111 65671
rect 18245 65637 18279 65671
rect 4629 65569 4663 65603
rect 11805 65501 11839 65535
rect 11897 65501 11931 65535
rect 12081 65501 12115 65535
rect 18061 65501 18095 65535
rect 4353 65433 4387 65467
rect 11253 65433 11287 65467
rect 12541 65433 12575 65467
rect 4537 65365 4571 65399
rect 7941 65161 7975 65195
rect 14381 65161 14415 65195
rect 13268 65093 13302 65127
rect 8309 65025 8343 65059
rect 18153 65025 18187 65059
rect 8401 64957 8435 64991
rect 8585 64957 8619 64991
rect 13001 64957 13035 64991
rect 18337 64889 18371 64923
rect 2605 64413 2639 64447
rect 11805 64413 11839 64447
rect 12050 64345 12084 64379
rect 2421 64277 2455 64311
rect 13185 64277 13219 64311
rect 12265 63937 12299 63971
rect 18061 63937 18095 63971
rect 12357 63869 12391 63903
rect 12541 63869 12575 63903
rect 11897 63801 11931 63835
rect 10701 63733 10735 63767
rect 11069 63733 11103 63767
rect 12909 63733 12943 63767
rect 13277 63733 13311 63767
rect 13645 63733 13679 63767
rect 18245 63733 18279 63767
rect 16313 63461 16347 63495
rect 14289 63325 14323 63359
rect 16497 63325 16531 63359
rect 6285 63257 6319 63291
rect 6377 63189 6411 63223
rect 14473 63189 14507 63223
rect 7941 62985 7975 63019
rect 6561 62849 6595 62883
rect 6817 62849 6851 62883
rect 5641 62781 5675 62815
rect 5917 62781 5951 62815
rect 8401 62645 8435 62679
rect 8769 62645 8803 62679
rect 18061 62237 18095 62271
rect 4261 62169 4295 62203
rect 4353 62101 4387 62135
rect 18245 62101 18279 62135
rect 11713 61897 11747 61931
rect 12081 61829 12115 61863
rect 12173 61693 12207 61727
rect 12265 61693 12299 61727
rect 15945 61149 15979 61183
rect 15669 61081 15703 61115
rect 16212 61081 16246 61115
rect 17601 61081 17635 61115
rect 17325 61013 17359 61047
rect 9505 60741 9539 60775
rect 6561 60673 6595 60707
rect 6817 60673 6851 60707
rect 8309 60673 8343 60707
rect 8677 60673 8711 60707
rect 5917 60605 5951 60639
rect 9413 60605 9447 60639
rect 9597 60605 9631 60639
rect 7941 60469 7975 60503
rect 9045 60469 9079 60503
rect 16129 60265 16163 60299
rect 9137 60197 9171 60231
rect 15669 60197 15703 60231
rect 8217 60129 8251 60163
rect 9781 60129 9815 60163
rect 16589 60129 16623 60163
rect 16681 60129 16715 60163
rect 8033 60061 8067 60095
rect 14289 60061 14323 60095
rect 18061 60061 18095 60095
rect 7941 59993 7975 60027
rect 9505 59993 9539 60027
rect 14556 59993 14590 60027
rect 7573 59925 7607 59959
rect 9597 59925 9631 59959
rect 16497 59925 16531 59959
rect 18245 59925 18279 59959
rect 4629 59721 4663 59755
rect 3249 59585 3283 59619
rect 3516 59585 3550 59619
rect 2237 59517 2271 59551
rect 2605 59517 2639 59551
rect 2973 59517 3007 59551
rect 4997 59381 5031 59415
rect 5273 59381 5307 59415
rect 15209 59041 15243 59075
rect 15393 59041 15427 59075
rect 7297 58973 7331 59007
rect 7573 58973 7607 59007
rect 15301 58905 15335 58939
rect 13737 58837 13771 58871
rect 14381 58837 14415 58871
rect 14823 58837 14857 58871
rect 15761 58837 15795 58871
rect 18061 58497 18095 58531
rect 18245 58293 18279 58327
rect 17325 57545 17359 57579
rect 16957 57477 16991 57511
rect 17693 57477 17727 57511
rect 2789 57409 2823 57443
rect 3056 57409 3090 57443
rect 15209 57409 15243 57443
rect 2513 57341 2547 57375
rect 17785 57341 17819 57375
rect 17877 57341 17911 57375
rect 4169 57205 4203 57239
rect 15025 57205 15059 57239
rect 1685 56933 1719 56967
rect 2237 56865 2271 56899
rect 1961 56797 1995 56831
rect 2145 56661 2179 56695
rect 2697 56661 2731 56695
rect 3402 56389 3436 56423
rect 2513 56321 2547 56355
rect 3157 56321 3191 56355
rect 18061 56321 18095 56355
rect 12449 56253 12483 56287
rect 12725 56253 12759 56287
rect 2789 56185 2823 56219
rect 2329 56117 2363 56151
rect 4537 56117 4571 56151
rect 18245 56117 18279 56151
rect 11805 55777 11839 55811
rect 1685 55709 1719 55743
rect 11529 55709 11563 55743
rect 1930 55641 1964 55675
rect 3065 55573 3099 55607
rect 3617 55369 3651 55403
rect 4077 55369 4111 55403
rect 4445 55369 4479 55403
rect 4813 55369 4847 55403
rect 5181 55369 5215 55403
rect 16865 55369 16899 55403
rect 17325 55301 17359 55335
rect 2237 55233 2271 55267
rect 2504 55233 2538 55267
rect 5549 55233 5583 55267
rect 5733 55233 5767 55267
rect 6561 55233 6595 55267
rect 17233 55233 17267 55267
rect 17417 55165 17451 55199
rect 18061 54621 18095 54655
rect 18245 54485 18279 54519
rect 9965 54145 9999 54179
rect 10609 54145 10643 54179
rect 10701 54145 10735 54179
rect 13001 54145 13035 54179
rect 10885 54077 10919 54111
rect 10241 54009 10275 54043
rect 12817 53941 12851 53975
rect 13737 53193 13771 53227
rect 1961 53125 1995 53159
rect 2145 53125 2179 53159
rect 9965 53125 9999 53159
rect 8585 53057 8619 53091
rect 12624 53057 12658 53091
rect 2237 52989 2271 53023
rect 9873 52989 9907 53023
rect 10057 52989 10091 53023
rect 12357 52989 12391 53023
rect 8769 52921 8803 52955
rect 1685 52853 1719 52887
rect 9505 52853 9539 52887
rect 18245 52581 18279 52615
rect 14289 52513 14323 52547
rect 14556 52445 14590 52479
rect 18061 52445 18095 52479
rect 15669 52309 15703 52343
rect 18061 52105 18095 52139
rect 18245 51969 18279 52003
rect 5365 51561 5399 51595
rect 3985 51425 4019 51459
rect 10425 51425 10459 51459
rect 14565 51425 14599 51459
rect 8585 51357 8619 51391
rect 14289 51357 14323 51391
rect 4252 51289 4286 51323
rect 10692 51289 10726 51323
rect 8401 51221 8435 51255
rect 11805 51221 11839 51255
rect 8401 50881 8435 50915
rect 8677 50881 8711 50915
rect 9312 50881 9346 50915
rect 18061 50881 18095 50915
rect 9045 50813 9079 50847
rect 10425 50677 10459 50711
rect 10701 50677 10735 50711
rect 18245 50677 18279 50711
rect 2789 50405 2823 50439
rect 3249 50337 3283 50371
rect 3341 50269 3375 50303
rect 14473 50269 14507 50303
rect 3249 50133 3283 50167
rect 14289 50133 14323 50167
rect 4445 49929 4479 49963
rect 3332 49861 3366 49895
rect 8300 49861 8334 49895
rect 3065 49725 3099 49759
rect 8033 49725 8067 49759
rect 9413 49657 9447 49691
rect 7389 49317 7423 49351
rect 6009 49181 6043 49215
rect 6276 49113 6310 49147
rect 7481 48841 7515 48875
rect 15853 48841 15887 48875
rect 10701 48773 10735 48807
rect 3157 48705 3191 48739
rect 3700 48705 3734 48739
rect 7665 48705 7699 48739
rect 14657 48705 14691 48739
rect 16037 48705 16071 48739
rect 18061 48705 18095 48739
rect 3433 48637 3467 48671
rect 10793 48637 10827 48671
rect 10885 48637 10919 48671
rect 14749 48637 14783 48671
rect 14933 48637 14967 48671
rect 4813 48569 4847 48603
rect 14289 48569 14323 48603
rect 10333 48501 10367 48535
rect 18245 48501 18279 48535
rect 2421 47753 2455 47787
rect 6561 47753 6595 47787
rect 11897 47753 11931 47787
rect 7021 47685 7055 47719
rect 13154 47685 13188 47719
rect 2329 47617 2363 47651
rect 3065 47617 3099 47651
rect 4997 47617 5031 47651
rect 6929 47617 6963 47651
rect 12081 47617 12115 47651
rect 7205 47549 7239 47583
rect 12909 47549 12943 47583
rect 3249 47481 3283 47515
rect 4813 47413 4847 47447
rect 14289 47413 14323 47447
rect 2789 47141 2823 47175
rect 7389 47141 7423 47175
rect 3065 47005 3099 47039
rect 7573 47005 7607 47039
rect 18061 47005 18095 47039
rect 3249 46937 3283 46971
rect 3341 46937 3375 46971
rect 18245 46869 18279 46903
rect 12532 46597 12566 46631
rect 12265 46461 12299 46495
rect 13645 46325 13679 46359
rect 16405 45033 16439 45067
rect 14289 44897 14323 44931
rect 14565 44897 14599 44931
rect 13093 44829 13127 44863
rect 16589 44829 16623 44863
rect 18061 44829 18095 44863
rect 13461 44761 13495 44795
rect 15669 44693 15703 44727
rect 18245 44693 18279 44727
rect 1961 44421 1995 44455
rect 2145 44421 2179 44455
rect 2237 44421 2271 44455
rect 4353 44353 4387 44387
rect 4609 44353 4643 44387
rect 1685 44149 1719 44183
rect 5733 44149 5767 44183
rect 7297 43809 7331 43843
rect 7205 43741 7239 43775
rect 7113 43673 7147 43707
rect 6745 43605 6779 43639
rect 18061 43265 18095 43299
rect 18245 43061 18279 43095
rect 13001 42857 13035 42891
rect 2145 42721 2179 42755
rect 2697 42721 2731 42755
rect 11069 42721 11103 42755
rect 13645 42721 13679 42755
rect 2237 42653 2271 42687
rect 2973 42653 3007 42687
rect 9965 42653 9999 42687
rect 2145 42585 2179 42619
rect 10885 42585 10919 42619
rect 13369 42585 13403 42619
rect 1675 42517 1709 42551
rect 2789 42517 2823 42551
rect 9781 42517 9815 42551
rect 10517 42517 10551 42551
rect 10977 42517 11011 42551
rect 13461 42517 13495 42551
rect 3525 42313 3559 42347
rect 8677 42313 8711 42347
rect 9137 42313 9171 42347
rect 2390 42245 2424 42279
rect 7564 42245 7598 42279
rect 9597 42245 9631 42279
rect 2145 42177 2179 42211
rect 7297 42177 7331 42211
rect 9505 42177 9539 42211
rect 9781 42109 9815 42143
rect 6377 41633 6411 41667
rect 5733 41429 5767 41463
rect 6101 41429 6135 41463
rect 6193 41429 6227 41463
rect 18061 41089 18095 41123
rect 18245 40885 18279 40919
rect 7849 40137 7883 40171
rect 10977 40137 11011 40171
rect 8217 40069 8251 40103
rect 9853 40001 9887 40035
rect 15761 40001 15795 40035
rect 8309 39933 8343 39967
rect 8493 39933 8527 39967
rect 9597 39933 9631 39967
rect 15485 39933 15519 39967
rect 13001 39457 13035 39491
rect 12725 39389 12759 39423
rect 18061 39389 18095 39423
rect 12817 39321 12851 39355
rect 12357 39253 12391 39287
rect 18245 39253 18279 39287
rect 3976 38981 4010 39015
rect 3709 38913 3743 38947
rect 17049 38913 17083 38947
rect 17693 38913 17727 38947
rect 18245 38845 18279 38879
rect 5089 38709 5123 38743
rect 16865 38709 16899 38743
rect 15485 38301 15519 38335
rect 15301 38165 15335 38199
rect 15945 37961 15979 37995
rect 16037 37825 16071 37859
rect 16129 37757 16163 37791
rect 15577 37621 15611 37655
rect 12633 37417 12667 37451
rect 13277 37281 13311 37315
rect 1961 37213 1995 37247
rect 13001 37213 13035 37247
rect 18061 37213 18095 37247
rect 2206 37145 2240 37179
rect 3341 37077 3375 37111
rect 13093 37077 13127 37111
rect 18245 37077 18279 37111
rect 8125 36873 8159 36907
rect 8585 36873 8619 36907
rect 8493 36737 8527 36771
rect 8677 36669 8711 36703
rect 2237 36329 2271 36363
rect 11437 36261 11471 36295
rect 2881 36193 2915 36227
rect 12357 36193 12391 36227
rect 2697 36125 2731 36159
rect 12173 36125 12207 36159
rect 2605 36057 2639 36091
rect 12265 36057 12299 36091
rect 11805 35989 11839 36023
rect 13338 35717 13372 35751
rect 12357 35649 12391 35683
rect 18061 35649 18095 35683
rect 13093 35581 13127 35615
rect 14473 35513 14507 35547
rect 12449 35445 12483 35479
rect 18245 35445 18279 35479
rect 10517 35241 10551 35275
rect 13001 35173 13035 35207
rect 8309 35105 8343 35139
rect 8493 35105 8527 35139
rect 13645 35105 13679 35139
rect 8217 35037 8251 35071
rect 9137 35037 9171 35071
rect 13369 35037 13403 35071
rect 9382 34969 9416 35003
rect 13461 34969 13495 35003
rect 7849 34901 7883 34935
rect 10149 34697 10183 34731
rect 12265 34697 12299 34731
rect 14749 34697 14783 34731
rect 15393 34697 15427 34731
rect 3065 34629 3099 34663
rect 3249 34629 3283 34663
rect 15853 34629 15887 34663
rect 2771 34561 2805 34595
rect 9025 34561 9059 34595
rect 12633 34561 12667 34595
rect 13369 34561 13403 34595
rect 13625 34561 13659 34595
rect 15025 34561 15059 34595
rect 15761 34561 15795 34595
rect 3341 34493 3375 34527
rect 8769 34493 8803 34527
rect 12725 34493 12759 34527
rect 12817 34493 12851 34527
rect 16037 34493 16071 34527
rect 16865 34085 16899 34119
rect 17417 34017 17451 34051
rect 16313 33949 16347 33983
rect 17141 33881 17175 33915
rect 16129 33813 16163 33847
rect 17325 33813 17359 33847
rect 15577 33609 15611 33643
rect 15761 33473 15795 33507
rect 18061 33473 18095 33507
rect 18245 33269 18279 33303
rect 16957 33065 16991 33099
rect 15577 32929 15611 32963
rect 15844 32793 15878 32827
rect 7297 32521 7331 32555
rect 17110 32453 17144 32487
rect 7205 32385 7239 32419
rect 11989 32385 12023 32419
rect 12256 32385 12290 32419
rect 16865 32385 16899 32419
rect 7389 32317 7423 32351
rect 6837 32181 6871 32215
rect 13369 32181 13403 32215
rect 18245 32181 18279 32215
rect 18061 31773 18095 31807
rect 18245 31637 18279 31671
rect 1593 31433 1627 31467
rect 18245 31433 18279 31467
rect 17110 31365 17144 31399
rect 1777 31297 1811 31331
rect 16865 31297 16899 31331
rect 6377 30753 6411 30787
rect 6101 30617 6135 30651
rect 5733 30549 5767 30583
rect 6193 30549 6227 30583
rect 7113 30277 7147 30311
rect 8013 30277 8047 30311
rect 14832 30277 14866 30311
rect 3249 30209 3283 30243
rect 3801 30209 3835 30243
rect 7757 30209 7791 30243
rect 14565 30209 14599 30243
rect 7113 30141 7147 30175
rect 7205 30141 7239 30175
rect 9137 30073 9171 30107
rect 6653 30005 6687 30039
rect 15945 30005 15979 30039
rect 15669 29801 15703 29835
rect 16313 29665 16347 29699
rect 18061 29597 18095 29631
rect 16037 29461 16071 29495
rect 16129 29461 16163 29495
rect 18245 29461 18279 29495
rect 9597 29257 9631 29291
rect 4629 29189 4663 29223
rect 4445 29121 4479 29155
rect 9965 29121 9999 29155
rect 10057 29053 10091 29087
rect 10241 29053 10275 29087
rect 9321 28713 9355 28747
rect 5365 28577 5399 28611
rect 9781 28577 9815 28611
rect 5641 28509 5675 28543
rect 9873 28441 9907 28475
rect 9781 28373 9815 28407
rect 4322 28101 4356 28135
rect 18061 28033 18095 28067
rect 4077 27965 4111 27999
rect 5457 27829 5491 27863
rect 18245 27829 18279 27863
rect 18245 27557 18279 27591
rect 4261 27489 4295 27523
rect 4077 27421 4111 27455
rect 18061 27421 18095 27455
rect 14657 27081 14691 27115
rect 13277 26945 13311 26979
rect 13533 26945 13567 26979
rect 3433 26537 3467 26571
rect 6929 26537 6963 26571
rect 5549 26401 5583 26435
rect 2053 26333 2087 26367
rect 2320 26265 2354 26299
rect 5816 26265 5850 26299
rect 10149 25993 10183 26027
rect 10517 25993 10551 26027
rect 18061 25857 18095 25891
rect 10609 25789 10643 25823
rect 10793 25789 10827 25823
rect 18245 25653 18279 25687
rect 5365 25449 5399 25483
rect 9873 25381 9907 25415
rect 6653 25313 6687 25347
rect 6929 25313 6963 25347
rect 10333 25313 10367 25347
rect 10425 25313 10459 25347
rect 12909 25313 12943 25347
rect 3985 25245 4019 25279
rect 10241 25245 10275 25279
rect 12725 25245 12759 25279
rect 4252 25177 4286 25211
rect 12817 25177 12851 25211
rect 12357 25109 12391 25143
rect 17969 24905 18003 24939
rect 9229 24769 9263 24803
rect 9781 24769 9815 24803
rect 9965 24769 9999 24803
rect 18061 24701 18095 24735
rect 18153 24701 18187 24735
rect 17601 24633 17635 24667
rect 9045 24565 9079 24599
rect 18061 24157 18095 24191
rect 18245 24021 18279 24055
rect 9321 23817 9355 23851
rect 17417 23817 17451 23851
rect 8186 23749 8220 23783
rect 17233 23749 17267 23783
rect 3433 23681 3467 23715
rect 7941 23681 7975 23715
rect 17509 23681 17543 23715
rect 16957 23545 16991 23579
rect 3249 23477 3283 23511
rect 17693 22729 17727 22763
rect 17785 22593 17819 22627
rect 17693 22525 17727 22559
rect 17233 22457 17267 22491
rect 2421 22117 2455 22151
rect 7021 22117 7055 22151
rect 2881 22049 2915 22083
rect 5181 21981 5215 22015
rect 7205 21981 7239 22015
rect 14565 21981 14599 22015
rect 18061 21981 18095 22015
rect 2973 21913 3007 21947
rect 3433 21913 3467 21947
rect 4169 21913 4203 21947
rect 4537 21913 4571 21947
rect 4905 21913 4939 21947
rect 5448 21913 5482 21947
rect 2881 21845 2915 21879
rect 6561 21845 6595 21879
rect 6929 21845 6963 21879
rect 14381 21845 14415 21879
rect 18245 21845 18279 21879
rect 11161 21641 11195 21675
rect 11897 21641 11931 21675
rect 12357 21641 12391 21675
rect 12725 21641 12759 21675
rect 11805 21505 11839 21539
rect 9137 21097 9171 21131
rect 17141 21097 17175 21131
rect 8309 21029 8343 21063
rect 6929 20961 6963 20995
rect 9597 20961 9631 20995
rect 9781 20961 9815 20995
rect 15761 20961 15795 20995
rect 6285 20893 6319 20927
rect 6653 20893 6687 20927
rect 7196 20893 7230 20927
rect 14657 20893 14691 20927
rect 15025 20825 15059 20859
rect 16028 20825 16062 20859
rect 9505 20757 9539 20791
rect 16957 20553 16991 20587
rect 17325 20553 17359 20587
rect 2145 20485 2179 20519
rect 14933 20485 14967 20519
rect 2237 20417 2271 20451
rect 11969 20417 12003 20451
rect 14841 20417 14875 20451
rect 2145 20349 2179 20383
rect 11713 20349 11747 20383
rect 15025 20349 15059 20383
rect 17417 20349 17451 20383
rect 17601 20349 17635 20383
rect 1685 20281 1719 20315
rect 13093 20281 13127 20315
rect 14473 20281 14507 20315
rect 2697 20213 2731 20247
rect 18245 19941 18279 19975
rect 18061 19805 18095 19839
rect 11989 19465 12023 19499
rect 12173 19329 12207 19363
rect 15301 18377 15335 18411
rect 14188 18309 14222 18343
rect 13921 18241 13955 18275
rect 18061 18241 18095 18275
rect 18245 18037 18279 18071
rect 11989 17833 12023 17867
rect 13001 17765 13035 17799
rect 10609 17697 10643 17731
rect 13461 17697 13495 17731
rect 13645 17697 13679 17731
rect 10876 17629 10910 17663
rect 13369 17629 13403 17663
rect 10701 17221 10735 17255
rect 10793 16949 10827 16983
rect 17969 16745 18003 16779
rect 6009 16609 6043 16643
rect 7113 16609 7147 16643
rect 5825 16541 5859 16575
rect 17877 16541 17911 16575
rect 7358 16473 7392 16507
rect 5457 16405 5491 16439
rect 5917 16405 5951 16439
rect 8493 16405 8527 16439
rect 7021 16201 7055 16235
rect 7389 16201 7423 16235
rect 7757 16201 7791 16235
rect 8217 16201 8251 16235
rect 8677 16201 8711 16235
rect 9045 16201 9079 16235
rect 9321 16201 9355 16235
rect 9781 16201 9815 16235
rect 18245 16201 18279 16235
rect 9229 16133 9263 16167
rect 8033 16065 8067 16099
rect 18061 16065 18095 16099
rect 8677 15657 8711 15691
rect 11897 15657 11931 15691
rect 12541 15589 12575 15623
rect 13001 15521 13035 15555
rect 13093 15521 13127 15555
rect 12081 15453 12115 15487
rect 16865 15453 16899 15487
rect 17110 15385 17144 15419
rect 12909 15317 12943 15351
rect 18245 15317 18279 15351
rect 1869 15113 1903 15147
rect 2421 15113 2455 15147
rect 18153 15113 18187 15147
rect 2329 15045 2363 15079
rect 17969 15045 18003 15079
rect 18245 14977 18279 15011
rect 17693 14841 17727 14875
rect 7665 14569 7699 14603
rect 16865 14569 16899 14603
rect 8585 14501 8619 14535
rect 7849 14365 7883 14399
rect 8401 14365 8435 14399
rect 15485 14365 15519 14399
rect 18061 14365 18095 14399
rect 15730 14297 15764 14331
rect 18245 14229 18279 14263
rect 6561 14025 6595 14059
rect 6745 13889 6779 13923
rect 16129 13481 16163 13515
rect 16405 13277 16439 13311
rect 16681 13209 16715 13243
rect 16589 13141 16623 13175
rect 4537 12937 4571 12971
rect 18245 12937 18279 12971
rect 2513 12869 2547 12903
rect 2881 12869 2915 12903
rect 3424 12869 3458 12903
rect 4997 12869 5031 12903
rect 5273 12869 5307 12903
rect 17132 12869 17166 12903
rect 16865 12801 16899 12835
rect 3157 12733 3191 12767
rect 7389 12393 7423 12427
rect 12173 12325 12207 12359
rect 18245 12325 18279 12359
rect 8585 12257 8619 12291
rect 9137 12257 9171 12291
rect 6009 12189 6043 12223
rect 9413 12189 9447 12223
rect 10333 12189 10367 12223
rect 10701 12189 10735 12223
rect 10793 12189 10827 12223
rect 11060 12189 11094 12223
rect 18061 12189 18095 12223
rect 6276 12121 6310 12155
rect 14565 11169 14599 11203
rect 15301 11169 15335 11203
rect 14657 11101 14691 11135
rect 14841 11101 14875 11135
rect 1869 10761 1903 10795
rect 2697 10761 2731 10795
rect 3157 10761 3191 10795
rect 2237 10693 2271 10727
rect 2605 10693 2639 10727
rect 18061 10625 18095 10659
rect 18245 10421 18279 10455
rect 1869 10217 1903 10251
rect 7665 10081 7699 10115
rect 7941 10081 7975 10115
rect 5181 10013 5215 10047
rect 6929 10013 6963 10047
rect 7021 10013 7055 10047
rect 7205 10013 7239 10047
rect 4997 9877 5031 9911
rect 6009 9877 6043 9911
rect 6285 9877 6319 9911
rect 6193 9605 6227 9639
rect 7481 9605 7515 9639
rect 7573 9605 7607 9639
rect 1777 9537 1811 9571
rect 2145 9537 2179 9571
rect 2513 9537 2547 9571
rect 4005 9537 4039 9571
rect 4261 9537 4295 9571
rect 4629 9537 4663 9571
rect 4997 9537 5031 9571
rect 5365 9537 5399 9571
rect 5733 9537 5767 9571
rect 6653 9537 6687 9571
rect 7481 9469 7515 9503
rect 7021 9401 7055 9435
rect 2881 9333 2915 9367
rect 4169 9129 4203 9163
rect 4537 9129 4571 9163
rect 4905 9129 4939 9163
rect 8033 9129 8067 9163
rect 17693 9129 17727 9163
rect 5733 8993 5767 9027
rect 5181 8925 5215 8959
rect 8217 8925 8251 8959
rect 18061 8925 18095 8959
rect 10149 8857 10183 8891
rect 8493 8789 8527 8823
rect 9321 8789 9355 8823
rect 9689 8789 9723 8823
rect 10241 8789 10275 8823
rect 10609 8789 10643 8823
rect 10977 8789 11011 8823
rect 18245 8789 18279 8823
rect 3709 8585 3743 8619
rect 17969 8585 18003 8619
rect 2053 8449 2087 8483
rect 9597 8449 9631 8483
rect 9864 8449 9898 8483
rect 14657 8449 14691 8483
rect 17785 8449 17819 8483
rect 2329 8381 2363 8415
rect 2605 8381 2639 8415
rect 14381 8381 14415 8415
rect 10977 8313 11011 8347
rect 2973 8041 3007 8075
rect 3341 8041 3375 8075
rect 4353 8041 4387 8075
rect 4721 8041 4755 8075
rect 5089 8041 5123 8075
rect 5457 8041 5491 8075
rect 11529 8041 11563 8075
rect 11897 8041 11931 8075
rect 9597 7905 9631 7939
rect 9781 7905 9815 7939
rect 4169 7837 4203 7871
rect 9505 7837 9539 7871
rect 12265 7837 12299 7871
rect 12909 7769 12943 7803
rect 13185 7769 13219 7803
rect 9137 7701 9171 7735
rect 12449 7701 12483 7735
rect 11989 7497 12023 7531
rect 14197 7429 14231 7463
rect 13829 7225 13863 7259
rect 14381 7225 14415 7259
rect 6929 6885 6963 6919
rect 9229 6885 9263 6919
rect 7389 6817 7423 6851
rect 7481 6817 7515 6851
rect 18061 6749 18095 6783
rect 9505 6681 9539 6715
rect 9689 6681 9723 6715
rect 9781 6681 9815 6715
rect 7389 6613 7423 6647
rect 18245 6613 18279 6647
rect 5089 5661 5123 5695
rect 5356 5661 5390 5695
rect 6469 5525 6503 5559
rect 13369 5253 13403 5287
rect 16957 5253 16991 5287
rect 5917 5185 5951 5219
rect 11713 5185 11747 5219
rect 16221 5185 16255 5219
rect 17141 5185 17175 5219
rect 17417 5185 17451 5219
rect 18061 5185 18095 5219
rect 11989 5117 12023 5151
rect 13645 5117 13679 5151
rect 14013 5117 14047 5151
rect 14381 5117 14415 5151
rect 17785 5117 17819 5151
rect 10701 5049 10735 5083
rect 11069 5049 11103 5083
rect 5733 4981 5767 5015
rect 18245 4981 18279 5015
rect 10333 4641 10367 4675
rect 10057 4573 10091 4607
rect 6561 4097 6595 4131
rect 6817 4097 6851 4131
rect 9781 4097 9815 4131
rect 10057 4029 10091 4063
rect 7941 3961 7975 3995
rect 13645 3689 13679 3723
rect 12265 3553 12299 3587
rect 12521 3485 12555 3519
rect 3893 3145 3927 3179
rect 2780 3077 2814 3111
rect 18061 3009 18095 3043
rect 2513 2941 2547 2975
rect 18245 2805 18279 2839
rect 7205 2601 7239 2635
rect 7573 2601 7607 2635
rect 7941 2601 7975 2635
rect 14473 2601 14507 2635
rect 18061 2465 18095 2499
rect 6561 2397 6595 2431
rect 10057 2397 10091 2431
rect 17877 2397 17911 2431
rect 14381 2329 14415 2363
rect 5641 2261 5675 2295
rect 5917 2261 5951 2295
rect 6745 2261 6779 2295
rect 10241 2261 10275 2295
<< metal1 >>
rect 1104 77818 18860 77840
rect 1104 77766 1950 77818
rect 2002 77766 2014 77818
rect 2066 77766 2078 77818
rect 2130 77766 2142 77818
rect 2194 77766 2206 77818
rect 2258 77766 6950 77818
rect 7002 77766 7014 77818
rect 7066 77766 7078 77818
rect 7130 77766 7142 77818
rect 7194 77766 7206 77818
rect 7258 77766 11950 77818
rect 12002 77766 12014 77818
rect 12066 77766 12078 77818
rect 12130 77766 12142 77818
rect 12194 77766 12206 77818
rect 12258 77766 16950 77818
rect 17002 77766 17014 77818
rect 17066 77766 17078 77818
rect 17130 77766 17142 77818
rect 17194 77766 17206 77818
rect 17258 77766 18860 77818
rect 1104 77744 18860 77766
rect 18049 77503 18107 77509
rect 18049 77469 18061 77503
rect 18095 77500 18107 77503
rect 18322 77500 18328 77512
rect 18095 77472 18328 77500
rect 18095 77469 18107 77472
rect 18049 77463 18107 77469
rect 18322 77460 18328 77472
rect 18380 77460 18386 77512
rect 16850 77324 16856 77376
rect 16908 77364 16914 77376
rect 16945 77367 17003 77373
rect 16945 77364 16957 77367
rect 16908 77336 16957 77364
rect 16908 77324 16914 77336
rect 16945 77333 16957 77336
rect 16991 77364 17003 77367
rect 17221 77367 17279 77373
rect 17221 77364 17233 77367
rect 16991 77336 17233 77364
rect 16991 77333 17003 77336
rect 16945 77327 17003 77333
rect 17221 77333 17233 77336
rect 17267 77333 17279 77367
rect 17221 77327 17279 77333
rect 18230 77324 18236 77376
rect 18288 77324 18294 77376
rect 1104 77274 18860 77296
rect 1104 77222 2610 77274
rect 2662 77222 2674 77274
rect 2726 77222 2738 77274
rect 2790 77222 2802 77274
rect 2854 77222 2866 77274
rect 2918 77222 7610 77274
rect 7662 77222 7674 77274
rect 7726 77222 7738 77274
rect 7790 77222 7802 77274
rect 7854 77222 7866 77274
rect 7918 77222 12610 77274
rect 12662 77222 12674 77274
rect 12726 77222 12738 77274
rect 12790 77222 12802 77274
rect 12854 77222 12866 77274
rect 12918 77222 17610 77274
rect 17662 77222 17674 77274
rect 17726 77222 17738 77274
rect 17790 77222 17802 77274
rect 17854 77222 17866 77274
rect 17918 77222 18860 77274
rect 1104 77200 18860 77222
rect 17129 76959 17187 76965
rect 17129 76956 17141 76959
rect 16546 76928 17141 76956
rect 16546 76832 16574 76928
rect 17129 76925 17141 76928
rect 17175 76956 17187 76959
rect 17405 76959 17463 76965
rect 17405 76956 17417 76959
rect 17175 76928 17417 76956
rect 17175 76925 17187 76928
rect 17129 76919 17187 76925
rect 17405 76925 17417 76928
rect 17451 76925 17463 76959
rect 17405 76919 17463 76925
rect 17494 76916 17500 76968
rect 17552 76956 17558 76968
rect 17681 76959 17739 76965
rect 17681 76956 17693 76959
rect 17552 76928 17693 76956
rect 17552 76916 17558 76928
rect 17681 76925 17693 76928
rect 17727 76925 17739 76959
rect 17681 76919 17739 76925
rect 13909 76823 13967 76829
rect 13909 76789 13921 76823
rect 13955 76820 13967 76823
rect 14277 76823 14335 76829
rect 14277 76820 14289 76823
rect 13955 76792 14289 76820
rect 13955 76789 13967 76792
rect 13909 76783 13967 76789
rect 14277 76789 14289 76792
rect 14323 76820 14335 76823
rect 14642 76820 14648 76832
rect 14323 76792 14648 76820
rect 14323 76789 14335 76792
rect 14277 76783 14335 76789
rect 14642 76780 14648 76792
rect 14700 76780 14706 76832
rect 15930 76780 15936 76832
rect 15988 76820 15994 76832
rect 16209 76823 16267 76829
rect 16209 76820 16221 76823
rect 15988 76792 16221 76820
rect 15988 76780 15994 76792
rect 16209 76789 16221 76792
rect 16255 76820 16267 76823
rect 16482 76820 16488 76832
rect 16255 76792 16488 76820
rect 16255 76789 16267 76792
rect 16209 76783 16267 76789
rect 16482 76780 16488 76792
rect 16540 76792 16574 76832
rect 16540 76780 16546 76792
rect 1104 76730 18860 76752
rect 1104 76678 1950 76730
rect 2002 76678 2014 76730
rect 2066 76678 2078 76730
rect 2130 76678 2142 76730
rect 2194 76678 2206 76730
rect 2258 76678 6950 76730
rect 7002 76678 7014 76730
rect 7066 76678 7078 76730
rect 7130 76678 7142 76730
rect 7194 76678 7206 76730
rect 7258 76678 11950 76730
rect 12002 76678 12014 76730
rect 12066 76678 12078 76730
rect 12130 76678 12142 76730
rect 12194 76678 12206 76730
rect 12258 76678 16950 76730
rect 17002 76678 17014 76730
rect 17066 76678 17078 76730
rect 17130 76678 17142 76730
rect 17194 76678 17206 76730
rect 17258 76678 18860 76730
rect 1104 76656 18860 76678
rect 16482 76576 16488 76628
rect 16540 76616 16546 76628
rect 17129 76619 17187 76625
rect 17129 76616 17141 76619
rect 16540 76588 17141 76616
rect 16540 76576 16546 76588
rect 17129 76585 17141 76588
rect 17175 76616 17187 76619
rect 17497 76619 17555 76625
rect 17497 76616 17509 76619
rect 17175 76588 17509 76616
rect 17175 76585 17187 76588
rect 17129 76579 17187 76585
rect 17497 76585 17509 76588
rect 17543 76616 17555 76619
rect 17865 76619 17923 76625
rect 17865 76616 17877 76619
rect 17543 76588 17877 76616
rect 17543 76585 17555 76588
rect 17497 76579 17555 76585
rect 17865 76585 17877 76588
rect 17911 76616 17923 76619
rect 18233 76619 18291 76625
rect 18233 76616 18245 76619
rect 17911 76588 18245 76616
rect 17911 76585 17923 76588
rect 17865 76579 17923 76585
rect 18233 76585 18245 76588
rect 18279 76585 18291 76619
rect 18233 76579 18291 76585
rect 7745 76483 7803 76489
rect 7745 76449 7757 76483
rect 7791 76480 7803 76483
rect 7926 76480 7932 76492
rect 7791 76452 7932 76480
rect 7791 76449 7803 76452
rect 7745 76443 7803 76449
rect 7926 76440 7932 76452
rect 7984 76440 7990 76492
rect 7837 76415 7895 76421
rect 7837 76381 7849 76415
rect 7883 76381 7895 76415
rect 7837 76375 7895 76381
rect 8021 76415 8079 76421
rect 8021 76381 8033 76415
rect 8067 76412 8079 76415
rect 8202 76412 8208 76424
rect 8067 76384 8208 76412
rect 8067 76381 8079 76384
rect 8021 76375 8079 76381
rect 2958 76236 2964 76288
rect 3016 76276 3022 76288
rect 7098 76276 7104 76288
rect 3016 76248 7104 76276
rect 3016 76236 3022 76248
rect 7098 76236 7104 76248
rect 7156 76236 7162 76288
rect 7193 76279 7251 76285
rect 7193 76245 7205 76279
rect 7239 76276 7251 76279
rect 7852 76276 7880 76375
rect 8202 76372 8208 76384
rect 8260 76372 8266 76424
rect 14918 76372 14924 76424
rect 14976 76372 14982 76424
rect 8478 76304 8484 76356
rect 8536 76304 8542 76356
rect 11609 76347 11667 76353
rect 11609 76313 11621 76347
rect 11655 76313 11667 76347
rect 11609 76307 11667 76313
rect 8938 76276 8944 76288
rect 7239 76248 8944 76276
rect 7239 76245 7251 76248
rect 7193 76239 7251 76245
rect 8938 76236 8944 76248
rect 8996 76236 9002 76288
rect 11238 76236 11244 76288
rect 11296 76276 11302 76288
rect 11624 76276 11652 76307
rect 14642 76304 14648 76356
rect 14700 76344 14706 76356
rect 15166 76347 15224 76353
rect 15166 76344 15178 76347
rect 14700 76316 15178 76344
rect 14700 76304 14706 76316
rect 15166 76313 15178 76316
rect 15212 76344 15224 76347
rect 16850 76344 16856 76356
rect 15212 76316 16856 76344
rect 15212 76313 15224 76316
rect 15166 76307 15224 76313
rect 16850 76304 16856 76316
rect 16908 76304 16914 76356
rect 11296 76248 11652 76276
rect 11296 76236 11302 76248
rect 11698 76236 11704 76288
rect 11756 76236 11762 76288
rect 16298 76236 16304 76288
rect 16356 76236 16362 76288
rect 1104 76186 18860 76208
rect 1104 76134 2610 76186
rect 2662 76134 2674 76186
rect 2726 76134 2738 76186
rect 2790 76134 2802 76186
rect 2854 76134 2866 76186
rect 2918 76134 7610 76186
rect 7662 76134 7674 76186
rect 7726 76134 7738 76186
rect 7790 76134 7802 76186
rect 7854 76134 7866 76186
rect 7918 76134 12610 76186
rect 12662 76134 12674 76186
rect 12726 76134 12738 76186
rect 12790 76134 12802 76186
rect 12854 76134 12866 76186
rect 12918 76134 17610 76186
rect 17662 76134 17674 76186
rect 17726 76134 17738 76186
rect 17790 76134 17802 76186
rect 17854 76134 17866 76186
rect 17918 76134 18860 76186
rect 1104 76112 18860 76134
rect 16666 76072 16672 76084
rect 5644 76044 16672 76072
rect 5534 76004 5540 76016
rect 3988 75976 5540 76004
rect 3988 75945 4016 75976
rect 5534 75964 5540 75976
rect 5592 75964 5598 76016
rect 3973 75939 4031 75945
rect 3973 75905 3985 75939
rect 4019 75905 4031 75939
rect 3973 75899 4031 75905
rect 4240 75939 4298 75945
rect 4240 75905 4252 75939
rect 4286 75936 4298 75939
rect 5644 75936 5672 76044
rect 16666 76032 16672 76044
rect 16724 76032 16730 76084
rect 4286 75908 5672 75936
rect 5736 75976 7512 76004
rect 4286 75905 4298 75908
rect 4240 75899 4298 75905
rect 5736 75868 5764 75976
rect 6917 75939 6975 75945
rect 6917 75905 6929 75939
rect 6963 75936 6975 75939
rect 6963 75908 7052 75936
rect 6963 75905 6975 75908
rect 6917 75899 6975 75905
rect 5368 75840 5764 75868
rect 5368 75809 5396 75840
rect 6638 75828 6644 75880
rect 6696 75868 6702 75880
rect 6825 75871 6883 75877
rect 6825 75868 6837 75871
rect 6696 75840 6837 75868
rect 6696 75828 6702 75840
rect 6825 75837 6837 75840
rect 6871 75837 6883 75871
rect 7024 75868 7052 75908
rect 7098 75896 7104 75948
rect 7156 75896 7162 75948
rect 7374 75936 7380 75948
rect 7208 75908 7380 75936
rect 7208 75868 7236 75908
rect 7374 75896 7380 75908
rect 7432 75896 7438 75948
rect 7484 75936 7512 75976
rect 7558 75964 7564 76016
rect 7616 75964 7622 76016
rect 8754 75964 8760 76016
rect 8812 75964 8818 76016
rect 12434 76004 12440 76016
rect 12406 75964 12440 76004
rect 12492 75964 12498 76016
rect 12406 75936 12434 75964
rect 7484 75908 12434 75936
rect 14090 75896 14096 75948
rect 14148 75896 14154 75948
rect 14182 75896 14188 75948
rect 14240 75896 14246 75948
rect 7024 75840 7236 75868
rect 14369 75871 14427 75877
rect 6825 75831 6883 75837
rect 14369 75837 14381 75871
rect 14415 75868 14427 75871
rect 14458 75868 14464 75880
rect 14415 75840 14464 75868
rect 14415 75837 14427 75840
rect 14369 75831 14427 75837
rect 14458 75828 14464 75840
rect 14516 75828 14522 75880
rect 5353 75803 5411 75809
rect 5353 75769 5365 75803
rect 5399 75769 5411 75803
rect 5353 75763 5411 75769
rect 8389 75735 8447 75741
rect 8389 75701 8401 75735
rect 8435 75732 8447 75735
rect 8849 75735 8907 75741
rect 8849 75732 8861 75735
rect 8435 75704 8861 75732
rect 8435 75701 8447 75704
rect 8389 75695 8447 75701
rect 8849 75701 8861 75704
rect 8895 75732 8907 75735
rect 9214 75732 9220 75744
rect 8895 75704 9220 75732
rect 8895 75701 8907 75704
rect 8849 75695 8907 75701
rect 9214 75692 9220 75704
rect 9272 75692 9278 75744
rect 13722 75692 13728 75744
rect 13780 75692 13786 75744
rect 1104 75642 18860 75664
rect 1104 75590 1950 75642
rect 2002 75590 2014 75642
rect 2066 75590 2078 75642
rect 2130 75590 2142 75642
rect 2194 75590 2206 75642
rect 2258 75590 6950 75642
rect 7002 75590 7014 75642
rect 7066 75590 7078 75642
rect 7130 75590 7142 75642
rect 7194 75590 7206 75642
rect 7258 75590 11950 75642
rect 12002 75590 12014 75642
rect 12066 75590 12078 75642
rect 12130 75590 12142 75642
rect 12194 75590 12206 75642
rect 12258 75590 16950 75642
rect 17002 75590 17014 75642
rect 17066 75590 17078 75642
rect 17130 75590 17142 75642
rect 17194 75590 17206 75642
rect 17258 75590 18860 75642
rect 1104 75568 18860 75590
rect 15194 75420 15200 75472
rect 15252 75420 15258 75472
rect 5721 75395 5779 75401
rect 5721 75361 5733 75395
rect 5767 75392 5779 75395
rect 11790 75392 11796 75404
rect 5767 75364 11796 75392
rect 5767 75361 5779 75364
rect 5721 75355 5779 75361
rect 11790 75352 11796 75364
rect 11848 75352 11854 75404
rect 5442 75284 5448 75336
rect 5500 75324 5506 75336
rect 5537 75327 5595 75333
rect 5537 75324 5549 75327
rect 5500 75296 5549 75324
rect 5500 75284 5506 75296
rect 5537 75293 5549 75296
rect 5583 75293 5595 75327
rect 5537 75287 5595 75293
rect 7282 75284 7288 75336
rect 7340 75324 7346 75336
rect 7561 75327 7619 75333
rect 7561 75324 7573 75327
rect 7340 75296 7573 75324
rect 7340 75284 7346 75296
rect 7561 75293 7573 75296
rect 7607 75293 7619 75327
rect 7561 75287 7619 75293
rect 8110 75284 8116 75336
rect 8168 75324 8174 75336
rect 15381 75327 15439 75333
rect 15381 75324 15393 75327
rect 8168 75296 15393 75324
rect 8168 75284 8174 75296
rect 15381 75293 15393 75296
rect 15427 75293 15439 75327
rect 18049 75327 18107 75333
rect 18049 75324 18061 75327
rect 15381 75287 15439 75293
rect 16546 75296 18061 75324
rect 4985 75259 5043 75265
rect 4985 75225 4997 75259
rect 5031 75256 5043 75259
rect 5031 75228 12434 75256
rect 5031 75225 5043 75228
rect 4985 75219 5043 75225
rect 5074 75148 5080 75200
rect 5132 75148 5138 75200
rect 5460 75197 5488 75228
rect 5445 75191 5503 75197
rect 5445 75157 5457 75191
rect 5491 75157 5503 75191
rect 5445 75151 5503 75157
rect 6181 75191 6239 75197
rect 6181 75157 6193 75191
rect 6227 75188 6239 75191
rect 6546 75188 6552 75200
rect 6227 75160 6552 75188
rect 6227 75157 6239 75160
rect 6181 75151 6239 75157
rect 6546 75148 6552 75160
rect 6604 75188 6610 75200
rect 6825 75191 6883 75197
rect 6825 75188 6837 75191
rect 6604 75160 6837 75188
rect 6604 75148 6610 75160
rect 6825 75157 6837 75160
rect 6871 75188 6883 75191
rect 7193 75191 7251 75197
rect 7193 75188 7205 75191
rect 6871 75160 7205 75188
rect 6871 75157 6883 75160
rect 6825 75151 6883 75157
rect 7193 75157 7205 75160
rect 7239 75188 7251 75191
rect 7745 75191 7803 75197
rect 7745 75188 7757 75191
rect 7239 75160 7757 75188
rect 7239 75157 7251 75160
rect 7193 75151 7251 75157
rect 7745 75157 7757 75160
rect 7791 75188 7803 75191
rect 8113 75191 8171 75197
rect 8113 75188 8125 75191
rect 7791 75160 8125 75188
rect 7791 75157 7803 75160
rect 7745 75151 7803 75157
rect 8113 75157 8125 75160
rect 8159 75188 8171 75191
rect 8481 75191 8539 75197
rect 8481 75188 8493 75191
rect 8159 75160 8493 75188
rect 8159 75157 8171 75160
rect 8113 75151 8171 75157
rect 8481 75157 8493 75160
rect 8527 75188 8539 75191
rect 9125 75191 9183 75197
rect 9125 75188 9137 75191
rect 8527 75160 9137 75188
rect 8527 75157 8539 75160
rect 8481 75151 8539 75157
rect 9125 75157 9137 75160
rect 9171 75157 9183 75191
rect 12406 75188 12434 75228
rect 14090 75216 14096 75268
rect 14148 75256 14154 75268
rect 16546 75256 16574 75296
rect 18049 75293 18061 75296
rect 18095 75293 18107 75327
rect 18049 75287 18107 75293
rect 14148 75228 16574 75256
rect 14148 75216 14154 75228
rect 16022 75188 16028 75200
rect 12406 75160 16028 75188
rect 9125 75151 9183 75157
rect 16022 75148 16028 75160
rect 16080 75148 16086 75200
rect 18230 75148 18236 75200
rect 18288 75148 18294 75200
rect 1104 75098 18860 75120
rect 1104 75046 2610 75098
rect 2662 75046 2674 75098
rect 2726 75046 2738 75098
rect 2790 75046 2802 75098
rect 2854 75046 2866 75098
rect 2918 75046 7610 75098
rect 7662 75046 7674 75098
rect 7726 75046 7738 75098
rect 7790 75046 7802 75098
rect 7854 75046 7866 75098
rect 7918 75046 12610 75098
rect 12662 75046 12674 75098
rect 12726 75046 12738 75098
rect 12790 75046 12802 75098
rect 12854 75046 12866 75098
rect 12918 75046 17610 75098
rect 17662 75046 17674 75098
rect 17726 75046 17738 75098
rect 17790 75046 17802 75098
rect 17854 75046 17866 75098
rect 17918 75046 18860 75098
rect 1104 75024 18860 75046
rect 4709 74987 4767 74993
rect 4709 74953 4721 74987
rect 4755 74984 4767 74987
rect 8110 74984 8116 74996
rect 4755 74956 8116 74984
rect 4755 74953 4767 74956
rect 4709 74947 4767 74953
rect 8110 74944 8116 74956
rect 8168 74944 8174 74996
rect 15286 74944 15292 74996
rect 15344 74984 15350 74996
rect 16209 74987 16267 74993
rect 16209 74984 16221 74987
rect 15344 74956 16221 74984
rect 15344 74944 15350 74956
rect 16209 74953 16221 74956
rect 16255 74953 16267 74987
rect 16209 74947 16267 74953
rect 5077 74919 5135 74925
rect 5077 74885 5089 74919
rect 5123 74916 5135 74919
rect 6546 74916 6552 74928
rect 5123 74888 6552 74916
rect 5123 74885 5135 74888
rect 5077 74879 5135 74885
rect 6546 74876 6552 74888
rect 6604 74876 6610 74928
rect 5169 74851 5227 74857
rect 5169 74817 5181 74851
rect 5215 74848 5227 74851
rect 5215 74820 6408 74848
rect 5215 74817 5227 74820
rect 5169 74811 5227 74817
rect 5261 74783 5319 74789
rect 5261 74749 5273 74783
rect 5307 74749 5319 74783
rect 6380 74780 6408 74820
rect 6454 74808 6460 74860
rect 6512 74848 6518 74860
rect 6641 74851 6699 74857
rect 6641 74848 6653 74851
rect 6512 74820 6653 74848
rect 6512 74808 6518 74820
rect 6641 74817 6653 74820
rect 6687 74817 6699 74851
rect 6641 74811 6699 74817
rect 14829 74851 14887 74857
rect 14829 74817 14841 74851
rect 14875 74848 14887 74851
rect 14918 74848 14924 74860
rect 14875 74820 14924 74848
rect 14875 74817 14887 74820
rect 14829 74811 14887 74817
rect 14918 74808 14924 74820
rect 14976 74808 14982 74860
rect 15102 74857 15108 74860
rect 15096 74811 15108 74857
rect 15102 74808 15108 74811
rect 15160 74808 15166 74860
rect 16850 74808 16856 74860
rect 16908 74808 16914 74860
rect 9398 74780 9404 74792
rect 6380 74752 9404 74780
rect 5261 74743 5319 74749
rect 4614 74672 4620 74724
rect 4672 74712 4678 74724
rect 5276 74712 5304 74743
rect 9398 74740 9404 74752
rect 9456 74740 9462 74792
rect 4672 74684 5304 74712
rect 4672 74672 4678 74684
rect 15838 74672 15844 74724
rect 15896 74712 15902 74724
rect 17494 74712 17500 74724
rect 15896 74684 17500 74712
rect 15896 74672 15902 74684
rect 17494 74672 17500 74684
rect 17552 74672 17558 74724
rect 6730 74604 6736 74656
rect 6788 74604 6794 74656
rect 17037 74647 17095 74653
rect 17037 74613 17049 74647
rect 17083 74644 17095 74647
rect 18782 74644 18788 74656
rect 17083 74616 18788 74644
rect 17083 74613 17095 74616
rect 17037 74607 17095 74613
rect 18782 74604 18788 74616
rect 18840 74604 18846 74656
rect 1104 74554 18860 74576
rect 1104 74502 1950 74554
rect 2002 74502 2014 74554
rect 2066 74502 2078 74554
rect 2130 74502 2142 74554
rect 2194 74502 2206 74554
rect 2258 74502 6950 74554
rect 7002 74502 7014 74554
rect 7066 74502 7078 74554
rect 7130 74502 7142 74554
rect 7194 74502 7206 74554
rect 7258 74502 11950 74554
rect 12002 74502 12014 74554
rect 12066 74502 12078 74554
rect 12130 74502 12142 74554
rect 12194 74502 12206 74554
rect 12258 74502 16950 74554
rect 17002 74502 17014 74554
rect 17066 74502 17078 74554
rect 17130 74502 17142 74554
rect 17194 74502 17206 74554
rect 17258 74502 18860 74554
rect 1104 74480 18860 74502
rect 7374 74400 7380 74452
rect 7432 74440 7438 74452
rect 10318 74440 10324 74452
rect 7432 74412 10324 74440
rect 7432 74400 7438 74412
rect 10318 74400 10324 74412
rect 10376 74400 10382 74452
rect 12069 74443 12127 74449
rect 12069 74409 12081 74443
rect 12115 74440 12127 74443
rect 16850 74440 16856 74452
rect 12115 74412 16856 74440
rect 12115 74409 12127 74412
rect 12069 74403 12127 74409
rect 16850 74400 16856 74412
rect 16908 74400 16914 74452
rect 12713 74307 12771 74313
rect 12713 74273 12725 74307
rect 12759 74304 12771 74307
rect 13722 74304 13728 74316
rect 12759 74276 13728 74304
rect 12759 74273 12771 74276
rect 12713 74267 12771 74273
rect 13722 74264 13728 74276
rect 13780 74264 13786 74316
rect 14274 74196 14280 74248
rect 14332 74236 14338 74248
rect 14918 74236 14924 74248
rect 14332 74208 14924 74236
rect 14332 74196 14338 74208
rect 14918 74196 14924 74208
rect 14976 74196 14982 74248
rect 10502 74128 10508 74180
rect 10560 74168 10566 74180
rect 12529 74171 12587 74177
rect 12529 74168 12541 74171
rect 10560 74140 12541 74168
rect 10560 74128 10566 74140
rect 12529 74137 12541 74140
rect 12575 74137 12587 74171
rect 14522 74171 14580 74177
rect 14522 74168 14534 74171
rect 12529 74131 12587 74137
rect 13648 74140 14534 74168
rect 12434 74060 12440 74112
rect 12492 74060 12498 74112
rect 13446 74060 13452 74112
rect 13504 74100 13510 74112
rect 13648 74109 13676 74140
rect 14522 74137 14534 74140
rect 14568 74168 14580 74171
rect 15933 74171 15991 74177
rect 15933 74168 15945 74171
rect 14568 74140 15945 74168
rect 14568 74137 14580 74140
rect 14522 74131 14580 74137
rect 15933 74137 15945 74140
rect 15979 74168 15991 74171
rect 16301 74171 16359 74177
rect 16301 74168 16313 74171
rect 15979 74140 16313 74168
rect 15979 74137 15991 74140
rect 15933 74131 15991 74137
rect 16301 74137 16313 74140
rect 16347 74137 16359 74171
rect 16301 74131 16359 74137
rect 13633 74103 13691 74109
rect 13633 74100 13645 74103
rect 13504 74072 13645 74100
rect 13504 74060 13510 74072
rect 13633 74069 13645 74072
rect 13679 74069 13691 74103
rect 13633 74063 13691 74069
rect 15562 74060 15568 74112
rect 15620 74100 15626 74112
rect 15657 74103 15715 74109
rect 15657 74100 15669 74103
rect 15620 74072 15669 74100
rect 15620 74060 15626 74072
rect 15657 74069 15669 74072
rect 15703 74069 15715 74103
rect 15657 74063 15715 74069
rect 1104 74010 18860 74032
rect 1104 73958 2610 74010
rect 2662 73958 2674 74010
rect 2726 73958 2738 74010
rect 2790 73958 2802 74010
rect 2854 73958 2866 74010
rect 2918 73958 7610 74010
rect 7662 73958 7674 74010
rect 7726 73958 7738 74010
rect 7790 73958 7802 74010
rect 7854 73958 7866 74010
rect 7918 73958 12610 74010
rect 12662 73958 12674 74010
rect 12726 73958 12738 74010
rect 12790 73958 12802 74010
rect 12854 73958 12866 74010
rect 12918 73958 17610 74010
rect 17662 73958 17674 74010
rect 17726 73958 17738 74010
rect 17790 73958 17802 74010
rect 17854 73958 17866 74010
rect 17918 73958 18860 74010
rect 1104 73936 18860 73958
rect 7282 73856 7288 73908
rect 7340 73856 7346 73908
rect 15930 73788 15936 73840
rect 15988 73828 15994 73840
rect 16298 73828 16304 73840
rect 15988 73800 16304 73828
rect 15988 73788 15994 73800
rect 16298 73788 16304 73800
rect 16356 73828 16362 73840
rect 16356 73800 16574 73828
rect 16356 73788 16362 73800
rect 7374 73720 7380 73772
rect 7432 73760 7438 73772
rect 7653 73763 7711 73769
rect 7653 73760 7665 73763
rect 7432 73732 7665 73760
rect 7432 73720 7438 73732
rect 7653 73729 7665 73732
rect 7699 73729 7711 73763
rect 7653 73723 7711 73729
rect 7745 73763 7803 73769
rect 7745 73729 7757 73763
rect 7791 73760 7803 73763
rect 16546 73760 16574 73800
rect 18049 73763 18107 73769
rect 18049 73760 18061 73763
rect 7791 73732 16160 73760
rect 16546 73732 18061 73760
rect 7791 73729 7803 73732
rect 7745 73723 7803 73729
rect 7929 73695 7987 73701
rect 7929 73661 7941 73695
rect 7975 73692 7987 73695
rect 8202 73692 8208 73704
rect 7975 73664 8208 73692
rect 7975 73661 7987 73664
rect 7929 73655 7987 73661
rect 8202 73652 8208 73664
rect 8260 73652 8266 73704
rect 16132 73692 16160 73732
rect 18049 73729 18061 73732
rect 18095 73729 18107 73763
rect 18049 73723 18107 73729
rect 17494 73692 17500 73704
rect 16132 73664 17500 73692
rect 17494 73652 17500 73664
rect 17552 73652 17558 73704
rect 18230 73516 18236 73568
rect 18288 73516 18294 73568
rect 1104 73466 18860 73488
rect 1104 73414 1950 73466
rect 2002 73414 2014 73466
rect 2066 73414 2078 73466
rect 2130 73414 2142 73466
rect 2194 73414 2206 73466
rect 2258 73414 6950 73466
rect 7002 73414 7014 73466
rect 7066 73414 7078 73466
rect 7130 73414 7142 73466
rect 7194 73414 7206 73466
rect 7258 73414 11950 73466
rect 12002 73414 12014 73466
rect 12066 73414 12078 73466
rect 12130 73414 12142 73466
rect 12194 73414 12206 73466
rect 12258 73414 16950 73466
rect 17002 73414 17014 73466
rect 17066 73414 17078 73466
rect 17130 73414 17142 73466
rect 17194 73414 17206 73466
rect 17258 73414 18860 73466
rect 1104 73392 18860 73414
rect 5534 73176 5540 73228
rect 5592 73216 5598 73228
rect 6641 73219 6699 73225
rect 6641 73216 6653 73219
rect 5592 73188 6653 73216
rect 5592 73176 5598 73188
rect 6641 73185 6653 73188
rect 6687 73185 6699 73219
rect 9125 73219 9183 73225
rect 9125 73216 9137 73219
rect 6641 73179 6699 73185
rect 8312 73188 9137 73216
rect 8312 73089 8340 73188
rect 9125 73185 9137 73188
rect 9171 73185 9183 73219
rect 9125 73179 9183 73185
rect 6886 73083 6944 73089
rect 6886 73080 6898 73083
rect 6288 73052 6898 73080
rect 1302 72972 1308 73024
rect 1360 73012 1366 73024
rect 6288 73021 6316 73052
rect 6886 73049 6898 73052
rect 6932 73080 6944 73083
rect 8297 73083 8355 73089
rect 8297 73080 8309 73083
rect 6932 73052 8309 73080
rect 6932 73049 6944 73052
rect 6886 73043 6944 73049
rect 8297 73049 8309 73052
rect 8343 73049 8355 73083
rect 8297 73043 8355 73049
rect 5537 73015 5595 73021
rect 5537 73012 5549 73015
rect 1360 72984 5549 73012
rect 1360 72972 1366 72984
rect 5537 72981 5549 72984
rect 5583 73012 5595 73015
rect 5905 73015 5963 73021
rect 5905 73012 5917 73015
rect 5583 72984 5917 73012
rect 5583 72981 5595 72984
rect 5537 72975 5595 72981
rect 5905 72981 5917 72984
rect 5951 73012 5963 73015
rect 6273 73015 6331 73021
rect 6273 73012 6285 73015
rect 5951 72984 6285 73012
rect 5951 72981 5963 72984
rect 5905 72975 5963 72981
rect 6273 72981 6285 72984
rect 6319 72981 6331 73015
rect 6273 72975 6331 72981
rect 8021 73015 8079 73021
rect 8021 72981 8033 73015
rect 8067 73012 8079 73015
rect 8110 73012 8116 73024
rect 8067 72984 8116 73012
rect 8067 72981 8079 72984
rect 8021 72975 8079 72981
rect 8110 72972 8116 72984
rect 8168 72972 8174 73024
rect 1104 72922 18860 72944
rect 1104 72870 2610 72922
rect 2662 72870 2674 72922
rect 2726 72870 2738 72922
rect 2790 72870 2802 72922
rect 2854 72870 2866 72922
rect 2918 72870 7610 72922
rect 7662 72870 7674 72922
rect 7726 72870 7738 72922
rect 7790 72870 7802 72922
rect 7854 72870 7866 72922
rect 7918 72870 12610 72922
rect 12662 72870 12674 72922
rect 12726 72870 12738 72922
rect 12790 72870 12802 72922
rect 12854 72870 12866 72922
rect 12918 72870 17610 72922
rect 17662 72870 17674 72922
rect 17726 72870 17738 72922
rect 17790 72870 17802 72922
rect 17854 72870 17866 72922
rect 17918 72870 18860 72922
rect 1104 72848 18860 72870
rect 8202 72700 8208 72752
rect 8260 72740 8266 72752
rect 8260 72712 13492 72740
rect 8260 72700 8266 72712
rect 12342 72632 12348 72684
rect 12400 72672 12406 72684
rect 13173 72675 13231 72681
rect 13173 72672 13185 72675
rect 12400 72644 13185 72672
rect 12400 72632 12406 72644
rect 13173 72641 13185 72644
rect 13219 72641 13231 72675
rect 13173 72635 13231 72641
rect 7374 72564 7380 72616
rect 7432 72604 7438 72616
rect 13464 72613 13492 72712
rect 13265 72607 13323 72613
rect 13265 72604 13277 72607
rect 7432 72576 13277 72604
rect 7432 72564 7438 72576
rect 13265 72573 13277 72576
rect 13311 72573 13323 72607
rect 13265 72567 13323 72573
rect 13449 72607 13507 72613
rect 13449 72573 13461 72607
rect 13495 72604 13507 72607
rect 16574 72604 16580 72616
rect 13495 72576 16580 72604
rect 13495 72573 13507 72576
rect 13449 72567 13507 72573
rect 16574 72564 16580 72576
rect 16632 72564 16638 72616
rect 12805 72471 12863 72477
rect 12805 72437 12817 72471
rect 12851 72468 12863 72471
rect 13262 72468 13268 72480
rect 12851 72440 13268 72468
rect 12851 72437 12863 72440
rect 12805 72431 12863 72437
rect 13262 72428 13268 72440
rect 13320 72428 13326 72480
rect 1104 72378 18860 72400
rect 1104 72326 1950 72378
rect 2002 72326 2014 72378
rect 2066 72326 2078 72378
rect 2130 72326 2142 72378
rect 2194 72326 2206 72378
rect 2258 72326 6950 72378
rect 7002 72326 7014 72378
rect 7066 72326 7078 72378
rect 7130 72326 7142 72378
rect 7194 72326 7206 72378
rect 7258 72326 11950 72378
rect 12002 72326 12014 72378
rect 12066 72326 12078 72378
rect 12130 72326 12142 72378
rect 12194 72326 12206 72378
rect 12258 72326 16950 72378
rect 17002 72326 17014 72378
rect 17066 72326 17078 72378
rect 17130 72326 17142 72378
rect 17194 72326 17206 72378
rect 17258 72326 18860 72378
rect 1104 72304 18860 72326
rect 16666 72224 16672 72276
rect 16724 72264 16730 72276
rect 17037 72267 17095 72273
rect 17037 72264 17049 72267
rect 16724 72236 17049 72264
rect 16724 72224 16730 72236
rect 17037 72233 17049 72236
rect 17083 72233 17095 72267
rect 17037 72227 17095 72233
rect 16850 72020 16856 72072
rect 16908 72060 16914 72072
rect 17221 72063 17279 72069
rect 17221 72060 17233 72063
rect 16908 72032 17233 72060
rect 16908 72020 16914 72032
rect 17221 72029 17233 72032
rect 17267 72029 17279 72063
rect 17221 72023 17279 72029
rect 16574 71884 16580 71936
rect 16632 71924 16638 71936
rect 16850 71924 16856 71936
rect 16632 71896 16856 71924
rect 16632 71884 16638 71896
rect 16850 71884 16856 71896
rect 16908 71884 16914 71936
rect 1104 71834 18860 71856
rect 1104 71782 2610 71834
rect 2662 71782 2674 71834
rect 2726 71782 2738 71834
rect 2790 71782 2802 71834
rect 2854 71782 2866 71834
rect 2918 71782 7610 71834
rect 7662 71782 7674 71834
rect 7726 71782 7738 71834
rect 7790 71782 7802 71834
rect 7854 71782 7866 71834
rect 7918 71782 12610 71834
rect 12662 71782 12674 71834
rect 12726 71782 12738 71834
rect 12790 71782 12802 71834
rect 12854 71782 12866 71834
rect 12918 71782 17610 71834
rect 17662 71782 17674 71834
rect 17726 71782 17738 71834
rect 17790 71782 17802 71834
rect 17854 71782 17866 71834
rect 17918 71782 18860 71834
rect 1104 71760 18860 71782
rect 12434 71680 12440 71732
rect 12492 71720 12498 71732
rect 18966 71720 18972 71732
rect 12492 71692 18972 71720
rect 12492 71680 12498 71692
rect 18966 71680 18972 71692
rect 19024 71680 19030 71732
rect 5534 71652 5540 71664
rect 3068 71624 5540 71652
rect 3068 71593 3096 71624
rect 5534 71612 5540 71624
rect 5592 71612 5598 71664
rect 3326 71593 3332 71596
rect 3053 71587 3111 71593
rect 3053 71553 3065 71587
rect 3099 71553 3111 71587
rect 3053 71547 3111 71553
rect 3320 71547 3332 71593
rect 3326 71544 3332 71547
rect 3384 71544 3390 71596
rect 15654 71544 15660 71596
rect 15712 71584 15718 71596
rect 18049 71587 18107 71593
rect 18049 71584 18061 71587
rect 15712 71556 18061 71584
rect 15712 71544 15718 71556
rect 18049 71553 18061 71556
rect 18095 71553 18107 71587
rect 18049 71547 18107 71553
rect 4433 71383 4491 71389
rect 4433 71349 4445 71383
rect 4479 71380 4491 71383
rect 8202 71380 8208 71392
rect 4479 71352 8208 71380
rect 4479 71349 4491 71352
rect 4433 71343 4491 71349
rect 8202 71340 8208 71352
rect 8260 71340 8266 71392
rect 18230 71340 18236 71392
rect 18288 71340 18294 71392
rect 1104 71290 18860 71312
rect 1104 71238 1950 71290
rect 2002 71238 2014 71290
rect 2066 71238 2078 71290
rect 2130 71238 2142 71290
rect 2194 71238 2206 71290
rect 2258 71238 6950 71290
rect 7002 71238 7014 71290
rect 7066 71238 7078 71290
rect 7130 71238 7142 71290
rect 7194 71238 7206 71290
rect 7258 71238 11950 71290
rect 12002 71238 12014 71290
rect 12066 71238 12078 71290
rect 12130 71238 12142 71290
rect 12194 71238 12206 71290
rect 12258 71238 16950 71290
rect 17002 71238 17014 71290
rect 17066 71238 17078 71290
rect 17130 71238 17142 71290
rect 17194 71238 17206 71290
rect 17258 71238 18860 71290
rect 1104 71216 18860 71238
rect 6270 71136 6276 71188
rect 6328 71176 6334 71188
rect 15194 71176 15200 71188
rect 6328 71148 15200 71176
rect 6328 71136 6334 71148
rect 15194 71136 15200 71148
rect 15252 71136 15258 71188
rect 10502 71068 10508 71120
rect 10560 71068 10566 71120
rect 5534 71000 5540 71052
rect 5592 71040 5598 71052
rect 5997 71043 6055 71049
rect 5997 71040 6009 71043
rect 5592 71012 6009 71040
rect 5592 71000 5598 71012
rect 5997 71009 6009 71012
rect 6043 71009 6055 71043
rect 5997 71003 6055 71009
rect 6012 70972 6040 71003
rect 6822 70972 6828 70984
rect 6012 70944 6828 70972
rect 6822 70932 6828 70944
rect 6880 70972 6886 70984
rect 9122 70972 9128 70984
rect 6880 70944 9128 70972
rect 6880 70932 6886 70944
rect 9122 70932 9128 70944
rect 9180 70932 9186 70984
rect 9858 70932 9864 70984
rect 9916 70972 9922 70984
rect 10520 70972 10548 71068
rect 9916 70944 10548 70972
rect 9916 70932 9922 70944
rect 14274 70932 14280 70984
rect 14332 70972 14338 70984
rect 15473 70975 15531 70981
rect 15473 70972 15485 70975
rect 14332 70944 15485 70972
rect 14332 70932 14338 70944
rect 15473 70941 15485 70944
rect 15519 70941 15531 70975
rect 15473 70935 15531 70941
rect 6270 70913 6276 70916
rect 6264 70867 6276 70913
rect 6270 70864 6276 70867
rect 6328 70864 6334 70916
rect 15746 70913 15752 70916
rect 9370 70907 9428 70913
rect 9370 70904 9382 70907
rect 6380 70876 9382 70904
rect 1118 70796 1124 70848
rect 1176 70836 1182 70848
rect 6380 70836 6408 70876
rect 9370 70873 9382 70876
rect 9416 70873 9428 70907
rect 9370 70867 9428 70873
rect 15740 70867 15752 70913
rect 15746 70864 15752 70867
rect 15804 70864 15810 70916
rect 1176 70808 6408 70836
rect 1176 70796 1182 70808
rect 6546 70796 6552 70848
rect 6604 70836 6610 70848
rect 7377 70839 7435 70845
rect 7377 70836 7389 70839
rect 6604 70808 7389 70836
rect 6604 70796 6610 70808
rect 7377 70805 7389 70808
rect 7423 70836 7435 70839
rect 9030 70836 9036 70848
rect 7423 70808 9036 70836
rect 7423 70805 7435 70808
rect 7377 70799 7435 70805
rect 9030 70796 9036 70808
rect 9088 70796 9094 70848
rect 16666 70796 16672 70848
rect 16724 70836 16730 70848
rect 16853 70839 16911 70845
rect 16853 70836 16865 70839
rect 16724 70808 16865 70836
rect 16724 70796 16730 70808
rect 16853 70805 16865 70808
rect 16899 70805 16911 70839
rect 16853 70799 16911 70805
rect 1104 70746 18860 70768
rect 1104 70694 2610 70746
rect 2662 70694 2674 70746
rect 2726 70694 2738 70746
rect 2790 70694 2802 70746
rect 2854 70694 2866 70746
rect 2918 70694 7610 70746
rect 7662 70694 7674 70746
rect 7726 70694 7738 70746
rect 7790 70694 7802 70746
rect 7854 70694 7866 70746
rect 7918 70694 12610 70746
rect 12662 70694 12674 70746
rect 12726 70694 12738 70746
rect 12790 70694 12802 70746
rect 12854 70694 12866 70746
rect 12918 70694 17610 70746
rect 17662 70694 17674 70746
rect 17726 70694 17738 70746
rect 17790 70694 17802 70746
rect 17854 70694 17866 70746
rect 17918 70694 18860 70746
rect 1104 70672 18860 70694
rect 1104 70202 18860 70224
rect 1104 70150 1950 70202
rect 2002 70150 2014 70202
rect 2066 70150 2078 70202
rect 2130 70150 2142 70202
rect 2194 70150 2206 70202
rect 2258 70150 6950 70202
rect 7002 70150 7014 70202
rect 7066 70150 7078 70202
rect 7130 70150 7142 70202
rect 7194 70150 7206 70202
rect 7258 70150 11950 70202
rect 12002 70150 12014 70202
rect 12066 70150 12078 70202
rect 12130 70150 12142 70202
rect 12194 70150 12206 70202
rect 12258 70150 16950 70202
rect 17002 70150 17014 70202
rect 17066 70150 17078 70202
rect 17130 70150 17142 70202
rect 17194 70150 17206 70202
rect 17258 70150 18860 70202
rect 1104 70128 18860 70150
rect 16666 70088 16672 70100
rect 6886 70060 16672 70088
rect 2038 69980 2044 70032
rect 2096 69980 2102 70032
rect 6886 70020 6914 70060
rect 16666 70048 16672 70060
rect 16724 70048 16730 70100
rect 2516 69992 6914 70020
rect 2516 69961 2544 69992
rect 2501 69955 2559 69961
rect 2501 69921 2513 69955
rect 2547 69921 2559 69955
rect 2501 69915 2559 69921
rect 12434 69912 12440 69964
rect 12492 69952 12498 69964
rect 13722 69952 13728 69964
rect 12492 69924 13728 69952
rect 12492 69912 12498 69924
rect 13722 69912 13728 69924
rect 13780 69952 13786 69964
rect 15289 69955 15347 69961
rect 15289 69952 15301 69955
rect 13780 69924 15301 69952
rect 13780 69912 13786 69924
rect 15289 69921 15301 69924
rect 15335 69921 15347 69955
rect 15289 69915 15347 69921
rect 2958 69844 2964 69896
rect 3016 69844 3022 69896
rect 3970 69844 3976 69896
rect 4028 69844 4034 69896
rect 7006 69844 7012 69896
rect 7064 69884 7070 69896
rect 7101 69887 7159 69893
rect 7101 69884 7113 69887
rect 7064 69856 7113 69884
rect 7064 69844 7070 69856
rect 7101 69853 7113 69856
rect 7147 69853 7159 69887
rect 7101 69847 7159 69853
rect 8294 69844 8300 69896
rect 8352 69884 8358 69896
rect 9125 69887 9183 69893
rect 9125 69884 9137 69887
rect 8352 69856 9137 69884
rect 8352 69844 8358 69856
rect 9125 69853 9137 69856
rect 9171 69853 9183 69887
rect 9125 69847 9183 69853
rect 9306 69844 9312 69896
rect 9364 69884 9370 69896
rect 9401 69887 9459 69893
rect 9401 69884 9413 69887
rect 9364 69856 9413 69884
rect 9364 69844 9370 69856
rect 9401 69853 9413 69856
rect 9447 69853 9459 69887
rect 9401 69847 9459 69853
rect 15010 69844 15016 69896
rect 15068 69844 15074 69896
rect 15102 69844 15108 69896
rect 15160 69884 15166 69896
rect 18049 69887 18107 69893
rect 18049 69884 18061 69887
rect 15160 69856 18061 69884
rect 15160 69844 15166 69856
rect 18049 69853 18061 69856
rect 18095 69853 18107 69887
rect 18049 69847 18107 69853
rect 2593 69819 2651 69825
rect 2593 69785 2605 69819
rect 2639 69816 2651 69819
rect 2976 69816 3004 69844
rect 3786 69816 3792 69828
rect 2639 69788 3792 69816
rect 2639 69785 2651 69788
rect 2593 69779 2651 69785
rect 3786 69776 3792 69788
rect 3844 69776 3850 69828
rect 6546 69776 6552 69828
rect 6604 69816 6610 69828
rect 7346 69819 7404 69825
rect 7346 69816 7358 69819
rect 6604 69788 7358 69816
rect 6604 69776 6610 69788
rect 7346 69785 7358 69788
rect 7392 69785 7404 69819
rect 7346 69779 7404 69785
rect 2498 69708 2504 69760
rect 2556 69708 2562 69760
rect 3053 69751 3111 69757
rect 3053 69717 3065 69751
rect 3099 69748 3111 69751
rect 3421 69751 3479 69757
rect 3421 69748 3433 69751
rect 3099 69720 3433 69748
rect 3099 69717 3111 69720
rect 3053 69711 3111 69717
rect 3421 69717 3433 69720
rect 3467 69748 3479 69751
rect 4157 69751 4215 69757
rect 4157 69748 4169 69751
rect 3467 69720 4169 69748
rect 3467 69717 3479 69720
rect 3421 69711 3479 69717
rect 4157 69717 4169 69720
rect 4203 69748 4215 69751
rect 4617 69751 4675 69757
rect 4617 69748 4629 69751
rect 4203 69720 4629 69748
rect 4203 69717 4215 69720
rect 4157 69711 4215 69717
rect 4617 69717 4629 69720
rect 4663 69748 4675 69751
rect 4985 69751 5043 69757
rect 4985 69748 4997 69751
rect 4663 69720 4997 69748
rect 4663 69717 4675 69720
rect 4617 69711 4675 69717
rect 4985 69717 4997 69720
rect 5031 69748 5043 69751
rect 5258 69748 5264 69760
rect 5031 69720 5264 69748
rect 5031 69717 5043 69720
rect 4985 69711 5043 69717
rect 5258 69708 5264 69720
rect 5316 69708 5322 69760
rect 6638 69708 6644 69760
rect 6696 69748 6702 69760
rect 6822 69748 6828 69760
rect 6696 69720 6828 69748
rect 6696 69708 6702 69720
rect 6822 69708 6828 69720
rect 6880 69708 6886 69760
rect 8481 69751 8539 69757
rect 8481 69717 8493 69751
rect 8527 69748 8539 69751
rect 15470 69748 15476 69760
rect 8527 69720 15476 69748
rect 8527 69717 8539 69720
rect 8481 69711 8539 69717
rect 15470 69708 15476 69720
rect 15528 69708 15534 69760
rect 18230 69708 18236 69760
rect 18288 69708 18294 69760
rect 1104 69658 18860 69680
rect 1104 69606 2610 69658
rect 2662 69606 2674 69658
rect 2726 69606 2738 69658
rect 2790 69606 2802 69658
rect 2854 69606 2866 69658
rect 2918 69606 7610 69658
rect 7662 69606 7674 69658
rect 7726 69606 7738 69658
rect 7790 69606 7802 69658
rect 7854 69606 7866 69658
rect 7918 69606 12610 69658
rect 12662 69606 12674 69658
rect 12726 69606 12738 69658
rect 12790 69606 12802 69658
rect 12854 69606 12866 69658
rect 12918 69606 17610 69658
rect 17662 69606 17674 69658
rect 17726 69606 17738 69658
rect 17790 69606 17802 69658
rect 17854 69606 17866 69658
rect 17918 69606 18860 69658
rect 1104 69584 18860 69606
rect 13170 69544 13176 69556
rect 6886 69516 13176 69544
rect 3970 69436 3976 69488
rect 4028 69476 4034 69488
rect 6886 69476 6914 69516
rect 13170 69504 13176 69516
rect 13228 69504 13234 69556
rect 4028 69448 6914 69476
rect 4028 69436 4034 69448
rect 7466 69436 7472 69488
rect 7524 69476 7530 69488
rect 9922 69479 9980 69485
rect 9922 69476 9934 69479
rect 7524 69448 9934 69476
rect 7524 69436 7530 69448
rect 9922 69445 9934 69448
rect 9968 69445 9980 69479
rect 9922 69439 9980 69445
rect 9122 69368 9128 69420
rect 9180 69408 9186 69420
rect 9677 69411 9735 69417
rect 9677 69408 9689 69411
rect 9180 69380 9689 69408
rect 9180 69368 9186 69380
rect 9677 69377 9689 69380
rect 9723 69377 9735 69411
rect 9677 69371 9735 69377
rect 11054 69164 11060 69216
rect 11112 69164 11118 69216
rect 1104 69114 18860 69136
rect 1104 69062 1950 69114
rect 2002 69062 2014 69114
rect 2066 69062 2078 69114
rect 2130 69062 2142 69114
rect 2194 69062 2206 69114
rect 2258 69062 6950 69114
rect 7002 69062 7014 69114
rect 7066 69062 7078 69114
rect 7130 69062 7142 69114
rect 7194 69062 7206 69114
rect 7258 69062 11950 69114
rect 12002 69062 12014 69114
rect 12066 69062 12078 69114
rect 12130 69062 12142 69114
rect 12194 69062 12206 69114
rect 12258 69062 16950 69114
rect 17002 69062 17014 69114
rect 17066 69062 17078 69114
rect 17130 69062 17142 69114
rect 17194 69062 17206 69114
rect 17258 69062 18860 69114
rect 1104 69040 18860 69062
rect 9122 68824 9128 68876
rect 9180 68824 9186 68876
rect 13814 68756 13820 68808
rect 13872 68796 13878 68808
rect 14274 68796 14280 68808
rect 13872 68768 14280 68796
rect 13872 68756 13878 68768
rect 14274 68756 14280 68768
rect 14332 68756 14338 68808
rect 9392 68731 9450 68737
rect 9392 68697 9404 68731
rect 9438 68728 9450 68731
rect 9582 68728 9588 68740
rect 9438 68700 9588 68728
rect 9438 68697 9450 68700
rect 9392 68691 9450 68697
rect 9582 68688 9588 68700
rect 9640 68688 9646 68740
rect 14550 68737 14556 68740
rect 14544 68691 14556 68737
rect 14550 68688 14556 68691
rect 14608 68688 14614 68740
rect 10502 68620 10508 68672
rect 10560 68620 10566 68672
rect 15654 68620 15660 68672
rect 15712 68620 15718 68672
rect 1104 68570 18860 68592
rect 1104 68518 2610 68570
rect 2662 68518 2674 68570
rect 2726 68518 2738 68570
rect 2790 68518 2802 68570
rect 2854 68518 2866 68570
rect 2918 68518 7610 68570
rect 7662 68518 7674 68570
rect 7726 68518 7738 68570
rect 7790 68518 7802 68570
rect 7854 68518 7866 68570
rect 7918 68518 12610 68570
rect 12662 68518 12674 68570
rect 12726 68518 12738 68570
rect 12790 68518 12802 68570
rect 12854 68518 12866 68570
rect 12918 68518 17610 68570
rect 17662 68518 17674 68570
rect 17726 68518 17738 68570
rect 17790 68518 17802 68570
rect 17854 68518 17866 68570
rect 17918 68518 18860 68570
rect 1104 68496 18860 68518
rect 6178 68280 6184 68332
rect 6236 68320 6242 68332
rect 14918 68320 14924 68332
rect 6236 68292 14924 68320
rect 6236 68280 6242 68292
rect 14918 68280 14924 68292
rect 14976 68280 14982 68332
rect 1104 68026 18860 68048
rect 1104 67974 1950 68026
rect 2002 67974 2014 68026
rect 2066 67974 2078 68026
rect 2130 67974 2142 68026
rect 2194 67974 2206 68026
rect 2258 67974 6950 68026
rect 7002 67974 7014 68026
rect 7066 67974 7078 68026
rect 7130 67974 7142 68026
rect 7194 67974 7206 68026
rect 7258 67974 11950 68026
rect 12002 67974 12014 68026
rect 12066 67974 12078 68026
rect 12130 67974 12142 68026
rect 12194 67974 12206 68026
rect 12258 67974 16950 68026
rect 17002 67974 17014 68026
rect 17066 67974 17078 68026
rect 17130 67974 17142 68026
rect 17194 67974 17206 68026
rect 17258 67974 18860 68026
rect 1104 67952 18860 67974
rect 10410 67804 10416 67856
rect 10468 67844 10474 67856
rect 12437 67847 12495 67853
rect 12437 67844 12449 67847
rect 10468 67816 12449 67844
rect 10468 67804 10474 67816
rect 12437 67813 12449 67816
rect 12483 67813 12495 67847
rect 12437 67807 12495 67813
rect 18230 67804 18236 67856
rect 18288 67804 18294 67856
rect 12621 67711 12679 67717
rect 12621 67708 12633 67711
rect 12084 67680 12633 67708
rect 12084 67652 12112 67680
rect 12621 67677 12633 67680
rect 12667 67677 12679 67711
rect 12621 67671 12679 67677
rect 17402 67668 17408 67720
rect 17460 67708 17466 67720
rect 18049 67711 18107 67717
rect 18049 67708 18061 67711
rect 17460 67680 18061 67708
rect 17460 67668 17466 67680
rect 18049 67677 18061 67680
rect 18095 67677 18107 67711
rect 18049 67671 18107 67677
rect 12066 67600 12072 67652
rect 12124 67600 12130 67652
rect 1104 67482 18860 67504
rect 1104 67430 2610 67482
rect 2662 67430 2674 67482
rect 2726 67430 2738 67482
rect 2790 67430 2802 67482
rect 2854 67430 2866 67482
rect 2918 67430 7610 67482
rect 7662 67430 7674 67482
rect 7726 67430 7738 67482
rect 7790 67430 7802 67482
rect 7854 67430 7866 67482
rect 7918 67430 12610 67482
rect 12662 67430 12674 67482
rect 12726 67430 12738 67482
rect 12790 67430 12802 67482
rect 12854 67430 12866 67482
rect 12918 67430 17610 67482
rect 17662 67430 17674 67482
rect 17726 67430 17738 67482
rect 17790 67430 17802 67482
rect 17854 67430 17866 67482
rect 17918 67430 18860 67482
rect 1104 67408 18860 67430
rect 11790 67260 11796 67312
rect 11848 67300 11854 67312
rect 11848 67272 18184 67300
rect 11848 67260 11854 67272
rect 3694 67192 3700 67244
rect 3752 67232 3758 67244
rect 7929 67235 7987 67241
rect 7929 67232 7941 67235
rect 3752 67204 7941 67232
rect 3752 67192 3758 67204
rect 7929 67201 7941 67204
rect 7975 67201 7987 67235
rect 7929 67195 7987 67201
rect 13998 67192 14004 67244
rect 14056 67232 14062 67244
rect 17957 67235 18015 67241
rect 17957 67232 17969 67235
rect 14056 67204 17969 67232
rect 14056 67192 14062 67204
rect 17957 67201 17969 67204
rect 18003 67201 18015 67235
rect 17957 67195 18015 67201
rect 16022 67124 16028 67176
rect 16080 67164 16086 67176
rect 16482 67164 16488 67176
rect 16080 67136 16488 67164
rect 16080 67124 16086 67136
rect 16482 67124 16488 67136
rect 16540 67164 16546 67176
rect 18156 67173 18184 67272
rect 17313 67167 17371 67173
rect 17313 67164 17325 67167
rect 16540 67136 17325 67164
rect 16540 67124 16546 67136
rect 17313 67133 17325 67136
rect 17359 67164 17371 67167
rect 18049 67167 18107 67173
rect 18049 67164 18061 67167
rect 17359 67136 18061 67164
rect 17359 67133 17371 67136
rect 17313 67127 17371 67133
rect 18049 67133 18061 67136
rect 18095 67133 18107 67167
rect 18049 67127 18107 67133
rect 18141 67167 18199 67173
rect 18141 67133 18153 67167
rect 18187 67133 18199 67167
rect 18141 67127 18199 67133
rect 1210 66988 1216 67040
rect 1268 67028 1274 67040
rect 8113 67031 8171 67037
rect 8113 67028 8125 67031
rect 1268 67000 8125 67028
rect 1268 66988 1274 67000
rect 8113 66997 8125 67000
rect 8159 66997 8171 67031
rect 8113 66991 8171 66997
rect 17310 66988 17316 67040
rect 17368 67028 17374 67040
rect 17589 67031 17647 67037
rect 17589 67028 17601 67031
rect 17368 67000 17601 67028
rect 17368 66988 17374 67000
rect 17589 66997 17601 67000
rect 17635 66997 17647 67031
rect 17589 66991 17647 66997
rect 1104 66938 18860 66960
rect 1104 66886 1950 66938
rect 2002 66886 2014 66938
rect 2066 66886 2078 66938
rect 2130 66886 2142 66938
rect 2194 66886 2206 66938
rect 2258 66886 6950 66938
rect 7002 66886 7014 66938
rect 7066 66886 7078 66938
rect 7130 66886 7142 66938
rect 7194 66886 7206 66938
rect 7258 66886 11950 66938
rect 12002 66886 12014 66938
rect 12066 66886 12078 66938
rect 12130 66886 12142 66938
rect 12194 66886 12206 66938
rect 12258 66886 16950 66938
rect 17002 66886 17014 66938
rect 17066 66886 17078 66938
rect 17130 66886 17142 66938
rect 17194 66886 17206 66938
rect 17258 66886 18860 66938
rect 1104 66864 18860 66886
rect 1104 66394 18860 66416
rect 1104 66342 2610 66394
rect 2662 66342 2674 66394
rect 2726 66342 2738 66394
rect 2790 66342 2802 66394
rect 2854 66342 2866 66394
rect 2918 66342 7610 66394
rect 7662 66342 7674 66394
rect 7726 66342 7738 66394
rect 7790 66342 7802 66394
rect 7854 66342 7866 66394
rect 7918 66342 12610 66394
rect 12662 66342 12674 66394
rect 12726 66342 12738 66394
rect 12790 66342 12802 66394
rect 12854 66342 12866 66394
rect 12918 66342 17610 66394
rect 17662 66342 17674 66394
rect 17726 66342 17738 66394
rect 17790 66342 17802 66394
rect 17854 66342 17866 66394
rect 17918 66342 18860 66394
rect 1104 66320 18860 66342
rect 13808 66215 13866 66221
rect 13808 66181 13820 66215
rect 13854 66212 13866 66215
rect 13906 66212 13912 66224
rect 13854 66184 13912 66212
rect 13854 66181 13866 66184
rect 13808 66175 13866 66181
rect 13906 66172 13912 66184
rect 13964 66172 13970 66224
rect 16574 66172 16580 66224
rect 16632 66212 16638 66224
rect 17494 66212 17500 66224
rect 16632 66184 17500 66212
rect 16632 66172 16638 66184
rect 17494 66172 17500 66184
rect 17552 66212 17558 66224
rect 17957 66215 18015 66221
rect 17957 66212 17969 66215
rect 17552 66184 17969 66212
rect 17552 66172 17558 66184
rect 17957 66181 17969 66184
rect 18003 66181 18015 66215
rect 17957 66175 18015 66181
rect 13541 66147 13599 66153
rect 13541 66113 13553 66147
rect 13587 66144 13599 66147
rect 13630 66144 13636 66156
rect 13587 66116 13636 66144
rect 13587 66113 13599 66116
rect 13541 66107 13599 66113
rect 13630 66104 13636 66116
rect 13688 66104 13694 66156
rect 17402 66104 17408 66156
rect 17460 66144 17466 66156
rect 17773 66147 17831 66153
rect 17773 66144 17785 66147
rect 17460 66116 17785 66144
rect 17460 66104 17466 66116
rect 17773 66113 17785 66116
rect 17819 66113 17831 66147
rect 17773 66107 17831 66113
rect 18049 66079 18107 66085
rect 18049 66045 18061 66079
rect 18095 66045 18107 66079
rect 18049 66039 18107 66045
rect 18064 66008 18092 66039
rect 14752 65980 18092 66008
rect 14274 65900 14280 65952
rect 14332 65940 14338 65952
rect 14752 65940 14780 65980
rect 14332 65912 14780 65940
rect 14332 65900 14338 65912
rect 14826 65900 14832 65952
rect 14884 65940 14890 65952
rect 14921 65943 14979 65949
rect 14921 65940 14933 65943
rect 14884 65912 14933 65940
rect 14884 65900 14890 65912
rect 14921 65909 14933 65912
rect 14967 65909 14979 65943
rect 14921 65903 14979 65909
rect 17494 65900 17500 65952
rect 17552 65900 17558 65952
rect 1104 65850 18860 65872
rect 1104 65798 1950 65850
rect 2002 65798 2014 65850
rect 2066 65798 2078 65850
rect 2130 65798 2142 65850
rect 2194 65798 2206 65850
rect 2258 65798 6950 65850
rect 7002 65798 7014 65850
rect 7066 65798 7078 65850
rect 7130 65798 7142 65850
rect 7194 65798 7206 65850
rect 7258 65798 11950 65850
rect 12002 65798 12014 65850
rect 12066 65798 12078 65850
rect 12130 65798 12142 65850
rect 12194 65798 12206 65850
rect 12258 65798 16950 65850
rect 17002 65798 17014 65850
rect 17066 65798 17078 65850
rect 17130 65798 17142 65850
rect 17194 65798 17206 65850
rect 17258 65798 18860 65850
rect 1104 65776 18860 65798
rect 4062 65628 4068 65680
rect 4120 65628 4126 65680
rect 11790 65628 11796 65680
rect 11848 65628 11854 65680
rect 18230 65628 18236 65680
rect 18288 65628 18294 65680
rect 4614 65560 4620 65612
rect 4672 65560 4678 65612
rect 11514 65560 11520 65612
rect 11572 65600 11578 65612
rect 11808 65600 11836 65628
rect 11572 65572 12112 65600
rect 11572 65560 11578 65572
rect 11790 65492 11796 65544
rect 11848 65492 11854 65544
rect 11882 65492 11888 65544
rect 11940 65492 11946 65544
rect 12084 65541 12112 65572
rect 12069 65535 12127 65541
rect 12069 65501 12081 65535
rect 12115 65501 12127 65535
rect 12069 65495 12127 65501
rect 15562 65492 15568 65544
rect 15620 65532 15626 65544
rect 16206 65532 16212 65544
rect 15620 65504 16212 65532
rect 15620 65492 15626 65504
rect 16206 65492 16212 65504
rect 16264 65532 16270 65544
rect 18049 65535 18107 65541
rect 18049 65532 18061 65535
rect 16264 65504 18061 65532
rect 16264 65492 16270 65504
rect 18049 65501 18061 65504
rect 18095 65501 18107 65535
rect 18049 65495 18107 65501
rect 4341 65467 4399 65473
rect 4341 65433 4353 65467
rect 4387 65464 4399 65467
rect 9490 65464 9496 65476
rect 4387 65436 9496 65464
rect 4387 65433 4399 65436
rect 4341 65427 4399 65433
rect 9490 65424 9496 65436
rect 9548 65424 9554 65476
rect 11241 65467 11299 65473
rect 11241 65433 11253 65467
rect 11287 65464 11299 65467
rect 11422 65464 11428 65476
rect 11287 65436 11428 65464
rect 11287 65433 11299 65436
rect 11241 65427 11299 65433
rect 11422 65424 11428 65436
rect 11480 65464 11486 65476
rect 12529 65467 12587 65473
rect 12529 65464 12541 65467
rect 11480 65436 12541 65464
rect 11480 65424 11486 65436
rect 12529 65433 12541 65436
rect 12575 65433 12587 65467
rect 12529 65427 12587 65433
rect 3602 65356 3608 65408
rect 3660 65396 3666 65408
rect 4525 65399 4583 65405
rect 4525 65396 4537 65399
rect 3660 65368 4537 65396
rect 3660 65356 3666 65368
rect 4525 65365 4537 65368
rect 4571 65365 4583 65399
rect 4525 65359 4583 65365
rect 1104 65306 18860 65328
rect 1104 65254 2610 65306
rect 2662 65254 2674 65306
rect 2726 65254 2738 65306
rect 2790 65254 2802 65306
rect 2854 65254 2866 65306
rect 2918 65254 7610 65306
rect 7662 65254 7674 65306
rect 7726 65254 7738 65306
rect 7790 65254 7802 65306
rect 7854 65254 7866 65306
rect 7918 65254 12610 65306
rect 12662 65254 12674 65306
rect 12726 65254 12738 65306
rect 12790 65254 12802 65306
rect 12854 65254 12866 65306
rect 12918 65254 17610 65306
rect 17662 65254 17674 65306
rect 17726 65254 17738 65306
rect 17790 65254 17802 65306
rect 17854 65254 17866 65306
rect 17918 65254 18860 65306
rect 1104 65232 18860 65254
rect 7929 65195 7987 65201
rect 7929 65161 7941 65195
rect 7975 65192 7987 65195
rect 8294 65192 8300 65204
rect 7975 65164 8300 65192
rect 7975 65161 7987 65164
rect 7929 65155 7987 65161
rect 8294 65152 8300 65164
rect 8352 65152 8358 65204
rect 14366 65152 14372 65204
rect 14424 65192 14430 65204
rect 15102 65192 15108 65204
rect 14424 65164 15108 65192
rect 14424 65152 14430 65164
rect 15102 65152 15108 65164
rect 15160 65152 15166 65204
rect 17402 65152 17408 65204
rect 17460 65192 17466 65204
rect 17586 65192 17592 65204
rect 17460 65164 17592 65192
rect 17460 65152 17466 65164
rect 17586 65152 17592 65164
rect 17644 65152 17650 65204
rect 13256 65127 13314 65133
rect 13256 65093 13268 65127
rect 13302 65124 13314 65127
rect 19150 65124 19156 65136
rect 13302 65096 19156 65124
rect 13302 65093 13314 65096
rect 13256 65087 13314 65093
rect 19150 65084 19156 65096
rect 19208 65084 19214 65136
rect 7926 65016 7932 65068
rect 7984 65016 7990 65068
rect 8297 65059 8355 65065
rect 8297 65025 8309 65059
rect 8343 65056 8355 65059
rect 8662 65056 8668 65068
rect 8343 65028 8668 65056
rect 8343 65025 8355 65028
rect 8297 65019 8355 65025
rect 8662 65016 8668 65028
rect 8720 65016 8726 65068
rect 18141 65059 18199 65065
rect 18141 65025 18153 65059
rect 18187 65056 18199 65059
rect 19334 65056 19340 65068
rect 18187 65028 19340 65056
rect 18187 65025 18199 65028
rect 18141 65019 18199 65025
rect 19334 65016 19340 65028
rect 19392 65016 19398 65068
rect 7944 64988 7972 65016
rect 8389 64991 8447 64997
rect 8389 64988 8401 64991
rect 7944 64960 8401 64988
rect 8220 64852 8248 64960
rect 8389 64957 8401 64960
rect 8435 64957 8447 64991
rect 8573 64991 8631 64997
rect 8573 64988 8585 64991
rect 8389 64951 8447 64957
rect 8496 64960 8585 64988
rect 8294 64880 8300 64932
rect 8352 64920 8358 64932
rect 8496 64920 8524 64960
rect 8573 64957 8585 64960
rect 8619 64988 8631 64991
rect 12434 64988 12440 65000
rect 8619 64960 12440 64988
rect 8619 64957 8631 64960
rect 8573 64951 8631 64957
rect 12434 64948 12440 64960
rect 12492 64948 12498 65000
rect 12989 64991 13047 64997
rect 12989 64957 13001 64991
rect 13035 64957 13047 64991
rect 12989 64951 13047 64957
rect 11882 64920 11888 64932
rect 8352 64892 8524 64920
rect 8588 64892 11888 64920
rect 8352 64880 8358 64892
rect 8588 64852 8616 64892
rect 11882 64880 11888 64892
rect 11940 64880 11946 64932
rect 8220 64824 8616 64852
rect 13004 64852 13032 64951
rect 17034 64880 17040 64932
rect 17092 64920 17098 64932
rect 17402 64920 17408 64932
rect 17092 64892 17408 64920
rect 17092 64880 17098 64892
rect 17402 64880 17408 64892
rect 17460 64880 17466 64932
rect 18325 64923 18383 64929
rect 18325 64889 18337 64923
rect 18371 64920 18383 64923
rect 18414 64920 18420 64932
rect 18371 64892 18420 64920
rect 18371 64889 18383 64892
rect 18325 64883 18383 64889
rect 18414 64880 18420 64892
rect 18472 64880 18478 64932
rect 13722 64852 13728 64864
rect 13004 64824 13728 64852
rect 13722 64812 13728 64824
rect 13780 64812 13786 64864
rect 16482 64812 16488 64864
rect 16540 64852 16546 64864
rect 16942 64852 16948 64864
rect 16540 64824 16948 64852
rect 16540 64812 16546 64824
rect 16942 64812 16948 64824
rect 17000 64812 17006 64864
rect 1104 64762 18860 64784
rect 1104 64710 1950 64762
rect 2002 64710 2014 64762
rect 2066 64710 2078 64762
rect 2130 64710 2142 64762
rect 2194 64710 2206 64762
rect 2258 64710 6950 64762
rect 7002 64710 7014 64762
rect 7066 64710 7078 64762
rect 7130 64710 7142 64762
rect 7194 64710 7206 64762
rect 7258 64710 11950 64762
rect 12002 64710 12014 64762
rect 12066 64710 12078 64762
rect 12130 64710 12142 64762
rect 12194 64710 12206 64762
rect 12258 64710 16950 64762
rect 17002 64710 17014 64762
rect 17066 64710 17078 64762
rect 17130 64710 17142 64762
rect 17194 64710 17206 64762
rect 17258 64710 18860 64762
rect 1104 64688 18860 64710
rect 13262 64648 13268 64660
rect 6886 64620 13268 64648
rect 2593 64447 2651 64453
rect 2593 64413 2605 64447
rect 2639 64444 2651 64447
rect 6886 64444 6914 64620
rect 13262 64608 13268 64620
rect 13320 64608 13326 64660
rect 8110 64472 8116 64524
rect 8168 64512 8174 64524
rect 8386 64512 8392 64524
rect 8168 64484 8392 64512
rect 8168 64472 8174 64484
rect 8386 64472 8392 64484
rect 8444 64472 8450 64524
rect 2639 64416 6914 64444
rect 2639 64413 2651 64416
rect 2593 64407 2651 64413
rect 7282 64404 7288 64456
rect 7340 64444 7346 64456
rect 11793 64447 11851 64453
rect 11793 64444 11805 64447
rect 7340 64416 11805 64444
rect 7340 64404 7346 64416
rect 11793 64413 11805 64416
rect 11839 64444 11851 64447
rect 13722 64444 13728 64456
rect 11839 64416 13728 64444
rect 11839 64413 11851 64416
rect 11793 64407 11851 64413
rect 13722 64404 13728 64416
rect 13780 64404 13786 64456
rect 11330 64336 11336 64388
rect 11388 64376 11394 64388
rect 12038 64379 12096 64385
rect 12038 64376 12050 64379
rect 11388 64348 12050 64376
rect 11388 64336 11394 64348
rect 12038 64345 12050 64348
rect 12084 64345 12096 64379
rect 12038 64339 12096 64345
rect 1762 64268 1768 64320
rect 1820 64308 1826 64320
rect 2409 64311 2467 64317
rect 2409 64308 2421 64311
rect 1820 64280 2421 64308
rect 1820 64268 1826 64280
rect 2409 64277 2421 64280
rect 2455 64277 2467 64311
rect 2409 64271 2467 64277
rect 7926 64268 7932 64320
rect 7984 64308 7990 64320
rect 8110 64308 8116 64320
rect 7984 64280 8116 64308
rect 7984 64268 7990 64280
rect 8110 64268 8116 64280
rect 8168 64268 8174 64320
rect 13173 64311 13231 64317
rect 13173 64277 13185 64311
rect 13219 64308 13231 64311
rect 13906 64308 13912 64320
rect 13219 64280 13912 64308
rect 13219 64277 13231 64280
rect 13173 64271 13231 64277
rect 13906 64268 13912 64280
rect 13964 64268 13970 64320
rect 1104 64218 18860 64240
rect 1104 64166 2610 64218
rect 2662 64166 2674 64218
rect 2726 64166 2738 64218
rect 2790 64166 2802 64218
rect 2854 64166 2866 64218
rect 2918 64166 7610 64218
rect 7662 64166 7674 64218
rect 7726 64166 7738 64218
rect 7790 64166 7802 64218
rect 7854 64166 7866 64218
rect 7918 64166 12610 64218
rect 12662 64166 12674 64218
rect 12726 64166 12738 64218
rect 12790 64166 12802 64218
rect 12854 64166 12866 64218
rect 12918 64166 17610 64218
rect 17662 64166 17674 64218
rect 17726 64166 17738 64218
rect 17790 64166 17802 64218
rect 17854 64166 17866 64218
rect 17918 64166 18860 64218
rect 1104 64144 18860 64166
rect 11238 63928 11244 63980
rect 11296 63968 11302 63980
rect 12253 63971 12311 63977
rect 12253 63968 12265 63971
rect 11296 63940 12265 63968
rect 11296 63928 11302 63940
rect 12253 63937 12265 63940
rect 12299 63937 12311 63971
rect 12253 63931 12311 63937
rect 18049 63971 18107 63977
rect 18049 63937 18061 63971
rect 18095 63968 18107 63971
rect 18506 63968 18512 63980
rect 18095 63940 18512 63968
rect 18095 63937 18107 63940
rect 18049 63931 18107 63937
rect 18506 63928 18512 63940
rect 18564 63928 18570 63980
rect 12345 63903 12403 63909
rect 12345 63869 12357 63903
rect 12391 63869 12403 63903
rect 12345 63863 12403 63869
rect 12529 63903 12587 63909
rect 12529 63869 12541 63903
rect 12575 63900 12587 63903
rect 15378 63900 15384 63912
rect 12575 63872 15384 63900
rect 12575 63869 12587 63872
rect 12529 63863 12587 63869
rect 9674 63792 9680 63844
rect 9732 63832 9738 63844
rect 11885 63835 11943 63841
rect 11885 63832 11897 63835
rect 9732 63804 11897 63832
rect 9732 63792 9738 63804
rect 11885 63801 11897 63804
rect 11931 63801 11943 63835
rect 11885 63795 11943 63801
rect 9950 63724 9956 63776
rect 10008 63764 10014 63776
rect 10689 63767 10747 63773
rect 10689 63764 10701 63767
rect 10008 63736 10701 63764
rect 10008 63724 10014 63736
rect 10689 63733 10701 63736
rect 10735 63764 10747 63767
rect 11057 63767 11115 63773
rect 11057 63764 11069 63767
rect 10735 63736 11069 63764
rect 10735 63733 10747 63736
rect 10689 63727 10747 63733
rect 11057 63733 11069 63736
rect 11103 63764 11115 63767
rect 12360 63764 12388 63863
rect 15378 63860 15384 63872
rect 15436 63860 15442 63912
rect 12897 63767 12955 63773
rect 12897 63764 12909 63767
rect 11103 63736 12909 63764
rect 11103 63733 11115 63736
rect 11057 63727 11115 63733
rect 12897 63733 12909 63736
rect 12943 63764 12955 63767
rect 13265 63767 13323 63773
rect 13265 63764 13277 63767
rect 12943 63736 13277 63764
rect 12943 63733 12955 63736
rect 12897 63727 12955 63733
rect 13265 63733 13277 63736
rect 13311 63764 13323 63767
rect 13633 63767 13691 63773
rect 13633 63764 13645 63767
rect 13311 63736 13645 63764
rect 13311 63733 13323 63736
rect 13265 63727 13323 63733
rect 13633 63733 13645 63736
rect 13679 63733 13691 63767
rect 13633 63727 13691 63733
rect 18230 63724 18236 63776
rect 18288 63724 18294 63776
rect 1104 63674 18860 63696
rect 1104 63622 1950 63674
rect 2002 63622 2014 63674
rect 2066 63622 2078 63674
rect 2130 63622 2142 63674
rect 2194 63622 2206 63674
rect 2258 63622 6950 63674
rect 7002 63622 7014 63674
rect 7066 63622 7078 63674
rect 7130 63622 7142 63674
rect 7194 63622 7206 63674
rect 7258 63622 11950 63674
rect 12002 63622 12014 63674
rect 12066 63622 12078 63674
rect 12130 63622 12142 63674
rect 12194 63622 12206 63674
rect 12258 63622 16950 63674
rect 17002 63622 17014 63674
rect 17066 63622 17078 63674
rect 17130 63622 17142 63674
rect 17194 63622 17206 63674
rect 17258 63622 18860 63674
rect 1104 63600 18860 63622
rect 13906 63520 13912 63572
rect 13964 63560 13970 63572
rect 14918 63560 14924 63572
rect 13964 63532 14924 63560
rect 13964 63520 13970 63532
rect 14918 63520 14924 63532
rect 14976 63520 14982 63572
rect 6546 63452 6552 63504
rect 6604 63492 6610 63504
rect 7282 63492 7288 63504
rect 6604 63464 7288 63492
rect 6604 63452 6610 63464
rect 7282 63452 7288 63464
rect 7340 63452 7346 63504
rect 14550 63452 14556 63504
rect 14608 63492 14614 63504
rect 16301 63495 16359 63501
rect 16301 63492 16313 63495
rect 14608 63464 16313 63492
rect 14608 63452 14614 63464
rect 16301 63461 16313 63464
rect 16347 63461 16359 63495
rect 16301 63455 16359 63461
rect 14277 63359 14335 63365
rect 14277 63325 14289 63359
rect 14323 63356 14335 63359
rect 15562 63356 15568 63368
rect 14323 63328 15568 63356
rect 14323 63325 14335 63328
rect 14277 63319 14335 63325
rect 15562 63316 15568 63328
rect 15620 63316 15626 63368
rect 16482 63316 16488 63368
rect 16540 63316 16546 63368
rect 6273 63291 6331 63297
rect 6273 63257 6285 63291
rect 6319 63288 6331 63291
rect 9674 63288 9680 63300
rect 6319 63260 9680 63288
rect 6319 63257 6331 63260
rect 6273 63251 6331 63257
rect 9674 63248 9680 63260
rect 9732 63248 9738 63300
rect 6362 63180 6368 63232
rect 6420 63180 6426 63232
rect 14458 63180 14464 63232
rect 14516 63180 14522 63232
rect 1104 63130 18860 63152
rect 1104 63078 2610 63130
rect 2662 63078 2674 63130
rect 2726 63078 2738 63130
rect 2790 63078 2802 63130
rect 2854 63078 2866 63130
rect 2918 63078 7610 63130
rect 7662 63078 7674 63130
rect 7726 63078 7738 63130
rect 7790 63078 7802 63130
rect 7854 63078 7866 63130
rect 7918 63078 12610 63130
rect 12662 63078 12674 63130
rect 12726 63078 12738 63130
rect 12790 63078 12802 63130
rect 12854 63078 12866 63130
rect 12918 63078 17610 63130
rect 17662 63078 17674 63130
rect 17726 63078 17738 63130
rect 17790 63078 17802 63130
rect 17854 63078 17866 63130
rect 17918 63078 18860 63130
rect 1104 63056 18860 63078
rect 5442 62976 5448 63028
rect 5500 63016 5506 63028
rect 7929 63019 7987 63025
rect 7929 63016 7941 63019
rect 5500 62988 7941 63016
rect 5500 62976 5506 62988
rect 7929 62985 7941 62988
rect 7975 63016 7987 63019
rect 11146 63016 11152 63028
rect 7975 62988 11152 63016
rect 7975 62985 7987 62988
rect 7929 62979 7987 62985
rect 11146 62976 11152 62988
rect 11204 62976 11210 63028
rect 6546 62840 6552 62892
rect 6604 62840 6610 62892
rect 6805 62883 6863 62889
rect 6805 62880 6817 62883
rect 6656 62852 6817 62880
rect 5629 62815 5687 62821
rect 5629 62781 5641 62815
rect 5675 62812 5687 62815
rect 5905 62815 5963 62821
rect 5905 62812 5917 62815
rect 5675 62784 5917 62812
rect 5675 62781 5687 62784
rect 5629 62775 5687 62781
rect 5905 62781 5917 62784
rect 5951 62812 5963 62815
rect 6656 62812 6684 62852
rect 6805 62849 6817 62852
rect 6851 62880 6863 62883
rect 6851 62852 8432 62880
rect 6851 62849 6863 62852
rect 6805 62843 6863 62849
rect 5951 62784 6684 62812
rect 5951 62781 5963 62784
rect 5905 62775 5963 62781
rect 8404 62685 8432 62852
rect 9582 62772 9588 62824
rect 9640 62812 9646 62824
rect 19058 62812 19064 62824
rect 9640 62784 19064 62812
rect 9640 62772 9646 62784
rect 19058 62772 19064 62784
rect 19116 62772 19122 62824
rect 8389 62679 8447 62685
rect 8389 62645 8401 62679
rect 8435 62676 8447 62679
rect 8754 62676 8760 62688
rect 8435 62648 8760 62676
rect 8435 62645 8447 62648
rect 8389 62639 8447 62645
rect 8754 62636 8760 62648
rect 8812 62636 8818 62688
rect 1104 62586 18860 62608
rect 1104 62534 1950 62586
rect 2002 62534 2014 62586
rect 2066 62534 2078 62586
rect 2130 62534 2142 62586
rect 2194 62534 2206 62586
rect 2258 62534 6950 62586
rect 7002 62534 7014 62586
rect 7066 62534 7078 62586
rect 7130 62534 7142 62586
rect 7194 62534 7206 62586
rect 7258 62534 11950 62586
rect 12002 62534 12014 62586
rect 12066 62534 12078 62586
rect 12130 62534 12142 62586
rect 12194 62534 12206 62586
rect 12258 62534 16950 62586
rect 17002 62534 17014 62586
rect 17066 62534 17078 62586
rect 17130 62534 17142 62586
rect 17194 62534 17206 62586
rect 17258 62534 18860 62586
rect 1104 62512 18860 62534
rect 4154 62432 4160 62484
rect 4212 62472 4218 62484
rect 13814 62472 13820 62484
rect 4212 62444 13820 62472
rect 4212 62432 4218 62444
rect 13814 62432 13820 62444
rect 13872 62432 13878 62484
rect 11146 62364 11152 62416
rect 11204 62404 11210 62416
rect 11790 62404 11796 62416
rect 11204 62376 11796 62404
rect 11204 62364 11210 62376
rect 11790 62364 11796 62376
rect 11848 62364 11854 62416
rect 18049 62271 18107 62277
rect 18049 62237 18061 62271
rect 18095 62268 18107 62271
rect 18598 62268 18604 62280
rect 18095 62240 18604 62268
rect 18095 62237 18107 62240
rect 18049 62231 18107 62237
rect 18598 62228 18604 62240
rect 18656 62228 18662 62280
rect 4246 62160 4252 62212
rect 4304 62160 4310 62212
rect 4338 62092 4344 62144
rect 4396 62092 4402 62144
rect 18230 62092 18236 62144
rect 18288 62092 18294 62144
rect 1104 62042 18860 62064
rect 1104 61990 2610 62042
rect 2662 61990 2674 62042
rect 2726 61990 2738 62042
rect 2790 61990 2802 62042
rect 2854 61990 2866 62042
rect 2918 61990 7610 62042
rect 7662 61990 7674 62042
rect 7726 61990 7738 62042
rect 7790 61990 7802 62042
rect 7854 61990 7866 62042
rect 7918 61990 12610 62042
rect 12662 61990 12674 62042
rect 12726 61990 12738 62042
rect 12790 61990 12802 62042
rect 12854 61990 12866 62042
rect 12918 61990 17610 62042
rect 17662 61990 17674 62042
rect 17726 61990 17738 62042
rect 17790 61990 17802 62042
rect 17854 61990 17866 62042
rect 17918 61990 18860 62042
rect 1104 61968 18860 61990
rect 11701 61931 11759 61937
rect 11701 61897 11713 61931
rect 11747 61928 11759 61931
rect 16482 61928 16488 61940
rect 11747 61900 16488 61928
rect 11747 61897 11759 61900
rect 11701 61891 11759 61897
rect 16482 61888 16488 61900
rect 16540 61888 16546 61940
rect 12069 61863 12127 61869
rect 12069 61829 12081 61863
rect 12115 61860 12127 61863
rect 15654 61860 15660 61872
rect 12115 61832 15660 61860
rect 12115 61829 12127 61832
rect 12069 61823 12127 61829
rect 15654 61820 15660 61832
rect 15712 61820 15718 61872
rect 12342 61792 12348 61804
rect 12176 61764 12348 61792
rect 11606 61684 11612 61736
rect 11664 61724 11670 61736
rect 12176 61733 12204 61764
rect 12342 61752 12348 61764
rect 12400 61752 12406 61804
rect 12161 61727 12219 61733
rect 12161 61724 12173 61727
rect 11664 61696 12173 61724
rect 11664 61684 11670 61696
rect 12161 61693 12173 61696
rect 12207 61693 12219 61727
rect 12161 61687 12219 61693
rect 12253 61727 12311 61733
rect 12253 61693 12265 61727
rect 12299 61724 12311 61727
rect 13538 61724 13544 61736
rect 12299 61696 13544 61724
rect 12299 61693 12311 61696
rect 12253 61687 12311 61693
rect 13538 61684 13544 61696
rect 13596 61724 13602 61736
rect 14274 61724 14280 61736
rect 13596 61696 14280 61724
rect 13596 61684 13602 61696
rect 14274 61684 14280 61696
rect 14332 61684 14338 61736
rect 1104 61498 18860 61520
rect 1104 61446 1950 61498
rect 2002 61446 2014 61498
rect 2066 61446 2078 61498
rect 2130 61446 2142 61498
rect 2194 61446 2206 61498
rect 2258 61446 6950 61498
rect 7002 61446 7014 61498
rect 7066 61446 7078 61498
rect 7130 61446 7142 61498
rect 7194 61446 7206 61498
rect 7258 61446 11950 61498
rect 12002 61446 12014 61498
rect 12066 61446 12078 61498
rect 12130 61446 12142 61498
rect 12194 61446 12206 61498
rect 12258 61446 16950 61498
rect 17002 61446 17014 61498
rect 17066 61446 17078 61498
rect 17130 61446 17142 61498
rect 17194 61446 17206 61498
rect 17258 61446 18860 61498
rect 1104 61424 18860 61446
rect 4798 61344 4804 61396
rect 4856 61384 4862 61396
rect 16206 61384 16212 61396
rect 4856 61356 16212 61384
rect 4856 61344 4862 61356
rect 16206 61344 16212 61356
rect 16264 61344 16270 61396
rect 13814 61140 13820 61192
rect 13872 61180 13878 61192
rect 14274 61180 14280 61192
rect 13872 61152 14280 61180
rect 13872 61140 13878 61152
rect 14274 61140 14280 61152
rect 14332 61180 14338 61192
rect 15933 61183 15991 61189
rect 15933 61180 15945 61183
rect 14332 61152 15945 61180
rect 14332 61140 14338 61152
rect 15933 61149 15945 61152
rect 15979 61149 15991 61183
rect 15933 61143 15991 61149
rect 16206 61121 16212 61124
rect 15657 61115 15715 61121
rect 15657 61081 15669 61115
rect 15703 61112 15715 61115
rect 16200 61112 16212 61121
rect 15703 61084 16212 61112
rect 15703 61081 15715 61084
rect 15657 61075 15715 61081
rect 16200 61075 16212 61084
rect 16264 61112 16270 61124
rect 17589 61115 17647 61121
rect 17589 61112 17601 61115
rect 16264 61084 17601 61112
rect 16206 61072 16212 61075
rect 16264 61072 16270 61084
rect 17589 61081 17601 61084
rect 17635 61081 17647 61115
rect 17589 61075 17647 61081
rect 17313 61047 17371 61053
rect 17313 61013 17325 61047
rect 17359 61044 17371 61047
rect 17954 61044 17960 61056
rect 17359 61016 17960 61044
rect 17359 61013 17371 61016
rect 17313 61007 17371 61013
rect 17954 61004 17960 61016
rect 18012 61004 18018 61056
rect 1104 60954 18860 60976
rect 1104 60902 2610 60954
rect 2662 60902 2674 60954
rect 2726 60902 2738 60954
rect 2790 60902 2802 60954
rect 2854 60902 2866 60954
rect 2918 60902 7610 60954
rect 7662 60902 7674 60954
rect 7726 60902 7738 60954
rect 7790 60902 7802 60954
rect 7854 60902 7866 60954
rect 7918 60902 12610 60954
rect 12662 60902 12674 60954
rect 12726 60902 12738 60954
rect 12790 60902 12802 60954
rect 12854 60902 12866 60954
rect 12918 60902 17610 60954
rect 17662 60902 17674 60954
rect 17726 60902 17738 60954
rect 17790 60902 17802 60954
rect 17854 60902 17866 60954
rect 17918 60902 18860 60954
rect 1104 60880 18860 60902
rect 8478 60732 8484 60784
rect 8536 60772 8542 60784
rect 9490 60772 9496 60784
rect 8536 60744 9496 60772
rect 8536 60732 8542 60744
rect 9490 60732 9496 60744
rect 9548 60732 9554 60784
rect 6546 60664 6552 60716
rect 6604 60664 6610 60716
rect 6805 60707 6863 60713
rect 6805 60704 6817 60707
rect 6656 60676 6817 60704
rect 5902 60596 5908 60648
rect 5960 60636 5966 60648
rect 6656 60636 6684 60676
rect 6805 60673 6817 60676
rect 6851 60704 6863 60707
rect 8297 60707 8355 60713
rect 8297 60704 8309 60707
rect 6851 60676 8309 60704
rect 6851 60673 6863 60676
rect 6805 60667 6863 60673
rect 8297 60673 8309 60676
rect 8343 60704 8355 60707
rect 8665 60707 8723 60713
rect 8665 60704 8677 60707
rect 8343 60676 8677 60704
rect 8343 60673 8355 60676
rect 8297 60667 8355 60673
rect 8665 60673 8677 60676
rect 8711 60673 8723 60707
rect 8665 60667 8723 60673
rect 5960 60608 6684 60636
rect 5960 60596 5966 60608
rect 9398 60596 9404 60648
rect 9456 60596 9462 60648
rect 9585 60639 9643 60645
rect 9585 60605 9597 60639
rect 9631 60605 9643 60639
rect 9585 60599 9643 60605
rect 9600 60568 9628 60599
rect 10962 60568 10968 60580
rect 7852 60540 10968 60568
rect 4614 60460 4620 60512
rect 4672 60500 4678 60512
rect 7852 60500 7880 60540
rect 10962 60528 10968 60540
rect 11020 60528 11026 60580
rect 4672 60472 7880 60500
rect 4672 60460 4678 60472
rect 7926 60460 7932 60512
rect 7984 60460 7990 60512
rect 8018 60460 8024 60512
rect 8076 60500 8082 60512
rect 9033 60503 9091 60509
rect 9033 60500 9045 60503
rect 8076 60472 9045 60500
rect 8076 60460 8082 60472
rect 9033 60469 9045 60472
rect 9079 60469 9091 60503
rect 9033 60463 9091 60469
rect 1104 60410 18860 60432
rect 1104 60358 1950 60410
rect 2002 60358 2014 60410
rect 2066 60358 2078 60410
rect 2130 60358 2142 60410
rect 2194 60358 2206 60410
rect 2258 60358 6950 60410
rect 7002 60358 7014 60410
rect 7066 60358 7078 60410
rect 7130 60358 7142 60410
rect 7194 60358 7206 60410
rect 7258 60358 11950 60410
rect 12002 60358 12014 60410
rect 12066 60358 12078 60410
rect 12130 60358 12142 60410
rect 12194 60358 12206 60410
rect 12258 60358 16950 60410
rect 17002 60358 17014 60410
rect 17066 60358 17078 60410
rect 17130 60358 17142 60410
rect 17194 60358 17206 60410
rect 17258 60358 18860 60410
rect 1104 60336 18860 60358
rect 1026 60256 1032 60308
rect 1084 60296 1090 60308
rect 8018 60296 8024 60308
rect 1084 60268 8024 60296
rect 1084 60256 1090 60268
rect 8018 60256 8024 60268
rect 8076 60256 8082 60308
rect 13170 60256 13176 60308
rect 13228 60296 13234 60308
rect 16117 60299 16175 60305
rect 16117 60296 16129 60299
rect 13228 60268 16129 60296
rect 13228 60256 13234 60268
rect 16117 60265 16129 60268
rect 16163 60265 16175 60299
rect 16117 60259 16175 60265
rect 9125 60231 9183 60237
rect 9125 60197 9137 60231
rect 9171 60228 9183 60231
rect 10502 60228 10508 60240
rect 9171 60200 10508 60228
rect 9171 60197 9183 60200
rect 9125 60191 9183 60197
rect 10502 60188 10508 60200
rect 10560 60188 10566 60240
rect 15657 60231 15715 60237
rect 15657 60197 15669 60231
rect 15703 60228 15715 60231
rect 16482 60228 16488 60240
rect 15703 60200 16488 60228
rect 15703 60197 15715 60200
rect 15657 60191 15715 60197
rect 16482 60188 16488 60200
rect 16540 60188 16546 60240
rect 7190 60120 7196 60172
rect 7248 60160 7254 60172
rect 8110 60160 8116 60172
rect 7248 60132 8116 60160
rect 7248 60120 7254 60132
rect 8110 60120 8116 60132
rect 8168 60120 8174 60172
rect 8205 60163 8263 60169
rect 8205 60129 8217 60163
rect 8251 60160 8263 60163
rect 9769 60163 9827 60169
rect 9769 60160 9781 60163
rect 8251 60132 9781 60160
rect 8251 60129 8263 60132
rect 8205 60123 8263 60129
rect 9769 60129 9781 60132
rect 9815 60160 9827 60163
rect 10778 60160 10784 60172
rect 9815 60132 10784 60160
rect 9815 60129 9827 60132
rect 9769 60123 9827 60129
rect 10778 60120 10784 60132
rect 10836 60120 10842 60172
rect 15470 60120 15476 60172
rect 15528 60160 15534 60172
rect 16390 60160 16396 60172
rect 15528 60132 16396 60160
rect 15528 60120 15534 60132
rect 16390 60120 16396 60132
rect 16448 60160 16454 60172
rect 16577 60163 16635 60169
rect 16577 60160 16589 60163
rect 16448 60132 16589 60160
rect 16448 60120 16454 60132
rect 16577 60129 16589 60132
rect 16623 60129 16635 60163
rect 16577 60123 16635 60129
rect 16669 60163 16727 60169
rect 16669 60129 16681 60163
rect 16715 60129 16727 60163
rect 16669 60123 16727 60129
rect 8021 60095 8079 60101
rect 8021 60061 8033 60095
rect 8067 60092 8079 60095
rect 8067 60064 13584 60092
rect 8067 60061 8079 60064
rect 8021 60055 8079 60061
rect 6270 59984 6276 60036
rect 6328 60024 6334 60036
rect 6822 60024 6828 60036
rect 6328 59996 6828 60024
rect 6328 59984 6334 59996
rect 6822 59984 6828 59996
rect 6880 59984 6886 60036
rect 7929 60027 7987 60033
rect 7929 59993 7941 60027
rect 7975 60024 7987 60027
rect 8110 60024 8116 60036
rect 7975 59996 8116 60024
rect 7975 59993 7987 59996
rect 7929 59987 7987 59993
rect 8110 59984 8116 59996
rect 8168 59984 8174 60036
rect 9493 60027 9551 60033
rect 9493 59993 9505 60027
rect 9539 60024 9551 60027
rect 13078 60024 13084 60036
rect 9539 59996 13084 60024
rect 9539 59993 9551 59996
rect 9493 59987 9551 59993
rect 13078 59984 13084 59996
rect 13136 59984 13142 60036
rect 7282 59916 7288 59968
rect 7340 59956 7346 59968
rect 7561 59959 7619 59965
rect 7561 59956 7573 59959
rect 7340 59928 7573 59956
rect 7340 59916 7346 59928
rect 7561 59925 7573 59928
rect 7607 59925 7619 59959
rect 7561 59919 7619 59925
rect 9582 59916 9588 59968
rect 9640 59916 9646 59968
rect 13556 59956 13584 60064
rect 14274 60052 14280 60104
rect 14332 60052 14338 60104
rect 15378 60052 15384 60104
rect 15436 60092 15442 60104
rect 16684 60092 16712 60123
rect 15436 60064 16712 60092
rect 18049 60095 18107 60101
rect 15436 60052 15442 60064
rect 18049 60061 18061 60095
rect 18095 60092 18107 60095
rect 19242 60092 19248 60104
rect 18095 60064 19248 60092
rect 18095 60061 18107 60064
rect 18049 60055 18107 60061
rect 19242 60052 19248 60064
rect 19300 60052 19306 60104
rect 14550 60033 14556 60036
rect 14544 59987 14556 60033
rect 14550 59984 14556 59987
rect 14608 59984 14614 60036
rect 16114 59956 16120 59968
rect 13556 59928 16120 59956
rect 16114 59916 16120 59928
rect 16172 59956 16178 59968
rect 16485 59959 16543 59965
rect 16485 59956 16497 59959
rect 16172 59928 16497 59956
rect 16172 59916 16178 59928
rect 16485 59925 16497 59928
rect 16531 59925 16543 59959
rect 16485 59919 16543 59925
rect 18230 59916 18236 59968
rect 18288 59916 18294 59968
rect 1104 59866 18860 59888
rect 1104 59814 2610 59866
rect 2662 59814 2674 59866
rect 2726 59814 2738 59866
rect 2790 59814 2802 59866
rect 2854 59814 2866 59866
rect 2918 59814 7610 59866
rect 7662 59814 7674 59866
rect 7726 59814 7738 59866
rect 7790 59814 7802 59866
rect 7854 59814 7866 59866
rect 7918 59814 12610 59866
rect 12662 59814 12674 59866
rect 12726 59814 12738 59866
rect 12790 59814 12802 59866
rect 12854 59814 12866 59866
rect 12918 59814 17610 59866
rect 17662 59814 17674 59866
rect 17726 59814 17738 59866
rect 17790 59814 17802 59866
rect 17854 59814 17866 59866
rect 17918 59814 18860 59866
rect 1104 59792 18860 59814
rect 4617 59755 4675 59761
rect 4617 59721 4629 59755
rect 4663 59752 4675 59755
rect 4663 59724 6914 59752
rect 4663 59721 4675 59724
rect 4617 59715 4675 59721
rect 6546 59684 6552 59696
rect 3252 59656 6552 59684
rect 3252 59628 3280 59656
rect 6546 59644 6552 59656
rect 6604 59644 6610 59696
rect 6886 59684 6914 59724
rect 7190 59684 7196 59696
rect 6886 59656 7196 59684
rect 7190 59644 7196 59656
rect 7248 59684 7254 59696
rect 8202 59684 8208 59696
rect 7248 59656 8208 59684
rect 7248 59644 7254 59656
rect 8202 59644 8208 59656
rect 8260 59644 8266 59696
rect 3234 59576 3240 59628
rect 3292 59576 3298 59628
rect 3504 59619 3562 59625
rect 3504 59616 3516 59619
rect 3344 59588 3516 59616
rect 2225 59551 2283 59557
rect 2225 59517 2237 59551
rect 2271 59548 2283 59551
rect 2593 59551 2651 59557
rect 2593 59548 2605 59551
rect 2271 59520 2605 59548
rect 2271 59517 2283 59520
rect 2225 59511 2283 59517
rect 2593 59517 2605 59520
rect 2639 59548 2651 59551
rect 2961 59551 3019 59557
rect 2961 59548 2973 59551
rect 2639 59520 2973 59548
rect 2639 59517 2651 59520
rect 2593 59511 2651 59517
rect 2961 59517 2973 59520
rect 3007 59548 3019 59551
rect 3344 59548 3372 59588
rect 3504 59585 3516 59588
rect 3550 59616 3562 59619
rect 3550 59588 5028 59616
rect 3550 59585 3562 59588
rect 3504 59579 3562 59585
rect 3007 59520 3372 59548
rect 3007 59517 3019 59520
rect 2961 59511 3019 59517
rect 5000 59421 5028 59588
rect 4985 59415 5043 59421
rect 4985 59381 4997 59415
rect 5031 59412 5043 59415
rect 5166 59412 5172 59424
rect 5031 59384 5172 59412
rect 5031 59381 5043 59384
rect 4985 59375 5043 59381
rect 5166 59372 5172 59384
rect 5224 59412 5230 59424
rect 5261 59415 5319 59421
rect 5261 59412 5273 59415
rect 5224 59384 5273 59412
rect 5224 59372 5230 59384
rect 5261 59381 5273 59384
rect 5307 59381 5319 59415
rect 5261 59375 5319 59381
rect 1104 59322 18860 59344
rect 1104 59270 1950 59322
rect 2002 59270 2014 59322
rect 2066 59270 2078 59322
rect 2130 59270 2142 59322
rect 2194 59270 2206 59322
rect 2258 59270 6950 59322
rect 7002 59270 7014 59322
rect 7066 59270 7078 59322
rect 7130 59270 7142 59322
rect 7194 59270 7206 59322
rect 7258 59270 11950 59322
rect 12002 59270 12014 59322
rect 12066 59270 12078 59322
rect 12130 59270 12142 59322
rect 12194 59270 12206 59322
rect 12258 59270 16950 59322
rect 17002 59270 17014 59322
rect 17066 59270 17078 59322
rect 17130 59270 17142 59322
rect 17194 59270 17206 59322
rect 17258 59270 18860 59322
rect 1104 59248 18860 59270
rect 15194 59032 15200 59084
rect 15252 59032 15258 59084
rect 15378 59032 15384 59084
rect 15436 59032 15442 59084
rect 4062 58964 4068 59016
rect 4120 59004 4126 59016
rect 7285 59007 7343 59013
rect 7285 59004 7297 59007
rect 4120 58976 7297 59004
rect 4120 58964 4126 58976
rect 7285 58973 7297 58976
rect 7331 58973 7343 59007
rect 7285 58967 7343 58973
rect 7561 59007 7619 59013
rect 7561 58973 7573 59007
rect 7607 59004 7619 59007
rect 18874 59004 18880 59016
rect 7607 58976 18880 59004
rect 7607 58973 7619 58976
rect 7561 58967 7619 58973
rect 18874 58964 18880 58976
rect 18932 58964 18938 59016
rect 15286 58896 15292 58948
rect 15344 58936 15350 58948
rect 15470 58936 15476 58948
rect 15344 58908 15476 58936
rect 15344 58896 15350 58908
rect 15470 58896 15476 58908
rect 15528 58896 15534 58948
rect 13722 58828 13728 58880
rect 13780 58868 13786 58880
rect 14369 58871 14427 58877
rect 14369 58868 14381 58871
rect 13780 58840 14381 58868
rect 13780 58828 13786 58840
rect 14369 58837 14381 58840
rect 14415 58868 14427 58871
rect 14811 58871 14869 58877
rect 14811 58868 14823 58871
rect 14415 58840 14823 58868
rect 14415 58837 14427 58840
rect 14369 58831 14427 58837
rect 14811 58837 14823 58840
rect 14857 58868 14869 58871
rect 15749 58871 15807 58877
rect 15749 58868 15761 58871
rect 14857 58840 15761 58868
rect 14857 58837 14869 58840
rect 14811 58831 14869 58837
rect 15749 58837 15761 58840
rect 15795 58837 15807 58871
rect 15749 58831 15807 58837
rect 1104 58778 18860 58800
rect 1104 58726 2610 58778
rect 2662 58726 2674 58778
rect 2726 58726 2738 58778
rect 2790 58726 2802 58778
rect 2854 58726 2866 58778
rect 2918 58726 7610 58778
rect 7662 58726 7674 58778
rect 7726 58726 7738 58778
rect 7790 58726 7802 58778
rect 7854 58726 7866 58778
rect 7918 58726 12610 58778
rect 12662 58726 12674 58778
rect 12726 58726 12738 58778
rect 12790 58726 12802 58778
rect 12854 58726 12866 58778
rect 12918 58726 17610 58778
rect 17662 58726 17674 58778
rect 17726 58726 17738 58778
rect 17790 58726 17802 58778
rect 17854 58726 17866 58778
rect 17918 58726 18860 58778
rect 1104 58704 18860 58726
rect 16666 58488 16672 58540
rect 16724 58528 16730 58540
rect 18049 58531 18107 58537
rect 18049 58528 18061 58531
rect 16724 58500 18061 58528
rect 16724 58488 16730 58500
rect 18049 58497 18061 58500
rect 18095 58497 18107 58531
rect 18049 58491 18107 58497
rect 18230 58284 18236 58336
rect 18288 58284 18294 58336
rect 1104 58234 18860 58256
rect 1104 58182 1950 58234
rect 2002 58182 2014 58234
rect 2066 58182 2078 58234
rect 2130 58182 2142 58234
rect 2194 58182 2206 58234
rect 2258 58182 6950 58234
rect 7002 58182 7014 58234
rect 7066 58182 7078 58234
rect 7130 58182 7142 58234
rect 7194 58182 7206 58234
rect 7258 58182 11950 58234
rect 12002 58182 12014 58234
rect 12066 58182 12078 58234
rect 12130 58182 12142 58234
rect 12194 58182 12206 58234
rect 12258 58182 16950 58234
rect 17002 58182 17014 58234
rect 17066 58182 17078 58234
rect 17130 58182 17142 58234
rect 17194 58182 17206 58234
rect 17258 58182 18860 58234
rect 1104 58160 18860 58182
rect 2314 57740 2320 57792
rect 2372 57780 2378 57792
rect 8110 57780 8116 57792
rect 2372 57752 8116 57780
rect 2372 57740 2378 57752
rect 8110 57740 8116 57752
rect 8168 57780 8174 57792
rect 10042 57780 10048 57792
rect 8168 57752 10048 57780
rect 8168 57740 8174 57752
rect 10042 57740 10048 57752
rect 10100 57740 10106 57792
rect 1104 57690 18860 57712
rect 1104 57638 2610 57690
rect 2662 57638 2674 57690
rect 2726 57638 2738 57690
rect 2790 57638 2802 57690
rect 2854 57638 2866 57690
rect 2918 57638 7610 57690
rect 7662 57638 7674 57690
rect 7726 57638 7738 57690
rect 7790 57638 7802 57690
rect 7854 57638 7866 57690
rect 7918 57638 12610 57690
rect 12662 57638 12674 57690
rect 12726 57638 12738 57690
rect 12790 57638 12802 57690
rect 12854 57638 12866 57690
rect 12918 57638 17610 57690
rect 17662 57638 17674 57690
rect 17726 57638 17738 57690
rect 17790 57638 17802 57690
rect 17854 57638 17866 57690
rect 17918 57638 18860 57690
rect 1104 57616 18860 57638
rect 8110 57536 8116 57588
rect 8168 57576 8174 57588
rect 8386 57576 8392 57588
rect 8168 57548 8392 57576
rect 8168 57536 8174 57548
rect 8386 57536 8392 57548
rect 8444 57536 8450 57588
rect 15562 57536 15568 57588
rect 15620 57576 15626 57588
rect 17313 57579 17371 57585
rect 17313 57576 17325 57579
rect 15620 57548 17325 57576
rect 15620 57536 15626 57548
rect 17313 57545 17325 57548
rect 17359 57545 17371 57579
rect 17313 57539 17371 57545
rect 3234 57508 3240 57520
rect 2792 57480 3240 57508
rect 2792 57449 2820 57480
rect 3234 57468 3240 57480
rect 3292 57468 3298 57520
rect 4982 57468 4988 57520
rect 5040 57508 5046 57520
rect 16574 57508 16580 57520
rect 5040 57480 16580 57508
rect 5040 57468 5046 57480
rect 16574 57468 16580 57480
rect 16632 57508 16638 57520
rect 16945 57511 17003 57517
rect 16945 57508 16957 57511
rect 16632 57480 16957 57508
rect 16632 57468 16638 57480
rect 16945 57477 16957 57480
rect 16991 57508 17003 57511
rect 17681 57511 17739 57517
rect 17681 57508 17693 57511
rect 16991 57480 17693 57508
rect 16991 57477 17003 57480
rect 16945 57471 17003 57477
rect 17681 57477 17693 57480
rect 17727 57477 17739 57511
rect 17681 57471 17739 57477
rect 3050 57449 3056 57452
rect 2777 57443 2835 57449
rect 2777 57409 2789 57443
rect 2823 57409 2835 57443
rect 3044 57440 3056 57449
rect 2777 57403 2835 57409
rect 2884 57412 3056 57440
rect 2501 57375 2559 57381
rect 2501 57341 2513 57375
rect 2547 57372 2559 57375
rect 2884 57372 2912 57412
rect 3044 57403 3056 57412
rect 3050 57400 3056 57403
rect 3108 57400 3114 57452
rect 15197 57443 15255 57449
rect 15197 57409 15209 57443
rect 15243 57440 15255 57443
rect 16850 57440 16856 57452
rect 15243 57412 16856 57440
rect 15243 57409 15255 57412
rect 15197 57403 15255 57409
rect 16850 57400 16856 57412
rect 16908 57400 16914 57452
rect 2547 57344 2912 57372
rect 2547 57341 2559 57344
rect 2501 57335 2559 57341
rect 15286 57332 15292 57384
rect 15344 57372 15350 57384
rect 17773 57375 17831 57381
rect 17773 57372 17785 57375
rect 15344 57344 17785 57372
rect 15344 57332 15350 57344
rect 17773 57341 17785 57344
rect 17819 57341 17831 57375
rect 17773 57335 17831 57341
rect 17865 57375 17923 57381
rect 17865 57341 17877 57375
rect 17911 57341 17923 57375
rect 17865 57335 17923 57341
rect 17402 57264 17408 57316
rect 17460 57304 17466 57316
rect 17880 57304 17908 57335
rect 17460 57276 17908 57304
rect 17460 57264 17466 57276
rect 4154 57196 4160 57248
rect 4212 57196 4218 57248
rect 8294 57196 8300 57248
rect 8352 57236 8358 57248
rect 15013 57239 15071 57245
rect 15013 57236 15025 57239
rect 8352 57208 15025 57236
rect 8352 57196 8358 57208
rect 15013 57205 15025 57208
rect 15059 57205 15071 57239
rect 15013 57199 15071 57205
rect 1104 57146 18860 57168
rect 1104 57094 1950 57146
rect 2002 57094 2014 57146
rect 2066 57094 2078 57146
rect 2130 57094 2142 57146
rect 2194 57094 2206 57146
rect 2258 57094 6950 57146
rect 7002 57094 7014 57146
rect 7066 57094 7078 57146
rect 7130 57094 7142 57146
rect 7194 57094 7206 57146
rect 7258 57094 11950 57146
rect 12002 57094 12014 57146
rect 12066 57094 12078 57146
rect 12130 57094 12142 57146
rect 12194 57094 12206 57146
rect 12258 57094 16950 57146
rect 17002 57094 17014 57146
rect 17066 57094 17078 57146
rect 17130 57094 17142 57146
rect 17194 57094 17206 57146
rect 17258 57094 18860 57146
rect 1104 57072 18860 57094
rect 4154 56992 4160 57044
rect 4212 57032 4218 57044
rect 13170 57032 13176 57044
rect 4212 57004 13176 57032
rect 4212 56992 4218 57004
rect 13170 56992 13176 57004
rect 13228 56992 13234 57044
rect 1673 56967 1731 56973
rect 1673 56933 1685 56967
rect 1719 56964 1731 56967
rect 3510 56964 3516 56976
rect 1719 56936 3516 56964
rect 1719 56933 1731 56936
rect 1673 56927 1731 56933
rect 3510 56924 3516 56936
rect 3568 56924 3574 56976
rect 1486 56856 1492 56908
rect 1544 56896 1550 56908
rect 2225 56899 2283 56905
rect 2225 56896 2237 56899
rect 1544 56868 2237 56896
rect 1544 56856 1550 56868
rect 2225 56865 2237 56868
rect 2271 56896 2283 56899
rect 2314 56896 2320 56908
rect 2271 56868 2320 56896
rect 2271 56865 2283 56868
rect 2225 56859 2283 56865
rect 2314 56856 2320 56868
rect 2372 56856 2378 56908
rect 1949 56831 2007 56837
rect 1949 56797 1961 56831
rect 1995 56828 2007 56831
rect 1995 56800 2728 56828
rect 1995 56797 2007 56800
rect 1949 56791 2007 56797
rect 2133 56695 2191 56701
rect 2133 56661 2145 56695
rect 2179 56692 2191 56695
rect 2406 56692 2412 56704
rect 2179 56664 2412 56692
rect 2179 56661 2191 56664
rect 2133 56655 2191 56661
rect 2406 56652 2412 56664
rect 2464 56652 2470 56704
rect 2700 56701 2728 56800
rect 2685 56695 2743 56701
rect 2685 56661 2697 56695
rect 2731 56692 2743 56695
rect 17954 56692 17960 56704
rect 2731 56664 17960 56692
rect 2731 56661 2743 56664
rect 2685 56655 2743 56661
rect 17954 56652 17960 56664
rect 18012 56652 18018 56704
rect 1104 56602 18860 56624
rect 1104 56550 2610 56602
rect 2662 56550 2674 56602
rect 2726 56550 2738 56602
rect 2790 56550 2802 56602
rect 2854 56550 2866 56602
rect 2918 56550 7610 56602
rect 7662 56550 7674 56602
rect 7726 56550 7738 56602
rect 7790 56550 7802 56602
rect 7854 56550 7866 56602
rect 7918 56550 12610 56602
rect 12662 56550 12674 56602
rect 12726 56550 12738 56602
rect 12790 56550 12802 56602
rect 12854 56550 12866 56602
rect 12918 56550 17610 56602
rect 17662 56550 17674 56602
rect 17726 56550 17738 56602
rect 17790 56550 17802 56602
rect 17854 56550 17866 56602
rect 17918 56550 18860 56602
rect 1104 56528 18860 56550
rect 3390 56423 3448 56429
rect 3390 56420 3402 56423
rect 2792 56392 3402 56420
rect 1670 56312 1676 56364
rect 1728 56352 1734 56364
rect 2501 56355 2559 56361
rect 2501 56352 2513 56355
rect 1728 56324 2513 56352
rect 1728 56312 1734 56324
rect 2501 56321 2513 56324
rect 2547 56321 2559 56355
rect 2501 56315 2559 56321
rect 934 56176 940 56228
rect 992 56216 998 56228
rect 2792 56225 2820 56392
rect 3390 56389 3402 56392
rect 3436 56389 3448 56423
rect 3390 56383 3448 56389
rect 2958 56312 2964 56364
rect 3016 56352 3022 56364
rect 3145 56355 3203 56361
rect 3145 56352 3157 56355
rect 3016 56324 3157 56352
rect 3016 56312 3022 56324
rect 3145 56321 3157 56324
rect 3191 56352 3203 56355
rect 3234 56352 3240 56364
rect 3191 56324 3240 56352
rect 3191 56321 3203 56324
rect 3145 56315 3203 56321
rect 3234 56312 3240 56324
rect 3292 56312 3298 56364
rect 8110 56312 8116 56364
rect 8168 56352 8174 56364
rect 18049 56355 18107 56361
rect 18049 56352 18061 56355
rect 8168 56324 18061 56352
rect 8168 56312 8174 56324
rect 18049 56321 18061 56324
rect 18095 56321 18107 56355
rect 18049 56315 18107 56321
rect 12434 56244 12440 56296
rect 12492 56244 12498 56296
rect 12713 56287 12771 56293
rect 12713 56253 12725 56287
rect 12759 56284 12771 56287
rect 12986 56284 12992 56296
rect 12759 56256 12992 56284
rect 12759 56253 12771 56256
rect 12713 56247 12771 56253
rect 12986 56244 12992 56256
rect 13044 56244 13050 56296
rect 2777 56219 2835 56225
rect 2777 56216 2789 56219
rect 992 56188 2789 56216
rect 992 56176 998 56188
rect 2777 56185 2789 56188
rect 2823 56185 2835 56219
rect 2777 56179 2835 56185
rect 2314 56108 2320 56160
rect 2372 56108 2378 56160
rect 4522 56108 4528 56160
rect 4580 56108 4586 56160
rect 18230 56108 18236 56160
rect 18288 56108 18294 56160
rect 1104 56058 18860 56080
rect 1104 56006 1950 56058
rect 2002 56006 2014 56058
rect 2066 56006 2078 56058
rect 2130 56006 2142 56058
rect 2194 56006 2206 56058
rect 2258 56006 6950 56058
rect 7002 56006 7014 56058
rect 7066 56006 7078 56058
rect 7130 56006 7142 56058
rect 7194 56006 7206 56058
rect 7258 56006 11950 56058
rect 12002 56006 12014 56058
rect 12066 56006 12078 56058
rect 12130 56006 12142 56058
rect 12194 56006 12206 56058
rect 12258 56006 16950 56058
rect 17002 56006 17014 56058
rect 17066 56006 17078 56058
rect 17130 56006 17142 56058
rect 17194 56006 17206 56058
rect 17258 56006 18860 56058
rect 1104 55984 18860 56006
rect 4890 55836 4896 55888
rect 4948 55876 4954 55888
rect 11698 55876 11704 55888
rect 4948 55848 11704 55876
rect 4948 55836 4954 55848
rect 11698 55836 11704 55848
rect 11756 55836 11762 55888
rect 10962 55768 10968 55820
rect 11020 55808 11026 55820
rect 11793 55811 11851 55817
rect 11793 55808 11805 55811
rect 11020 55780 11805 55808
rect 11020 55768 11026 55780
rect 11793 55777 11805 55780
rect 11839 55808 11851 55811
rect 11839 55780 16574 55808
rect 11839 55777 11851 55780
rect 11793 55771 11851 55777
rect 1673 55743 1731 55749
rect 1673 55709 1685 55743
rect 1719 55740 1731 55743
rect 2958 55740 2964 55752
rect 1719 55712 2964 55740
rect 1719 55709 1731 55712
rect 1673 55703 1731 55709
rect 2958 55700 2964 55712
rect 3016 55700 3022 55752
rect 11517 55743 11575 55749
rect 11517 55709 11529 55743
rect 11563 55740 11575 55743
rect 11698 55740 11704 55752
rect 11563 55712 11704 55740
rect 11563 55709 11575 55712
rect 11517 55703 11575 55709
rect 11698 55700 11704 55712
rect 11756 55700 11762 55752
rect 842 55632 848 55684
rect 900 55672 906 55684
rect 1918 55675 1976 55681
rect 1918 55672 1930 55675
rect 900 55644 1930 55672
rect 900 55632 906 55644
rect 1918 55641 1930 55644
rect 1964 55641 1976 55675
rect 16546 55672 16574 55780
rect 17126 55672 17132 55684
rect 16546 55644 17132 55672
rect 1918 55635 1976 55641
rect 17126 55632 17132 55644
rect 17184 55632 17190 55684
rect 3053 55607 3111 55613
rect 3053 55573 3065 55607
rect 3099 55604 3111 55607
rect 10226 55604 10232 55616
rect 3099 55576 10232 55604
rect 3099 55573 3111 55576
rect 3053 55567 3111 55573
rect 10226 55564 10232 55576
rect 10284 55564 10290 55616
rect 1104 55514 18860 55536
rect 1104 55462 2610 55514
rect 2662 55462 2674 55514
rect 2726 55462 2738 55514
rect 2790 55462 2802 55514
rect 2854 55462 2866 55514
rect 2918 55462 7610 55514
rect 7662 55462 7674 55514
rect 7726 55462 7738 55514
rect 7790 55462 7802 55514
rect 7854 55462 7866 55514
rect 7918 55462 12610 55514
rect 12662 55462 12674 55514
rect 12726 55462 12738 55514
rect 12790 55462 12802 55514
rect 12854 55462 12866 55514
rect 12918 55462 17610 55514
rect 17662 55462 17674 55514
rect 17726 55462 17738 55514
rect 17790 55462 17802 55514
rect 17854 55462 17866 55514
rect 17918 55462 18860 55514
rect 1104 55440 18860 55462
rect 3602 55360 3608 55412
rect 3660 55360 3666 55412
rect 4065 55403 4123 55409
rect 4065 55369 4077 55403
rect 4111 55400 4123 55403
rect 4433 55403 4491 55409
rect 4433 55400 4445 55403
rect 4111 55372 4445 55400
rect 4111 55369 4123 55372
rect 4065 55363 4123 55369
rect 4433 55369 4445 55372
rect 4479 55400 4491 55403
rect 4801 55403 4859 55409
rect 4801 55400 4813 55403
rect 4479 55372 4813 55400
rect 4479 55369 4491 55372
rect 4433 55363 4491 55369
rect 4801 55369 4813 55372
rect 4847 55400 4859 55403
rect 5169 55403 5227 55409
rect 5169 55400 5181 55403
rect 4847 55372 5181 55400
rect 4847 55369 4859 55372
rect 4801 55363 4859 55369
rect 5169 55369 5181 55372
rect 5215 55400 5227 55403
rect 5718 55400 5724 55412
rect 5215 55372 5724 55400
rect 5215 55369 5227 55372
rect 5169 55363 5227 55369
rect 5718 55360 5724 55372
rect 5776 55360 5782 55412
rect 16850 55360 16856 55412
rect 16908 55360 16914 55412
rect 2958 55332 2964 55344
rect 2240 55304 2964 55332
rect 2240 55273 2268 55304
rect 2958 55292 2964 55304
rect 3016 55292 3022 55344
rect 10410 55332 10416 55344
rect 3896 55304 10416 55332
rect 2225 55267 2283 55273
rect 2225 55233 2237 55267
rect 2271 55233 2283 55267
rect 2225 55227 2283 55233
rect 2492 55267 2550 55273
rect 2492 55233 2504 55267
rect 2538 55264 2550 55267
rect 3896 55264 3924 55304
rect 10410 55292 10416 55304
rect 10468 55292 10474 55344
rect 16574 55292 16580 55344
rect 16632 55332 16638 55344
rect 17313 55335 17371 55341
rect 17313 55332 17325 55335
rect 16632 55304 17325 55332
rect 16632 55292 16638 55304
rect 17313 55301 17325 55304
rect 17359 55301 17371 55335
rect 17313 55295 17371 55301
rect 2538 55236 3924 55264
rect 2538 55233 2550 55236
rect 2492 55227 2550 55233
rect 5534 55224 5540 55276
rect 5592 55224 5598 55276
rect 5718 55224 5724 55276
rect 5776 55264 5782 55276
rect 6546 55264 6552 55276
rect 5776 55236 6552 55264
rect 5776 55224 5782 55236
rect 6546 55224 6552 55236
rect 6604 55224 6610 55276
rect 16850 55224 16856 55276
rect 16908 55264 16914 55276
rect 17221 55267 17279 55273
rect 17221 55264 17233 55267
rect 16908 55236 17233 55264
rect 16908 55224 16914 55236
rect 17221 55233 17233 55236
rect 17267 55233 17279 55267
rect 17221 55227 17279 55233
rect 17126 55156 17132 55208
rect 17184 55196 17190 55208
rect 17405 55199 17463 55205
rect 17405 55196 17417 55199
rect 17184 55168 17417 55196
rect 17184 55156 17190 55168
rect 17405 55165 17417 55168
rect 17451 55165 17463 55199
rect 17405 55159 17463 55165
rect 1104 54970 18860 54992
rect 1104 54918 1950 54970
rect 2002 54918 2014 54970
rect 2066 54918 2078 54970
rect 2130 54918 2142 54970
rect 2194 54918 2206 54970
rect 2258 54918 6950 54970
rect 7002 54918 7014 54970
rect 7066 54918 7078 54970
rect 7130 54918 7142 54970
rect 7194 54918 7206 54970
rect 7258 54918 11950 54970
rect 12002 54918 12014 54970
rect 12066 54918 12078 54970
rect 12130 54918 12142 54970
rect 12194 54918 12206 54970
rect 12258 54918 16950 54970
rect 17002 54918 17014 54970
rect 17066 54918 17078 54970
rect 17130 54918 17142 54970
rect 17194 54918 17206 54970
rect 17258 54918 18860 54970
rect 1104 54896 18860 54918
rect 18049 54655 18107 54661
rect 18049 54621 18061 54655
rect 18095 54652 18107 54655
rect 18138 54652 18144 54664
rect 18095 54624 18144 54652
rect 18095 54621 18107 54624
rect 18049 54615 18107 54621
rect 18138 54612 18144 54624
rect 18196 54612 18202 54664
rect 18230 54476 18236 54528
rect 18288 54476 18294 54528
rect 1104 54426 18860 54448
rect 1104 54374 2610 54426
rect 2662 54374 2674 54426
rect 2726 54374 2738 54426
rect 2790 54374 2802 54426
rect 2854 54374 2866 54426
rect 2918 54374 7610 54426
rect 7662 54374 7674 54426
rect 7726 54374 7738 54426
rect 7790 54374 7802 54426
rect 7854 54374 7866 54426
rect 7918 54374 12610 54426
rect 12662 54374 12674 54426
rect 12726 54374 12738 54426
rect 12790 54374 12802 54426
rect 12854 54374 12866 54426
rect 12918 54374 17610 54426
rect 17662 54374 17674 54426
rect 17726 54374 17738 54426
rect 17790 54374 17802 54426
rect 17854 54374 17866 54426
rect 17918 54374 18860 54426
rect 1104 54352 18860 54374
rect 8110 54272 8116 54324
rect 8168 54312 8174 54324
rect 8386 54312 8392 54324
rect 8168 54284 8392 54312
rect 8168 54272 8174 54284
rect 8386 54272 8392 54284
rect 8444 54272 8450 54324
rect 11054 54272 11060 54324
rect 11112 54312 11118 54324
rect 11422 54312 11428 54324
rect 11112 54284 11428 54312
rect 11112 54272 11118 54284
rect 11422 54272 11428 54284
rect 11480 54272 11486 54324
rect 7374 54136 7380 54188
rect 7432 54176 7438 54188
rect 8110 54176 8116 54188
rect 7432 54148 8116 54176
rect 7432 54136 7438 54148
rect 8110 54136 8116 54148
rect 8168 54136 8174 54188
rect 9953 54179 10011 54185
rect 9953 54145 9965 54179
rect 9999 54176 10011 54179
rect 10594 54176 10600 54188
rect 9999 54148 10600 54176
rect 9999 54145 10011 54148
rect 9953 54139 10011 54145
rect 10594 54136 10600 54148
rect 10652 54136 10658 54188
rect 10689 54179 10747 54185
rect 10689 54145 10701 54179
rect 10735 54176 10747 54179
rect 11054 54176 11060 54188
rect 10735 54148 11060 54176
rect 10735 54145 10747 54148
rect 10689 54139 10747 54145
rect 11054 54136 11060 54148
rect 11112 54176 11118 54188
rect 11238 54176 11244 54188
rect 11112 54148 11244 54176
rect 11112 54136 11118 54148
rect 11238 54136 11244 54148
rect 11296 54136 11302 54188
rect 12434 54136 12440 54188
rect 12492 54176 12498 54188
rect 12989 54179 13047 54185
rect 12989 54176 13001 54179
rect 12492 54148 13001 54176
rect 12492 54136 12498 54148
rect 12989 54145 13001 54148
rect 13035 54145 13047 54179
rect 12989 54139 13047 54145
rect 10778 54068 10784 54120
rect 10836 54108 10842 54120
rect 10873 54111 10931 54117
rect 10873 54108 10885 54111
rect 10836 54080 10885 54108
rect 10836 54068 10842 54080
rect 10873 54077 10885 54080
rect 10919 54108 10931 54111
rect 10962 54108 10968 54120
rect 10919 54080 10968 54108
rect 10919 54077 10931 54080
rect 10873 54071 10931 54077
rect 10962 54068 10968 54080
rect 11020 54068 11026 54120
rect 7374 54000 7380 54052
rect 7432 54040 7438 54052
rect 10229 54043 10287 54049
rect 10229 54040 10241 54043
rect 7432 54012 10241 54040
rect 7432 54000 7438 54012
rect 10229 54009 10241 54012
rect 10275 54009 10287 54043
rect 10229 54003 10287 54009
rect 12526 53932 12532 53984
rect 12584 53972 12590 53984
rect 12805 53975 12863 53981
rect 12805 53972 12817 53975
rect 12584 53944 12817 53972
rect 12584 53932 12590 53944
rect 12805 53941 12817 53944
rect 12851 53941 12863 53975
rect 12805 53935 12863 53941
rect 1104 53882 18860 53904
rect 1104 53830 1950 53882
rect 2002 53830 2014 53882
rect 2066 53830 2078 53882
rect 2130 53830 2142 53882
rect 2194 53830 2206 53882
rect 2258 53830 6950 53882
rect 7002 53830 7014 53882
rect 7066 53830 7078 53882
rect 7130 53830 7142 53882
rect 7194 53830 7206 53882
rect 7258 53830 11950 53882
rect 12002 53830 12014 53882
rect 12066 53830 12078 53882
rect 12130 53830 12142 53882
rect 12194 53830 12206 53882
rect 12258 53830 16950 53882
rect 17002 53830 17014 53882
rect 17066 53830 17078 53882
rect 17130 53830 17142 53882
rect 17194 53830 17206 53882
rect 17258 53830 18860 53882
rect 1104 53808 18860 53830
rect 1946 53388 1952 53440
rect 2004 53428 2010 53440
rect 15930 53428 15936 53440
rect 2004 53400 15936 53428
rect 2004 53388 2010 53400
rect 15930 53388 15936 53400
rect 15988 53388 15994 53440
rect 1104 53338 18860 53360
rect 1104 53286 2610 53338
rect 2662 53286 2674 53338
rect 2726 53286 2738 53338
rect 2790 53286 2802 53338
rect 2854 53286 2866 53338
rect 2918 53286 7610 53338
rect 7662 53286 7674 53338
rect 7726 53286 7738 53338
rect 7790 53286 7802 53338
rect 7854 53286 7866 53338
rect 7918 53286 12610 53338
rect 12662 53286 12674 53338
rect 12726 53286 12738 53338
rect 12790 53286 12802 53338
rect 12854 53286 12866 53338
rect 12918 53286 17610 53338
rect 17662 53286 17674 53338
rect 17726 53286 17738 53338
rect 17790 53286 17802 53338
rect 17854 53286 17866 53338
rect 17918 53286 18860 53338
rect 1104 53264 18860 53286
rect 7834 53184 7840 53236
rect 7892 53224 7898 53236
rect 13725 53227 13783 53233
rect 13725 53224 13737 53227
rect 7892 53196 13737 53224
rect 7892 53184 7898 53196
rect 13725 53193 13737 53196
rect 13771 53224 13783 53227
rect 15286 53224 15292 53236
rect 13771 53196 15292 53224
rect 13771 53193 13783 53196
rect 13725 53187 13783 53193
rect 15286 53184 15292 53196
rect 15344 53184 15350 53236
rect 1946 53116 1952 53168
rect 2004 53116 2010 53168
rect 2133 53159 2191 53165
rect 2133 53125 2145 53159
rect 2179 53156 2191 53159
rect 9953 53159 10011 53165
rect 2179 53128 9904 53156
rect 2179 53125 2191 53128
rect 2133 53119 2191 53125
rect 8573 53091 8631 53097
rect 8573 53057 8585 53091
rect 8619 53088 8631 53091
rect 9122 53088 9128 53100
rect 8619 53060 9128 53088
rect 8619 53057 8631 53060
rect 8573 53051 8631 53057
rect 9122 53048 9128 53060
rect 9180 53048 9186 53100
rect 9876 53088 9904 53128
rect 9953 53125 9965 53159
rect 9999 53156 10011 53159
rect 10134 53156 10140 53168
rect 9999 53128 10140 53156
rect 9999 53125 10011 53128
rect 9953 53119 10011 53125
rect 10134 53116 10140 53128
rect 10192 53116 10198 53168
rect 14274 53156 14280 53168
rect 12360 53128 14280 53156
rect 11422 53088 11428 53100
rect 9876 53060 11428 53088
rect 11422 53048 11428 53060
rect 11480 53048 11486 53100
rect 2225 53023 2283 53029
rect 2225 52989 2237 53023
rect 2271 53020 2283 53023
rect 3326 53020 3332 53032
rect 2271 52992 3332 53020
rect 2271 52989 2283 52992
rect 2225 52983 2283 52989
rect 3326 52980 3332 52992
rect 3384 52980 3390 53032
rect 9858 52980 9864 53032
rect 9916 52980 9922 53032
rect 10045 53023 10103 53029
rect 10045 52989 10057 53023
rect 10091 52989 10103 53023
rect 10045 52983 10103 52989
rect 750 52912 756 52964
rect 808 52952 814 52964
rect 8757 52955 8815 52961
rect 8757 52952 8769 52955
rect 808 52924 8769 52952
rect 808 52912 814 52924
rect 8757 52921 8769 52924
rect 8803 52921 8815 52955
rect 8757 52915 8815 52921
rect 1673 52887 1731 52893
rect 1673 52853 1685 52887
rect 1719 52884 1731 52887
rect 1762 52884 1768 52896
rect 1719 52856 1768 52884
rect 1719 52853 1731 52856
rect 1673 52847 1731 52853
rect 1762 52844 1768 52856
rect 1820 52844 1826 52896
rect 8018 52844 8024 52896
rect 8076 52884 8082 52896
rect 8570 52884 8576 52896
rect 8076 52856 8576 52884
rect 8076 52844 8082 52856
rect 8570 52844 8576 52856
rect 8628 52844 8634 52896
rect 9490 52844 9496 52896
rect 9548 52844 9554 52896
rect 10060 52884 10088 52983
rect 10410 52980 10416 53032
rect 10468 53020 10474 53032
rect 12360 53029 12388 53128
rect 14274 53116 14280 53128
rect 14332 53116 14338 53168
rect 12612 53091 12670 53097
rect 12612 53057 12624 53091
rect 12658 53088 12670 53091
rect 15838 53088 15844 53100
rect 12658 53060 15844 53088
rect 12658 53057 12670 53060
rect 12612 53051 12670 53057
rect 15838 53048 15844 53060
rect 15896 53048 15902 53100
rect 12345 53023 12403 53029
rect 12345 53020 12357 53023
rect 10468 52992 12357 53020
rect 10468 52980 10474 52992
rect 12345 52989 12357 52992
rect 12391 52989 12403 53023
rect 12345 52983 12403 52989
rect 10870 52884 10876 52896
rect 10060 52856 10876 52884
rect 10870 52844 10876 52856
rect 10928 52884 10934 52896
rect 13262 52884 13268 52896
rect 10928 52856 13268 52884
rect 10928 52844 10934 52856
rect 13262 52844 13268 52856
rect 13320 52844 13326 52896
rect 1104 52794 18860 52816
rect 1104 52742 1950 52794
rect 2002 52742 2014 52794
rect 2066 52742 2078 52794
rect 2130 52742 2142 52794
rect 2194 52742 2206 52794
rect 2258 52742 6950 52794
rect 7002 52742 7014 52794
rect 7066 52742 7078 52794
rect 7130 52742 7142 52794
rect 7194 52742 7206 52794
rect 7258 52742 11950 52794
rect 12002 52742 12014 52794
rect 12066 52742 12078 52794
rect 12130 52742 12142 52794
rect 12194 52742 12206 52794
rect 12258 52742 16950 52794
rect 17002 52742 17014 52794
rect 17066 52742 17078 52794
rect 17130 52742 17142 52794
rect 17194 52742 17206 52794
rect 17258 52742 18860 52794
rect 1104 52720 18860 52742
rect 6914 52640 6920 52692
rect 6972 52680 6978 52692
rect 7834 52680 7840 52692
rect 6972 52652 7840 52680
rect 6972 52640 6978 52652
rect 7834 52640 7840 52652
rect 7892 52640 7898 52692
rect 18230 52572 18236 52624
rect 18288 52572 18294 52624
rect 14274 52504 14280 52556
rect 14332 52504 14338 52556
rect 8754 52436 8760 52488
rect 8812 52476 8818 52488
rect 9306 52476 9312 52488
rect 8812 52448 9312 52476
rect 8812 52436 8818 52448
rect 9306 52436 9312 52448
rect 9364 52436 9370 52488
rect 14544 52479 14602 52485
rect 14544 52445 14556 52479
rect 14590 52476 14602 52479
rect 15562 52476 15568 52488
rect 14590 52448 15568 52476
rect 14590 52445 14602 52448
rect 14544 52439 14602 52445
rect 15562 52436 15568 52448
rect 15620 52436 15626 52488
rect 17954 52436 17960 52488
rect 18012 52476 18018 52488
rect 18049 52479 18107 52485
rect 18049 52476 18061 52479
rect 18012 52448 18061 52476
rect 18012 52436 18018 52448
rect 18049 52445 18061 52448
rect 18095 52445 18107 52479
rect 18049 52439 18107 52445
rect 15654 52300 15660 52352
rect 15712 52300 15718 52352
rect 1104 52250 18860 52272
rect 1104 52198 2610 52250
rect 2662 52198 2674 52250
rect 2726 52198 2738 52250
rect 2790 52198 2802 52250
rect 2854 52198 2866 52250
rect 2918 52198 7610 52250
rect 7662 52198 7674 52250
rect 7726 52198 7738 52250
rect 7790 52198 7802 52250
rect 7854 52198 7866 52250
rect 7918 52198 12610 52250
rect 12662 52198 12674 52250
rect 12726 52198 12738 52250
rect 12790 52198 12802 52250
rect 12854 52198 12866 52250
rect 12918 52198 17610 52250
rect 17662 52198 17674 52250
rect 17726 52198 17738 52250
rect 17790 52198 17802 52250
rect 17854 52198 17866 52250
rect 17918 52198 18860 52250
rect 1104 52176 18860 52198
rect 14550 52096 14556 52148
rect 14608 52136 14614 52148
rect 18049 52139 18107 52145
rect 18049 52136 18061 52139
rect 14608 52108 18061 52136
rect 14608 52096 14614 52108
rect 18049 52105 18061 52108
rect 18095 52105 18107 52139
rect 18049 52099 18107 52105
rect 18233 52003 18291 52009
rect 18233 51969 18245 52003
rect 18279 52000 18291 52003
rect 18690 52000 18696 52012
rect 18279 51972 18696 52000
rect 18279 51969 18291 51972
rect 18233 51963 18291 51969
rect 18690 51960 18696 51972
rect 18748 51960 18754 52012
rect 1104 51706 18860 51728
rect 1104 51654 1950 51706
rect 2002 51654 2014 51706
rect 2066 51654 2078 51706
rect 2130 51654 2142 51706
rect 2194 51654 2206 51706
rect 2258 51654 6950 51706
rect 7002 51654 7014 51706
rect 7066 51654 7078 51706
rect 7130 51654 7142 51706
rect 7194 51654 7206 51706
rect 7258 51654 11950 51706
rect 12002 51654 12014 51706
rect 12066 51654 12078 51706
rect 12130 51654 12142 51706
rect 12194 51654 12206 51706
rect 12258 51654 16950 51706
rect 17002 51654 17014 51706
rect 17066 51654 17078 51706
rect 17130 51654 17142 51706
rect 17194 51654 17206 51706
rect 17258 51654 18860 51706
rect 1104 51632 18860 51654
rect 5353 51595 5411 51601
rect 5353 51561 5365 51595
rect 5399 51592 5411 51595
rect 7834 51592 7840 51604
rect 5399 51564 7840 51592
rect 5399 51561 5411 51564
rect 5353 51555 5411 51561
rect 7834 51552 7840 51564
rect 7892 51552 7898 51604
rect 2958 51416 2964 51468
rect 3016 51456 3022 51468
rect 3973 51459 4031 51465
rect 3973 51456 3985 51459
rect 3016 51428 3985 51456
rect 3016 51416 3022 51428
rect 3973 51425 3985 51428
rect 4019 51425 4031 51459
rect 3973 51419 4031 51425
rect 10410 51416 10416 51468
rect 10468 51416 10474 51468
rect 13354 51416 13360 51468
rect 13412 51456 13418 51468
rect 14553 51459 14611 51465
rect 14553 51456 14565 51459
rect 13412 51428 14565 51456
rect 13412 51416 13418 51428
rect 14553 51425 14565 51428
rect 14599 51425 14611 51459
rect 14553 51419 14611 51425
rect 1394 51348 1400 51400
rect 1452 51388 1458 51400
rect 8573 51391 8631 51397
rect 8573 51388 8585 51391
rect 1452 51360 8585 51388
rect 1452 51348 1458 51360
rect 8573 51357 8585 51360
rect 8619 51357 8631 51391
rect 14090 51388 14096 51400
rect 8573 51351 8631 51357
rect 10612 51360 14096 51388
rect 4240 51323 4298 51329
rect 4240 51289 4252 51323
rect 4286 51320 4298 51323
rect 10612 51320 10640 51360
rect 14090 51348 14096 51360
rect 14148 51348 14154 51400
rect 14274 51348 14280 51400
rect 14332 51348 14338 51400
rect 4286 51292 10640 51320
rect 10680 51323 10738 51329
rect 4286 51289 4298 51292
rect 4240 51283 4298 51289
rect 10680 51289 10692 51323
rect 10726 51289 10738 51323
rect 10680 51283 10738 51289
rect 4154 51212 4160 51264
rect 4212 51252 4218 51264
rect 8389 51255 8447 51261
rect 8389 51252 8401 51255
rect 4212 51224 8401 51252
rect 4212 51212 4218 51224
rect 8389 51221 8401 51224
rect 8435 51221 8447 51255
rect 8389 51215 8447 51221
rect 10594 51212 10600 51264
rect 10652 51252 10658 51264
rect 10704 51252 10732 51283
rect 10652 51224 10732 51252
rect 10652 51212 10658 51224
rect 11238 51212 11244 51264
rect 11296 51252 11302 51264
rect 11793 51255 11851 51261
rect 11793 51252 11805 51255
rect 11296 51224 11805 51252
rect 11296 51212 11302 51224
rect 11793 51221 11805 51224
rect 11839 51221 11851 51255
rect 11793 51215 11851 51221
rect 1104 51162 18860 51184
rect 1104 51110 2610 51162
rect 2662 51110 2674 51162
rect 2726 51110 2738 51162
rect 2790 51110 2802 51162
rect 2854 51110 2866 51162
rect 2918 51110 7610 51162
rect 7662 51110 7674 51162
rect 7726 51110 7738 51162
rect 7790 51110 7802 51162
rect 7854 51110 7866 51162
rect 7918 51110 12610 51162
rect 12662 51110 12674 51162
rect 12726 51110 12738 51162
rect 12790 51110 12802 51162
rect 12854 51110 12866 51162
rect 12918 51110 17610 51162
rect 17662 51110 17674 51162
rect 17726 51110 17738 51162
rect 17790 51110 17802 51162
rect 17854 51110 17866 51162
rect 17918 51110 18860 51162
rect 1104 51088 18860 51110
rect 6086 50940 6092 50992
rect 6144 50980 6150 50992
rect 8018 50980 8024 50992
rect 6144 50952 8024 50980
rect 6144 50940 6150 50952
rect 8018 50940 8024 50952
rect 8076 50940 8082 50992
rect 8389 50915 8447 50921
rect 8389 50881 8401 50915
rect 8435 50912 8447 50915
rect 8665 50915 8723 50921
rect 8665 50912 8677 50915
rect 8435 50884 8677 50912
rect 8435 50881 8447 50884
rect 8389 50875 8447 50881
rect 8665 50881 8677 50884
rect 8711 50912 8723 50915
rect 9300 50915 9358 50921
rect 9300 50912 9312 50915
rect 8711 50884 9312 50912
rect 8711 50881 8723 50884
rect 8665 50875 8723 50881
rect 9300 50881 9312 50884
rect 9346 50912 9358 50915
rect 10686 50912 10692 50924
rect 9346 50884 10692 50912
rect 9346 50881 9358 50884
rect 9300 50875 9358 50881
rect 10686 50872 10692 50884
rect 10744 50872 10750 50924
rect 13170 50872 13176 50924
rect 13228 50912 13234 50924
rect 18049 50915 18107 50921
rect 18049 50912 18061 50915
rect 13228 50884 18061 50912
rect 13228 50872 13234 50884
rect 18049 50881 18061 50884
rect 18095 50881 18107 50915
rect 18049 50875 18107 50881
rect 8018 50804 8024 50856
rect 8076 50844 8082 50856
rect 9033 50847 9091 50853
rect 9033 50844 9045 50847
rect 8076 50816 9045 50844
rect 8076 50804 8082 50816
rect 9033 50813 9045 50816
rect 9079 50813 9091 50847
rect 9033 50807 9091 50813
rect 8110 50736 8116 50788
rect 8168 50776 8174 50788
rect 8754 50776 8760 50788
rect 8168 50748 8760 50776
rect 8168 50736 8174 50748
rect 8754 50736 8760 50748
rect 8812 50736 8818 50788
rect 2314 50668 2320 50720
rect 2372 50708 2378 50720
rect 2590 50708 2596 50720
rect 2372 50680 2596 50708
rect 2372 50668 2378 50680
rect 2590 50668 2596 50680
rect 2648 50668 2654 50720
rect 9306 50668 9312 50720
rect 9364 50708 9370 50720
rect 10413 50711 10471 50717
rect 10413 50708 10425 50711
rect 9364 50680 10425 50708
rect 9364 50668 9370 50680
rect 10413 50677 10425 50680
rect 10459 50677 10471 50711
rect 10413 50671 10471 50677
rect 10686 50668 10692 50720
rect 10744 50668 10750 50720
rect 18230 50668 18236 50720
rect 18288 50668 18294 50720
rect 1104 50618 18860 50640
rect 1104 50566 1950 50618
rect 2002 50566 2014 50618
rect 2066 50566 2078 50618
rect 2130 50566 2142 50618
rect 2194 50566 2206 50618
rect 2258 50566 6950 50618
rect 7002 50566 7014 50618
rect 7066 50566 7078 50618
rect 7130 50566 7142 50618
rect 7194 50566 7206 50618
rect 7258 50566 11950 50618
rect 12002 50566 12014 50618
rect 12066 50566 12078 50618
rect 12130 50566 12142 50618
rect 12194 50566 12206 50618
rect 12258 50566 16950 50618
rect 17002 50566 17014 50618
rect 17066 50566 17078 50618
rect 17130 50566 17142 50618
rect 17194 50566 17206 50618
rect 17258 50566 18860 50618
rect 1104 50544 18860 50566
rect 2777 50439 2835 50445
rect 2777 50405 2789 50439
rect 2823 50436 2835 50439
rect 3142 50436 3148 50448
rect 2823 50408 3148 50436
rect 2823 50405 2835 50408
rect 2777 50399 2835 50405
rect 3142 50396 3148 50408
rect 3200 50396 3206 50448
rect 3237 50371 3295 50377
rect 3237 50337 3249 50371
rect 3283 50368 3295 50371
rect 4798 50368 4804 50380
rect 3283 50340 4804 50368
rect 3283 50337 3295 50340
rect 3237 50331 3295 50337
rect 4798 50328 4804 50340
rect 4856 50328 4862 50380
rect 3326 50260 3332 50312
rect 3384 50260 3390 50312
rect 5074 50260 5080 50312
rect 5132 50300 5138 50312
rect 14461 50303 14519 50309
rect 14461 50300 14473 50303
rect 5132 50272 14473 50300
rect 5132 50260 5138 50272
rect 14461 50269 14473 50272
rect 14507 50269 14519 50303
rect 14461 50263 14519 50269
rect 3237 50167 3295 50173
rect 3237 50133 3249 50167
rect 3283 50164 3295 50167
rect 7558 50164 7564 50176
rect 3283 50136 7564 50164
rect 3283 50133 3295 50136
rect 3237 50127 3295 50133
rect 7558 50124 7564 50136
rect 7616 50124 7622 50176
rect 14277 50167 14335 50173
rect 14277 50133 14289 50167
rect 14323 50164 14335 50167
rect 14550 50164 14556 50176
rect 14323 50136 14556 50164
rect 14323 50133 14335 50136
rect 14277 50127 14335 50133
rect 14550 50124 14556 50136
rect 14608 50124 14614 50176
rect 1104 50074 18860 50096
rect 1104 50022 2610 50074
rect 2662 50022 2674 50074
rect 2726 50022 2738 50074
rect 2790 50022 2802 50074
rect 2854 50022 2866 50074
rect 2918 50022 7610 50074
rect 7662 50022 7674 50074
rect 7726 50022 7738 50074
rect 7790 50022 7802 50074
rect 7854 50022 7866 50074
rect 7918 50022 12610 50074
rect 12662 50022 12674 50074
rect 12726 50022 12738 50074
rect 12790 50022 12802 50074
rect 12854 50022 12866 50074
rect 12918 50022 17610 50074
rect 17662 50022 17674 50074
rect 17726 50022 17738 50074
rect 17790 50022 17802 50074
rect 17854 50022 17866 50074
rect 17918 50022 18860 50074
rect 1104 50000 18860 50022
rect 1854 49920 1860 49972
rect 1912 49960 1918 49972
rect 3694 49960 3700 49972
rect 1912 49932 3700 49960
rect 1912 49920 1918 49932
rect 3694 49920 3700 49932
rect 3752 49920 3758 49972
rect 4430 49920 4436 49972
rect 4488 49920 4494 49972
rect 3320 49895 3378 49901
rect 3320 49861 3332 49895
rect 3366 49892 3378 49895
rect 4154 49892 4160 49904
rect 3366 49864 4160 49892
rect 3366 49861 3378 49864
rect 3320 49855 3378 49861
rect 4154 49852 4160 49864
rect 4212 49852 4218 49904
rect 8294 49901 8300 49904
rect 8288 49892 8300 49901
rect 8255 49864 8300 49892
rect 8288 49855 8300 49864
rect 8294 49852 8300 49855
rect 8352 49852 8358 49904
rect 2958 49716 2964 49768
rect 3016 49756 3022 49768
rect 3053 49759 3111 49765
rect 3053 49756 3065 49759
rect 3016 49728 3065 49756
rect 3016 49716 3022 49728
rect 3053 49725 3065 49728
rect 3099 49725 3111 49759
rect 3053 49719 3111 49725
rect 3068 49620 3096 49719
rect 8018 49716 8024 49768
rect 8076 49716 8082 49768
rect 9582 49756 9588 49768
rect 9416 49728 9588 49756
rect 9416 49697 9444 49728
rect 9582 49716 9588 49728
rect 9640 49756 9646 49768
rect 16850 49756 16856 49768
rect 9640 49728 16856 49756
rect 9640 49716 9646 49728
rect 16850 49716 16856 49728
rect 16908 49716 16914 49768
rect 9401 49691 9459 49697
rect 9401 49657 9413 49691
rect 9447 49657 9459 49691
rect 9401 49651 9459 49657
rect 3418 49620 3424 49632
rect 3068 49592 3424 49620
rect 3418 49580 3424 49592
rect 3476 49580 3482 49632
rect 1104 49530 18860 49552
rect 1104 49478 1950 49530
rect 2002 49478 2014 49530
rect 2066 49478 2078 49530
rect 2130 49478 2142 49530
rect 2194 49478 2206 49530
rect 2258 49478 6950 49530
rect 7002 49478 7014 49530
rect 7066 49478 7078 49530
rect 7130 49478 7142 49530
rect 7194 49478 7206 49530
rect 7258 49478 11950 49530
rect 12002 49478 12014 49530
rect 12066 49478 12078 49530
rect 12130 49478 12142 49530
rect 12194 49478 12206 49530
rect 12258 49478 16950 49530
rect 17002 49478 17014 49530
rect 17066 49478 17078 49530
rect 17130 49478 17142 49530
rect 17194 49478 17206 49530
rect 17258 49478 18860 49530
rect 1104 49456 18860 49478
rect 7377 49351 7435 49357
rect 7377 49317 7389 49351
rect 7423 49348 7435 49351
rect 13998 49348 14004 49360
rect 7423 49320 14004 49348
rect 7423 49317 7435 49320
rect 7377 49311 7435 49317
rect 13998 49308 14004 49320
rect 14056 49308 14062 49360
rect 3418 49172 3424 49224
rect 3476 49212 3482 49224
rect 5997 49215 6055 49221
rect 5997 49212 6009 49215
rect 3476 49184 6009 49212
rect 3476 49172 3482 49184
rect 5997 49181 6009 49184
rect 6043 49212 6055 49215
rect 8018 49212 8024 49224
rect 6043 49184 8024 49212
rect 6043 49181 6055 49184
rect 5997 49175 6055 49181
rect 8018 49172 8024 49184
rect 8076 49172 8082 49224
rect 6264 49147 6322 49153
rect 6264 49113 6276 49147
rect 6310 49144 6322 49147
rect 16390 49144 16396 49156
rect 6310 49116 16396 49144
rect 6310 49113 6322 49116
rect 6264 49107 6322 49113
rect 16390 49104 16396 49116
rect 16448 49104 16454 49156
rect 8018 49036 8024 49088
rect 8076 49076 8082 49088
rect 8570 49076 8576 49088
rect 8076 49048 8576 49076
rect 8076 49036 8082 49048
rect 8570 49036 8576 49048
rect 8628 49036 8634 49088
rect 1104 48986 18860 49008
rect 1104 48934 2610 48986
rect 2662 48934 2674 48986
rect 2726 48934 2738 48986
rect 2790 48934 2802 48986
rect 2854 48934 2866 48986
rect 2918 48934 7610 48986
rect 7662 48934 7674 48986
rect 7726 48934 7738 48986
rect 7790 48934 7802 48986
rect 7854 48934 7866 48986
rect 7918 48934 12610 48986
rect 12662 48934 12674 48986
rect 12726 48934 12738 48986
rect 12790 48934 12802 48986
rect 12854 48934 12866 48986
rect 12918 48934 17610 48986
rect 17662 48934 17674 48986
rect 17726 48934 17738 48986
rect 17790 48934 17802 48986
rect 17854 48934 17866 48986
rect 17918 48934 18860 48986
rect 1104 48912 18860 48934
rect 7466 48832 7472 48884
rect 7524 48832 7530 48884
rect 14090 48832 14096 48884
rect 14148 48872 14154 48884
rect 15841 48875 15899 48881
rect 15841 48872 15853 48875
rect 14148 48844 15853 48872
rect 14148 48832 14154 48844
rect 15841 48841 15853 48844
rect 15887 48841 15899 48875
rect 15841 48835 15899 48841
rect 10226 48764 10232 48816
rect 10284 48804 10290 48816
rect 10689 48807 10747 48813
rect 10689 48804 10701 48807
rect 10284 48776 10701 48804
rect 10284 48764 10290 48776
rect 10689 48773 10701 48776
rect 10735 48804 10747 48807
rect 10778 48804 10784 48816
rect 10735 48776 10784 48804
rect 10735 48773 10747 48776
rect 10689 48767 10747 48773
rect 10778 48764 10784 48776
rect 10836 48764 10842 48816
rect 12406 48776 16574 48804
rect 3694 48745 3700 48748
rect 3145 48739 3203 48745
rect 3145 48705 3157 48739
rect 3191 48736 3203 48739
rect 3688 48736 3700 48745
rect 3191 48708 3700 48736
rect 3191 48705 3203 48708
rect 3145 48699 3203 48705
rect 3688 48699 3700 48708
rect 3694 48696 3700 48699
rect 3752 48696 3758 48748
rect 7653 48739 7711 48745
rect 7653 48705 7665 48739
rect 7699 48736 7711 48739
rect 8570 48736 8576 48748
rect 7699 48708 8576 48736
rect 7699 48705 7711 48708
rect 7653 48699 7711 48705
rect 8570 48696 8576 48708
rect 8628 48696 8634 48748
rect 12406 48736 12434 48776
rect 8680 48708 12434 48736
rect 3418 48628 3424 48680
rect 3476 48628 3482 48680
rect 4801 48603 4859 48609
rect 4801 48569 4813 48603
rect 4847 48600 4859 48603
rect 6270 48600 6276 48612
rect 4847 48572 6276 48600
rect 4847 48569 4859 48572
rect 4801 48563 4859 48569
rect 6270 48560 6276 48572
rect 6328 48600 6334 48612
rect 8680 48600 8708 48708
rect 14642 48696 14648 48748
rect 14700 48696 14706 48748
rect 16022 48696 16028 48748
rect 16080 48696 16086 48748
rect 16546 48736 16574 48776
rect 18049 48739 18107 48745
rect 18049 48736 18061 48739
rect 16546 48708 18061 48736
rect 18049 48705 18061 48708
rect 18095 48705 18107 48739
rect 18049 48699 18107 48705
rect 10686 48628 10692 48680
rect 10744 48668 10750 48680
rect 10781 48671 10839 48677
rect 10781 48668 10793 48671
rect 10744 48640 10793 48668
rect 10744 48628 10750 48640
rect 10781 48637 10793 48640
rect 10827 48637 10839 48671
rect 10781 48631 10839 48637
rect 10873 48671 10931 48677
rect 10873 48637 10885 48671
rect 10919 48637 10931 48671
rect 10873 48631 10931 48637
rect 6328 48572 8708 48600
rect 6328 48560 6334 48572
rect 10042 48560 10048 48612
rect 10100 48600 10106 48612
rect 10226 48600 10232 48612
rect 10100 48572 10232 48600
rect 10100 48560 10106 48572
rect 10226 48560 10232 48572
rect 10284 48600 10290 48612
rect 10888 48600 10916 48631
rect 11054 48628 11060 48680
rect 11112 48668 11118 48680
rect 14734 48668 14740 48680
rect 11112 48640 14740 48668
rect 11112 48628 11118 48640
rect 14734 48628 14740 48640
rect 14792 48628 14798 48680
rect 14921 48671 14979 48677
rect 14921 48637 14933 48671
rect 14967 48668 14979 48671
rect 15010 48668 15016 48680
rect 14967 48640 15016 48668
rect 14967 48637 14979 48640
rect 14921 48631 14979 48637
rect 15010 48628 15016 48640
rect 15068 48668 15074 48680
rect 15378 48668 15384 48680
rect 15068 48640 15384 48668
rect 15068 48628 15074 48640
rect 15378 48628 15384 48640
rect 15436 48628 15442 48680
rect 10284 48572 10916 48600
rect 14277 48603 14335 48609
rect 10284 48560 10290 48572
rect 14277 48569 14289 48603
rect 14323 48600 14335 48603
rect 16666 48600 16672 48612
rect 14323 48572 16672 48600
rect 14323 48569 14335 48572
rect 14277 48563 14335 48569
rect 16666 48560 16672 48572
rect 16724 48560 16730 48612
rect 6638 48492 6644 48544
rect 6696 48532 6702 48544
rect 10321 48535 10379 48541
rect 10321 48532 10333 48535
rect 6696 48504 10333 48532
rect 6696 48492 6702 48504
rect 10321 48501 10333 48504
rect 10367 48501 10379 48535
rect 10321 48495 10379 48501
rect 10686 48492 10692 48544
rect 10744 48532 10750 48544
rect 15654 48532 15660 48544
rect 10744 48504 15660 48532
rect 10744 48492 10750 48504
rect 15654 48492 15660 48504
rect 15712 48492 15718 48544
rect 18230 48492 18236 48544
rect 18288 48492 18294 48544
rect 1104 48442 18860 48464
rect 1104 48390 1950 48442
rect 2002 48390 2014 48442
rect 2066 48390 2078 48442
rect 2130 48390 2142 48442
rect 2194 48390 2206 48442
rect 2258 48390 6950 48442
rect 7002 48390 7014 48442
rect 7066 48390 7078 48442
rect 7130 48390 7142 48442
rect 7194 48390 7206 48442
rect 7258 48390 11950 48442
rect 12002 48390 12014 48442
rect 12066 48390 12078 48442
rect 12130 48390 12142 48442
rect 12194 48390 12206 48442
rect 12258 48390 16950 48442
rect 17002 48390 17014 48442
rect 17066 48390 17078 48442
rect 17130 48390 17142 48442
rect 17194 48390 17206 48442
rect 17258 48390 18860 48442
rect 1104 48368 18860 48390
rect 1578 48288 1584 48340
rect 1636 48328 1642 48340
rect 6638 48328 6644 48340
rect 1636 48300 6644 48328
rect 1636 48288 1642 48300
rect 6638 48288 6644 48300
rect 6696 48288 6702 48340
rect 10042 48288 10048 48340
rect 10100 48328 10106 48340
rect 10686 48328 10692 48340
rect 10100 48300 10692 48328
rect 10100 48288 10106 48300
rect 10686 48288 10692 48300
rect 10744 48288 10750 48340
rect 1104 47898 18860 47920
rect 1104 47846 2610 47898
rect 2662 47846 2674 47898
rect 2726 47846 2738 47898
rect 2790 47846 2802 47898
rect 2854 47846 2866 47898
rect 2918 47846 7610 47898
rect 7662 47846 7674 47898
rect 7726 47846 7738 47898
rect 7790 47846 7802 47898
rect 7854 47846 7866 47898
rect 7918 47846 12610 47898
rect 12662 47846 12674 47898
rect 12726 47846 12738 47898
rect 12790 47846 12802 47898
rect 12854 47846 12866 47898
rect 12918 47846 17610 47898
rect 17662 47846 17674 47898
rect 17726 47846 17738 47898
rect 17790 47846 17802 47898
rect 17854 47846 17866 47898
rect 17918 47846 18860 47898
rect 1104 47824 18860 47846
rect 2409 47787 2467 47793
rect 2409 47753 2421 47787
rect 2455 47784 2467 47787
rect 6178 47784 6184 47796
rect 2455 47756 6184 47784
rect 2455 47753 2467 47756
rect 2409 47747 2467 47753
rect 6178 47744 6184 47756
rect 6236 47744 6242 47796
rect 6454 47744 6460 47796
rect 6512 47784 6518 47796
rect 6549 47787 6607 47793
rect 6549 47784 6561 47787
rect 6512 47756 6561 47784
rect 6512 47744 6518 47756
rect 6549 47753 6561 47756
rect 6595 47753 6607 47787
rect 6549 47747 6607 47753
rect 7650 47744 7656 47796
rect 7708 47784 7714 47796
rect 8386 47784 8392 47796
rect 7708 47756 8392 47784
rect 7708 47744 7714 47756
rect 8386 47744 8392 47756
rect 8444 47744 8450 47796
rect 11885 47787 11943 47793
rect 11885 47753 11897 47787
rect 11931 47784 11943 47787
rect 11931 47756 12434 47784
rect 11931 47753 11943 47756
rect 11885 47747 11943 47753
rect 7009 47719 7067 47725
rect 7009 47685 7021 47719
rect 7055 47716 7067 47719
rect 8846 47716 8852 47728
rect 7055 47688 8852 47716
rect 7055 47685 7067 47688
rect 7009 47679 7067 47685
rect 8846 47676 8852 47688
rect 8904 47676 8910 47728
rect 12406 47716 12434 47756
rect 13142 47719 13200 47725
rect 13142 47716 13154 47719
rect 12406 47688 13154 47716
rect 13142 47685 13154 47688
rect 13188 47685 13200 47719
rect 13142 47679 13200 47685
rect 2317 47651 2375 47657
rect 2317 47617 2329 47651
rect 2363 47648 2375 47651
rect 2958 47648 2964 47660
rect 2363 47620 2964 47648
rect 2363 47617 2375 47620
rect 2317 47611 2375 47617
rect 2958 47608 2964 47620
rect 3016 47608 3022 47660
rect 3050 47608 3056 47660
rect 3108 47608 3114 47660
rect 4985 47651 5043 47657
rect 4985 47617 4997 47651
rect 5031 47617 5043 47651
rect 4985 47611 5043 47617
rect 6917 47651 6975 47657
rect 6917 47617 6929 47651
rect 6963 47648 6975 47651
rect 7374 47648 7380 47660
rect 6963 47620 7380 47648
rect 6963 47617 6975 47620
rect 6917 47611 6975 47617
rect 3237 47515 3295 47521
rect 3237 47481 3249 47515
rect 3283 47512 3295 47515
rect 3970 47512 3976 47524
rect 3283 47484 3976 47512
rect 3283 47481 3295 47484
rect 3237 47475 3295 47481
rect 3970 47472 3976 47484
rect 4028 47472 4034 47524
rect 5000 47512 5028 47611
rect 7374 47608 7380 47620
rect 7432 47608 7438 47660
rect 7466 47608 7472 47660
rect 7524 47648 7530 47660
rect 7742 47648 7748 47660
rect 7524 47620 7748 47648
rect 7524 47608 7530 47620
rect 7742 47608 7748 47620
rect 7800 47608 7806 47660
rect 10502 47608 10508 47660
rect 10560 47648 10566 47660
rect 12069 47651 12127 47657
rect 12069 47648 12081 47651
rect 10560 47620 12081 47648
rect 10560 47608 10566 47620
rect 12069 47617 12081 47620
rect 12115 47617 12127 47651
rect 12069 47611 12127 47617
rect 7193 47583 7251 47589
rect 7193 47549 7205 47583
rect 7239 47580 7251 47583
rect 11514 47580 11520 47592
rect 7239 47552 11520 47580
rect 7239 47549 7251 47552
rect 7193 47543 7251 47549
rect 11514 47540 11520 47552
rect 11572 47540 11578 47592
rect 12434 47540 12440 47592
rect 12492 47580 12498 47592
rect 12897 47583 12955 47589
rect 12897 47580 12909 47583
rect 12492 47552 12909 47580
rect 12492 47540 12498 47552
rect 12897 47549 12909 47552
rect 12943 47549 12955 47583
rect 12897 47543 12955 47549
rect 7558 47512 7564 47524
rect 5000 47484 7564 47512
rect 7558 47472 7564 47484
rect 7616 47472 7622 47524
rect 4798 47404 4804 47456
rect 4856 47404 4862 47456
rect 13078 47404 13084 47456
rect 13136 47444 13142 47456
rect 14277 47447 14335 47453
rect 14277 47444 14289 47447
rect 13136 47416 14289 47444
rect 13136 47404 13142 47416
rect 14277 47413 14289 47416
rect 14323 47444 14335 47447
rect 19242 47444 19248 47456
rect 14323 47416 19248 47444
rect 14323 47413 14335 47416
rect 14277 47407 14335 47413
rect 19242 47404 19248 47416
rect 19300 47404 19306 47456
rect 1104 47354 18860 47376
rect 1104 47302 1950 47354
rect 2002 47302 2014 47354
rect 2066 47302 2078 47354
rect 2130 47302 2142 47354
rect 2194 47302 2206 47354
rect 2258 47302 6950 47354
rect 7002 47302 7014 47354
rect 7066 47302 7078 47354
rect 7130 47302 7142 47354
rect 7194 47302 7206 47354
rect 7258 47302 11950 47354
rect 12002 47302 12014 47354
rect 12066 47302 12078 47354
rect 12130 47302 12142 47354
rect 12194 47302 12206 47354
rect 12258 47302 16950 47354
rect 17002 47302 17014 47354
rect 17066 47302 17078 47354
rect 17130 47302 17142 47354
rect 17194 47302 17206 47354
rect 17258 47302 18860 47354
rect 1104 47280 18860 47302
rect 2777 47175 2835 47181
rect 2777 47141 2789 47175
rect 2823 47172 2835 47175
rect 3050 47172 3056 47184
rect 2823 47144 3056 47172
rect 2823 47141 2835 47144
rect 2777 47135 2835 47141
rect 3050 47132 3056 47144
rect 3108 47132 3114 47184
rect 7377 47175 7435 47181
rect 7377 47141 7389 47175
rect 7423 47172 7435 47175
rect 11422 47172 11428 47184
rect 7423 47144 11428 47172
rect 7423 47141 7435 47144
rect 7377 47135 7435 47141
rect 11422 47132 11428 47144
rect 11480 47132 11486 47184
rect 2958 47064 2964 47116
rect 3016 47104 3022 47116
rect 15102 47104 15108 47116
rect 3016 47076 15108 47104
rect 3016 47064 3022 47076
rect 15102 47064 15108 47076
rect 15160 47064 15166 47116
rect 3053 47039 3111 47045
rect 3053 47005 3065 47039
rect 3099 47036 3111 47039
rect 7561 47039 7619 47045
rect 3099 47008 5764 47036
rect 3099 47005 3111 47008
rect 3053 46999 3111 47005
rect 3234 46928 3240 46980
rect 3292 46928 3298 46980
rect 3329 46971 3387 46977
rect 3329 46937 3341 46971
rect 3375 46968 3387 46971
rect 3786 46968 3792 46980
rect 3375 46940 3792 46968
rect 3375 46937 3387 46940
rect 3329 46931 3387 46937
rect 3786 46928 3792 46940
rect 3844 46928 3850 46980
rect 5736 46968 5764 47008
rect 7561 47005 7573 47039
rect 7607 47036 7619 47039
rect 7742 47036 7748 47048
rect 7607 47008 7748 47036
rect 7607 47005 7619 47008
rect 7561 46999 7619 47005
rect 7742 46996 7748 47008
rect 7800 46996 7806 47048
rect 15838 46996 15844 47048
rect 15896 47036 15902 47048
rect 16482 47036 16488 47048
rect 15896 47008 16488 47036
rect 15896 46996 15902 47008
rect 16482 46996 16488 47008
rect 16540 47036 16546 47048
rect 18049 47039 18107 47045
rect 18049 47036 18061 47039
rect 16540 47008 18061 47036
rect 16540 46996 16546 47008
rect 18049 47005 18061 47008
rect 18095 47005 18107 47039
rect 18049 46999 18107 47005
rect 7650 46968 7656 46980
rect 5736 46940 7656 46968
rect 7650 46928 7656 46940
rect 7708 46928 7714 46980
rect 18230 46860 18236 46912
rect 18288 46860 18294 46912
rect 1104 46810 18860 46832
rect 1104 46758 2610 46810
rect 2662 46758 2674 46810
rect 2726 46758 2738 46810
rect 2790 46758 2802 46810
rect 2854 46758 2866 46810
rect 2918 46758 7610 46810
rect 7662 46758 7674 46810
rect 7726 46758 7738 46810
rect 7790 46758 7802 46810
rect 7854 46758 7866 46810
rect 7918 46758 12610 46810
rect 12662 46758 12674 46810
rect 12726 46758 12738 46810
rect 12790 46758 12802 46810
rect 12854 46758 12866 46810
rect 12918 46758 17610 46810
rect 17662 46758 17674 46810
rect 17726 46758 17738 46810
rect 17790 46758 17802 46810
rect 17854 46758 17866 46810
rect 17918 46758 18860 46810
rect 1104 46736 18860 46758
rect 3970 46656 3976 46708
rect 4028 46696 4034 46708
rect 4028 46668 16574 46696
rect 4028 46656 4034 46668
rect 12526 46637 12532 46640
rect 12520 46628 12532 46637
rect 12487 46600 12532 46628
rect 12520 46591 12532 46600
rect 12526 46588 12532 46591
rect 12584 46588 12590 46640
rect 16546 46560 16574 46668
rect 16850 46560 16856 46572
rect 16546 46532 16856 46560
rect 16850 46520 16856 46532
rect 16908 46520 16914 46572
rect 12253 46495 12311 46501
rect 12253 46461 12265 46495
rect 12299 46461 12311 46495
rect 12253 46455 12311 46461
rect 6454 46316 6460 46368
rect 6512 46356 6518 46368
rect 8018 46356 8024 46368
rect 6512 46328 8024 46356
rect 6512 46316 6518 46328
rect 8018 46316 8024 46328
rect 8076 46316 8082 46368
rect 12268 46356 12296 46455
rect 12434 46356 12440 46368
rect 12268 46328 12440 46356
rect 12434 46316 12440 46328
rect 12492 46316 12498 46368
rect 13630 46316 13636 46368
rect 13688 46316 13694 46368
rect 1104 46266 18860 46288
rect 1104 46214 1950 46266
rect 2002 46214 2014 46266
rect 2066 46214 2078 46266
rect 2130 46214 2142 46266
rect 2194 46214 2206 46266
rect 2258 46214 6950 46266
rect 7002 46214 7014 46266
rect 7066 46214 7078 46266
rect 7130 46214 7142 46266
rect 7194 46214 7206 46266
rect 7258 46214 11950 46266
rect 12002 46214 12014 46266
rect 12066 46214 12078 46266
rect 12130 46214 12142 46266
rect 12194 46214 12206 46266
rect 12258 46214 16950 46266
rect 17002 46214 17014 46266
rect 17066 46214 17078 46266
rect 17130 46214 17142 46266
rect 17194 46214 17206 46266
rect 17258 46214 18860 46266
rect 1104 46192 18860 46214
rect 7282 46112 7288 46164
rect 7340 46152 7346 46164
rect 8018 46152 8024 46164
rect 7340 46124 8024 46152
rect 7340 46112 7346 46124
rect 8018 46112 8024 46124
rect 8076 46112 8082 46164
rect 1104 45722 18860 45744
rect 1104 45670 2610 45722
rect 2662 45670 2674 45722
rect 2726 45670 2738 45722
rect 2790 45670 2802 45722
rect 2854 45670 2866 45722
rect 2918 45670 7610 45722
rect 7662 45670 7674 45722
rect 7726 45670 7738 45722
rect 7790 45670 7802 45722
rect 7854 45670 7866 45722
rect 7918 45670 12610 45722
rect 12662 45670 12674 45722
rect 12726 45670 12738 45722
rect 12790 45670 12802 45722
rect 12854 45670 12866 45722
rect 12918 45670 17610 45722
rect 17662 45670 17674 45722
rect 17726 45670 17738 45722
rect 17790 45670 17802 45722
rect 17854 45670 17866 45722
rect 17918 45670 18860 45722
rect 1104 45648 18860 45670
rect 7282 45568 7288 45620
rect 7340 45608 7346 45620
rect 12434 45608 12440 45620
rect 7340 45580 12440 45608
rect 7340 45568 7346 45580
rect 12434 45568 12440 45580
rect 12492 45568 12498 45620
rect 1104 45178 18860 45200
rect 1104 45126 1950 45178
rect 2002 45126 2014 45178
rect 2066 45126 2078 45178
rect 2130 45126 2142 45178
rect 2194 45126 2206 45178
rect 2258 45126 6950 45178
rect 7002 45126 7014 45178
rect 7066 45126 7078 45178
rect 7130 45126 7142 45178
rect 7194 45126 7206 45178
rect 7258 45126 11950 45178
rect 12002 45126 12014 45178
rect 12066 45126 12078 45178
rect 12130 45126 12142 45178
rect 12194 45126 12206 45178
rect 12258 45126 16950 45178
rect 17002 45126 17014 45178
rect 17066 45126 17078 45178
rect 17130 45126 17142 45178
rect 17194 45126 17206 45178
rect 17258 45126 18860 45178
rect 1104 45104 18860 45126
rect 13538 45024 13544 45076
rect 13596 45064 13602 45076
rect 13814 45064 13820 45076
rect 13596 45036 13820 45064
rect 13596 45024 13602 45036
rect 13814 45024 13820 45036
rect 13872 45024 13878 45076
rect 16390 45024 16396 45076
rect 16448 45024 16454 45076
rect 12434 44888 12440 44940
rect 12492 44928 12498 44940
rect 14277 44931 14335 44937
rect 14277 44928 14289 44931
rect 12492 44900 14289 44928
rect 12492 44888 12498 44900
rect 14277 44897 14289 44900
rect 14323 44897 14335 44931
rect 14277 44891 14335 44897
rect 14550 44888 14556 44940
rect 14608 44888 14614 44940
rect 11698 44820 11704 44872
rect 11756 44860 11762 44872
rect 13081 44863 13139 44869
rect 13081 44860 13093 44863
rect 11756 44832 13093 44860
rect 11756 44820 11762 44832
rect 13081 44829 13093 44832
rect 13127 44860 13139 44863
rect 13127 44832 13676 44860
rect 13127 44829 13139 44832
rect 13081 44823 13139 44829
rect 2498 44752 2504 44804
rect 2556 44792 2562 44804
rect 4430 44792 4436 44804
rect 2556 44764 4436 44792
rect 2556 44752 2562 44764
rect 4430 44752 4436 44764
rect 4488 44752 4494 44804
rect 11514 44752 11520 44804
rect 11572 44792 11578 44804
rect 13446 44792 13452 44804
rect 11572 44764 13452 44792
rect 11572 44752 11578 44764
rect 13446 44752 13452 44764
rect 13504 44752 13510 44804
rect 13648 44792 13676 44832
rect 13722 44820 13728 44872
rect 13780 44860 13786 44872
rect 16577 44863 16635 44869
rect 16577 44860 16589 44863
rect 13780 44832 16589 44860
rect 13780 44820 13786 44832
rect 16577 44829 16589 44832
rect 16623 44829 16635 44863
rect 16577 44823 16635 44829
rect 18049 44863 18107 44869
rect 18049 44829 18061 44863
rect 18095 44860 18107 44863
rect 19518 44860 19524 44872
rect 18095 44832 19524 44860
rect 18095 44829 18107 44832
rect 18049 44823 18107 44829
rect 19518 44820 19524 44832
rect 19576 44820 19582 44872
rect 13998 44792 14004 44804
rect 13648 44764 14004 44792
rect 13998 44752 14004 44764
rect 14056 44752 14062 44804
rect 2130 44684 2136 44736
rect 2188 44724 2194 44736
rect 3878 44724 3884 44736
rect 2188 44696 3884 44724
rect 2188 44684 2194 44696
rect 3878 44684 3884 44696
rect 3936 44724 3942 44736
rect 6086 44724 6092 44736
rect 3936 44696 6092 44724
rect 3936 44684 3942 44696
rect 6086 44684 6092 44696
rect 6144 44684 6150 44736
rect 15286 44684 15292 44736
rect 15344 44724 15350 44736
rect 15657 44727 15715 44733
rect 15657 44724 15669 44727
rect 15344 44696 15669 44724
rect 15344 44684 15350 44696
rect 15657 44693 15669 44696
rect 15703 44724 15715 44727
rect 16758 44724 16764 44736
rect 15703 44696 16764 44724
rect 15703 44693 15715 44696
rect 15657 44687 15715 44693
rect 16758 44684 16764 44696
rect 16816 44684 16822 44736
rect 18230 44684 18236 44736
rect 18288 44684 18294 44736
rect 1104 44634 18860 44656
rect 1104 44582 2610 44634
rect 2662 44582 2674 44634
rect 2726 44582 2738 44634
rect 2790 44582 2802 44634
rect 2854 44582 2866 44634
rect 2918 44582 7610 44634
rect 7662 44582 7674 44634
rect 7726 44582 7738 44634
rect 7790 44582 7802 44634
rect 7854 44582 7866 44634
rect 7918 44582 12610 44634
rect 12662 44582 12674 44634
rect 12726 44582 12738 44634
rect 12790 44582 12802 44634
rect 12854 44582 12866 44634
rect 12918 44582 17610 44634
rect 17662 44582 17674 44634
rect 17726 44582 17738 44634
rect 17790 44582 17802 44634
rect 17854 44582 17866 44634
rect 17918 44582 18860 44634
rect 1104 44560 18860 44582
rect 14366 44520 14372 44532
rect 1964 44492 14372 44520
rect 1964 44461 1992 44492
rect 14366 44480 14372 44492
rect 14424 44480 14430 44532
rect 1949 44455 2007 44461
rect 1949 44421 1961 44455
rect 1995 44421 2007 44455
rect 1949 44415 2007 44421
rect 2130 44412 2136 44464
rect 2188 44412 2194 44464
rect 2225 44455 2283 44461
rect 2225 44421 2237 44455
rect 2271 44452 2283 44455
rect 3326 44452 3332 44464
rect 2271 44424 3332 44452
rect 2271 44421 2283 44424
rect 2225 44415 2283 44421
rect 3326 44412 3332 44424
rect 3384 44412 3390 44464
rect 7282 44452 7288 44464
rect 4356 44424 7288 44452
rect 4356 44393 4384 44424
rect 7282 44412 7288 44424
rect 7340 44412 7346 44464
rect 4341 44387 4399 44393
rect 4341 44353 4353 44387
rect 4387 44353 4399 44387
rect 4341 44347 4399 44353
rect 2314 44276 2320 44328
rect 2372 44316 2378 44328
rect 3418 44316 3424 44328
rect 2372 44288 3424 44316
rect 2372 44276 2378 44288
rect 3418 44276 3424 44288
rect 3476 44316 3482 44328
rect 4356 44316 4384 44347
rect 4430 44344 4436 44396
rect 4488 44384 4494 44396
rect 4597 44387 4655 44393
rect 4597 44384 4609 44387
rect 4488 44356 4609 44384
rect 4488 44344 4494 44356
rect 4597 44353 4609 44356
rect 4643 44353 4655 44387
rect 4597 44347 4655 44353
rect 18322 44344 18328 44396
rect 18380 44384 18386 44396
rect 18380 44356 18920 44384
rect 18380 44344 18386 44356
rect 3476 44288 4384 44316
rect 3476 44276 3482 44288
rect 2222 44208 2228 44260
rect 2280 44248 2286 44260
rect 2498 44248 2504 44260
rect 2280 44220 2504 44248
rect 2280 44208 2286 44220
rect 2498 44208 2504 44220
rect 2556 44208 2562 44260
rect 5644 44220 12434 44248
rect 1673 44183 1731 44189
rect 1673 44149 1685 44183
rect 1719 44180 1731 44183
rect 5644 44180 5672 44220
rect 1719 44152 5672 44180
rect 1719 44149 1731 44152
rect 1673 44143 1731 44149
rect 5718 44140 5724 44192
rect 5776 44140 5782 44192
rect 8386 44140 8392 44192
rect 8444 44180 8450 44192
rect 10594 44180 10600 44192
rect 8444 44152 10600 44180
rect 8444 44140 8450 44152
rect 10594 44140 10600 44152
rect 10652 44140 10658 44192
rect 12406 44180 12434 44220
rect 18138 44180 18144 44192
rect 12406 44152 18144 44180
rect 18138 44140 18144 44152
rect 18196 44140 18202 44192
rect 18892 44112 18920 44356
rect 19426 44112 19432 44124
rect 1104 44090 18860 44112
rect 1104 44038 1950 44090
rect 2002 44038 2014 44090
rect 2066 44038 2078 44090
rect 2130 44038 2142 44090
rect 2194 44038 2206 44090
rect 2258 44038 6950 44090
rect 7002 44038 7014 44090
rect 7066 44038 7078 44090
rect 7130 44038 7142 44090
rect 7194 44038 7206 44090
rect 7258 44038 11950 44090
rect 12002 44038 12014 44090
rect 12066 44038 12078 44090
rect 12130 44038 12142 44090
rect 12194 44038 12206 44090
rect 12258 44038 16950 44090
rect 17002 44038 17014 44090
rect 17066 44038 17078 44090
rect 17130 44038 17142 44090
rect 17194 44038 17206 44090
rect 17258 44038 18860 44090
rect 18892 44084 19432 44112
rect 19426 44072 19432 44084
rect 19484 44072 19490 44124
rect 1104 44016 18860 44038
rect 3326 43800 3332 43852
rect 3384 43840 3390 43852
rect 7285 43843 7343 43849
rect 7285 43840 7297 43843
rect 3384 43812 7297 43840
rect 3384 43800 3390 43812
rect 7285 43809 7297 43812
rect 7331 43840 7343 43843
rect 9766 43840 9772 43852
rect 7331 43812 9772 43840
rect 7331 43809 7343 43812
rect 7285 43803 7343 43809
rect 9766 43800 9772 43812
rect 9824 43800 9830 43852
rect 7193 43775 7251 43781
rect 7193 43741 7205 43775
rect 7239 43772 7251 43775
rect 8754 43772 8760 43784
rect 7239 43744 8760 43772
rect 7239 43741 7251 43744
rect 7193 43735 7251 43741
rect 8754 43732 8760 43744
rect 8812 43772 8818 43784
rect 14826 43772 14832 43784
rect 8812 43744 14832 43772
rect 8812 43732 8818 43744
rect 14826 43732 14832 43744
rect 14884 43732 14890 43784
rect 7101 43707 7159 43713
rect 7101 43673 7113 43707
rect 7147 43704 7159 43707
rect 19426 43704 19432 43716
rect 7147 43676 19432 43704
rect 7147 43673 7159 43676
rect 7101 43667 7159 43673
rect 19426 43664 19432 43676
rect 19484 43664 19490 43716
rect 6730 43596 6736 43648
rect 6788 43596 6794 43648
rect 1104 43546 18860 43568
rect 1104 43494 2610 43546
rect 2662 43494 2674 43546
rect 2726 43494 2738 43546
rect 2790 43494 2802 43546
rect 2854 43494 2866 43546
rect 2918 43494 7610 43546
rect 7662 43494 7674 43546
rect 7726 43494 7738 43546
rect 7790 43494 7802 43546
rect 7854 43494 7866 43546
rect 7918 43494 12610 43546
rect 12662 43494 12674 43546
rect 12726 43494 12738 43546
rect 12790 43494 12802 43546
rect 12854 43494 12866 43546
rect 12918 43494 17610 43546
rect 17662 43494 17674 43546
rect 17726 43494 17738 43546
rect 17790 43494 17802 43546
rect 17854 43494 17866 43546
rect 17918 43494 18860 43546
rect 1104 43472 18860 43494
rect 13722 43392 13728 43444
rect 13780 43432 13786 43444
rect 18506 43432 18512 43444
rect 13780 43404 18512 43432
rect 13780 43392 13786 43404
rect 18506 43392 18512 43404
rect 18564 43392 18570 43444
rect 18049 43299 18107 43305
rect 18049 43265 18061 43299
rect 18095 43296 18107 43299
rect 18506 43296 18512 43308
rect 18095 43268 18512 43296
rect 18095 43265 18107 43268
rect 18049 43259 18107 43265
rect 18506 43256 18512 43268
rect 18564 43256 18570 43308
rect 8938 43188 8944 43240
rect 8996 43228 9002 43240
rect 12526 43228 12532 43240
rect 8996 43200 12532 43228
rect 8996 43188 9002 43200
rect 12526 43188 12532 43200
rect 12584 43188 12590 43240
rect 18230 43052 18236 43104
rect 18288 43052 18294 43104
rect 1104 43002 18860 43024
rect 1104 42950 1950 43002
rect 2002 42950 2014 43002
rect 2066 42950 2078 43002
rect 2130 42950 2142 43002
rect 2194 42950 2206 43002
rect 2258 42950 6950 43002
rect 7002 42950 7014 43002
rect 7066 42950 7078 43002
rect 7130 42950 7142 43002
rect 7194 42950 7206 43002
rect 7258 42950 11950 43002
rect 12002 42950 12014 43002
rect 12066 42950 12078 43002
rect 12130 42950 12142 43002
rect 12194 42950 12206 43002
rect 12258 42950 16950 43002
rect 17002 42950 17014 43002
rect 17066 42950 17078 43002
rect 17130 42950 17142 43002
rect 17194 42950 17206 43002
rect 17258 42950 18860 43002
rect 1104 42928 18860 42950
rect 12989 42891 13047 42897
rect 12989 42857 13001 42891
rect 13035 42857 13047 42891
rect 12989 42851 13047 42857
rect 6454 42780 6460 42832
rect 6512 42820 6518 42832
rect 6730 42820 6736 42832
rect 6512 42792 6736 42820
rect 6512 42780 6518 42792
rect 6730 42780 6736 42792
rect 6788 42780 6794 42832
rect 10962 42780 10968 42832
rect 11020 42820 11026 42832
rect 11020 42792 11100 42820
rect 11020 42780 11026 42792
rect 1670 42712 1676 42764
rect 1728 42752 1734 42764
rect 1946 42752 1952 42764
rect 1728 42724 1952 42752
rect 1728 42712 1734 42724
rect 1946 42712 1952 42724
rect 2004 42712 2010 42764
rect 2133 42755 2191 42761
rect 2133 42721 2145 42755
rect 2179 42752 2191 42755
rect 2685 42755 2743 42761
rect 2685 42752 2697 42755
rect 2179 42724 2697 42752
rect 2179 42721 2191 42724
rect 2133 42715 2191 42721
rect 2685 42721 2697 42724
rect 2731 42752 2743 42755
rect 2731 42724 6408 42752
rect 2731 42721 2743 42724
rect 2685 42715 2743 42721
rect 1486 42644 1492 42696
rect 1544 42684 1550 42696
rect 2225 42687 2283 42693
rect 2225 42684 2237 42687
rect 1544 42656 2237 42684
rect 1544 42644 1550 42656
rect 2225 42653 2237 42656
rect 2271 42653 2283 42687
rect 2225 42647 2283 42653
rect 2961 42687 3019 42693
rect 2961 42653 2973 42687
rect 3007 42684 3019 42687
rect 5442 42684 5448 42696
rect 3007 42656 5448 42684
rect 3007 42653 3019 42656
rect 2961 42647 3019 42653
rect 5442 42644 5448 42656
rect 5500 42644 5506 42696
rect 2133 42619 2191 42625
rect 2133 42585 2145 42619
rect 2179 42616 2191 42619
rect 3602 42616 3608 42628
rect 2179 42588 3608 42616
rect 2179 42585 2191 42588
rect 2133 42579 2191 42585
rect 3602 42576 3608 42588
rect 3660 42576 3666 42628
rect 1670 42557 1676 42560
rect 1663 42551 1676 42557
rect 1663 42517 1675 42551
rect 1663 42511 1676 42517
rect 1670 42508 1676 42511
rect 1728 42508 1734 42560
rect 2777 42551 2835 42557
rect 2777 42517 2789 42551
rect 2823 42548 2835 42551
rect 3326 42548 3332 42560
rect 2823 42520 3332 42548
rect 2823 42517 2835 42520
rect 2777 42511 2835 42517
rect 3326 42508 3332 42520
rect 3384 42508 3390 42560
rect 6380 42548 6408 42724
rect 7466 42712 7472 42764
rect 7524 42752 7530 42764
rect 11072 42761 11100 42792
rect 11057 42755 11115 42761
rect 7524 42724 11008 42752
rect 7524 42712 7530 42724
rect 6454 42644 6460 42696
rect 6512 42684 6518 42696
rect 9953 42687 10011 42693
rect 9953 42684 9965 42687
rect 6512 42656 9965 42684
rect 6512 42644 6518 42656
rect 9953 42653 9965 42656
rect 9999 42653 10011 42687
rect 10980 42684 11008 42724
rect 11057 42721 11069 42755
rect 11103 42721 11115 42755
rect 13004 42752 13032 42851
rect 13354 42780 13360 42832
rect 13412 42820 13418 42832
rect 13906 42820 13912 42832
rect 13412 42792 13912 42820
rect 13412 42780 13418 42792
rect 13906 42780 13912 42792
rect 13964 42780 13970 42832
rect 11057 42715 11115 42721
rect 11164 42724 13032 42752
rect 13633 42755 13691 42761
rect 11164 42684 11192 42724
rect 13633 42721 13645 42755
rect 13679 42752 13691 42755
rect 13814 42752 13820 42764
rect 13679 42724 13820 42752
rect 13679 42721 13691 42724
rect 13633 42715 13691 42721
rect 13814 42712 13820 42724
rect 13872 42712 13878 42764
rect 15194 42684 15200 42696
rect 10980 42656 11192 42684
rect 12406 42656 15200 42684
rect 9953 42647 10011 42653
rect 10410 42616 10416 42628
rect 9600 42588 10416 42616
rect 9306 42548 9312 42560
rect 6380 42520 9312 42548
rect 9306 42508 9312 42520
rect 9364 42548 9370 42560
rect 9600 42548 9628 42588
rect 10410 42576 10416 42588
rect 10468 42576 10474 42628
rect 10873 42619 10931 42625
rect 10873 42585 10885 42619
rect 10919 42616 10931 42619
rect 11698 42616 11704 42628
rect 10919 42588 11704 42616
rect 10919 42585 10931 42588
rect 10873 42579 10931 42585
rect 11698 42576 11704 42588
rect 11756 42576 11762 42628
rect 9364 42520 9628 42548
rect 9364 42508 9370 42520
rect 9674 42508 9680 42560
rect 9732 42548 9738 42560
rect 9769 42551 9827 42557
rect 9769 42548 9781 42551
rect 9732 42520 9781 42548
rect 9732 42508 9738 42520
rect 9769 42517 9781 42520
rect 9815 42517 9827 42551
rect 9769 42511 9827 42517
rect 10502 42508 10508 42560
rect 10560 42508 10566 42560
rect 10686 42508 10692 42560
rect 10744 42548 10750 42560
rect 10965 42551 11023 42557
rect 10965 42548 10977 42551
rect 10744 42520 10977 42548
rect 10744 42508 10750 42520
rect 10965 42517 10977 42520
rect 11011 42548 11023 42551
rect 12406 42548 12434 42656
rect 15194 42644 15200 42656
rect 15252 42644 15258 42696
rect 13357 42619 13415 42625
rect 13357 42585 13369 42619
rect 13403 42616 13415 42619
rect 13722 42616 13728 42628
rect 13403 42588 13728 42616
rect 13403 42585 13415 42588
rect 13357 42579 13415 42585
rect 13722 42576 13728 42588
rect 13780 42576 13786 42628
rect 11011 42520 12434 42548
rect 11011 42517 11023 42520
rect 10965 42511 11023 42517
rect 13170 42508 13176 42560
rect 13228 42548 13234 42560
rect 13449 42551 13507 42557
rect 13449 42548 13461 42551
rect 13228 42520 13461 42548
rect 13228 42508 13234 42520
rect 13449 42517 13461 42520
rect 13495 42517 13507 42551
rect 13449 42511 13507 42517
rect 16758 42508 16764 42560
rect 16816 42548 16822 42560
rect 17310 42548 17316 42560
rect 16816 42520 17316 42548
rect 16816 42508 16822 42520
rect 17310 42508 17316 42520
rect 17368 42508 17374 42560
rect 17402 42508 17408 42560
rect 17460 42548 17466 42560
rect 17586 42548 17592 42560
rect 17460 42520 17592 42548
rect 17460 42508 17466 42520
rect 17586 42508 17592 42520
rect 17644 42508 17650 42560
rect 1104 42458 18860 42480
rect 1104 42406 2610 42458
rect 2662 42406 2674 42458
rect 2726 42406 2738 42458
rect 2790 42406 2802 42458
rect 2854 42406 2866 42458
rect 2918 42406 7610 42458
rect 7662 42406 7674 42458
rect 7726 42406 7738 42458
rect 7790 42406 7802 42458
rect 7854 42406 7866 42458
rect 7918 42406 12610 42458
rect 12662 42406 12674 42458
rect 12726 42406 12738 42458
rect 12790 42406 12802 42458
rect 12854 42406 12866 42458
rect 12918 42406 17610 42458
rect 17662 42406 17674 42458
rect 17726 42406 17738 42458
rect 17790 42406 17802 42458
rect 17854 42406 17866 42458
rect 17918 42406 18860 42458
rect 1104 42384 18860 42406
rect 3513 42347 3571 42353
rect 3513 42313 3525 42347
rect 3559 42344 3571 42347
rect 3559 42316 8248 42344
rect 3559 42313 3571 42316
rect 3513 42307 3571 42313
rect 1946 42236 1952 42288
rect 2004 42276 2010 42288
rect 2378 42279 2436 42285
rect 2378 42276 2390 42279
rect 2004 42248 2390 42276
rect 2004 42236 2010 42248
rect 2378 42245 2390 42248
rect 2424 42245 2436 42279
rect 2378 42239 2436 42245
rect 7552 42279 7610 42285
rect 7552 42245 7564 42279
rect 7598 42276 7610 42279
rect 8110 42276 8116 42288
rect 7598 42248 8116 42276
rect 7598 42245 7610 42248
rect 7552 42239 7610 42245
rect 8110 42236 8116 42248
rect 8168 42236 8174 42288
rect 2133 42211 2191 42217
rect 2133 42177 2145 42211
rect 2179 42208 2191 42211
rect 2222 42208 2228 42220
rect 2179 42180 2228 42208
rect 2179 42177 2191 42180
rect 2133 42171 2191 42177
rect 2222 42168 2228 42180
rect 2280 42168 2286 42220
rect 7282 42168 7288 42220
rect 7340 42168 7346 42220
rect 8220 42208 8248 42316
rect 8662 42304 8668 42356
rect 8720 42304 8726 42356
rect 9122 42304 9128 42356
rect 9180 42304 9186 42356
rect 13170 42344 13176 42356
rect 9232 42316 13176 42344
rect 8294 42236 8300 42288
rect 8352 42276 8358 42288
rect 9232 42276 9260 42316
rect 13170 42304 13176 42316
rect 13228 42304 13234 42356
rect 8352 42248 9260 42276
rect 8352 42236 8358 42248
rect 9306 42236 9312 42288
rect 9364 42276 9370 42288
rect 9585 42279 9643 42285
rect 9585 42276 9597 42279
rect 9364 42248 9597 42276
rect 9364 42236 9370 42248
rect 9585 42245 9597 42248
rect 9631 42245 9643 42279
rect 9585 42239 9643 42245
rect 10502 42236 10508 42288
rect 10560 42276 10566 42288
rect 17310 42276 17316 42288
rect 10560 42248 17316 42276
rect 10560 42236 10566 42248
rect 17310 42236 17316 42248
rect 17368 42236 17374 42288
rect 9493 42211 9551 42217
rect 8220 42180 9076 42208
rect 9048 42004 9076 42180
rect 9493 42177 9505 42211
rect 9539 42177 9551 42211
rect 9493 42171 9551 42177
rect 9508 42084 9536 42171
rect 9766 42100 9772 42152
rect 9824 42140 9830 42152
rect 13814 42140 13820 42152
rect 9824 42112 13820 42140
rect 9824 42100 9830 42112
rect 13814 42100 13820 42112
rect 13872 42100 13878 42152
rect 18598 42140 18604 42152
rect 17926 42112 18604 42140
rect 9490 42032 9496 42084
rect 9548 42072 9554 42084
rect 17926 42072 17954 42112
rect 18598 42100 18604 42112
rect 18656 42100 18662 42152
rect 9548 42044 17954 42072
rect 9548 42032 9554 42044
rect 11606 42004 11612 42016
rect 9048 41976 11612 42004
rect 11606 41964 11612 41976
rect 11664 41964 11670 42016
rect 1104 41914 18860 41936
rect 1104 41862 1950 41914
rect 2002 41862 2014 41914
rect 2066 41862 2078 41914
rect 2130 41862 2142 41914
rect 2194 41862 2206 41914
rect 2258 41862 6950 41914
rect 7002 41862 7014 41914
rect 7066 41862 7078 41914
rect 7130 41862 7142 41914
rect 7194 41862 7206 41914
rect 7258 41862 11950 41914
rect 12002 41862 12014 41914
rect 12066 41862 12078 41914
rect 12130 41862 12142 41914
rect 12194 41862 12206 41914
rect 12258 41862 16950 41914
rect 17002 41862 17014 41914
rect 17066 41862 17078 41914
rect 17130 41862 17142 41914
rect 17194 41862 17206 41914
rect 17258 41862 18860 41914
rect 1104 41840 18860 41862
rect 7190 41760 7196 41812
rect 7248 41800 7254 41812
rect 7374 41800 7380 41812
rect 7248 41772 7380 41800
rect 7248 41760 7254 41772
rect 7374 41760 7380 41772
rect 7432 41760 7438 41812
rect 8110 41760 8116 41812
rect 8168 41800 8174 41812
rect 8386 41800 8392 41812
rect 8168 41772 8392 41800
rect 8168 41760 8174 41772
rect 8386 41760 8392 41772
rect 8444 41760 8450 41812
rect 6270 41624 6276 41676
rect 6328 41664 6334 41676
rect 6365 41667 6423 41673
rect 6365 41664 6377 41667
rect 6328 41636 6377 41664
rect 6328 41624 6334 41636
rect 6365 41633 6377 41636
rect 6411 41664 6423 41667
rect 10962 41664 10968 41676
rect 6411 41636 10968 41664
rect 6411 41633 6423 41636
rect 6365 41627 6423 41633
rect 10962 41624 10968 41636
rect 11020 41624 11026 41676
rect 658 41556 664 41608
rect 716 41596 722 41608
rect 6454 41596 6460 41608
rect 716 41568 6460 41596
rect 716 41556 722 41568
rect 6454 41556 6460 41568
rect 6512 41556 6518 41608
rect 6730 41556 6736 41608
rect 6788 41596 6794 41608
rect 7466 41596 7472 41608
rect 6788 41568 7472 41596
rect 6788 41556 6794 41568
rect 7466 41556 7472 41568
rect 7524 41596 7530 41608
rect 9306 41596 9312 41608
rect 7524 41568 9312 41596
rect 7524 41556 7530 41568
rect 9306 41556 9312 41568
rect 9364 41556 9370 41608
rect 15194 41528 15200 41540
rect 5736 41500 15200 41528
rect 5736 41469 5764 41500
rect 15194 41488 15200 41500
rect 15252 41488 15258 41540
rect 5721 41463 5779 41469
rect 5721 41429 5733 41463
rect 5767 41429 5779 41463
rect 5721 41423 5779 41429
rect 6086 41420 6092 41472
rect 6144 41420 6150 41472
rect 6178 41420 6184 41472
rect 6236 41420 6242 41472
rect 1104 41370 18860 41392
rect 1104 41318 2610 41370
rect 2662 41318 2674 41370
rect 2726 41318 2738 41370
rect 2790 41318 2802 41370
rect 2854 41318 2866 41370
rect 2918 41318 7610 41370
rect 7662 41318 7674 41370
rect 7726 41318 7738 41370
rect 7790 41318 7802 41370
rect 7854 41318 7866 41370
rect 7918 41318 12610 41370
rect 12662 41318 12674 41370
rect 12726 41318 12738 41370
rect 12790 41318 12802 41370
rect 12854 41318 12866 41370
rect 12918 41318 17610 41370
rect 17662 41318 17674 41370
rect 17726 41318 17738 41370
rect 17790 41318 17802 41370
rect 17854 41318 17866 41370
rect 17918 41318 18860 41370
rect 1104 41296 18860 41318
rect 18049 41123 18107 41129
rect 18049 41089 18061 41123
rect 18095 41120 18107 41123
rect 19794 41120 19800 41132
rect 18095 41092 19800 41120
rect 18095 41089 18107 41092
rect 18049 41083 18107 41089
rect 19794 41080 19800 41092
rect 19852 41080 19858 41132
rect 7190 40876 7196 40928
rect 7248 40916 7254 40928
rect 7650 40916 7656 40928
rect 7248 40888 7656 40916
rect 7248 40876 7254 40888
rect 7650 40876 7656 40888
rect 7708 40876 7714 40928
rect 18230 40876 18236 40928
rect 18288 40876 18294 40928
rect 1104 40826 18860 40848
rect 1104 40774 1950 40826
rect 2002 40774 2014 40826
rect 2066 40774 2078 40826
rect 2130 40774 2142 40826
rect 2194 40774 2206 40826
rect 2258 40774 6950 40826
rect 7002 40774 7014 40826
rect 7066 40774 7078 40826
rect 7130 40774 7142 40826
rect 7194 40774 7206 40826
rect 7258 40774 11950 40826
rect 12002 40774 12014 40826
rect 12066 40774 12078 40826
rect 12130 40774 12142 40826
rect 12194 40774 12206 40826
rect 12258 40774 16950 40826
rect 17002 40774 17014 40826
rect 17066 40774 17078 40826
rect 17130 40774 17142 40826
rect 17194 40774 17206 40826
rect 17258 40774 18860 40826
rect 1104 40752 18860 40774
rect 8662 40468 8668 40520
rect 8720 40508 8726 40520
rect 8938 40508 8944 40520
rect 8720 40480 8944 40508
rect 8720 40468 8726 40480
rect 8938 40468 8944 40480
rect 8996 40468 9002 40520
rect 6638 40332 6644 40384
rect 6696 40372 6702 40384
rect 7650 40372 7656 40384
rect 6696 40344 7656 40372
rect 6696 40332 6702 40344
rect 7650 40332 7656 40344
rect 7708 40372 7714 40384
rect 10962 40372 10968 40384
rect 7708 40344 10968 40372
rect 7708 40332 7714 40344
rect 10962 40332 10968 40344
rect 11020 40332 11026 40384
rect 1104 40282 18860 40304
rect 1104 40230 2610 40282
rect 2662 40230 2674 40282
rect 2726 40230 2738 40282
rect 2790 40230 2802 40282
rect 2854 40230 2866 40282
rect 2918 40230 7610 40282
rect 7662 40230 7674 40282
rect 7726 40230 7738 40282
rect 7790 40230 7802 40282
rect 7854 40230 7866 40282
rect 7918 40230 12610 40282
rect 12662 40230 12674 40282
rect 12726 40230 12738 40282
rect 12790 40230 12802 40282
rect 12854 40230 12866 40282
rect 12918 40230 17610 40282
rect 17662 40230 17674 40282
rect 17726 40230 17738 40282
rect 17790 40230 17802 40282
rect 17854 40230 17866 40282
rect 17918 40230 18860 40282
rect 1104 40208 18860 40230
rect 5074 40128 5080 40180
rect 5132 40168 5138 40180
rect 7837 40171 7895 40177
rect 7837 40168 7849 40171
rect 5132 40140 7849 40168
rect 5132 40128 5138 40140
rect 7837 40137 7849 40140
rect 7883 40137 7895 40171
rect 7837 40131 7895 40137
rect 8478 40128 8484 40180
rect 8536 40168 8542 40180
rect 9306 40168 9312 40180
rect 8536 40140 9312 40168
rect 8536 40128 8542 40140
rect 9306 40128 9312 40140
rect 9364 40128 9370 40180
rect 10962 40128 10968 40180
rect 11020 40128 11026 40180
rect 8205 40103 8263 40109
rect 8205 40069 8217 40103
rect 8251 40100 8263 40103
rect 8846 40100 8852 40112
rect 8251 40072 8852 40100
rect 8251 40069 8263 40072
rect 8205 40063 8263 40069
rect 8846 40060 8852 40072
rect 8904 40060 8910 40112
rect 6822 39992 6828 40044
rect 6880 40032 6886 40044
rect 9841 40035 9899 40041
rect 9841 40032 9853 40035
rect 6880 40004 9853 40032
rect 6880 39992 6886 40004
rect 9841 40001 9853 40004
rect 9887 40001 9899 40035
rect 9841 39995 9899 40001
rect 11330 39992 11336 40044
rect 11388 40032 11394 40044
rect 15749 40035 15807 40041
rect 15749 40032 15761 40035
rect 11388 40004 15761 40032
rect 11388 39992 11394 40004
rect 15749 40001 15761 40004
rect 15795 40001 15807 40035
rect 15749 39995 15807 40001
rect 8297 39967 8355 39973
rect 8297 39933 8309 39967
rect 8343 39964 8355 39967
rect 8386 39964 8392 39976
rect 8343 39936 8392 39964
rect 8343 39933 8355 39936
rect 8297 39927 8355 39933
rect 8386 39924 8392 39936
rect 8444 39924 8450 39976
rect 8478 39924 8484 39976
rect 8536 39924 8542 39976
rect 8754 39924 8760 39976
rect 8812 39964 8818 39976
rect 9585 39967 9643 39973
rect 9585 39964 9597 39967
rect 8812 39936 9597 39964
rect 8812 39924 8818 39936
rect 9585 39933 9597 39936
rect 9631 39933 9643 39967
rect 9585 39927 9643 39933
rect 15473 39967 15531 39973
rect 15473 39933 15485 39967
rect 15519 39964 15531 39967
rect 16758 39964 16764 39976
rect 15519 39936 16764 39964
rect 15519 39933 15531 39936
rect 15473 39927 15531 39933
rect 16758 39924 16764 39936
rect 16816 39924 16822 39976
rect 7282 39856 7288 39908
rect 7340 39896 7346 39908
rect 8772 39896 8800 39924
rect 7340 39868 8800 39896
rect 10520 39868 12434 39896
rect 7340 39856 7346 39868
rect 8478 39788 8484 39840
rect 8536 39828 8542 39840
rect 8662 39828 8668 39840
rect 8536 39800 8668 39828
rect 8536 39788 8542 39800
rect 8662 39788 8668 39800
rect 8720 39828 8726 39840
rect 10520 39828 10548 39868
rect 8720 39800 10548 39828
rect 12406 39828 12434 39868
rect 15010 39828 15016 39840
rect 12406 39800 15016 39828
rect 8720 39788 8726 39800
rect 15010 39788 15016 39800
rect 15068 39788 15074 39840
rect 16758 39788 16764 39840
rect 16816 39828 16822 39840
rect 16942 39828 16948 39840
rect 16816 39800 16948 39828
rect 16816 39788 16822 39800
rect 16942 39788 16948 39800
rect 17000 39788 17006 39840
rect 1104 39738 18860 39760
rect 1104 39686 1950 39738
rect 2002 39686 2014 39738
rect 2066 39686 2078 39738
rect 2130 39686 2142 39738
rect 2194 39686 2206 39738
rect 2258 39686 6950 39738
rect 7002 39686 7014 39738
rect 7066 39686 7078 39738
rect 7130 39686 7142 39738
rect 7194 39686 7206 39738
rect 7258 39686 11950 39738
rect 12002 39686 12014 39738
rect 12066 39686 12078 39738
rect 12130 39686 12142 39738
rect 12194 39686 12206 39738
rect 12258 39686 16950 39738
rect 17002 39686 17014 39738
rect 17066 39686 17078 39738
rect 17130 39686 17142 39738
rect 17194 39686 17206 39738
rect 17258 39686 18860 39738
rect 1104 39664 18860 39686
rect 2498 39584 2504 39636
rect 2556 39624 2562 39636
rect 2556 39596 2774 39624
rect 2556 39584 2562 39596
rect 2746 39420 2774 39596
rect 8386 39584 8392 39636
rect 8444 39624 8450 39636
rect 11790 39624 11796 39636
rect 8444 39596 11796 39624
rect 8444 39584 8450 39596
rect 11790 39584 11796 39596
rect 11848 39624 11854 39636
rect 14182 39624 14188 39636
rect 11848 39596 14188 39624
rect 11848 39584 11854 39596
rect 14182 39584 14188 39596
rect 14240 39584 14246 39636
rect 8938 39516 8944 39568
rect 8996 39556 9002 39568
rect 8996 39528 18092 39556
rect 8996 39516 9002 39528
rect 12526 39448 12532 39500
rect 12584 39488 12590 39500
rect 12989 39491 13047 39497
rect 12989 39488 13001 39491
rect 12584 39460 13001 39488
rect 12584 39448 12590 39460
rect 12989 39457 13001 39460
rect 13035 39488 13047 39491
rect 13446 39488 13452 39500
rect 13035 39460 13452 39488
rect 13035 39457 13047 39460
rect 12989 39451 13047 39457
rect 13446 39448 13452 39460
rect 13504 39448 13510 39500
rect 8478 39420 8484 39432
rect 2746 39392 8484 39420
rect 8478 39380 8484 39392
rect 8536 39420 8542 39432
rect 18064 39429 18092 39528
rect 12713 39423 12771 39429
rect 12713 39420 12725 39423
rect 8536 39392 12725 39420
rect 8536 39380 8542 39392
rect 12713 39389 12725 39392
rect 12759 39389 12771 39423
rect 12713 39383 12771 39389
rect 18049 39423 18107 39429
rect 18049 39389 18061 39423
rect 18095 39389 18107 39423
rect 18049 39383 18107 39389
rect 9122 39312 9128 39364
rect 9180 39352 9186 39364
rect 10502 39352 10508 39364
rect 9180 39324 10508 39352
rect 9180 39312 9186 39324
rect 10502 39312 10508 39324
rect 10560 39352 10566 39364
rect 12805 39355 12863 39361
rect 12805 39352 12817 39355
rect 10560 39324 12817 39352
rect 10560 39312 10566 39324
rect 12805 39321 12817 39324
rect 12851 39321 12863 39355
rect 12805 39315 12863 39321
rect 12342 39244 12348 39296
rect 12400 39244 12406 39296
rect 18230 39244 18236 39296
rect 18288 39244 18294 39296
rect 1104 39194 18860 39216
rect 1104 39142 2610 39194
rect 2662 39142 2674 39194
rect 2726 39142 2738 39194
rect 2790 39142 2802 39194
rect 2854 39142 2866 39194
rect 2918 39142 7610 39194
rect 7662 39142 7674 39194
rect 7726 39142 7738 39194
rect 7790 39142 7802 39194
rect 7854 39142 7866 39194
rect 7918 39142 12610 39194
rect 12662 39142 12674 39194
rect 12726 39142 12738 39194
rect 12790 39142 12802 39194
rect 12854 39142 12866 39194
rect 12918 39142 17610 39194
rect 17662 39142 17674 39194
rect 17726 39142 17738 39194
rect 17790 39142 17802 39194
rect 17854 39142 17866 39194
rect 17918 39142 18860 39194
rect 1104 39120 18860 39142
rect 3964 39015 4022 39021
rect 3964 38981 3976 39015
rect 4010 39012 4022 39015
rect 4890 39012 4896 39024
rect 4010 38984 4896 39012
rect 4010 38981 4022 38984
rect 3964 38975 4022 38981
rect 4890 38972 4896 38984
rect 4948 38972 4954 39024
rect 2314 38904 2320 38956
rect 2372 38944 2378 38956
rect 3697 38947 3755 38953
rect 3697 38944 3709 38947
rect 2372 38916 3709 38944
rect 2372 38904 2378 38916
rect 3697 38913 3709 38916
rect 3743 38913 3755 38947
rect 3697 38907 3755 38913
rect 17037 38947 17095 38953
rect 17037 38913 17049 38947
rect 17083 38944 17095 38947
rect 17310 38944 17316 38956
rect 17083 38916 17316 38944
rect 17083 38913 17095 38916
rect 17037 38907 17095 38913
rect 17310 38904 17316 38916
rect 17368 38904 17374 38956
rect 17681 38947 17739 38953
rect 17681 38913 17693 38947
rect 17727 38913 17739 38947
rect 17681 38907 17739 38913
rect 17696 38876 17724 38907
rect 14476 38848 17724 38876
rect 18233 38879 18291 38885
rect 7282 38808 7288 38820
rect 4632 38780 7288 38808
rect 2958 38700 2964 38752
rect 3016 38740 3022 38752
rect 4632 38740 4660 38780
rect 7282 38768 7288 38780
rect 7340 38768 7346 38820
rect 14476 38752 14504 38848
rect 18233 38845 18245 38879
rect 18279 38876 18291 38879
rect 19610 38876 19616 38888
rect 18279 38848 19616 38876
rect 18279 38845 18291 38848
rect 18233 38839 18291 38845
rect 15010 38768 15016 38820
rect 15068 38808 15074 38820
rect 18248 38808 18276 38839
rect 19610 38836 19616 38848
rect 19668 38836 19674 38888
rect 15068 38780 18276 38808
rect 15068 38768 15074 38780
rect 3016 38712 4660 38740
rect 5077 38743 5135 38749
rect 3016 38700 3022 38712
rect 5077 38709 5089 38743
rect 5123 38740 5135 38743
rect 6822 38740 6828 38752
rect 5123 38712 6828 38740
rect 5123 38709 5135 38712
rect 5077 38703 5135 38709
rect 6822 38700 6828 38712
rect 6880 38700 6886 38752
rect 13998 38700 14004 38752
rect 14056 38740 14062 38752
rect 14458 38740 14464 38752
rect 14056 38712 14464 38740
rect 14056 38700 14062 38712
rect 14458 38700 14464 38712
rect 14516 38700 14522 38752
rect 16853 38743 16911 38749
rect 16853 38709 16865 38743
rect 16899 38740 16911 38743
rect 17310 38740 17316 38752
rect 16899 38712 17316 38740
rect 16899 38709 16911 38712
rect 16853 38703 16911 38709
rect 17310 38700 17316 38712
rect 17368 38700 17374 38752
rect 1104 38650 18860 38672
rect 1104 38598 1950 38650
rect 2002 38598 2014 38650
rect 2066 38598 2078 38650
rect 2130 38598 2142 38650
rect 2194 38598 2206 38650
rect 2258 38598 6950 38650
rect 7002 38598 7014 38650
rect 7066 38598 7078 38650
rect 7130 38598 7142 38650
rect 7194 38598 7206 38650
rect 7258 38598 11950 38650
rect 12002 38598 12014 38650
rect 12066 38598 12078 38650
rect 12130 38598 12142 38650
rect 12194 38598 12206 38650
rect 12258 38598 16950 38650
rect 17002 38598 17014 38650
rect 17066 38598 17078 38650
rect 17130 38598 17142 38650
rect 17194 38598 17206 38650
rect 17258 38598 18860 38650
rect 1104 38576 18860 38598
rect 6638 38496 6644 38548
rect 6696 38536 6702 38548
rect 7282 38536 7288 38548
rect 6696 38508 7288 38536
rect 6696 38496 6702 38508
rect 7282 38496 7288 38508
rect 7340 38496 7346 38548
rect 15194 38292 15200 38344
rect 15252 38332 15258 38344
rect 15473 38335 15531 38341
rect 15473 38332 15485 38335
rect 15252 38304 15485 38332
rect 15252 38292 15258 38304
rect 15473 38301 15485 38304
rect 15519 38301 15531 38335
rect 15473 38295 15531 38301
rect 13538 38224 13544 38276
rect 13596 38264 13602 38276
rect 19886 38264 19892 38276
rect 13596 38236 19892 38264
rect 13596 38224 13602 38236
rect 19886 38224 19892 38236
rect 19944 38224 19950 38276
rect 11330 38156 11336 38208
rect 11388 38196 11394 38208
rect 15289 38199 15347 38205
rect 15289 38196 15301 38199
rect 11388 38168 15301 38196
rect 11388 38156 11394 38168
rect 15289 38165 15301 38168
rect 15335 38165 15347 38199
rect 15289 38159 15347 38165
rect 1104 38106 18860 38128
rect 1104 38054 2610 38106
rect 2662 38054 2674 38106
rect 2726 38054 2738 38106
rect 2790 38054 2802 38106
rect 2854 38054 2866 38106
rect 2918 38054 7610 38106
rect 7662 38054 7674 38106
rect 7726 38054 7738 38106
rect 7790 38054 7802 38106
rect 7854 38054 7866 38106
rect 7918 38054 12610 38106
rect 12662 38054 12674 38106
rect 12726 38054 12738 38106
rect 12790 38054 12802 38106
rect 12854 38054 12866 38106
rect 12918 38054 17610 38106
rect 17662 38054 17674 38106
rect 17726 38054 17738 38106
rect 17790 38054 17802 38106
rect 17854 38054 17866 38106
rect 17918 38054 18860 38106
rect 1104 38032 18860 38054
rect 15930 37952 15936 38004
rect 15988 37992 15994 38004
rect 18322 37992 18328 38004
rect 15988 37964 18328 37992
rect 15988 37952 15994 37964
rect 18322 37952 18328 37964
rect 18380 37952 18386 38004
rect 5534 37884 5540 37936
rect 5592 37924 5598 37936
rect 15378 37924 15384 37936
rect 5592 37896 15384 37924
rect 5592 37884 5598 37896
rect 15378 37884 15384 37896
rect 15436 37884 15442 37936
rect 16025 37859 16083 37865
rect 16025 37825 16037 37859
rect 16071 37856 16083 37859
rect 16482 37856 16488 37868
rect 16071 37828 16488 37856
rect 16071 37825 16083 37828
rect 16025 37819 16083 37825
rect 16482 37816 16488 37828
rect 16540 37816 16546 37868
rect 13538 37748 13544 37800
rect 13596 37788 13602 37800
rect 16117 37791 16175 37797
rect 16117 37788 16129 37791
rect 13596 37760 16129 37788
rect 13596 37748 13602 37760
rect 16117 37757 16129 37760
rect 16163 37757 16175 37791
rect 16117 37751 16175 37757
rect 15194 37612 15200 37664
rect 15252 37652 15258 37664
rect 15565 37655 15623 37661
rect 15565 37652 15577 37655
rect 15252 37624 15577 37652
rect 15252 37612 15258 37624
rect 15565 37621 15577 37624
rect 15611 37621 15623 37655
rect 15565 37615 15623 37621
rect 1104 37562 18860 37584
rect 1104 37510 1950 37562
rect 2002 37510 2014 37562
rect 2066 37510 2078 37562
rect 2130 37510 2142 37562
rect 2194 37510 2206 37562
rect 2258 37510 6950 37562
rect 7002 37510 7014 37562
rect 7066 37510 7078 37562
rect 7130 37510 7142 37562
rect 7194 37510 7206 37562
rect 7258 37510 11950 37562
rect 12002 37510 12014 37562
rect 12066 37510 12078 37562
rect 12130 37510 12142 37562
rect 12194 37510 12206 37562
rect 12258 37510 16950 37562
rect 17002 37510 17014 37562
rect 17066 37510 17078 37562
rect 17130 37510 17142 37562
rect 17194 37510 17206 37562
rect 17258 37510 18860 37562
rect 1104 37488 18860 37510
rect 9582 37408 9588 37460
rect 9640 37448 9646 37460
rect 9766 37448 9772 37460
rect 9640 37420 9772 37448
rect 9640 37408 9646 37420
rect 9766 37408 9772 37420
rect 9824 37408 9830 37460
rect 12618 37408 12624 37460
rect 12676 37408 12682 37460
rect 12434 37340 12440 37392
rect 12492 37380 12498 37392
rect 15010 37380 15016 37392
rect 12492 37352 15016 37380
rect 12492 37340 12498 37352
rect 15010 37340 15016 37352
rect 15068 37340 15074 37392
rect 13265 37315 13323 37321
rect 13265 37281 13277 37315
rect 13311 37312 13323 37315
rect 13538 37312 13544 37324
rect 13311 37284 13544 37312
rect 13311 37281 13323 37284
rect 13265 37275 13323 37281
rect 13538 37272 13544 37284
rect 13596 37272 13602 37324
rect 14826 37272 14832 37324
rect 14884 37312 14890 37324
rect 15746 37312 15752 37324
rect 14884 37284 15752 37312
rect 14884 37272 14890 37284
rect 15746 37272 15752 37284
rect 15804 37272 15810 37324
rect 1949 37247 2007 37253
rect 1949 37213 1961 37247
rect 1995 37244 2007 37247
rect 2958 37244 2964 37256
rect 1995 37216 2964 37244
rect 1995 37213 2007 37216
rect 1949 37207 2007 37213
rect 2958 37204 2964 37216
rect 3016 37204 3022 37256
rect 12989 37247 13047 37253
rect 12989 37213 13001 37247
rect 13035 37244 13047 37247
rect 13078 37244 13084 37256
rect 13035 37216 13084 37244
rect 13035 37213 13047 37216
rect 12989 37207 13047 37213
rect 13078 37204 13084 37216
rect 13136 37204 13142 37256
rect 18046 37204 18052 37256
rect 18104 37204 18110 37256
rect 1854 37136 1860 37188
rect 1912 37176 1918 37188
rect 2194 37179 2252 37185
rect 2194 37176 2206 37179
rect 1912 37148 2206 37176
rect 1912 37136 1918 37148
rect 2194 37145 2206 37148
rect 2240 37145 2252 37179
rect 2194 37139 2252 37145
rect 12618 37136 12624 37188
rect 12676 37176 12682 37188
rect 13446 37176 13452 37188
rect 12676 37148 13452 37176
rect 12676 37136 12682 37148
rect 13446 37136 13452 37148
rect 13504 37136 13510 37188
rect 3329 37111 3387 37117
rect 3329 37077 3341 37111
rect 3375 37108 3387 37111
rect 8386 37108 8392 37120
rect 3375 37080 8392 37108
rect 3375 37077 3387 37080
rect 3329 37071 3387 37077
rect 8386 37068 8392 37080
rect 8444 37068 8450 37120
rect 9030 37068 9036 37120
rect 9088 37108 9094 37120
rect 13081 37111 13139 37117
rect 13081 37108 13093 37111
rect 9088 37080 13093 37108
rect 9088 37068 9094 37080
rect 13081 37077 13093 37080
rect 13127 37108 13139 37111
rect 13170 37108 13176 37120
rect 13127 37080 13176 37108
rect 13127 37077 13139 37080
rect 13081 37071 13139 37077
rect 13170 37068 13176 37080
rect 13228 37068 13234 37120
rect 18230 37068 18236 37120
rect 18288 37068 18294 37120
rect 1104 37018 18860 37040
rect 1104 36966 2610 37018
rect 2662 36966 2674 37018
rect 2726 36966 2738 37018
rect 2790 36966 2802 37018
rect 2854 36966 2866 37018
rect 2918 36966 7610 37018
rect 7662 36966 7674 37018
rect 7726 36966 7738 37018
rect 7790 36966 7802 37018
rect 7854 36966 7866 37018
rect 7918 36966 12610 37018
rect 12662 36966 12674 37018
rect 12726 36966 12738 37018
rect 12790 36966 12802 37018
rect 12854 36966 12866 37018
rect 12918 36966 17610 37018
rect 17662 36966 17674 37018
rect 17726 36966 17738 37018
rect 17790 36966 17802 37018
rect 17854 36966 17866 37018
rect 17918 36966 18860 37018
rect 1104 36944 18860 36966
rect 4062 36864 4068 36916
rect 4120 36904 4126 36916
rect 8113 36907 8171 36913
rect 8113 36904 8125 36907
rect 4120 36876 8125 36904
rect 4120 36864 4126 36876
rect 8113 36873 8125 36876
rect 8159 36873 8171 36907
rect 8113 36867 8171 36873
rect 8386 36864 8392 36916
rect 8444 36904 8450 36916
rect 8573 36907 8631 36913
rect 8573 36904 8585 36907
rect 8444 36876 8585 36904
rect 8444 36864 8450 36876
rect 8573 36873 8585 36876
rect 8619 36904 8631 36907
rect 10686 36904 10692 36916
rect 8619 36876 10692 36904
rect 8619 36873 8631 36876
rect 8573 36867 8631 36873
rect 10686 36864 10692 36876
rect 10744 36864 10750 36916
rect 11606 36864 11612 36916
rect 11664 36904 11670 36916
rect 11664 36876 12848 36904
rect 11664 36864 11670 36876
rect 8481 36771 8539 36777
rect 8481 36737 8493 36771
rect 8527 36768 8539 36771
rect 9122 36768 9128 36780
rect 8527 36740 9128 36768
rect 8527 36737 8539 36740
rect 8481 36731 8539 36737
rect 9122 36728 9128 36740
rect 9180 36728 9186 36780
rect 12820 36768 12848 36876
rect 12986 36864 12992 36916
rect 13044 36904 13050 36916
rect 13354 36904 13360 36916
rect 13044 36876 13360 36904
rect 13044 36864 13050 36876
rect 13354 36864 13360 36876
rect 13412 36864 13418 36916
rect 17494 36864 17500 36916
rect 17552 36864 17558 36916
rect 15930 36768 15936 36780
rect 12820 36740 15936 36768
rect 15930 36728 15936 36740
rect 15988 36728 15994 36780
rect 17512 36768 17540 36864
rect 17420 36740 17540 36768
rect 17420 36712 17448 36740
rect 8662 36660 8668 36712
rect 8720 36660 8726 36712
rect 9766 36660 9772 36712
rect 9824 36700 9830 36712
rect 10410 36700 10416 36712
rect 9824 36672 10416 36700
rect 9824 36660 9830 36672
rect 10410 36660 10416 36672
rect 10468 36700 10474 36712
rect 13262 36700 13268 36712
rect 10468 36672 13268 36700
rect 10468 36660 10474 36672
rect 13262 36660 13268 36672
rect 13320 36660 13326 36712
rect 17402 36660 17408 36712
rect 17460 36660 17466 36712
rect 6638 36592 6644 36644
rect 6696 36632 6702 36644
rect 13998 36632 14004 36644
rect 6696 36604 14004 36632
rect 6696 36592 6702 36604
rect 13998 36592 14004 36604
rect 14056 36592 14062 36644
rect 15102 36524 15108 36576
rect 15160 36564 15166 36576
rect 15654 36564 15660 36576
rect 15160 36536 15660 36564
rect 15160 36524 15166 36536
rect 15654 36524 15660 36536
rect 15712 36524 15718 36576
rect 18322 36524 18328 36576
rect 18380 36564 18386 36576
rect 19426 36564 19432 36576
rect 18380 36536 19432 36564
rect 18380 36524 18386 36536
rect 19426 36524 19432 36536
rect 19484 36524 19490 36576
rect 1104 36474 18860 36496
rect 1104 36422 1950 36474
rect 2002 36422 2014 36474
rect 2066 36422 2078 36474
rect 2130 36422 2142 36474
rect 2194 36422 2206 36474
rect 2258 36422 6950 36474
rect 7002 36422 7014 36474
rect 7066 36422 7078 36474
rect 7130 36422 7142 36474
rect 7194 36422 7206 36474
rect 7258 36422 11950 36474
rect 12002 36422 12014 36474
rect 12066 36422 12078 36474
rect 12130 36422 12142 36474
rect 12194 36422 12206 36474
rect 12258 36422 16950 36474
rect 17002 36422 17014 36474
rect 17066 36422 17078 36474
rect 17130 36422 17142 36474
rect 17194 36422 17206 36474
rect 17258 36422 18860 36474
rect 1104 36400 18860 36422
rect 2225 36363 2283 36369
rect 2225 36329 2237 36363
rect 2271 36360 2283 36363
rect 6638 36360 6644 36372
rect 2271 36332 6644 36360
rect 2271 36329 2283 36332
rect 2225 36323 2283 36329
rect 6638 36320 6644 36332
rect 6696 36320 6702 36372
rect 10226 36320 10232 36372
rect 10284 36360 10290 36372
rect 10594 36360 10600 36372
rect 10284 36332 10600 36360
rect 10284 36320 10290 36332
rect 10594 36320 10600 36332
rect 10652 36360 10658 36372
rect 10652 36332 12388 36360
rect 10652 36320 10658 36332
rect 4522 36252 4528 36304
rect 4580 36292 4586 36304
rect 11425 36295 11483 36301
rect 11425 36292 11437 36295
rect 4580 36264 11437 36292
rect 4580 36252 4586 36264
rect 11425 36261 11437 36264
rect 11471 36292 11483 36295
rect 11471 36264 12204 36292
rect 11471 36261 11483 36264
rect 11425 36255 11483 36261
rect 2869 36227 2927 36233
rect 2869 36193 2881 36227
rect 2915 36224 2927 36227
rect 9766 36224 9772 36236
rect 2915 36196 9772 36224
rect 2915 36193 2927 36196
rect 2869 36187 2927 36193
rect 9766 36184 9772 36196
rect 9824 36184 9830 36236
rect 2685 36159 2743 36165
rect 2685 36125 2697 36159
rect 2731 36156 2743 36159
rect 9858 36156 9864 36168
rect 2731 36128 9864 36156
rect 2731 36125 2743 36128
rect 2685 36119 2743 36125
rect 9858 36116 9864 36128
rect 9916 36116 9922 36168
rect 12176 36165 12204 36264
rect 12360 36233 12388 36332
rect 12345 36227 12403 36233
rect 12345 36193 12357 36227
rect 12391 36193 12403 36227
rect 12345 36187 12403 36193
rect 12161 36159 12219 36165
rect 12161 36125 12173 36159
rect 12207 36156 12219 36159
rect 12207 36128 12434 36156
rect 12207 36125 12219 36128
rect 12161 36119 12219 36125
rect 2593 36091 2651 36097
rect 2593 36057 2605 36091
rect 2639 36088 2651 36091
rect 2639 36060 2774 36088
rect 2639 36057 2651 36060
rect 2593 36051 2651 36057
rect 2746 36020 2774 36060
rect 9306 36048 9312 36100
rect 9364 36088 9370 36100
rect 12253 36091 12311 36097
rect 12253 36088 12265 36091
rect 9364 36060 12265 36088
rect 9364 36048 9370 36060
rect 12253 36057 12265 36060
rect 12299 36057 12311 36091
rect 12406 36088 12434 36128
rect 18046 36088 18052 36100
rect 12406 36060 18052 36088
rect 12253 36051 12311 36057
rect 18046 36048 18052 36060
rect 18104 36048 18110 36100
rect 10042 36020 10048 36032
rect 2746 35992 10048 36020
rect 10042 35980 10048 35992
rect 10100 35980 10106 36032
rect 11514 35980 11520 36032
rect 11572 36020 11578 36032
rect 11793 36023 11851 36029
rect 11793 36020 11805 36023
rect 11572 35992 11805 36020
rect 11572 35980 11578 35992
rect 11793 35989 11805 35992
rect 11839 35989 11851 36023
rect 11793 35983 11851 35989
rect 1104 35930 18860 35952
rect 1104 35878 2610 35930
rect 2662 35878 2674 35930
rect 2726 35878 2738 35930
rect 2790 35878 2802 35930
rect 2854 35878 2866 35930
rect 2918 35878 7610 35930
rect 7662 35878 7674 35930
rect 7726 35878 7738 35930
rect 7790 35878 7802 35930
rect 7854 35878 7866 35930
rect 7918 35878 12610 35930
rect 12662 35878 12674 35930
rect 12726 35878 12738 35930
rect 12790 35878 12802 35930
rect 12854 35878 12866 35930
rect 12918 35878 17610 35930
rect 17662 35878 17674 35930
rect 17726 35878 17738 35930
rect 17790 35878 17802 35930
rect 17854 35878 17866 35930
rect 17918 35878 18860 35930
rect 1104 35856 18860 35878
rect 3694 35776 3700 35828
rect 3752 35816 3758 35828
rect 4982 35816 4988 35828
rect 3752 35788 4988 35816
rect 3752 35776 3758 35788
rect 4982 35776 4988 35788
rect 5040 35776 5046 35828
rect 6822 35776 6828 35828
rect 6880 35816 6886 35828
rect 9766 35816 9772 35828
rect 6880 35788 9772 35816
rect 6880 35776 6886 35788
rect 9766 35776 9772 35788
rect 9824 35816 9830 35828
rect 11882 35816 11888 35828
rect 9824 35788 11888 35816
rect 9824 35776 9830 35788
rect 11882 35776 11888 35788
rect 11940 35776 11946 35828
rect 11422 35708 11428 35760
rect 11480 35748 11486 35760
rect 13326 35751 13384 35757
rect 13326 35748 13338 35751
rect 11480 35720 13338 35748
rect 11480 35708 11486 35720
rect 13326 35717 13338 35720
rect 13372 35717 13384 35751
rect 13326 35711 13384 35717
rect 8018 35640 8024 35692
rect 8076 35680 8082 35692
rect 12345 35683 12403 35689
rect 12345 35680 12357 35683
rect 8076 35652 12357 35680
rect 8076 35640 8082 35652
rect 12345 35649 12357 35652
rect 12391 35649 12403 35683
rect 18049 35683 18107 35689
rect 18049 35680 18061 35683
rect 12345 35643 12403 35649
rect 13004 35652 18061 35680
rect 11422 35572 11428 35624
rect 11480 35612 11486 35624
rect 11790 35612 11796 35624
rect 11480 35584 11796 35612
rect 11480 35572 11486 35584
rect 11790 35572 11796 35584
rect 11848 35572 11854 35624
rect 11882 35572 11888 35624
rect 11940 35612 11946 35624
rect 13004 35612 13032 35652
rect 18049 35649 18061 35652
rect 18095 35649 18107 35683
rect 18049 35643 18107 35649
rect 11940 35584 13032 35612
rect 13081 35615 13139 35621
rect 11940 35572 11946 35584
rect 13081 35581 13093 35615
rect 13127 35581 13139 35615
rect 13081 35575 13139 35581
rect 5718 35504 5724 35556
rect 5776 35544 5782 35556
rect 12986 35544 12992 35556
rect 5776 35516 12992 35544
rect 5776 35504 5782 35516
rect 12986 35504 12992 35516
rect 13044 35504 13050 35556
rect 12434 35436 12440 35488
rect 12492 35436 12498 35488
rect 13096 35476 13124 35575
rect 14090 35504 14096 35556
rect 14148 35544 14154 35556
rect 14461 35547 14519 35553
rect 14461 35544 14473 35547
rect 14148 35516 14473 35544
rect 14148 35504 14154 35516
rect 14461 35513 14473 35516
rect 14507 35544 14519 35547
rect 19702 35544 19708 35556
rect 14507 35516 19708 35544
rect 14507 35513 14519 35516
rect 14461 35507 14519 35513
rect 19702 35504 19708 35516
rect 19760 35504 19766 35556
rect 13814 35476 13820 35488
rect 13096 35448 13820 35476
rect 13814 35436 13820 35448
rect 13872 35436 13878 35488
rect 18230 35436 18236 35488
rect 18288 35436 18294 35488
rect 1104 35386 18860 35408
rect 1104 35334 1950 35386
rect 2002 35334 2014 35386
rect 2066 35334 2078 35386
rect 2130 35334 2142 35386
rect 2194 35334 2206 35386
rect 2258 35334 6950 35386
rect 7002 35334 7014 35386
rect 7066 35334 7078 35386
rect 7130 35334 7142 35386
rect 7194 35334 7206 35386
rect 7258 35334 11950 35386
rect 12002 35334 12014 35386
rect 12066 35334 12078 35386
rect 12130 35334 12142 35386
rect 12194 35334 12206 35386
rect 12258 35334 16950 35386
rect 17002 35334 17014 35386
rect 17066 35334 17078 35386
rect 17130 35334 17142 35386
rect 17194 35334 17206 35386
rect 17258 35334 18860 35386
rect 1104 35312 18860 35334
rect 10505 35275 10563 35281
rect 10505 35241 10517 35275
rect 10551 35272 10563 35275
rect 13722 35272 13728 35284
rect 10551 35244 13728 35272
rect 10551 35241 10563 35244
rect 10505 35235 10563 35241
rect 13722 35232 13728 35244
rect 13780 35232 13786 35284
rect 12989 35207 13047 35213
rect 12989 35173 13001 35207
rect 13035 35204 13047 35207
rect 18690 35204 18696 35216
rect 13035 35176 18696 35204
rect 13035 35173 13047 35176
rect 12989 35167 13047 35173
rect 18690 35164 18696 35176
rect 18748 35164 18754 35216
rect 8297 35139 8355 35145
rect 8297 35105 8309 35139
rect 8343 35136 8355 35139
rect 8386 35136 8392 35148
rect 8343 35108 8392 35136
rect 8343 35105 8355 35108
rect 8297 35099 8355 35105
rect 8386 35096 8392 35108
rect 8444 35096 8450 35148
rect 8481 35139 8539 35145
rect 8481 35105 8493 35139
rect 8527 35136 8539 35139
rect 8527 35108 9260 35136
rect 8527 35105 8539 35108
rect 8481 35099 8539 35105
rect 8202 35028 8208 35080
rect 8260 35028 8266 35080
rect 8754 35028 8760 35080
rect 8812 35068 8818 35080
rect 9125 35071 9183 35077
rect 9125 35068 9137 35071
rect 8812 35040 9137 35068
rect 8812 35028 8818 35040
rect 9125 35037 9137 35040
rect 9171 35037 9183 35071
rect 9232 35068 9260 35108
rect 13538 35096 13544 35148
rect 13596 35136 13602 35148
rect 13633 35139 13691 35145
rect 13633 35136 13645 35139
rect 13596 35108 13645 35136
rect 13596 35096 13602 35108
rect 13633 35105 13645 35108
rect 13679 35136 13691 35139
rect 13722 35136 13728 35148
rect 13679 35108 13728 35136
rect 13679 35105 13691 35108
rect 13633 35099 13691 35105
rect 13722 35096 13728 35108
rect 13780 35096 13786 35148
rect 12526 35068 12532 35080
rect 9232 35040 12532 35068
rect 9125 35031 9183 35037
rect 12526 35028 12532 35040
rect 12584 35068 12590 35080
rect 12986 35068 12992 35080
rect 12584 35040 12992 35068
rect 12584 35028 12590 35040
rect 12986 35028 12992 35040
rect 13044 35028 13050 35080
rect 13357 35071 13415 35077
rect 13357 35037 13369 35071
rect 13403 35068 13415 35071
rect 15838 35068 15844 35080
rect 13403 35040 15844 35068
rect 13403 35037 13415 35040
rect 13357 35031 13415 35037
rect 15838 35028 15844 35040
rect 15896 35028 15902 35080
rect 4798 34960 4804 35012
rect 4856 35000 4862 35012
rect 9370 35003 9428 35009
rect 9370 35000 9382 35003
rect 4856 34972 9382 35000
rect 4856 34960 4862 34972
rect 9370 34969 9382 34972
rect 9416 34969 9428 35003
rect 9370 34963 9428 34969
rect 10318 34960 10324 35012
rect 10376 35000 10382 35012
rect 12434 35000 12440 35012
rect 10376 34972 12440 35000
rect 10376 34960 10382 34972
rect 12434 34960 12440 34972
rect 12492 34960 12498 35012
rect 13078 34960 13084 35012
rect 13136 35000 13142 35012
rect 13449 35003 13507 35009
rect 13449 35000 13461 35003
rect 13136 34972 13461 35000
rect 13136 34960 13142 34972
rect 13449 34969 13461 34972
rect 13495 34969 13507 35003
rect 13449 34963 13507 34969
rect 7837 34935 7895 34941
rect 7837 34901 7849 34935
rect 7883 34932 7895 34935
rect 8202 34932 8208 34944
rect 7883 34904 8208 34932
rect 7883 34901 7895 34904
rect 7837 34895 7895 34901
rect 8202 34892 8208 34904
rect 8260 34892 8266 34944
rect 9674 34892 9680 34944
rect 9732 34932 9738 34944
rect 13262 34932 13268 34944
rect 9732 34904 13268 34932
rect 9732 34892 9738 34904
rect 13262 34892 13268 34904
rect 13320 34892 13326 34944
rect 13538 34892 13544 34944
rect 13596 34932 13602 34944
rect 15010 34932 15016 34944
rect 13596 34904 15016 34932
rect 13596 34892 13602 34904
rect 15010 34892 15016 34904
rect 15068 34892 15074 34944
rect 1104 34842 18860 34864
rect 1104 34790 2610 34842
rect 2662 34790 2674 34842
rect 2726 34790 2738 34842
rect 2790 34790 2802 34842
rect 2854 34790 2866 34842
rect 2918 34790 7610 34842
rect 7662 34790 7674 34842
rect 7726 34790 7738 34842
rect 7790 34790 7802 34842
rect 7854 34790 7866 34842
rect 7918 34790 12610 34842
rect 12662 34790 12674 34842
rect 12726 34790 12738 34842
rect 12790 34790 12802 34842
rect 12854 34790 12866 34842
rect 12918 34790 17610 34842
rect 17662 34790 17674 34842
rect 17726 34790 17738 34842
rect 17790 34790 17802 34842
rect 17854 34790 17866 34842
rect 17918 34790 18860 34842
rect 1104 34768 18860 34790
rect 5350 34728 5356 34740
rect 3068 34700 5356 34728
rect 2406 34620 2412 34672
rect 2464 34660 2470 34672
rect 3068 34669 3096 34700
rect 5350 34688 5356 34700
rect 5408 34728 5414 34740
rect 5408 34700 9168 34728
rect 5408 34688 5414 34700
rect 3053 34663 3111 34669
rect 3053 34660 3065 34663
rect 2464 34632 3065 34660
rect 2464 34620 2470 34632
rect 3053 34629 3065 34632
rect 3099 34629 3111 34663
rect 3053 34623 3111 34629
rect 3234 34620 3240 34672
rect 3292 34620 3298 34672
rect 2759 34595 2817 34601
rect 2759 34561 2771 34595
rect 2805 34592 2817 34595
rect 4890 34592 4896 34604
rect 2805 34564 4896 34592
rect 2805 34561 2817 34564
rect 2759 34555 2817 34561
rect 4890 34552 4896 34564
rect 4948 34552 4954 34604
rect 8018 34552 8024 34604
rect 8076 34592 8082 34604
rect 9013 34595 9071 34601
rect 9013 34592 9025 34595
rect 8076 34564 9025 34592
rect 8076 34552 8082 34564
rect 9013 34561 9025 34564
rect 9059 34561 9071 34595
rect 9140 34592 9168 34700
rect 10134 34688 10140 34740
rect 10192 34688 10198 34740
rect 12253 34731 12311 34737
rect 12253 34697 12265 34731
rect 12299 34697 12311 34731
rect 14737 34731 14795 34737
rect 12253 34691 12311 34697
rect 12406 34700 14136 34728
rect 9490 34620 9496 34672
rect 9548 34660 9554 34672
rect 12268 34660 12296 34691
rect 9548 34632 12296 34660
rect 9548 34620 9554 34632
rect 12406 34592 12434 34700
rect 13814 34660 13820 34672
rect 13372 34632 13820 34660
rect 9140 34564 12434 34592
rect 12621 34595 12679 34601
rect 9013 34555 9071 34561
rect 12621 34561 12633 34595
rect 12667 34592 12679 34595
rect 13170 34592 13176 34604
rect 12667 34564 13176 34592
rect 12667 34561 12679 34564
rect 12621 34555 12679 34561
rect 13170 34552 13176 34564
rect 13228 34552 13234 34604
rect 13262 34552 13268 34604
rect 13320 34552 13326 34604
rect 13372 34601 13400 34632
rect 13814 34620 13820 34632
rect 13872 34620 13878 34672
rect 14108 34660 14136 34700
rect 14737 34697 14749 34731
rect 14783 34728 14795 34731
rect 15102 34728 15108 34740
rect 14783 34700 15108 34728
rect 14783 34697 14795 34700
rect 14737 34691 14795 34697
rect 15102 34688 15108 34700
rect 15160 34688 15166 34740
rect 15378 34688 15384 34740
rect 15436 34688 15442 34740
rect 15841 34663 15899 34669
rect 15841 34660 15853 34663
rect 14108 34632 15853 34660
rect 15841 34629 15853 34632
rect 15887 34629 15899 34663
rect 15841 34623 15899 34629
rect 13357 34595 13415 34601
rect 13357 34561 13369 34595
rect 13403 34561 13415 34595
rect 13613 34595 13671 34601
rect 13613 34592 13625 34595
rect 13357 34555 13415 34561
rect 13464 34564 13625 34592
rect 3329 34527 3387 34533
rect 3329 34493 3341 34527
rect 3375 34524 3387 34527
rect 7282 34524 7288 34536
rect 3375 34496 7288 34524
rect 3375 34493 3387 34496
rect 3329 34487 3387 34493
rect 7282 34484 7288 34496
rect 7340 34484 7346 34536
rect 8754 34484 8760 34536
rect 8812 34484 8818 34536
rect 12434 34484 12440 34536
rect 12492 34524 12498 34536
rect 12713 34527 12771 34533
rect 12713 34524 12725 34527
rect 12492 34496 12725 34524
rect 12492 34484 12498 34496
rect 12713 34493 12725 34496
rect 12759 34493 12771 34527
rect 12713 34487 12771 34493
rect 12805 34527 12863 34533
rect 12805 34493 12817 34527
rect 12851 34493 12863 34527
rect 13280 34524 13308 34552
rect 13464 34524 13492 34564
rect 13613 34561 13625 34564
rect 13659 34561 13671 34595
rect 13613 34555 13671 34561
rect 15010 34552 15016 34604
rect 15068 34592 15074 34604
rect 15749 34595 15807 34601
rect 15749 34592 15761 34595
rect 15068 34564 15761 34592
rect 15068 34552 15074 34564
rect 15749 34561 15761 34564
rect 15795 34561 15807 34595
rect 15749 34555 15807 34561
rect 13280 34496 13492 34524
rect 16025 34527 16083 34533
rect 12805 34487 12863 34493
rect 16025 34493 16037 34527
rect 16071 34493 16083 34527
rect 16025 34487 16083 34493
rect 12820 34456 12848 34487
rect 12986 34456 12992 34468
rect 12820 34428 12992 34456
rect 12986 34416 12992 34428
rect 13044 34456 13050 34468
rect 13262 34456 13268 34468
rect 13044 34428 13268 34456
rect 13044 34416 13050 34428
rect 13262 34416 13268 34428
rect 13320 34416 13326 34468
rect 16040 34456 16068 34487
rect 17402 34456 17408 34468
rect 16040 34428 17408 34456
rect 7282 34348 7288 34400
rect 7340 34388 7346 34400
rect 16040 34388 16068 34428
rect 17402 34416 17408 34428
rect 17460 34416 17466 34468
rect 7340 34360 16068 34388
rect 7340 34348 7346 34360
rect 1104 34298 18860 34320
rect 1104 34246 1950 34298
rect 2002 34246 2014 34298
rect 2066 34246 2078 34298
rect 2130 34246 2142 34298
rect 2194 34246 2206 34298
rect 2258 34246 6950 34298
rect 7002 34246 7014 34298
rect 7066 34246 7078 34298
rect 7130 34246 7142 34298
rect 7194 34246 7206 34298
rect 7258 34246 11950 34298
rect 12002 34246 12014 34298
rect 12066 34246 12078 34298
rect 12130 34246 12142 34298
rect 12194 34246 12206 34298
rect 12258 34246 16950 34298
rect 17002 34246 17014 34298
rect 17066 34246 17078 34298
rect 17130 34246 17142 34298
rect 17194 34246 17206 34298
rect 17258 34246 18860 34298
rect 1104 34224 18860 34246
rect 16758 34076 16764 34128
rect 16816 34116 16822 34128
rect 16853 34119 16911 34125
rect 16853 34116 16865 34119
rect 16816 34088 16865 34116
rect 16816 34076 16822 34088
rect 16853 34085 16865 34088
rect 16899 34085 16911 34119
rect 16853 34079 16911 34085
rect 17402 34008 17408 34060
rect 17460 34008 17466 34060
rect 16298 33940 16304 33992
rect 16356 33940 16362 33992
rect 7006 33872 7012 33924
rect 7064 33912 7070 33924
rect 17129 33915 17187 33921
rect 17129 33912 17141 33915
rect 7064 33884 17141 33912
rect 7064 33872 7070 33884
rect 17129 33881 17141 33884
rect 17175 33881 17187 33915
rect 17129 33875 17187 33881
rect 16114 33804 16120 33856
rect 16172 33804 16178 33856
rect 16482 33804 16488 33856
rect 16540 33844 16546 33856
rect 17313 33847 17371 33853
rect 17313 33844 17325 33847
rect 16540 33816 17325 33844
rect 16540 33804 16546 33816
rect 17313 33813 17325 33816
rect 17359 33813 17371 33847
rect 17313 33807 17371 33813
rect 1104 33754 18860 33776
rect 1104 33702 2610 33754
rect 2662 33702 2674 33754
rect 2726 33702 2738 33754
rect 2790 33702 2802 33754
rect 2854 33702 2866 33754
rect 2918 33702 7610 33754
rect 7662 33702 7674 33754
rect 7726 33702 7738 33754
rect 7790 33702 7802 33754
rect 7854 33702 7866 33754
rect 7918 33702 12610 33754
rect 12662 33702 12674 33754
rect 12726 33702 12738 33754
rect 12790 33702 12802 33754
rect 12854 33702 12866 33754
rect 12918 33702 17610 33754
rect 17662 33702 17674 33754
rect 17726 33702 17738 33754
rect 17790 33702 17802 33754
rect 17854 33702 17866 33754
rect 17918 33702 18860 33754
rect 1104 33680 18860 33702
rect 15562 33600 15568 33652
rect 15620 33600 15626 33652
rect 15746 33600 15752 33652
rect 15804 33640 15810 33652
rect 16482 33640 16488 33652
rect 15804 33612 16488 33640
rect 15804 33600 15810 33612
rect 16482 33600 16488 33612
rect 16540 33600 16546 33652
rect 13998 33464 14004 33516
rect 14056 33504 14062 33516
rect 15749 33507 15807 33513
rect 15749 33504 15761 33507
rect 14056 33476 15761 33504
rect 14056 33464 14062 33476
rect 15749 33473 15761 33476
rect 15795 33473 15807 33507
rect 15749 33467 15807 33473
rect 18049 33507 18107 33513
rect 18049 33473 18061 33507
rect 18095 33473 18107 33507
rect 18049 33467 18107 33473
rect 9030 33396 9036 33448
rect 9088 33436 9094 33448
rect 18064 33436 18092 33467
rect 9088 33408 18092 33436
rect 9088 33396 9094 33408
rect 3234 33260 3240 33312
rect 3292 33300 3298 33312
rect 6638 33300 6644 33312
rect 3292 33272 6644 33300
rect 3292 33260 3298 33272
rect 6638 33260 6644 33272
rect 6696 33300 6702 33312
rect 7006 33300 7012 33312
rect 6696 33272 7012 33300
rect 6696 33260 6702 33272
rect 7006 33260 7012 33272
rect 7064 33260 7070 33312
rect 18230 33260 18236 33312
rect 18288 33260 18294 33312
rect 1104 33210 18860 33232
rect 1104 33158 1950 33210
rect 2002 33158 2014 33210
rect 2066 33158 2078 33210
rect 2130 33158 2142 33210
rect 2194 33158 2206 33210
rect 2258 33158 6950 33210
rect 7002 33158 7014 33210
rect 7066 33158 7078 33210
rect 7130 33158 7142 33210
rect 7194 33158 7206 33210
rect 7258 33158 11950 33210
rect 12002 33158 12014 33210
rect 12066 33158 12078 33210
rect 12130 33158 12142 33210
rect 12194 33158 12206 33210
rect 12258 33158 16950 33210
rect 17002 33158 17014 33210
rect 17066 33158 17078 33210
rect 17130 33158 17142 33210
rect 17194 33158 17206 33210
rect 17258 33158 18860 33210
rect 1104 33136 18860 33158
rect 4614 33056 4620 33108
rect 4672 33096 4678 33108
rect 6730 33096 6736 33108
rect 4672 33068 6736 33096
rect 4672 33056 4678 33068
rect 6730 33056 6736 33068
rect 6788 33056 6794 33108
rect 16482 33056 16488 33108
rect 16540 33096 16546 33108
rect 16945 33099 17003 33105
rect 16945 33096 16957 33099
rect 16540 33068 16957 33096
rect 16540 33056 16546 33068
rect 16945 33065 16957 33068
rect 16991 33096 17003 33099
rect 19518 33096 19524 33108
rect 16991 33068 19524 33096
rect 16991 33065 17003 33068
rect 16945 33059 17003 33065
rect 19518 33056 19524 33068
rect 19576 33056 19582 33108
rect 13814 32920 13820 32972
rect 13872 32960 13878 32972
rect 15565 32963 15623 32969
rect 15565 32960 15577 32963
rect 13872 32932 15577 32960
rect 13872 32920 13878 32932
rect 15565 32929 15577 32932
rect 15611 32929 15623 32963
rect 15565 32923 15623 32929
rect 15580 32892 15608 32923
rect 16850 32892 16856 32904
rect 15580 32864 16856 32892
rect 16850 32852 16856 32864
rect 16908 32852 16914 32904
rect 15832 32827 15890 32833
rect 15832 32793 15844 32827
rect 15878 32824 15890 32827
rect 16114 32824 16120 32836
rect 15878 32796 16120 32824
rect 15878 32793 15890 32796
rect 15832 32787 15890 32793
rect 16114 32784 16120 32796
rect 16172 32784 16178 32836
rect 1104 32666 18860 32688
rect 1104 32614 2610 32666
rect 2662 32614 2674 32666
rect 2726 32614 2738 32666
rect 2790 32614 2802 32666
rect 2854 32614 2866 32666
rect 2918 32614 7610 32666
rect 7662 32614 7674 32666
rect 7726 32614 7738 32666
rect 7790 32614 7802 32666
rect 7854 32614 7866 32666
rect 7918 32614 12610 32666
rect 12662 32614 12674 32666
rect 12726 32614 12738 32666
rect 12790 32614 12802 32666
rect 12854 32614 12866 32666
rect 12918 32614 17610 32666
rect 17662 32614 17674 32666
rect 17726 32614 17738 32666
rect 17790 32614 17802 32666
rect 17854 32614 17866 32666
rect 17918 32614 18860 32666
rect 1104 32592 18860 32614
rect 7285 32555 7343 32561
rect 7285 32521 7297 32555
rect 7331 32552 7343 32555
rect 7466 32552 7472 32564
rect 7331 32524 7472 32552
rect 7331 32521 7343 32524
rect 7285 32515 7343 32521
rect 7466 32512 7472 32524
rect 7524 32512 7530 32564
rect 13354 32512 13360 32564
rect 13412 32552 13418 32564
rect 13412 32524 17141 32552
rect 13412 32512 13418 32524
rect 13814 32484 13820 32496
rect 11992 32456 13820 32484
rect 7193 32419 7251 32425
rect 7193 32385 7205 32419
rect 7239 32416 7251 32419
rect 7466 32416 7472 32428
rect 7239 32388 7472 32416
rect 7239 32385 7251 32388
rect 7193 32379 7251 32385
rect 7466 32376 7472 32388
rect 7524 32416 7530 32428
rect 8294 32416 8300 32428
rect 7524 32388 8300 32416
rect 7524 32376 7530 32388
rect 8294 32376 8300 32388
rect 8352 32376 8358 32428
rect 11992 32425 12020 32456
rect 13814 32444 13820 32456
rect 13872 32444 13878 32496
rect 17113 32493 17141 32524
rect 17098 32487 17156 32493
rect 15396 32456 16988 32484
rect 11977 32419 12035 32425
rect 11977 32385 11989 32419
rect 12023 32385 12035 32419
rect 11977 32379 12035 32385
rect 12244 32419 12302 32425
rect 12244 32385 12256 32419
rect 12290 32416 12302 32419
rect 15396 32416 15424 32456
rect 12290 32388 15424 32416
rect 12290 32385 12302 32388
rect 12244 32379 12302 32385
rect 16850 32376 16856 32428
rect 16908 32376 16914 32428
rect 16960 32416 16988 32456
rect 17098 32453 17110 32487
rect 17144 32453 17156 32487
rect 17098 32447 17156 32453
rect 18414 32416 18420 32428
rect 16960 32388 18420 32416
rect 18414 32376 18420 32388
rect 18472 32376 18478 32428
rect 7282 32308 7288 32360
rect 7340 32348 7346 32360
rect 7377 32351 7435 32357
rect 7377 32348 7389 32351
rect 7340 32320 7389 32348
rect 7340 32308 7346 32320
rect 7377 32317 7389 32320
rect 7423 32348 7435 32351
rect 8386 32348 8392 32360
rect 7423 32320 8392 32348
rect 7423 32317 7435 32320
rect 7377 32311 7435 32317
rect 8386 32308 8392 32320
rect 8444 32308 8450 32360
rect 2406 32240 2412 32292
rect 2464 32280 2470 32292
rect 11514 32280 11520 32292
rect 2464 32252 11520 32280
rect 2464 32240 2470 32252
rect 11514 32240 11520 32252
rect 11572 32240 11578 32292
rect 6730 32172 6736 32224
rect 6788 32212 6794 32224
rect 6825 32215 6883 32221
rect 6825 32212 6837 32215
rect 6788 32184 6837 32212
rect 6788 32172 6794 32184
rect 6825 32181 6837 32184
rect 6871 32181 6883 32215
rect 6825 32175 6883 32181
rect 6914 32172 6920 32224
rect 6972 32212 6978 32224
rect 7282 32212 7288 32224
rect 6972 32184 7288 32212
rect 6972 32172 6978 32184
rect 7282 32172 7288 32184
rect 7340 32172 7346 32224
rect 11790 32172 11796 32224
rect 11848 32212 11854 32224
rect 13357 32215 13415 32221
rect 13357 32212 13369 32215
rect 11848 32184 13369 32212
rect 11848 32172 11854 32184
rect 13357 32181 13369 32184
rect 13403 32212 13415 32215
rect 17954 32212 17960 32224
rect 13403 32184 17960 32212
rect 13403 32181 13415 32184
rect 13357 32175 13415 32181
rect 17954 32172 17960 32184
rect 18012 32172 18018 32224
rect 18233 32215 18291 32221
rect 18233 32181 18245 32215
rect 18279 32212 18291 32215
rect 18414 32212 18420 32224
rect 18279 32184 18420 32212
rect 18279 32181 18291 32184
rect 18233 32175 18291 32181
rect 18414 32172 18420 32184
rect 18472 32172 18478 32224
rect 1104 32122 18860 32144
rect 1104 32070 1950 32122
rect 2002 32070 2014 32122
rect 2066 32070 2078 32122
rect 2130 32070 2142 32122
rect 2194 32070 2206 32122
rect 2258 32070 6950 32122
rect 7002 32070 7014 32122
rect 7066 32070 7078 32122
rect 7130 32070 7142 32122
rect 7194 32070 7206 32122
rect 7258 32070 11950 32122
rect 12002 32070 12014 32122
rect 12066 32070 12078 32122
rect 12130 32070 12142 32122
rect 12194 32070 12206 32122
rect 12258 32070 16950 32122
rect 17002 32070 17014 32122
rect 17066 32070 17078 32122
rect 17130 32070 17142 32122
rect 17194 32070 17206 32122
rect 17258 32070 18860 32122
rect 1104 32048 18860 32070
rect 11330 31968 11336 32020
rect 11388 32008 11394 32020
rect 11514 32008 11520 32020
rect 11388 31980 11520 32008
rect 11388 31968 11394 31980
rect 11514 31968 11520 31980
rect 11572 31968 11578 32020
rect 16482 31968 16488 32020
rect 16540 31968 16546 32020
rect 6454 31832 6460 31884
rect 6512 31872 6518 31884
rect 9490 31872 9496 31884
rect 6512 31844 9496 31872
rect 6512 31832 6518 31844
rect 9490 31832 9496 31844
rect 9548 31832 9554 31884
rect 16500 31816 16528 31968
rect 16758 31872 16764 31884
rect 16592 31844 16764 31872
rect 16592 31816 16620 31844
rect 16758 31832 16764 31844
rect 16816 31832 16822 31884
rect 16482 31764 16488 31816
rect 16540 31764 16546 31816
rect 16574 31764 16580 31816
rect 16632 31764 16638 31816
rect 18046 31764 18052 31816
rect 18104 31764 18110 31816
rect 8018 31696 8024 31748
rect 8076 31696 8082 31748
rect 6914 31628 6920 31680
rect 6972 31668 6978 31680
rect 8036 31668 8064 31696
rect 6972 31640 8064 31668
rect 6972 31628 6978 31640
rect 8110 31628 8116 31680
rect 8168 31668 8174 31680
rect 8294 31668 8300 31680
rect 8168 31640 8300 31668
rect 8168 31628 8174 31640
rect 8294 31628 8300 31640
rect 8352 31628 8358 31680
rect 18230 31628 18236 31680
rect 18288 31628 18294 31680
rect 1104 31578 18860 31600
rect 1104 31526 2610 31578
rect 2662 31526 2674 31578
rect 2726 31526 2738 31578
rect 2790 31526 2802 31578
rect 2854 31526 2866 31578
rect 2918 31526 7610 31578
rect 7662 31526 7674 31578
rect 7726 31526 7738 31578
rect 7790 31526 7802 31578
rect 7854 31526 7866 31578
rect 7918 31526 12610 31578
rect 12662 31526 12674 31578
rect 12726 31526 12738 31578
rect 12790 31526 12802 31578
rect 12854 31526 12866 31578
rect 12918 31526 17610 31578
rect 17662 31526 17674 31578
rect 17726 31526 17738 31578
rect 17790 31526 17802 31578
rect 17854 31526 17866 31578
rect 17918 31526 18860 31578
rect 1104 31504 18860 31526
rect 1581 31467 1639 31473
rect 1581 31433 1593 31467
rect 1627 31464 1639 31467
rect 6914 31464 6920 31476
rect 1627 31436 6920 31464
rect 1627 31433 1639 31436
rect 1581 31427 1639 31433
rect 6914 31424 6920 31436
rect 6972 31424 6978 31476
rect 14734 31424 14740 31476
rect 14792 31464 14798 31476
rect 18233 31467 18291 31473
rect 18233 31464 18245 31467
rect 14792 31436 18245 31464
rect 14792 31424 14798 31436
rect 18233 31433 18245 31436
rect 18279 31433 18291 31467
rect 18233 31427 18291 31433
rect 6362 31356 6368 31408
rect 6420 31396 6426 31408
rect 17098 31399 17156 31405
rect 17098 31396 17110 31399
rect 6420 31368 17110 31396
rect 6420 31356 6426 31368
rect 17098 31365 17110 31368
rect 17144 31365 17156 31399
rect 17098 31359 17156 31365
rect 1762 31288 1768 31340
rect 1820 31288 1826 31340
rect 7282 31288 7288 31340
rect 7340 31288 7346 31340
rect 7374 31288 7380 31340
rect 7432 31328 7438 31340
rect 8202 31328 8208 31340
rect 7432 31300 8208 31328
rect 7432 31288 7438 31300
rect 8202 31288 8208 31300
rect 8260 31288 8266 31340
rect 16850 31288 16856 31340
rect 16908 31288 16914 31340
rect 7300 31136 7328 31288
rect 7282 31084 7288 31136
rect 7340 31084 7346 31136
rect 1104 31034 18860 31056
rect 1104 30982 1950 31034
rect 2002 30982 2014 31034
rect 2066 30982 2078 31034
rect 2130 30982 2142 31034
rect 2194 30982 2206 31034
rect 2258 30982 6950 31034
rect 7002 30982 7014 31034
rect 7066 30982 7078 31034
rect 7130 30982 7142 31034
rect 7194 30982 7206 31034
rect 7258 30982 11950 31034
rect 12002 30982 12014 31034
rect 12066 30982 12078 31034
rect 12130 30982 12142 31034
rect 12194 30982 12206 31034
rect 12258 30982 16950 31034
rect 17002 30982 17014 31034
rect 17066 30982 17078 31034
rect 17130 30982 17142 31034
rect 17194 30982 17206 31034
rect 17258 30982 18860 31034
rect 1104 30960 18860 30982
rect 6362 30744 6368 30796
rect 6420 30744 6426 30796
rect 6089 30651 6147 30657
rect 6089 30617 6101 30651
rect 6135 30648 6147 30651
rect 11238 30648 11244 30660
rect 6135 30620 11244 30648
rect 6135 30617 6147 30620
rect 6089 30611 6147 30617
rect 11238 30608 11244 30620
rect 11296 30648 11302 30660
rect 11296 30620 12434 30648
rect 11296 30608 11302 30620
rect 5718 30540 5724 30592
rect 5776 30540 5782 30592
rect 6181 30583 6239 30589
rect 6181 30549 6193 30583
rect 6227 30580 6239 30583
rect 9122 30580 9128 30592
rect 6227 30552 9128 30580
rect 6227 30549 6239 30552
rect 6181 30543 6239 30549
rect 9122 30540 9128 30552
rect 9180 30540 9186 30592
rect 12406 30580 12434 30620
rect 13262 30608 13268 30660
rect 13320 30648 13326 30660
rect 13722 30648 13728 30660
rect 13320 30620 13728 30648
rect 13320 30608 13326 30620
rect 13722 30608 13728 30620
rect 13780 30608 13786 30660
rect 19518 30580 19524 30592
rect 12406 30552 19524 30580
rect 19518 30540 19524 30552
rect 19576 30540 19582 30592
rect 1104 30490 18860 30512
rect 1104 30438 2610 30490
rect 2662 30438 2674 30490
rect 2726 30438 2738 30490
rect 2790 30438 2802 30490
rect 2854 30438 2866 30490
rect 2918 30438 7610 30490
rect 7662 30438 7674 30490
rect 7726 30438 7738 30490
rect 7790 30438 7802 30490
rect 7854 30438 7866 30490
rect 7918 30438 12610 30490
rect 12662 30438 12674 30490
rect 12726 30438 12738 30490
rect 12790 30438 12802 30490
rect 12854 30438 12866 30490
rect 12918 30438 17610 30490
rect 17662 30438 17674 30490
rect 17726 30438 17738 30490
rect 17790 30438 17802 30490
rect 17854 30438 17866 30490
rect 17918 30438 18860 30490
rect 1104 30416 18860 30438
rect 7101 30311 7159 30317
rect 7101 30277 7113 30311
rect 7147 30308 7159 30311
rect 7282 30308 7288 30320
rect 7147 30280 7288 30308
rect 7147 30277 7159 30280
rect 7101 30271 7159 30277
rect 7282 30268 7288 30280
rect 7340 30308 7346 30320
rect 7558 30308 7564 30320
rect 7340 30280 7564 30308
rect 7340 30268 7346 30280
rect 7558 30268 7564 30280
rect 7616 30268 7622 30320
rect 8018 30317 8024 30320
rect 8001 30311 8024 30317
rect 8001 30277 8013 30311
rect 8001 30271 8024 30277
rect 8018 30268 8024 30271
rect 8076 30268 8082 30320
rect 13262 30308 13268 30320
rect 12406 30280 13268 30308
rect 3234 30200 3240 30252
rect 3292 30200 3298 30252
rect 3786 30200 3792 30252
rect 3844 30240 3850 30252
rect 3844 30212 7236 30240
rect 3844 30200 3850 30212
rect 7208 30181 7236 30212
rect 7742 30200 7748 30252
rect 7800 30200 7806 30252
rect 12406 30240 12434 30280
rect 13262 30268 13268 30280
rect 13320 30308 13326 30320
rect 13630 30308 13636 30320
rect 13320 30280 13636 30308
rect 13320 30268 13326 30280
rect 13630 30268 13636 30280
rect 13688 30268 13694 30320
rect 14820 30311 14878 30317
rect 14820 30277 14832 30311
rect 14866 30308 14878 30311
rect 18874 30308 18880 30320
rect 14866 30280 18880 30308
rect 14866 30277 14878 30280
rect 14820 30271 14878 30277
rect 18874 30268 18880 30280
rect 18932 30268 18938 30320
rect 7852 30212 12434 30240
rect 7101 30175 7159 30181
rect 7101 30141 7113 30175
rect 7147 30141 7159 30175
rect 7101 30135 7159 30141
rect 7193 30175 7251 30181
rect 7193 30141 7205 30175
rect 7239 30172 7251 30175
rect 7852 30172 7880 30212
rect 13814 30200 13820 30252
rect 13872 30240 13878 30252
rect 14553 30243 14611 30249
rect 14553 30240 14565 30243
rect 13872 30212 14565 30240
rect 13872 30200 13878 30212
rect 14553 30209 14565 30212
rect 14599 30209 14611 30243
rect 17494 30240 17500 30252
rect 14553 30203 14611 30209
rect 14660 30212 17500 30240
rect 11790 30172 11796 30184
rect 7239 30144 7880 30172
rect 9048 30144 11796 30172
rect 7239 30141 7251 30144
rect 7193 30135 7251 30141
rect 6638 29996 6644 30048
rect 6696 29996 6702 30048
rect 7116 30036 7144 30135
rect 9048 30036 9076 30144
rect 11790 30132 11796 30144
rect 11848 30132 11854 30184
rect 14660 30172 14688 30212
rect 17494 30200 17500 30212
rect 17552 30200 17558 30252
rect 13556 30144 14688 30172
rect 9125 30107 9183 30113
rect 9125 30073 9137 30107
rect 9171 30104 9183 30107
rect 13556 30104 13584 30144
rect 16390 30104 16396 30116
rect 9171 30076 13584 30104
rect 15488 30076 16396 30104
rect 9171 30073 9183 30076
rect 9125 30067 9183 30073
rect 7116 30008 9076 30036
rect 10042 29996 10048 30048
rect 10100 30036 10106 30048
rect 15488 30036 15516 30076
rect 16390 30064 16396 30076
rect 16448 30064 16454 30116
rect 10100 30008 15516 30036
rect 10100 29996 10106 30008
rect 15930 29996 15936 30048
rect 15988 29996 15994 30048
rect 1104 29946 18860 29968
rect 1104 29894 1950 29946
rect 2002 29894 2014 29946
rect 2066 29894 2078 29946
rect 2130 29894 2142 29946
rect 2194 29894 2206 29946
rect 2258 29894 6950 29946
rect 7002 29894 7014 29946
rect 7066 29894 7078 29946
rect 7130 29894 7142 29946
rect 7194 29894 7206 29946
rect 7258 29894 11950 29946
rect 12002 29894 12014 29946
rect 12066 29894 12078 29946
rect 12130 29894 12142 29946
rect 12194 29894 12206 29946
rect 12258 29894 16950 29946
rect 17002 29894 17014 29946
rect 17066 29894 17078 29946
rect 17130 29894 17142 29946
rect 17194 29894 17206 29946
rect 17258 29894 18860 29946
rect 1104 29872 18860 29894
rect 3234 29792 3240 29844
rect 3292 29832 3298 29844
rect 14182 29832 14188 29844
rect 3292 29804 14188 29832
rect 3292 29792 3298 29804
rect 14182 29792 14188 29804
rect 14240 29792 14246 29844
rect 15654 29792 15660 29844
rect 15712 29792 15718 29844
rect 6638 29724 6644 29776
rect 6696 29764 6702 29776
rect 19334 29764 19340 29776
rect 6696 29736 19340 29764
rect 6696 29724 6702 29736
rect 19334 29724 19340 29736
rect 19392 29724 19398 29776
rect 7282 29656 7288 29708
rect 7340 29696 7346 29708
rect 7742 29696 7748 29708
rect 7340 29668 7748 29696
rect 7340 29656 7346 29668
rect 7742 29656 7748 29668
rect 7800 29696 7806 29708
rect 8754 29696 8760 29708
rect 7800 29668 8760 29696
rect 7800 29656 7806 29668
rect 8754 29656 8760 29668
rect 8812 29656 8818 29708
rect 9122 29656 9128 29708
rect 9180 29696 9186 29708
rect 15930 29696 15936 29708
rect 9180 29668 15936 29696
rect 9180 29656 9186 29668
rect 15930 29656 15936 29668
rect 15988 29656 15994 29708
rect 16301 29699 16359 29705
rect 16301 29665 16313 29699
rect 16347 29696 16359 29699
rect 17954 29696 17960 29708
rect 16347 29668 17960 29696
rect 16347 29665 16359 29668
rect 16301 29659 16359 29665
rect 17954 29656 17960 29668
rect 18012 29696 18018 29708
rect 19610 29696 19616 29708
rect 18012 29668 19616 29696
rect 18012 29656 18018 29668
rect 19610 29656 19616 29668
rect 19668 29656 19674 29708
rect 18049 29631 18107 29637
rect 18049 29597 18061 29631
rect 18095 29628 18107 29631
rect 18598 29628 18604 29640
rect 18095 29600 18604 29628
rect 18095 29597 18107 29600
rect 18049 29591 18107 29597
rect 18598 29588 18604 29600
rect 18656 29588 18662 29640
rect 7558 29452 7564 29504
rect 7616 29492 7622 29504
rect 9398 29492 9404 29504
rect 7616 29464 9404 29492
rect 7616 29452 7622 29464
rect 9398 29452 9404 29464
rect 9456 29452 9462 29504
rect 15470 29452 15476 29504
rect 15528 29492 15534 29504
rect 16022 29492 16028 29504
rect 15528 29464 16028 29492
rect 15528 29452 15534 29464
rect 16022 29452 16028 29464
rect 16080 29452 16086 29504
rect 16114 29452 16120 29504
rect 16172 29452 16178 29504
rect 18230 29452 18236 29504
rect 18288 29452 18294 29504
rect 1104 29402 18860 29424
rect 1104 29350 2610 29402
rect 2662 29350 2674 29402
rect 2726 29350 2738 29402
rect 2790 29350 2802 29402
rect 2854 29350 2866 29402
rect 2918 29350 7610 29402
rect 7662 29350 7674 29402
rect 7726 29350 7738 29402
rect 7790 29350 7802 29402
rect 7854 29350 7866 29402
rect 7918 29350 12610 29402
rect 12662 29350 12674 29402
rect 12726 29350 12738 29402
rect 12790 29350 12802 29402
rect 12854 29350 12866 29402
rect 12918 29350 17610 29402
rect 17662 29350 17674 29402
rect 17726 29350 17738 29402
rect 17790 29350 17802 29402
rect 17854 29350 17866 29402
rect 17918 29350 18860 29402
rect 1104 29328 18860 29350
rect 5442 29248 5448 29300
rect 5500 29288 5506 29300
rect 9585 29291 9643 29297
rect 9585 29288 9597 29291
rect 5500 29260 9597 29288
rect 5500 29248 5506 29260
rect 9585 29257 9597 29260
rect 9631 29257 9643 29291
rect 9585 29251 9643 29257
rect 4614 29180 4620 29232
rect 4672 29180 4678 29232
rect 7926 29180 7932 29232
rect 7984 29220 7990 29232
rect 8386 29220 8392 29232
rect 7984 29192 8392 29220
rect 7984 29180 7990 29192
rect 8386 29180 8392 29192
rect 8444 29180 8450 29232
rect 4430 29112 4436 29164
rect 4488 29112 4494 29164
rect 9953 29155 10011 29161
rect 9953 29121 9965 29155
rect 9999 29152 10011 29155
rect 10962 29152 10968 29164
rect 9999 29124 10968 29152
rect 9999 29121 10011 29124
rect 9953 29115 10011 29121
rect 10962 29112 10968 29124
rect 11020 29112 11026 29164
rect 8754 29044 8760 29096
rect 8812 29084 8818 29096
rect 9122 29084 9128 29096
rect 8812 29056 9128 29084
rect 8812 29044 8818 29056
rect 9122 29044 9128 29056
rect 9180 29044 9186 29096
rect 10042 29044 10048 29096
rect 10100 29044 10106 29096
rect 10229 29087 10287 29093
rect 10229 29053 10241 29087
rect 10275 29084 10287 29087
rect 10686 29084 10692 29096
rect 10275 29056 10692 29084
rect 10275 29053 10287 29056
rect 10229 29047 10287 29053
rect 6362 28976 6368 29028
rect 6420 29016 6426 29028
rect 10244 29016 10272 29047
rect 10686 29044 10692 29056
rect 10744 29044 10750 29096
rect 6420 28988 10272 29016
rect 6420 28976 6426 28988
rect 1104 28858 18860 28880
rect 1104 28806 1950 28858
rect 2002 28806 2014 28858
rect 2066 28806 2078 28858
rect 2130 28806 2142 28858
rect 2194 28806 2206 28858
rect 2258 28806 6950 28858
rect 7002 28806 7014 28858
rect 7066 28806 7078 28858
rect 7130 28806 7142 28858
rect 7194 28806 7206 28858
rect 7258 28806 11950 28858
rect 12002 28806 12014 28858
rect 12066 28806 12078 28858
rect 12130 28806 12142 28858
rect 12194 28806 12206 28858
rect 12258 28806 16950 28858
rect 17002 28806 17014 28858
rect 17066 28806 17078 28858
rect 17130 28806 17142 28858
rect 17194 28806 17206 28858
rect 17258 28806 18860 28858
rect 1104 28784 18860 28806
rect 9309 28747 9367 28753
rect 9309 28713 9321 28747
rect 9355 28744 9367 28747
rect 11054 28744 11060 28756
rect 9355 28716 11060 28744
rect 9355 28713 9367 28716
rect 9309 28707 9367 28713
rect 11054 28704 11060 28716
rect 11112 28704 11118 28756
rect 5353 28611 5411 28617
rect 5353 28577 5365 28611
rect 5399 28608 5411 28611
rect 9122 28608 9128 28620
rect 5399 28580 9128 28608
rect 5399 28577 5411 28580
rect 5353 28571 5411 28577
rect 9122 28568 9128 28580
rect 9180 28568 9186 28620
rect 9766 28568 9772 28620
rect 9824 28568 9830 28620
rect 5626 28500 5632 28552
rect 5684 28500 5690 28552
rect 9858 28432 9864 28484
rect 9916 28472 9922 28484
rect 10594 28472 10600 28484
rect 9916 28444 10600 28472
rect 9916 28432 9922 28444
rect 10594 28432 10600 28444
rect 10652 28432 10658 28484
rect 9769 28407 9827 28413
rect 9769 28373 9781 28407
rect 9815 28404 9827 28407
rect 10502 28404 10508 28416
rect 9815 28376 10508 28404
rect 9815 28373 9827 28376
rect 9769 28367 9827 28373
rect 10502 28364 10508 28376
rect 10560 28364 10566 28416
rect 1104 28314 18860 28336
rect 1104 28262 2610 28314
rect 2662 28262 2674 28314
rect 2726 28262 2738 28314
rect 2790 28262 2802 28314
rect 2854 28262 2866 28314
rect 2918 28262 7610 28314
rect 7662 28262 7674 28314
rect 7726 28262 7738 28314
rect 7790 28262 7802 28314
rect 7854 28262 7866 28314
rect 7918 28262 12610 28314
rect 12662 28262 12674 28314
rect 12726 28262 12738 28314
rect 12790 28262 12802 28314
rect 12854 28262 12866 28314
rect 12918 28262 17610 28314
rect 17662 28262 17674 28314
rect 17726 28262 17738 28314
rect 17790 28262 17802 28314
rect 17854 28262 17866 28314
rect 17918 28262 18860 28314
rect 1104 28240 18860 28262
rect 3326 28092 3332 28144
rect 3384 28132 3390 28144
rect 4310 28135 4368 28141
rect 4310 28132 4322 28135
rect 3384 28104 4322 28132
rect 3384 28092 3390 28104
rect 4310 28101 4322 28104
rect 4356 28101 4368 28135
rect 4310 28095 4368 28101
rect 10778 28024 10784 28076
rect 10836 28064 10842 28076
rect 18049 28067 18107 28073
rect 18049 28064 18061 28067
rect 10836 28036 18061 28064
rect 10836 28024 10842 28036
rect 18049 28033 18061 28036
rect 18095 28033 18107 28067
rect 18049 28027 18107 28033
rect 4062 27956 4068 28008
rect 4120 27956 4126 28008
rect 5445 27863 5503 27869
rect 5445 27829 5457 27863
rect 5491 27860 5503 27863
rect 10962 27860 10968 27872
rect 5491 27832 10968 27860
rect 5491 27829 5503 27832
rect 5445 27823 5503 27829
rect 10962 27820 10968 27832
rect 11020 27820 11026 27872
rect 17862 27820 17868 27872
rect 17920 27860 17926 27872
rect 18233 27863 18291 27869
rect 18233 27860 18245 27863
rect 17920 27832 18245 27860
rect 17920 27820 17926 27832
rect 18233 27829 18245 27832
rect 18279 27829 18291 27863
rect 18233 27823 18291 27829
rect 1104 27770 18860 27792
rect 1104 27718 1950 27770
rect 2002 27718 2014 27770
rect 2066 27718 2078 27770
rect 2130 27718 2142 27770
rect 2194 27718 2206 27770
rect 2258 27718 6950 27770
rect 7002 27718 7014 27770
rect 7066 27718 7078 27770
rect 7130 27718 7142 27770
rect 7194 27718 7206 27770
rect 7258 27718 11950 27770
rect 12002 27718 12014 27770
rect 12066 27718 12078 27770
rect 12130 27718 12142 27770
rect 12194 27718 12206 27770
rect 12258 27718 16950 27770
rect 17002 27718 17014 27770
rect 17066 27718 17078 27770
rect 17130 27718 17142 27770
rect 17194 27718 17206 27770
rect 17258 27718 18860 27770
rect 1104 27696 18860 27718
rect 4062 27548 4068 27600
rect 4120 27588 4126 27600
rect 7282 27588 7288 27600
rect 4120 27560 7288 27588
rect 4120 27548 4126 27560
rect 7282 27548 7288 27560
rect 7340 27548 7346 27600
rect 10870 27548 10876 27600
rect 10928 27588 10934 27600
rect 13906 27588 13912 27600
rect 10928 27560 13912 27588
rect 10928 27548 10934 27560
rect 13906 27548 13912 27560
rect 13964 27548 13970 27600
rect 18233 27591 18291 27597
rect 18233 27557 18245 27591
rect 18279 27588 18291 27591
rect 19150 27588 19156 27600
rect 18279 27560 19156 27588
rect 18279 27557 18291 27560
rect 18233 27551 18291 27557
rect 19150 27548 19156 27560
rect 19208 27548 19214 27600
rect 4154 27480 4160 27532
rect 4212 27520 4218 27532
rect 4249 27523 4307 27529
rect 4249 27520 4261 27523
rect 4212 27492 4261 27520
rect 4212 27480 4218 27492
rect 4249 27489 4261 27492
rect 4295 27489 4307 27523
rect 4249 27483 4307 27489
rect 4065 27455 4123 27461
rect 4065 27421 4077 27455
rect 4111 27452 4123 27455
rect 5074 27452 5080 27464
rect 4111 27424 5080 27452
rect 4111 27421 4123 27424
rect 4065 27415 4123 27421
rect 5074 27412 5080 27424
rect 5132 27412 5138 27464
rect 18049 27455 18107 27461
rect 18049 27421 18061 27455
rect 18095 27452 18107 27455
rect 18138 27452 18144 27464
rect 18095 27424 18144 27452
rect 18095 27421 18107 27424
rect 18049 27415 18107 27421
rect 18138 27412 18144 27424
rect 18196 27412 18202 27464
rect 1104 27226 18860 27248
rect 1104 27174 2610 27226
rect 2662 27174 2674 27226
rect 2726 27174 2738 27226
rect 2790 27174 2802 27226
rect 2854 27174 2866 27226
rect 2918 27174 7610 27226
rect 7662 27174 7674 27226
rect 7726 27174 7738 27226
rect 7790 27174 7802 27226
rect 7854 27174 7866 27226
rect 7918 27174 12610 27226
rect 12662 27174 12674 27226
rect 12726 27174 12738 27226
rect 12790 27174 12802 27226
rect 12854 27174 12866 27226
rect 12918 27174 17610 27226
rect 17662 27174 17674 27226
rect 17726 27174 17738 27226
rect 17790 27174 17802 27226
rect 17854 27174 17866 27226
rect 17918 27174 18860 27226
rect 1104 27152 18860 27174
rect 8386 27072 8392 27124
rect 8444 27112 8450 27124
rect 9490 27112 9496 27124
rect 8444 27084 9496 27112
rect 8444 27072 8450 27084
rect 9490 27072 9496 27084
rect 9548 27112 9554 27124
rect 14645 27115 14703 27121
rect 14645 27112 14657 27115
rect 9548 27084 14657 27112
rect 9548 27072 9554 27084
rect 14645 27081 14657 27084
rect 14691 27081 14703 27115
rect 14645 27075 14703 27081
rect 13814 27044 13820 27056
rect 13280 27016 13820 27044
rect 13280 26988 13308 27016
rect 13814 27004 13820 27016
rect 13872 27004 13878 27056
rect 1578 26936 1584 26988
rect 1636 26936 1642 26988
rect 13262 26936 13268 26988
rect 13320 26936 13326 26988
rect 13521 26979 13579 26985
rect 13521 26976 13533 26979
rect 13372 26948 13533 26976
rect 1486 26732 1492 26784
rect 1544 26772 1550 26784
rect 1596 26772 1624 26936
rect 8662 26868 8668 26920
rect 8720 26908 8726 26920
rect 9030 26908 9036 26920
rect 8720 26880 9036 26908
rect 8720 26868 8726 26880
rect 9030 26868 9036 26880
rect 9088 26868 9094 26920
rect 11790 26868 11796 26920
rect 11848 26908 11854 26920
rect 13372 26908 13400 26948
rect 13521 26945 13533 26948
rect 13567 26945 13579 26979
rect 13521 26939 13579 26945
rect 11848 26880 13400 26908
rect 11848 26868 11854 26880
rect 1544 26744 1624 26772
rect 1544 26732 1550 26744
rect 1104 26682 18860 26704
rect 1104 26630 1950 26682
rect 2002 26630 2014 26682
rect 2066 26630 2078 26682
rect 2130 26630 2142 26682
rect 2194 26630 2206 26682
rect 2258 26630 6950 26682
rect 7002 26630 7014 26682
rect 7066 26630 7078 26682
rect 7130 26630 7142 26682
rect 7194 26630 7206 26682
rect 7258 26630 11950 26682
rect 12002 26630 12014 26682
rect 12066 26630 12078 26682
rect 12130 26630 12142 26682
rect 12194 26630 12206 26682
rect 12258 26630 16950 26682
rect 17002 26630 17014 26682
rect 17066 26630 17078 26682
rect 17130 26630 17142 26682
rect 17194 26630 17206 26682
rect 17258 26630 18860 26682
rect 1104 26608 18860 26630
rect 3421 26571 3479 26577
rect 3421 26537 3433 26571
rect 3467 26568 3479 26571
rect 6178 26568 6184 26580
rect 3467 26540 6184 26568
rect 3467 26537 3479 26540
rect 3421 26531 3479 26537
rect 6178 26528 6184 26540
rect 6236 26528 6242 26580
rect 6917 26571 6975 26577
rect 6917 26537 6929 26571
rect 6963 26568 6975 26571
rect 7374 26568 7380 26580
rect 6963 26540 7380 26568
rect 6963 26537 6975 26540
rect 6917 26531 6975 26537
rect 7374 26528 7380 26540
rect 7432 26528 7438 26580
rect 4062 26392 4068 26444
rect 4120 26432 4126 26444
rect 5537 26435 5595 26441
rect 5537 26432 5549 26435
rect 4120 26404 5549 26432
rect 4120 26392 4126 26404
rect 5537 26401 5549 26404
rect 5583 26401 5595 26435
rect 5537 26395 5595 26401
rect 2041 26367 2099 26373
rect 2041 26333 2053 26367
rect 2087 26364 2099 26367
rect 4080 26364 4108 26392
rect 11514 26364 11520 26376
rect 2087 26336 4108 26364
rect 5184 26336 11520 26364
rect 2087 26333 2099 26336
rect 2041 26327 2099 26333
rect 2308 26299 2366 26305
rect 2308 26265 2320 26299
rect 2354 26296 2366 26299
rect 5184 26296 5212 26336
rect 11514 26324 11520 26336
rect 11572 26324 11578 26376
rect 5810 26305 5816 26308
rect 2354 26268 5212 26296
rect 2354 26265 2366 26268
rect 2308 26259 2366 26265
rect 5804 26259 5816 26305
rect 5810 26256 5816 26259
rect 5868 26256 5874 26308
rect 7282 26256 7288 26308
rect 7340 26296 7346 26308
rect 13262 26296 13268 26308
rect 7340 26268 13268 26296
rect 7340 26256 7346 26268
rect 13262 26256 13268 26268
rect 13320 26256 13326 26308
rect 7374 26188 7380 26240
rect 7432 26228 7438 26240
rect 8294 26228 8300 26240
rect 7432 26200 8300 26228
rect 7432 26188 7438 26200
rect 8294 26188 8300 26200
rect 8352 26188 8358 26240
rect 1104 26138 18860 26160
rect 1104 26086 2610 26138
rect 2662 26086 2674 26138
rect 2726 26086 2738 26138
rect 2790 26086 2802 26138
rect 2854 26086 2866 26138
rect 2918 26086 7610 26138
rect 7662 26086 7674 26138
rect 7726 26086 7738 26138
rect 7790 26086 7802 26138
rect 7854 26086 7866 26138
rect 7918 26086 12610 26138
rect 12662 26086 12674 26138
rect 12726 26086 12738 26138
rect 12790 26086 12802 26138
rect 12854 26086 12866 26138
rect 12918 26086 17610 26138
rect 17662 26086 17674 26138
rect 17726 26086 17738 26138
rect 17790 26086 17802 26138
rect 17854 26086 17866 26138
rect 17918 26086 18860 26138
rect 1104 26064 18860 26086
rect 10134 25984 10140 26036
rect 10192 25984 10198 26036
rect 10505 26027 10563 26033
rect 10505 25993 10517 26027
rect 10551 26024 10563 26027
rect 13722 26024 13728 26036
rect 10551 25996 13728 26024
rect 10551 25993 10563 25996
rect 10505 25987 10563 25993
rect 13722 25984 13728 25996
rect 13780 26024 13786 26036
rect 17494 26024 17500 26036
rect 13780 25996 17500 26024
rect 13780 25984 13786 25996
rect 17494 25984 17500 25996
rect 17552 25984 17558 26036
rect 14642 25888 14648 25900
rect 10612 25860 14648 25888
rect 9674 25780 9680 25832
rect 9732 25820 9738 25832
rect 10612 25829 10640 25860
rect 14642 25848 14648 25860
rect 14700 25848 14706 25900
rect 18049 25891 18107 25897
rect 18049 25857 18061 25891
rect 18095 25888 18107 25891
rect 18966 25888 18972 25900
rect 18095 25860 18972 25888
rect 18095 25857 18107 25860
rect 18049 25851 18107 25857
rect 18966 25848 18972 25860
rect 19024 25848 19030 25900
rect 10597 25823 10655 25829
rect 10597 25820 10609 25823
rect 9732 25792 10609 25820
rect 9732 25780 9738 25792
rect 10597 25789 10609 25792
rect 10643 25789 10655 25823
rect 10597 25783 10655 25789
rect 10778 25780 10784 25832
rect 10836 25780 10842 25832
rect 18230 25644 18236 25696
rect 18288 25644 18294 25696
rect 1104 25594 18860 25616
rect 1104 25542 1950 25594
rect 2002 25542 2014 25594
rect 2066 25542 2078 25594
rect 2130 25542 2142 25594
rect 2194 25542 2206 25594
rect 2258 25542 6950 25594
rect 7002 25542 7014 25594
rect 7066 25542 7078 25594
rect 7130 25542 7142 25594
rect 7194 25542 7206 25594
rect 7258 25542 11950 25594
rect 12002 25542 12014 25594
rect 12066 25542 12078 25594
rect 12130 25542 12142 25594
rect 12194 25542 12206 25594
rect 12258 25542 16950 25594
rect 17002 25542 17014 25594
rect 17066 25542 17078 25594
rect 17130 25542 17142 25594
rect 17194 25542 17206 25594
rect 17258 25542 18860 25594
rect 1104 25520 18860 25542
rect 1762 25440 1768 25492
rect 1820 25480 1826 25492
rect 1820 25452 5304 25480
rect 1820 25440 1826 25452
rect 5276 25412 5304 25452
rect 5350 25440 5356 25492
rect 5408 25440 5414 25492
rect 9861 25415 9919 25421
rect 9861 25412 9873 25415
rect 5276 25384 9873 25412
rect 9861 25381 9873 25384
rect 9907 25381 9919 25415
rect 9861 25375 9919 25381
rect 1486 25304 1492 25356
rect 1544 25344 1550 25356
rect 1762 25344 1768 25356
rect 1544 25316 1768 25344
rect 1544 25304 1550 25316
rect 1762 25304 1768 25316
rect 1820 25304 1826 25356
rect 5718 25304 5724 25356
rect 5776 25344 5782 25356
rect 6641 25347 6699 25353
rect 6641 25344 6653 25347
rect 5776 25316 6653 25344
rect 5776 25304 5782 25316
rect 6641 25313 6653 25316
rect 6687 25313 6699 25347
rect 6641 25307 6699 25313
rect 6917 25347 6975 25353
rect 6917 25313 6929 25347
rect 6963 25344 6975 25347
rect 7374 25344 7380 25356
rect 6963 25316 7380 25344
rect 6963 25313 6975 25316
rect 6917 25307 6975 25313
rect 7374 25304 7380 25316
rect 7432 25304 7438 25356
rect 10318 25304 10324 25356
rect 10376 25304 10382 25356
rect 10410 25304 10416 25356
rect 10468 25344 10474 25356
rect 12526 25344 12532 25356
rect 10468 25316 12532 25344
rect 10468 25304 10474 25316
rect 12526 25304 12532 25316
rect 12584 25304 12590 25356
rect 12897 25347 12955 25353
rect 12897 25313 12909 25347
rect 12943 25344 12955 25347
rect 13354 25344 13360 25356
rect 12943 25316 13360 25344
rect 12943 25313 12955 25316
rect 12897 25307 12955 25313
rect 13354 25304 13360 25316
rect 13412 25304 13418 25356
rect 3973 25279 4031 25285
rect 3973 25245 3985 25279
rect 4019 25276 4031 25279
rect 4062 25276 4068 25288
rect 4019 25248 4068 25276
rect 4019 25245 4031 25248
rect 3973 25239 4031 25245
rect 4062 25236 4068 25248
rect 4120 25236 4126 25288
rect 10226 25236 10232 25288
rect 10284 25236 10290 25288
rect 12434 25236 12440 25288
rect 12492 25276 12498 25288
rect 12713 25279 12771 25285
rect 12713 25276 12725 25279
rect 12492 25248 12725 25276
rect 12492 25236 12498 25248
rect 12713 25245 12725 25248
rect 12759 25276 12771 25279
rect 12986 25276 12992 25288
rect 12759 25248 12992 25276
rect 12759 25245 12771 25248
rect 12713 25239 12771 25245
rect 12986 25236 12992 25248
rect 13044 25236 13050 25288
rect 1486 25168 1492 25220
rect 1544 25208 1550 25220
rect 2314 25208 2320 25220
rect 1544 25180 2320 25208
rect 1544 25168 1550 25180
rect 2314 25168 2320 25180
rect 2372 25168 2378 25220
rect 4240 25211 4298 25217
rect 4240 25177 4252 25211
rect 4286 25208 4298 25211
rect 11514 25208 11520 25220
rect 4286 25180 11520 25208
rect 4286 25177 4298 25180
rect 4240 25171 4298 25177
rect 11514 25168 11520 25180
rect 11572 25168 11578 25220
rect 12805 25211 12863 25217
rect 12805 25177 12817 25211
rect 12851 25208 12863 25211
rect 13078 25208 13084 25220
rect 12851 25180 13084 25208
rect 12851 25177 12863 25180
rect 12805 25171 12863 25177
rect 13078 25168 13084 25180
rect 13136 25208 13142 25220
rect 15838 25208 15844 25220
rect 13136 25180 15844 25208
rect 13136 25168 13142 25180
rect 15838 25168 15844 25180
rect 15896 25168 15902 25220
rect 10502 25100 10508 25152
rect 10560 25140 10566 25152
rect 12345 25143 12403 25149
rect 12345 25140 12357 25143
rect 10560 25112 12357 25140
rect 10560 25100 10566 25112
rect 12345 25109 12357 25112
rect 12391 25109 12403 25143
rect 12345 25103 12403 25109
rect 1104 25050 18860 25072
rect 1104 24998 2610 25050
rect 2662 24998 2674 25050
rect 2726 24998 2738 25050
rect 2790 24998 2802 25050
rect 2854 24998 2866 25050
rect 2918 24998 7610 25050
rect 7662 24998 7674 25050
rect 7726 24998 7738 25050
rect 7790 24998 7802 25050
rect 7854 24998 7866 25050
rect 7918 24998 12610 25050
rect 12662 24998 12674 25050
rect 12726 24998 12738 25050
rect 12790 24998 12802 25050
rect 12854 24998 12866 25050
rect 12918 24998 17610 25050
rect 17662 24998 17674 25050
rect 17726 24998 17738 25050
rect 17790 24998 17802 25050
rect 17854 24998 17866 25050
rect 17918 24998 18860 25050
rect 1104 24976 18860 24998
rect 11422 24896 11428 24948
rect 11480 24936 11486 24948
rect 13814 24936 13820 24948
rect 11480 24908 13820 24936
rect 11480 24896 11486 24908
rect 13814 24896 13820 24908
rect 13872 24936 13878 24948
rect 17957 24939 18015 24945
rect 17957 24936 17969 24939
rect 13872 24908 17969 24936
rect 13872 24896 13878 24908
rect 17957 24905 17969 24908
rect 18003 24905 18015 24939
rect 17957 24899 18015 24905
rect 6730 24760 6736 24812
rect 6788 24800 6794 24812
rect 9217 24803 9275 24809
rect 9217 24800 9229 24803
rect 6788 24772 9229 24800
rect 6788 24760 6794 24772
rect 9217 24769 9229 24772
rect 9263 24769 9275 24803
rect 9217 24763 9275 24769
rect 9766 24760 9772 24812
rect 9824 24760 9830 24812
rect 9953 24803 10011 24809
rect 9953 24769 9965 24803
rect 9999 24800 10011 24803
rect 14826 24800 14832 24812
rect 9999 24772 14832 24800
rect 9999 24769 10011 24772
rect 9953 24763 10011 24769
rect 14826 24760 14832 24772
rect 14884 24760 14890 24812
rect 17954 24760 17960 24812
rect 18012 24800 18018 24812
rect 18012 24772 18184 24800
rect 18012 24760 18018 24772
rect 18156 24744 18184 24772
rect 14734 24692 14740 24744
rect 14792 24732 14798 24744
rect 15102 24732 15108 24744
rect 14792 24704 15108 24732
rect 14792 24692 14798 24704
rect 15102 24692 15108 24704
rect 15160 24692 15166 24744
rect 16390 24692 16396 24744
rect 16448 24732 16454 24744
rect 18049 24735 18107 24741
rect 18049 24732 18061 24735
rect 16448 24704 18061 24732
rect 16448 24692 16454 24704
rect 18049 24701 18061 24704
rect 18095 24701 18107 24735
rect 18049 24695 18107 24701
rect 18138 24692 18144 24744
rect 18196 24692 18202 24744
rect 14274 24624 14280 24676
rect 14332 24664 14338 24676
rect 17589 24667 17647 24673
rect 17589 24664 17601 24667
rect 14332 24636 17601 24664
rect 14332 24624 14338 24636
rect 17589 24633 17601 24636
rect 17635 24633 17647 24667
rect 17589 24627 17647 24633
rect 8938 24556 8944 24608
rect 8996 24596 9002 24608
rect 9033 24599 9091 24605
rect 9033 24596 9045 24599
rect 8996 24568 9045 24596
rect 8996 24556 9002 24568
rect 9033 24565 9045 24568
rect 9079 24565 9091 24599
rect 9033 24559 9091 24565
rect 1104 24506 18860 24528
rect 1104 24454 1950 24506
rect 2002 24454 2014 24506
rect 2066 24454 2078 24506
rect 2130 24454 2142 24506
rect 2194 24454 2206 24506
rect 2258 24454 6950 24506
rect 7002 24454 7014 24506
rect 7066 24454 7078 24506
rect 7130 24454 7142 24506
rect 7194 24454 7206 24506
rect 7258 24454 11950 24506
rect 12002 24454 12014 24506
rect 12066 24454 12078 24506
rect 12130 24454 12142 24506
rect 12194 24454 12206 24506
rect 12258 24454 16950 24506
rect 17002 24454 17014 24506
rect 17066 24454 17078 24506
rect 17130 24454 17142 24506
rect 17194 24454 17206 24506
rect 17258 24454 18860 24506
rect 1104 24432 18860 24454
rect 14734 24148 14740 24200
rect 14792 24188 14798 24200
rect 18049 24191 18107 24197
rect 18049 24188 18061 24191
rect 14792 24160 18061 24188
rect 14792 24148 14798 24160
rect 18049 24157 18061 24160
rect 18095 24157 18107 24191
rect 18049 24151 18107 24157
rect 6270 24080 6276 24132
rect 6328 24120 6334 24132
rect 13078 24120 13084 24132
rect 6328 24092 13084 24120
rect 6328 24080 6334 24092
rect 13078 24080 13084 24092
rect 13136 24120 13142 24132
rect 13722 24120 13728 24132
rect 13136 24092 13728 24120
rect 13136 24080 13142 24092
rect 13722 24080 13728 24092
rect 13780 24080 13786 24132
rect 18230 24012 18236 24064
rect 18288 24012 18294 24064
rect 1104 23962 18860 23984
rect 1104 23910 2610 23962
rect 2662 23910 2674 23962
rect 2726 23910 2738 23962
rect 2790 23910 2802 23962
rect 2854 23910 2866 23962
rect 2918 23910 7610 23962
rect 7662 23910 7674 23962
rect 7726 23910 7738 23962
rect 7790 23910 7802 23962
rect 7854 23910 7866 23962
rect 7918 23910 12610 23962
rect 12662 23910 12674 23962
rect 12726 23910 12738 23962
rect 12790 23910 12802 23962
rect 12854 23910 12866 23962
rect 12918 23910 17610 23962
rect 17662 23910 17674 23962
rect 17726 23910 17738 23962
rect 17790 23910 17802 23962
rect 17854 23910 17866 23962
rect 17918 23910 18860 23962
rect 1104 23888 18860 23910
rect 9306 23808 9312 23860
rect 9364 23808 9370 23860
rect 16666 23808 16672 23860
rect 16724 23848 16730 23860
rect 17405 23851 17463 23857
rect 17405 23848 17417 23851
rect 16724 23820 17417 23848
rect 16724 23808 16730 23820
rect 17405 23817 17417 23820
rect 17451 23817 17463 23851
rect 17405 23811 17463 23817
rect 7374 23740 7380 23792
rect 7432 23780 7438 23792
rect 8174 23783 8232 23789
rect 8174 23780 8186 23783
rect 7432 23752 8186 23780
rect 7432 23740 7438 23752
rect 8174 23749 8186 23752
rect 8220 23749 8232 23783
rect 8174 23743 8232 23749
rect 13722 23740 13728 23792
rect 13780 23780 13786 23792
rect 17221 23783 17279 23789
rect 17221 23780 17233 23783
rect 13780 23752 17233 23780
rect 13780 23740 13786 23752
rect 17221 23749 17233 23752
rect 17267 23749 17279 23783
rect 17221 23743 17279 23749
rect 3421 23715 3479 23721
rect 3421 23681 3433 23715
rect 3467 23712 3479 23715
rect 6454 23712 6460 23724
rect 3467 23684 6460 23712
rect 3467 23681 3479 23684
rect 3421 23675 3479 23681
rect 6454 23672 6460 23684
rect 6512 23672 6518 23724
rect 7282 23672 7288 23724
rect 7340 23712 7346 23724
rect 7929 23715 7987 23721
rect 7929 23712 7941 23715
rect 7340 23684 7941 23712
rect 7340 23672 7346 23684
rect 7929 23681 7941 23684
rect 7975 23681 7987 23715
rect 7929 23675 7987 23681
rect 12526 23672 12532 23724
rect 12584 23712 12590 23724
rect 17497 23715 17555 23721
rect 17497 23712 17509 23715
rect 12584 23684 17509 23712
rect 12584 23672 12590 23684
rect 17497 23681 17509 23684
rect 17543 23681 17555 23715
rect 17497 23675 17555 23681
rect 16574 23604 16580 23656
rect 16632 23604 16638 23656
rect 3237 23511 3295 23517
rect 3237 23477 3249 23511
rect 3283 23508 3295 23511
rect 11330 23508 11336 23520
rect 3283 23480 11336 23508
rect 3283 23477 3295 23480
rect 3237 23471 3295 23477
rect 11330 23468 11336 23480
rect 11388 23468 11394 23520
rect 16592 23508 16620 23604
rect 16942 23536 16948 23588
rect 17000 23536 17006 23588
rect 16758 23508 16764 23520
rect 16592 23480 16764 23508
rect 16758 23468 16764 23480
rect 16816 23468 16822 23520
rect 1104 23418 18860 23440
rect 1104 23366 1950 23418
rect 2002 23366 2014 23418
rect 2066 23366 2078 23418
rect 2130 23366 2142 23418
rect 2194 23366 2206 23418
rect 2258 23366 6950 23418
rect 7002 23366 7014 23418
rect 7066 23366 7078 23418
rect 7130 23366 7142 23418
rect 7194 23366 7206 23418
rect 7258 23366 11950 23418
rect 12002 23366 12014 23418
rect 12066 23366 12078 23418
rect 12130 23366 12142 23418
rect 12194 23366 12206 23418
rect 12258 23366 16950 23418
rect 17002 23366 17014 23418
rect 17066 23366 17078 23418
rect 17130 23366 17142 23418
rect 17194 23366 17206 23418
rect 17258 23366 18860 23418
rect 1104 23344 18860 23366
rect 18046 23264 18052 23316
rect 18104 23304 18110 23316
rect 18414 23304 18420 23316
rect 18104 23276 18420 23304
rect 18104 23264 18110 23276
rect 18414 23264 18420 23276
rect 18472 23264 18478 23316
rect 1104 22874 18860 22896
rect 1104 22822 2610 22874
rect 2662 22822 2674 22874
rect 2726 22822 2738 22874
rect 2790 22822 2802 22874
rect 2854 22822 2866 22874
rect 2918 22822 7610 22874
rect 7662 22822 7674 22874
rect 7726 22822 7738 22874
rect 7790 22822 7802 22874
rect 7854 22822 7866 22874
rect 7918 22822 12610 22874
rect 12662 22822 12674 22874
rect 12726 22822 12738 22874
rect 12790 22822 12802 22874
rect 12854 22822 12866 22874
rect 12918 22822 17610 22874
rect 17662 22822 17674 22874
rect 17726 22822 17738 22874
rect 17790 22822 17802 22874
rect 17854 22822 17866 22874
rect 17918 22822 18860 22874
rect 1104 22800 18860 22822
rect 7926 22720 7932 22772
rect 7984 22760 7990 22772
rect 8202 22760 8208 22772
rect 7984 22732 8208 22760
rect 7984 22720 7990 22732
rect 8202 22720 8208 22732
rect 8260 22720 8266 22772
rect 10318 22720 10324 22772
rect 10376 22760 10382 22772
rect 13354 22760 13360 22772
rect 10376 22732 13360 22760
rect 10376 22720 10382 22732
rect 13354 22720 13360 22732
rect 13412 22760 13418 22772
rect 17681 22763 17739 22769
rect 17681 22760 17693 22763
rect 13412 22732 17693 22760
rect 13412 22720 13418 22732
rect 17681 22729 17693 22732
rect 17727 22729 17739 22763
rect 17681 22723 17739 22729
rect 5534 22584 5540 22636
rect 5592 22624 5598 22636
rect 9858 22624 9864 22636
rect 5592 22596 9864 22624
rect 5592 22584 5598 22596
rect 9858 22584 9864 22596
rect 9916 22624 9922 22636
rect 17773 22627 17831 22633
rect 17773 22624 17785 22627
rect 9916 22596 17785 22624
rect 9916 22584 9922 22596
rect 17773 22593 17785 22596
rect 17819 22593 17831 22627
rect 17773 22587 17831 22593
rect 17681 22559 17739 22565
rect 17681 22525 17693 22559
rect 17727 22556 17739 22559
rect 18046 22556 18052 22568
rect 17727 22528 18052 22556
rect 17727 22525 17739 22528
rect 17681 22519 17739 22525
rect 18046 22516 18052 22528
rect 18104 22516 18110 22568
rect 17218 22448 17224 22500
rect 17276 22448 17282 22500
rect 1104 22330 18860 22352
rect 1104 22278 1950 22330
rect 2002 22278 2014 22330
rect 2066 22278 2078 22330
rect 2130 22278 2142 22330
rect 2194 22278 2206 22330
rect 2258 22278 6950 22330
rect 7002 22278 7014 22330
rect 7066 22278 7078 22330
rect 7130 22278 7142 22330
rect 7194 22278 7206 22330
rect 7258 22278 11950 22330
rect 12002 22278 12014 22330
rect 12066 22278 12078 22330
rect 12130 22278 12142 22330
rect 12194 22278 12206 22330
rect 12258 22278 16950 22330
rect 17002 22278 17014 22330
rect 17066 22278 17078 22330
rect 17130 22278 17142 22330
rect 17194 22278 17206 22330
rect 17258 22278 18860 22330
rect 1104 22256 18860 22278
rect 2409 22151 2467 22157
rect 2409 22117 2421 22151
rect 2455 22148 2467 22151
rect 7009 22151 7067 22157
rect 2455 22120 2489 22148
rect 2455 22117 2467 22120
rect 2409 22111 2467 22117
rect 7009 22117 7021 22151
rect 7055 22148 7067 22151
rect 9214 22148 9220 22160
rect 7055 22120 7089 22148
rect 7300 22120 9220 22148
rect 7055 22117 7067 22120
rect 7009 22111 7067 22117
rect 1394 22040 1400 22092
rect 1452 22080 1458 22092
rect 2424 22080 2452 22111
rect 1452 22052 2452 22080
rect 2869 22083 2927 22089
rect 1452 22040 1458 22052
rect 2869 22049 2881 22083
rect 2915 22080 2927 22083
rect 4154 22080 4160 22092
rect 2915 22052 4160 22080
rect 2915 22049 2927 22052
rect 2869 22043 2927 22049
rect 4154 22040 4160 22052
rect 4212 22040 4218 22092
rect 6178 22040 6184 22092
rect 6236 22080 6242 22092
rect 7024 22080 7052 22111
rect 7300 22094 7328 22120
rect 9214 22108 9220 22120
rect 9272 22108 9278 22160
rect 9766 22108 9772 22160
rect 9824 22148 9830 22160
rect 16206 22148 16212 22160
rect 9824 22120 16212 22148
rect 9824 22108 9830 22120
rect 16206 22108 16212 22120
rect 16264 22108 16270 22160
rect 7116 22092 7328 22094
rect 6236 22052 7052 22080
rect 6236 22040 6242 22052
rect 7098 22040 7104 22092
rect 7156 22066 7328 22092
rect 7156 22040 7162 22066
rect 5169 22015 5227 22021
rect 5169 21981 5181 22015
rect 5215 22012 5227 22015
rect 6914 22012 6920 22024
rect 5215 21984 6920 22012
rect 5215 21981 5227 21984
rect 5169 21975 5227 21981
rect 6914 21972 6920 21984
rect 6972 21972 6978 22024
rect 7193 22015 7251 22021
rect 7193 21981 7205 22015
rect 7239 22012 7251 22015
rect 9490 22012 9496 22024
rect 7239 21984 9496 22012
rect 7239 21981 7251 21984
rect 7193 21975 7251 21981
rect 9490 21972 9496 21984
rect 9548 21972 9554 22024
rect 14553 22015 14611 22021
rect 14553 21981 14565 22015
rect 14599 22012 14611 22015
rect 15194 22012 15200 22024
rect 14599 21984 15200 22012
rect 14599 21981 14611 21984
rect 14553 21975 14611 21981
rect 15194 21972 15200 21984
rect 15252 21972 15258 22024
rect 18046 21972 18052 22024
rect 18104 21972 18110 22024
rect 2961 21947 3019 21953
rect 2961 21913 2973 21947
rect 3007 21944 3019 21947
rect 3326 21944 3332 21956
rect 3007 21916 3332 21944
rect 3007 21913 3019 21916
rect 2961 21907 3019 21913
rect 3326 21904 3332 21916
rect 3384 21904 3390 21956
rect 3421 21947 3479 21953
rect 3421 21913 3433 21947
rect 3467 21944 3479 21947
rect 4157 21947 4215 21953
rect 4157 21944 4169 21947
rect 3467 21916 4169 21944
rect 3467 21913 3479 21916
rect 3421 21907 3479 21913
rect 4157 21913 4169 21916
rect 4203 21944 4215 21947
rect 4525 21947 4583 21953
rect 4525 21944 4537 21947
rect 4203 21916 4537 21944
rect 4203 21913 4215 21916
rect 4157 21907 4215 21913
rect 4525 21913 4537 21916
rect 4571 21944 4583 21947
rect 4893 21947 4951 21953
rect 4893 21944 4905 21947
rect 4571 21916 4905 21944
rect 4571 21913 4583 21916
rect 4525 21907 4583 21913
rect 4893 21913 4905 21916
rect 4939 21944 4951 21947
rect 5436 21947 5494 21953
rect 5436 21944 5448 21947
rect 4939 21916 5448 21944
rect 4939 21913 4951 21916
rect 4893 21907 4951 21913
rect 5436 21913 5448 21916
rect 5482 21944 5494 21947
rect 6932 21944 6960 21972
rect 7282 21944 7288 21956
rect 5482 21916 6776 21944
rect 6932 21916 7288 21944
rect 5482 21913 5494 21916
rect 5436 21907 5494 21913
rect 2869 21879 2927 21885
rect 2869 21845 2881 21879
rect 2915 21876 2927 21879
rect 6454 21876 6460 21888
rect 2915 21848 6460 21876
rect 2915 21845 2927 21848
rect 2869 21839 2927 21845
rect 6454 21836 6460 21848
rect 6512 21836 6518 21888
rect 6549 21879 6607 21885
rect 6549 21845 6561 21879
rect 6595 21876 6607 21879
rect 6638 21876 6644 21888
rect 6595 21848 6644 21876
rect 6595 21845 6607 21848
rect 6549 21839 6607 21845
rect 6638 21836 6644 21848
rect 6696 21836 6702 21888
rect 6748 21876 6776 21916
rect 7282 21904 7288 21916
rect 7340 21904 7346 21956
rect 6917 21879 6975 21885
rect 6917 21876 6929 21879
rect 6748 21848 6929 21876
rect 6917 21845 6929 21848
rect 6963 21876 6975 21879
rect 7098 21876 7104 21888
rect 6963 21848 7104 21876
rect 6963 21845 6975 21848
rect 6917 21839 6975 21845
rect 7098 21836 7104 21848
rect 7156 21836 7162 21888
rect 7926 21836 7932 21888
rect 7984 21876 7990 21888
rect 8202 21876 8208 21888
rect 7984 21848 8208 21876
rect 7984 21836 7990 21848
rect 8202 21836 8208 21848
rect 8260 21836 8266 21888
rect 11238 21836 11244 21888
rect 11296 21876 11302 21888
rect 12342 21876 12348 21888
rect 11296 21848 12348 21876
rect 11296 21836 11302 21848
rect 12342 21836 12348 21848
rect 12400 21836 12406 21888
rect 14090 21836 14096 21888
rect 14148 21876 14154 21888
rect 14369 21879 14427 21885
rect 14369 21876 14381 21879
rect 14148 21848 14381 21876
rect 14148 21836 14154 21848
rect 14369 21845 14381 21848
rect 14415 21845 14427 21879
rect 14369 21839 14427 21845
rect 18230 21836 18236 21888
rect 18288 21836 18294 21888
rect 1104 21786 18860 21808
rect 1104 21734 2610 21786
rect 2662 21734 2674 21786
rect 2726 21734 2738 21786
rect 2790 21734 2802 21786
rect 2854 21734 2866 21786
rect 2918 21734 7610 21786
rect 7662 21734 7674 21786
rect 7726 21734 7738 21786
rect 7790 21734 7802 21786
rect 7854 21734 7866 21786
rect 7918 21734 12610 21786
rect 12662 21734 12674 21786
rect 12726 21734 12738 21786
rect 12790 21734 12802 21786
rect 12854 21734 12866 21786
rect 12918 21734 17610 21786
rect 17662 21734 17674 21786
rect 17726 21734 17738 21786
rect 17790 21734 17802 21786
rect 17854 21734 17866 21786
rect 17918 21734 18860 21786
rect 1104 21712 18860 21734
rect 3326 21632 3332 21684
rect 3384 21672 3390 21684
rect 10778 21672 10784 21684
rect 3384 21644 10784 21672
rect 3384 21632 3390 21644
rect 10778 21632 10784 21644
rect 10836 21632 10842 21684
rect 11149 21675 11207 21681
rect 11149 21641 11161 21675
rect 11195 21672 11207 21675
rect 11885 21675 11943 21681
rect 11885 21672 11897 21675
rect 11195 21644 11897 21672
rect 11195 21641 11207 21644
rect 11149 21635 11207 21641
rect 11885 21641 11897 21644
rect 11931 21672 11943 21675
rect 12345 21675 12403 21681
rect 12345 21672 12357 21675
rect 11931 21644 12357 21672
rect 11931 21641 11943 21644
rect 11885 21635 11943 21641
rect 12345 21641 12357 21644
rect 12391 21672 12403 21675
rect 12713 21675 12771 21681
rect 12713 21672 12725 21675
rect 12391 21644 12725 21672
rect 12391 21641 12403 21644
rect 12345 21635 12403 21641
rect 12713 21641 12725 21644
rect 12759 21672 12771 21675
rect 19886 21672 19892 21684
rect 12759 21644 19892 21672
rect 12759 21641 12771 21644
rect 12713 21635 12771 21641
rect 19886 21632 19892 21644
rect 19944 21632 19950 21684
rect 3142 21496 3148 21548
rect 3200 21536 3206 21548
rect 11793 21539 11851 21545
rect 11793 21536 11805 21539
rect 3200 21508 11805 21536
rect 3200 21496 3206 21508
rect 11793 21505 11805 21508
rect 11839 21505 11851 21539
rect 11793 21499 11851 21505
rect 6454 21428 6460 21480
rect 6512 21468 6518 21480
rect 11422 21468 11428 21480
rect 6512 21440 11428 21468
rect 6512 21428 6518 21440
rect 11422 21428 11428 21440
rect 11480 21428 11486 21480
rect 12342 21292 12348 21344
rect 12400 21332 12406 21344
rect 18782 21332 18788 21344
rect 12400 21304 18788 21332
rect 12400 21292 12406 21304
rect 18782 21292 18788 21304
rect 18840 21292 18846 21344
rect 1104 21242 18860 21264
rect 1104 21190 1950 21242
rect 2002 21190 2014 21242
rect 2066 21190 2078 21242
rect 2130 21190 2142 21242
rect 2194 21190 2206 21242
rect 2258 21190 6950 21242
rect 7002 21190 7014 21242
rect 7066 21190 7078 21242
rect 7130 21190 7142 21242
rect 7194 21190 7206 21242
rect 7258 21190 11950 21242
rect 12002 21190 12014 21242
rect 12066 21190 12078 21242
rect 12130 21190 12142 21242
rect 12194 21190 12206 21242
rect 12258 21190 16950 21242
rect 17002 21190 17014 21242
rect 17066 21190 17078 21242
rect 17130 21190 17142 21242
rect 17194 21190 17206 21242
rect 17258 21190 18860 21242
rect 1104 21168 18860 21190
rect 9122 21088 9128 21140
rect 9180 21088 9186 21140
rect 12986 21088 12992 21140
rect 13044 21128 13050 21140
rect 17129 21131 17187 21137
rect 17129 21128 17141 21131
rect 13044 21100 17141 21128
rect 13044 21088 13050 21100
rect 17129 21097 17141 21100
rect 17175 21097 17187 21131
rect 17129 21091 17187 21097
rect 8297 21063 8355 21069
rect 8297 21029 8309 21063
rect 8343 21060 8355 21063
rect 9674 21060 9680 21072
rect 8343 21032 9680 21060
rect 8343 21029 8355 21032
rect 8297 21023 8355 21029
rect 9674 21020 9680 21032
rect 9732 21020 9738 21072
rect 13262 21060 13268 21072
rect 9784 21032 13268 21060
rect 6822 20952 6828 21004
rect 6880 20992 6886 21004
rect 6917 20995 6975 21001
rect 6917 20992 6929 20995
rect 6880 20964 6929 20992
rect 6880 20952 6886 20964
rect 6917 20961 6929 20964
rect 6963 20961 6975 20995
rect 6917 20955 6975 20961
rect 9398 20952 9404 21004
rect 9456 20992 9462 21004
rect 9784 21001 9812 21032
rect 13262 21020 13268 21032
rect 13320 21060 13326 21072
rect 15010 21060 15016 21072
rect 13320 21032 15016 21060
rect 13320 21020 13326 21032
rect 15010 21020 15016 21032
rect 15068 21020 15074 21072
rect 9585 20995 9643 21001
rect 9585 20992 9597 20995
rect 9456 20964 9597 20992
rect 9456 20952 9462 20964
rect 9585 20961 9597 20964
rect 9631 20961 9643 20995
rect 9585 20955 9643 20961
rect 9769 20995 9827 21001
rect 9769 20961 9781 20995
rect 9815 20961 9827 20995
rect 9769 20955 9827 20961
rect 13722 20952 13728 21004
rect 13780 20992 13786 21004
rect 15749 20995 15807 21001
rect 15749 20992 15761 20995
rect 13780 20964 15761 20992
rect 13780 20952 13786 20964
rect 15749 20961 15761 20964
rect 15795 20961 15807 20995
rect 15749 20955 15807 20961
rect 6273 20927 6331 20933
rect 6273 20893 6285 20927
rect 6319 20924 6331 20927
rect 6641 20927 6699 20933
rect 6641 20924 6653 20927
rect 6319 20896 6653 20924
rect 6319 20893 6331 20896
rect 6273 20887 6331 20893
rect 6641 20893 6653 20896
rect 6687 20924 6699 20927
rect 7184 20927 7242 20933
rect 7184 20924 7196 20927
rect 6687 20896 7196 20924
rect 6687 20893 6699 20896
rect 6641 20887 6699 20893
rect 7184 20893 7196 20896
rect 7230 20924 7242 20927
rect 12342 20924 12348 20936
rect 7230 20896 12348 20924
rect 7230 20893 7242 20896
rect 7184 20887 7242 20893
rect 12342 20884 12348 20896
rect 12400 20884 12406 20936
rect 14182 20884 14188 20936
rect 14240 20924 14246 20936
rect 14642 20924 14648 20936
rect 14240 20896 14648 20924
rect 14240 20884 14246 20896
rect 14642 20884 14648 20896
rect 14700 20884 14706 20936
rect 10778 20816 10784 20868
rect 10836 20856 10842 20868
rect 14826 20856 14832 20868
rect 10836 20828 14832 20856
rect 10836 20816 10842 20828
rect 14826 20816 14832 20828
rect 14884 20856 14890 20868
rect 15013 20859 15071 20865
rect 15013 20856 15025 20859
rect 14884 20828 15025 20856
rect 14884 20816 14890 20828
rect 15013 20825 15025 20828
rect 15059 20825 15071 20859
rect 15013 20819 15071 20825
rect 16016 20859 16074 20865
rect 16016 20825 16028 20859
rect 16062 20825 16074 20859
rect 16016 20819 16074 20825
rect 9306 20748 9312 20800
rect 9364 20788 9370 20800
rect 9493 20791 9551 20797
rect 9493 20788 9505 20791
rect 9364 20760 9505 20788
rect 9364 20748 9370 20760
rect 9493 20757 9505 20760
rect 9539 20788 9551 20791
rect 15654 20788 15660 20800
rect 9539 20760 15660 20788
rect 9539 20757 9551 20760
rect 9493 20751 9551 20757
rect 15654 20748 15660 20760
rect 15712 20748 15718 20800
rect 15930 20748 15936 20800
rect 15988 20788 15994 20800
rect 16040 20788 16068 20819
rect 15988 20760 16068 20788
rect 15988 20748 15994 20760
rect 1104 20698 18860 20720
rect 1104 20646 2610 20698
rect 2662 20646 2674 20698
rect 2726 20646 2738 20698
rect 2790 20646 2802 20698
rect 2854 20646 2866 20698
rect 2918 20646 7610 20698
rect 7662 20646 7674 20698
rect 7726 20646 7738 20698
rect 7790 20646 7802 20698
rect 7854 20646 7866 20698
rect 7918 20646 12610 20698
rect 12662 20646 12674 20698
rect 12726 20646 12738 20698
rect 12790 20646 12802 20698
rect 12854 20646 12866 20698
rect 12918 20646 17610 20698
rect 17662 20646 17674 20698
rect 17726 20646 17738 20698
rect 17790 20646 17802 20698
rect 17854 20646 17866 20698
rect 17918 20646 18860 20698
rect 1104 20624 18860 20646
rect 4338 20544 4344 20596
rect 4396 20584 4402 20596
rect 4396 20556 9674 20584
rect 4396 20544 4402 20556
rect 2133 20519 2191 20525
rect 2133 20485 2145 20519
rect 2179 20516 2191 20519
rect 8386 20516 8392 20528
rect 2179 20488 8392 20516
rect 2179 20485 2191 20488
rect 2133 20479 2191 20485
rect 8386 20476 8392 20488
rect 8444 20476 8450 20528
rect 2225 20451 2283 20457
rect 2225 20417 2237 20451
rect 2271 20448 2283 20451
rect 5534 20448 5540 20460
rect 2271 20420 5540 20448
rect 2271 20417 2283 20420
rect 2225 20411 2283 20417
rect 5534 20408 5540 20420
rect 5592 20408 5598 20460
rect 9646 20448 9674 20556
rect 11974 20544 11980 20596
rect 12032 20584 12038 20596
rect 16945 20587 17003 20593
rect 16945 20584 16957 20587
rect 12032 20556 16957 20584
rect 12032 20544 12038 20556
rect 16945 20553 16957 20556
rect 16991 20553 17003 20587
rect 16945 20547 17003 20553
rect 17218 20544 17224 20596
rect 17276 20584 17282 20596
rect 17313 20587 17371 20593
rect 17313 20584 17325 20587
rect 17276 20556 17325 20584
rect 17276 20544 17282 20556
rect 17313 20553 17325 20556
rect 17359 20553 17371 20587
rect 17313 20547 17371 20553
rect 14918 20476 14924 20528
rect 14976 20476 14982 20528
rect 11957 20451 12015 20457
rect 11957 20448 11969 20451
rect 9646 20420 11969 20448
rect 11957 20417 11969 20420
rect 12003 20417 12015 20451
rect 11957 20411 12015 20417
rect 14829 20451 14887 20457
rect 14829 20417 14841 20451
rect 14875 20448 14887 20451
rect 16482 20448 16488 20460
rect 14875 20420 16488 20448
rect 14875 20417 14887 20420
rect 14829 20411 14887 20417
rect 16482 20408 16488 20420
rect 16540 20408 16546 20460
rect 2133 20383 2191 20389
rect 2133 20349 2145 20383
rect 2179 20349 2191 20383
rect 2133 20343 2191 20349
rect 1673 20315 1731 20321
rect 1673 20281 1685 20315
rect 1719 20312 1731 20315
rect 1854 20312 1860 20324
rect 1719 20284 1860 20312
rect 1719 20281 1731 20284
rect 1673 20275 1731 20281
rect 1854 20272 1860 20284
rect 1912 20272 1918 20324
rect 2148 20312 2176 20343
rect 11422 20340 11428 20392
rect 11480 20380 11486 20392
rect 11701 20383 11759 20389
rect 11701 20380 11713 20383
rect 11480 20352 11713 20380
rect 11480 20340 11486 20352
rect 11701 20349 11713 20352
rect 11747 20349 11759 20383
rect 11701 20343 11759 20349
rect 13538 20340 13544 20392
rect 13596 20380 13602 20392
rect 15013 20383 15071 20389
rect 15013 20380 15025 20383
rect 13596 20352 15025 20380
rect 13596 20340 13602 20352
rect 15013 20349 15025 20352
rect 15059 20349 15071 20383
rect 15013 20343 15071 20349
rect 17405 20383 17463 20389
rect 17405 20349 17417 20383
rect 17451 20349 17463 20383
rect 17405 20343 17463 20349
rect 17589 20383 17647 20389
rect 17589 20349 17601 20383
rect 17635 20380 17647 20383
rect 18138 20380 18144 20392
rect 17635 20352 18144 20380
rect 17635 20349 17647 20352
rect 17589 20343 17647 20349
rect 8662 20312 8668 20324
rect 2148 20284 2728 20312
rect 2700 20253 2728 20284
rect 4356 20284 8668 20312
rect 2685 20247 2743 20253
rect 2685 20213 2697 20247
rect 2731 20244 2743 20247
rect 4356 20244 4384 20284
rect 8662 20272 8668 20284
rect 8720 20272 8726 20324
rect 13078 20272 13084 20324
rect 13136 20272 13142 20324
rect 14461 20315 14519 20321
rect 14461 20281 14473 20315
rect 14507 20312 14519 20315
rect 16298 20312 16304 20324
rect 14507 20284 16304 20312
rect 14507 20281 14519 20284
rect 14461 20275 14519 20281
rect 16298 20272 16304 20284
rect 16356 20272 16362 20324
rect 16850 20272 16856 20324
rect 16908 20312 16914 20324
rect 17420 20312 17448 20343
rect 16908 20284 17448 20312
rect 16908 20272 16914 20284
rect 2731 20216 4384 20244
rect 2731 20213 2743 20216
rect 2685 20207 2743 20213
rect 4430 20204 4436 20256
rect 4488 20244 4494 20256
rect 11974 20244 11980 20256
rect 4488 20216 11980 20244
rect 4488 20204 4494 20216
rect 11974 20204 11980 20216
rect 12032 20204 12038 20256
rect 13262 20204 13268 20256
rect 13320 20244 13326 20256
rect 17604 20244 17632 20343
rect 18138 20340 18144 20352
rect 18196 20340 18202 20392
rect 13320 20216 17632 20244
rect 13320 20204 13326 20216
rect 1104 20154 18860 20176
rect 1104 20102 1950 20154
rect 2002 20102 2014 20154
rect 2066 20102 2078 20154
rect 2130 20102 2142 20154
rect 2194 20102 2206 20154
rect 2258 20102 6950 20154
rect 7002 20102 7014 20154
rect 7066 20102 7078 20154
rect 7130 20102 7142 20154
rect 7194 20102 7206 20154
rect 7258 20102 11950 20154
rect 12002 20102 12014 20154
rect 12066 20102 12078 20154
rect 12130 20102 12142 20154
rect 12194 20102 12206 20154
rect 12258 20102 16950 20154
rect 17002 20102 17014 20154
rect 17066 20102 17078 20154
rect 17130 20102 17142 20154
rect 17194 20102 17206 20154
rect 17258 20102 18860 20154
rect 1104 20080 18860 20102
rect 10594 20000 10600 20052
rect 10652 20040 10658 20052
rect 11422 20040 11428 20052
rect 10652 20012 11428 20040
rect 10652 20000 10658 20012
rect 11422 20000 11428 20012
rect 11480 20040 11486 20052
rect 13722 20040 13728 20052
rect 11480 20012 13728 20040
rect 11480 20000 11486 20012
rect 13722 20000 13728 20012
rect 13780 20000 13786 20052
rect 14550 20000 14556 20052
rect 14608 20040 14614 20052
rect 16850 20040 16856 20052
rect 14608 20012 16856 20040
rect 14608 20000 14614 20012
rect 16850 20000 16856 20012
rect 16908 20000 16914 20052
rect 18230 19932 18236 19984
rect 18288 19932 18294 19984
rect 5994 19796 6000 19848
rect 6052 19836 6058 19848
rect 18049 19839 18107 19845
rect 18049 19836 18061 19839
rect 6052 19808 18061 19836
rect 6052 19796 6058 19808
rect 18049 19805 18061 19808
rect 18095 19805 18107 19839
rect 18049 19799 18107 19805
rect 1104 19610 18860 19632
rect 1104 19558 2610 19610
rect 2662 19558 2674 19610
rect 2726 19558 2738 19610
rect 2790 19558 2802 19610
rect 2854 19558 2866 19610
rect 2918 19558 7610 19610
rect 7662 19558 7674 19610
rect 7726 19558 7738 19610
rect 7790 19558 7802 19610
rect 7854 19558 7866 19610
rect 7918 19558 12610 19610
rect 12662 19558 12674 19610
rect 12726 19558 12738 19610
rect 12790 19558 12802 19610
rect 12854 19558 12866 19610
rect 12918 19558 17610 19610
rect 17662 19558 17674 19610
rect 17726 19558 17738 19610
rect 17790 19558 17802 19610
rect 17854 19558 17866 19610
rect 17918 19558 18860 19610
rect 1104 19536 18860 19558
rect 11977 19499 12035 19505
rect 11977 19465 11989 19499
rect 12023 19496 12035 19499
rect 14182 19496 14188 19508
rect 12023 19468 14188 19496
rect 12023 19465 12035 19468
rect 11977 19459 12035 19465
rect 14182 19456 14188 19468
rect 14240 19456 14246 19508
rect 12158 19320 12164 19372
rect 12216 19320 12222 19372
rect 1104 19066 18860 19088
rect 1104 19014 1950 19066
rect 2002 19014 2014 19066
rect 2066 19014 2078 19066
rect 2130 19014 2142 19066
rect 2194 19014 2206 19066
rect 2258 19014 6950 19066
rect 7002 19014 7014 19066
rect 7066 19014 7078 19066
rect 7130 19014 7142 19066
rect 7194 19014 7206 19066
rect 7258 19014 11950 19066
rect 12002 19014 12014 19066
rect 12066 19014 12078 19066
rect 12130 19014 12142 19066
rect 12194 19014 12206 19066
rect 12258 19014 16950 19066
rect 17002 19014 17014 19066
rect 17066 19014 17078 19066
rect 17130 19014 17142 19066
rect 17194 19014 17206 19066
rect 17258 19014 18860 19066
rect 1104 18992 18860 19014
rect 1104 18522 18860 18544
rect 1104 18470 2610 18522
rect 2662 18470 2674 18522
rect 2726 18470 2738 18522
rect 2790 18470 2802 18522
rect 2854 18470 2866 18522
rect 2918 18470 7610 18522
rect 7662 18470 7674 18522
rect 7726 18470 7738 18522
rect 7790 18470 7802 18522
rect 7854 18470 7866 18522
rect 7918 18470 12610 18522
rect 12662 18470 12674 18522
rect 12726 18470 12738 18522
rect 12790 18470 12802 18522
rect 12854 18470 12866 18522
rect 12918 18470 17610 18522
rect 17662 18470 17674 18522
rect 17726 18470 17738 18522
rect 17790 18470 17802 18522
rect 17854 18470 17866 18522
rect 17918 18470 18860 18522
rect 1104 18448 18860 18470
rect 15289 18411 15347 18417
rect 15289 18377 15301 18411
rect 15335 18408 15347 18411
rect 18322 18408 18328 18420
rect 15335 18380 18328 18408
rect 15335 18377 15347 18380
rect 15289 18371 15347 18377
rect 18322 18368 18328 18380
rect 18380 18368 18386 18420
rect 14182 18349 14188 18352
rect 14176 18340 14188 18349
rect 14143 18312 14188 18340
rect 14176 18303 14188 18312
rect 14182 18300 14188 18303
rect 14240 18300 14246 18352
rect 13722 18232 13728 18284
rect 13780 18272 13786 18284
rect 13909 18275 13967 18281
rect 13909 18272 13921 18275
rect 13780 18244 13921 18272
rect 13780 18232 13786 18244
rect 13909 18241 13921 18244
rect 13955 18241 13967 18275
rect 13909 18235 13967 18241
rect 18049 18275 18107 18281
rect 18049 18241 18061 18275
rect 18095 18272 18107 18275
rect 19242 18272 19248 18284
rect 18095 18244 19248 18272
rect 18095 18241 18107 18244
rect 18049 18235 18107 18241
rect 19242 18232 19248 18244
rect 19300 18232 19306 18284
rect 10318 18028 10324 18080
rect 10376 18068 10382 18080
rect 11054 18068 11060 18080
rect 10376 18040 11060 18068
rect 10376 18028 10382 18040
rect 11054 18028 11060 18040
rect 11112 18028 11118 18080
rect 18230 18028 18236 18080
rect 18288 18028 18294 18080
rect 1104 17978 18860 18000
rect 1104 17926 1950 17978
rect 2002 17926 2014 17978
rect 2066 17926 2078 17978
rect 2130 17926 2142 17978
rect 2194 17926 2206 17978
rect 2258 17926 6950 17978
rect 7002 17926 7014 17978
rect 7066 17926 7078 17978
rect 7130 17926 7142 17978
rect 7194 17926 7206 17978
rect 7258 17926 11950 17978
rect 12002 17926 12014 17978
rect 12066 17926 12078 17978
rect 12130 17926 12142 17978
rect 12194 17926 12206 17978
rect 12258 17926 16950 17978
rect 17002 17926 17014 17978
rect 17066 17926 17078 17978
rect 17130 17926 17142 17978
rect 17194 17926 17206 17978
rect 17258 17926 18860 17978
rect 1104 17904 18860 17926
rect 11977 17867 12035 17873
rect 11977 17833 11989 17867
rect 12023 17864 12035 17867
rect 13814 17864 13820 17876
rect 12023 17836 13820 17864
rect 12023 17833 12035 17836
rect 11977 17827 12035 17833
rect 13814 17824 13820 17836
rect 13872 17824 13878 17876
rect 12989 17799 13047 17805
rect 12989 17765 13001 17799
rect 13035 17796 13047 17799
rect 14550 17796 14556 17808
rect 13035 17768 14556 17796
rect 13035 17765 13047 17768
rect 12989 17759 13047 17765
rect 14550 17756 14556 17768
rect 14608 17756 14614 17808
rect 7282 17688 7288 17740
rect 7340 17728 7346 17740
rect 10594 17728 10600 17740
rect 7340 17700 10600 17728
rect 7340 17688 7346 17700
rect 10594 17688 10600 17700
rect 10652 17688 10658 17740
rect 13078 17688 13084 17740
rect 13136 17728 13142 17740
rect 13449 17731 13507 17737
rect 13449 17728 13461 17731
rect 13136 17700 13461 17728
rect 13136 17688 13142 17700
rect 13449 17697 13461 17700
rect 13495 17697 13507 17731
rect 13449 17691 13507 17697
rect 13633 17731 13691 17737
rect 13633 17697 13645 17731
rect 13679 17697 13691 17731
rect 13633 17691 13691 17697
rect 10870 17669 10876 17672
rect 10864 17623 10876 17669
rect 10870 17620 10876 17623
rect 10928 17620 10934 17672
rect 13354 17620 13360 17672
rect 13412 17620 13418 17672
rect 12526 17552 12532 17604
rect 12584 17592 12590 17604
rect 13538 17592 13544 17604
rect 12584 17564 13544 17592
rect 12584 17552 12590 17564
rect 13538 17552 13544 17564
rect 13596 17592 13602 17604
rect 13648 17592 13676 17691
rect 13596 17564 13676 17592
rect 13596 17552 13602 17564
rect 1104 17434 18860 17456
rect 1104 17382 2610 17434
rect 2662 17382 2674 17434
rect 2726 17382 2738 17434
rect 2790 17382 2802 17434
rect 2854 17382 2866 17434
rect 2918 17382 7610 17434
rect 7662 17382 7674 17434
rect 7726 17382 7738 17434
rect 7790 17382 7802 17434
rect 7854 17382 7866 17434
rect 7918 17382 12610 17434
rect 12662 17382 12674 17434
rect 12726 17382 12738 17434
rect 12790 17382 12802 17434
rect 12854 17382 12866 17434
rect 12918 17382 17610 17434
rect 17662 17382 17674 17434
rect 17726 17382 17738 17434
rect 17790 17382 17802 17434
rect 17854 17382 17866 17434
rect 17918 17382 18860 17434
rect 1104 17360 18860 17382
rect 5718 17280 5724 17332
rect 5776 17320 5782 17332
rect 5902 17320 5908 17332
rect 5776 17292 5908 17320
rect 5776 17280 5782 17292
rect 5902 17280 5908 17292
rect 5960 17280 5966 17332
rect 1578 17212 1584 17264
rect 1636 17252 1642 17264
rect 10689 17255 10747 17261
rect 10689 17252 10701 17255
rect 1636 17224 10701 17252
rect 1636 17212 1642 17224
rect 10689 17221 10701 17224
rect 10735 17221 10747 17255
rect 10689 17215 10747 17221
rect 5902 17008 5908 17060
rect 5960 17048 5966 17060
rect 10226 17048 10232 17060
rect 5960 17020 10232 17048
rect 5960 17008 5966 17020
rect 10226 17008 10232 17020
rect 10284 17008 10290 17060
rect 842 16940 848 16992
rect 900 16980 906 16992
rect 10781 16983 10839 16989
rect 10781 16980 10793 16983
rect 900 16952 10793 16980
rect 900 16940 906 16952
rect 10781 16949 10793 16952
rect 10827 16949 10839 16983
rect 10781 16943 10839 16949
rect 1104 16890 18860 16912
rect 1104 16838 1950 16890
rect 2002 16838 2014 16890
rect 2066 16838 2078 16890
rect 2130 16838 2142 16890
rect 2194 16838 2206 16890
rect 2258 16838 6950 16890
rect 7002 16838 7014 16890
rect 7066 16838 7078 16890
rect 7130 16838 7142 16890
rect 7194 16838 7206 16890
rect 7258 16838 11950 16890
rect 12002 16838 12014 16890
rect 12066 16838 12078 16890
rect 12130 16838 12142 16890
rect 12194 16838 12206 16890
rect 12258 16838 16950 16890
rect 17002 16838 17014 16890
rect 17066 16838 17078 16890
rect 17130 16838 17142 16890
rect 17194 16838 17206 16890
rect 17258 16838 18860 16890
rect 1104 16816 18860 16838
rect 7282 16776 7288 16788
rect 7116 16748 7288 16776
rect 5534 16600 5540 16652
rect 5592 16640 5598 16652
rect 7116 16649 7144 16748
rect 7282 16736 7288 16748
rect 7340 16736 7346 16788
rect 17954 16736 17960 16788
rect 18012 16736 18018 16788
rect 5997 16643 6055 16649
rect 5997 16640 6009 16643
rect 5592 16612 6009 16640
rect 5592 16600 5598 16612
rect 5997 16609 6009 16612
rect 6043 16609 6055 16643
rect 5997 16603 6055 16609
rect 7101 16643 7159 16649
rect 7101 16609 7113 16643
rect 7147 16609 7159 16643
rect 7101 16603 7159 16609
rect 5813 16575 5871 16581
rect 5813 16541 5825 16575
rect 5859 16572 5871 16575
rect 5859 16544 12434 16572
rect 5859 16541 5871 16544
rect 5813 16535 5871 16541
rect 750 16464 756 16516
rect 808 16504 814 16516
rect 7346 16507 7404 16513
rect 7346 16504 7358 16507
rect 808 16476 7358 16504
rect 808 16464 814 16476
rect 7346 16473 7358 16476
rect 7392 16473 7404 16507
rect 12406 16504 12434 16544
rect 13446 16532 13452 16584
rect 13504 16572 13510 16584
rect 17865 16575 17923 16581
rect 17865 16572 17877 16575
rect 13504 16544 17877 16572
rect 13504 16532 13510 16544
rect 17865 16541 17877 16544
rect 17911 16541 17923 16575
rect 17865 16535 17923 16541
rect 14734 16504 14740 16516
rect 12406 16476 14740 16504
rect 7346 16467 7404 16473
rect 14734 16464 14740 16476
rect 14792 16464 14798 16516
rect 658 16396 664 16448
rect 716 16436 722 16448
rect 5445 16439 5503 16445
rect 5445 16436 5457 16439
rect 716 16408 5457 16436
rect 716 16396 722 16408
rect 5445 16405 5457 16408
rect 5491 16405 5503 16439
rect 5445 16399 5503 16405
rect 5902 16396 5908 16448
rect 5960 16396 5966 16448
rect 8478 16396 8484 16448
rect 8536 16396 8542 16448
rect 1104 16346 18860 16368
rect 1104 16294 2610 16346
rect 2662 16294 2674 16346
rect 2726 16294 2738 16346
rect 2790 16294 2802 16346
rect 2854 16294 2866 16346
rect 2918 16294 7610 16346
rect 7662 16294 7674 16346
rect 7726 16294 7738 16346
rect 7790 16294 7802 16346
rect 7854 16294 7866 16346
rect 7918 16294 12610 16346
rect 12662 16294 12674 16346
rect 12726 16294 12738 16346
rect 12790 16294 12802 16346
rect 12854 16294 12866 16346
rect 12918 16294 17610 16346
rect 17662 16294 17674 16346
rect 17726 16294 17738 16346
rect 17790 16294 17802 16346
rect 17854 16294 17866 16346
rect 17918 16294 18860 16346
rect 1104 16272 18860 16294
rect 7009 16235 7067 16241
rect 7009 16201 7021 16235
rect 7055 16232 7067 16235
rect 7377 16235 7435 16241
rect 7377 16232 7389 16235
rect 7055 16204 7389 16232
rect 7055 16201 7067 16204
rect 7009 16195 7067 16201
rect 7377 16201 7389 16204
rect 7423 16232 7435 16235
rect 7745 16235 7803 16241
rect 7745 16232 7757 16235
rect 7423 16204 7757 16232
rect 7423 16201 7435 16204
rect 7377 16195 7435 16201
rect 7745 16201 7757 16204
rect 7791 16232 7803 16235
rect 8205 16235 8263 16241
rect 8205 16232 8217 16235
rect 7791 16204 8217 16232
rect 7791 16201 7803 16204
rect 7745 16195 7803 16201
rect 8205 16201 8217 16204
rect 8251 16232 8263 16235
rect 8665 16235 8723 16241
rect 8665 16232 8677 16235
rect 8251 16204 8677 16232
rect 8251 16201 8263 16204
rect 8205 16195 8263 16201
rect 8665 16201 8677 16204
rect 8711 16232 8723 16235
rect 9030 16232 9036 16244
rect 8711 16204 9036 16232
rect 8711 16201 8723 16204
rect 8665 16195 8723 16201
rect 9030 16192 9036 16204
rect 9088 16192 9094 16244
rect 9309 16235 9367 16241
rect 9309 16201 9321 16235
rect 9355 16232 9367 16235
rect 9766 16232 9772 16244
rect 9355 16204 9772 16232
rect 9355 16201 9367 16204
rect 9309 16195 9367 16201
rect 9766 16192 9772 16204
rect 9824 16192 9830 16244
rect 18230 16192 18236 16244
rect 18288 16192 18294 16244
rect 3510 16124 3516 16176
rect 3568 16164 3574 16176
rect 9217 16167 9275 16173
rect 9217 16164 9229 16167
rect 3568 16136 9229 16164
rect 3568 16124 3574 16136
rect 9217 16133 9229 16136
rect 9263 16133 9275 16167
rect 9217 16127 9275 16133
rect 1762 16056 1768 16108
rect 1820 16096 1826 16108
rect 8021 16099 8079 16105
rect 8021 16096 8033 16099
rect 1820 16068 8033 16096
rect 1820 16056 1826 16068
rect 8021 16065 8033 16068
rect 8067 16065 8079 16099
rect 8021 16059 8079 16065
rect 10962 16056 10968 16108
rect 11020 16096 11026 16108
rect 18049 16099 18107 16105
rect 18049 16096 18061 16099
rect 11020 16068 18061 16096
rect 11020 16056 11026 16068
rect 18049 16065 18061 16068
rect 18095 16065 18107 16099
rect 18049 16059 18107 16065
rect 7282 15988 7288 16040
rect 7340 16028 7346 16040
rect 8294 16028 8300 16040
rect 7340 16000 8300 16028
rect 7340 15988 7346 16000
rect 8294 15988 8300 16000
rect 8352 15988 8358 16040
rect 1104 15802 18860 15824
rect 1104 15750 1950 15802
rect 2002 15750 2014 15802
rect 2066 15750 2078 15802
rect 2130 15750 2142 15802
rect 2194 15750 2206 15802
rect 2258 15750 6950 15802
rect 7002 15750 7014 15802
rect 7066 15750 7078 15802
rect 7130 15750 7142 15802
rect 7194 15750 7206 15802
rect 7258 15750 11950 15802
rect 12002 15750 12014 15802
rect 12066 15750 12078 15802
rect 12130 15750 12142 15802
rect 12194 15750 12206 15802
rect 12258 15750 16950 15802
rect 17002 15750 17014 15802
rect 17066 15750 17078 15802
rect 17130 15750 17142 15802
rect 17194 15750 17206 15802
rect 17258 15750 18860 15802
rect 1104 15728 18860 15750
rect 8665 15691 8723 15697
rect 8665 15657 8677 15691
rect 8711 15688 8723 15691
rect 9766 15688 9772 15700
rect 8711 15660 9772 15688
rect 8711 15657 8723 15660
rect 8665 15651 8723 15657
rect 9766 15648 9772 15660
rect 9824 15648 9830 15700
rect 11790 15648 11796 15700
rect 11848 15688 11854 15700
rect 11885 15691 11943 15697
rect 11885 15688 11897 15691
rect 11848 15660 11897 15688
rect 11848 15648 11854 15660
rect 11885 15657 11897 15660
rect 11931 15657 11943 15691
rect 11885 15651 11943 15657
rect 9490 15580 9496 15632
rect 9548 15620 9554 15632
rect 12529 15623 12587 15629
rect 12529 15620 12541 15623
rect 9548 15592 12541 15620
rect 9548 15580 9554 15592
rect 12529 15589 12541 15592
rect 12575 15589 12587 15623
rect 12529 15583 12587 15589
rect 12986 15512 12992 15564
rect 13044 15512 13050 15564
rect 13078 15512 13084 15564
rect 13136 15552 13142 15564
rect 13630 15552 13636 15564
rect 13136 15524 13636 15552
rect 13136 15512 13142 15524
rect 13630 15512 13636 15524
rect 13688 15512 13694 15564
rect 1026 15444 1032 15496
rect 1084 15484 1090 15496
rect 12069 15487 12127 15493
rect 12069 15484 12081 15487
rect 1084 15456 12081 15484
rect 1084 15444 1090 15456
rect 12069 15453 12081 15456
rect 12115 15453 12127 15487
rect 12069 15447 12127 15453
rect 16850 15444 16856 15496
rect 16908 15444 16914 15496
rect 16574 15376 16580 15428
rect 16632 15416 16638 15428
rect 17098 15419 17156 15425
rect 17098 15416 17110 15419
rect 16632 15388 17110 15416
rect 16632 15376 16638 15388
rect 17098 15385 17110 15388
rect 17144 15385 17156 15419
rect 19794 15416 19800 15428
rect 17098 15379 17156 15385
rect 18156 15388 19800 15416
rect 11422 15308 11428 15360
rect 11480 15348 11486 15360
rect 12897 15351 12955 15357
rect 12897 15348 12909 15351
rect 11480 15320 12909 15348
rect 11480 15308 11486 15320
rect 12897 15317 12909 15320
rect 12943 15348 12955 15351
rect 18156 15348 18184 15388
rect 19794 15376 19800 15388
rect 19852 15376 19858 15428
rect 12943 15320 18184 15348
rect 12943 15317 12955 15320
rect 12897 15311 12955 15317
rect 18230 15308 18236 15360
rect 18288 15348 18294 15360
rect 18506 15348 18512 15360
rect 18288 15320 18512 15348
rect 18288 15308 18294 15320
rect 18506 15308 18512 15320
rect 18564 15308 18570 15360
rect 1104 15258 18860 15280
rect 1104 15206 2610 15258
rect 2662 15206 2674 15258
rect 2726 15206 2738 15258
rect 2790 15206 2802 15258
rect 2854 15206 2866 15258
rect 2918 15206 7610 15258
rect 7662 15206 7674 15258
rect 7726 15206 7738 15258
rect 7790 15206 7802 15258
rect 7854 15206 7866 15258
rect 7918 15206 12610 15258
rect 12662 15206 12674 15258
rect 12726 15206 12738 15258
rect 12790 15206 12802 15258
rect 12854 15206 12866 15258
rect 12918 15206 17610 15258
rect 17662 15206 17674 15258
rect 17726 15206 17738 15258
rect 17790 15206 17802 15258
rect 17854 15206 17866 15258
rect 17918 15206 18860 15258
rect 1104 15184 18860 15206
rect 934 15104 940 15156
rect 992 15144 998 15156
rect 1857 15147 1915 15153
rect 1857 15144 1869 15147
rect 992 15116 1869 15144
rect 992 15104 998 15116
rect 1857 15113 1869 15116
rect 1903 15144 1915 15147
rect 2409 15147 2467 15153
rect 2409 15144 2421 15147
rect 1903 15116 2421 15144
rect 1903 15113 1915 15116
rect 1857 15107 1915 15113
rect 2409 15113 2421 15116
rect 2455 15113 2467 15147
rect 2409 15107 2467 15113
rect 14918 15104 14924 15156
rect 14976 15144 14982 15156
rect 18141 15147 18199 15153
rect 18141 15144 18153 15147
rect 14976 15116 18153 15144
rect 14976 15104 14982 15116
rect 18141 15113 18153 15116
rect 18187 15113 18199 15147
rect 18141 15107 18199 15113
rect 2314 15036 2320 15088
rect 2372 15036 2378 15088
rect 15838 15036 15844 15088
rect 15896 15076 15902 15088
rect 17957 15079 18015 15085
rect 17957 15076 17969 15079
rect 15896 15048 17969 15076
rect 15896 15036 15902 15048
rect 17957 15045 17969 15048
rect 18003 15045 18015 15079
rect 17957 15039 18015 15045
rect 15010 14968 15016 15020
rect 15068 15008 15074 15020
rect 18233 15011 18291 15017
rect 18233 15008 18245 15011
rect 15068 14980 18245 15008
rect 15068 14968 15074 14980
rect 18233 14977 18245 14980
rect 18279 14977 18291 15011
rect 18233 14971 18291 14977
rect 17678 14832 17684 14884
rect 17736 14832 17742 14884
rect 1104 14714 18860 14736
rect 1104 14662 1950 14714
rect 2002 14662 2014 14714
rect 2066 14662 2078 14714
rect 2130 14662 2142 14714
rect 2194 14662 2206 14714
rect 2258 14662 6950 14714
rect 7002 14662 7014 14714
rect 7066 14662 7078 14714
rect 7130 14662 7142 14714
rect 7194 14662 7206 14714
rect 7258 14662 11950 14714
rect 12002 14662 12014 14714
rect 12066 14662 12078 14714
rect 12130 14662 12142 14714
rect 12194 14662 12206 14714
rect 12258 14662 16950 14714
rect 17002 14662 17014 14714
rect 17066 14662 17078 14714
rect 17130 14662 17142 14714
rect 17194 14662 17206 14714
rect 17258 14662 18860 14714
rect 1104 14640 18860 14662
rect 7374 14560 7380 14612
rect 7432 14600 7438 14612
rect 7653 14603 7711 14609
rect 7653 14600 7665 14603
rect 7432 14572 7665 14600
rect 7432 14560 7438 14572
rect 7653 14569 7665 14572
rect 7699 14569 7711 14603
rect 7653 14563 7711 14569
rect 13170 14560 13176 14612
rect 13228 14600 13234 14612
rect 16853 14603 16911 14609
rect 16853 14600 16865 14603
rect 13228 14572 16865 14600
rect 13228 14560 13234 14572
rect 16853 14569 16865 14572
rect 16899 14569 16911 14603
rect 16853 14563 16911 14569
rect 1118 14492 1124 14544
rect 1176 14532 1182 14544
rect 8573 14535 8631 14541
rect 8573 14532 8585 14535
rect 1176 14504 8585 14532
rect 1176 14492 1182 14504
rect 8573 14501 8585 14504
rect 8619 14501 8631 14535
rect 8573 14495 8631 14501
rect 7834 14356 7840 14408
rect 7892 14356 7898 14408
rect 8386 14356 8392 14408
rect 8444 14356 8450 14408
rect 15470 14356 15476 14408
rect 15528 14356 15534 14408
rect 18049 14399 18107 14405
rect 18049 14365 18061 14399
rect 18095 14396 18107 14399
rect 19518 14396 19524 14408
rect 18095 14368 19524 14396
rect 18095 14365 18107 14368
rect 18049 14359 18107 14365
rect 19518 14356 19524 14368
rect 19576 14356 19582 14408
rect 11330 14288 11336 14340
rect 11388 14328 11394 14340
rect 15718 14331 15776 14337
rect 15718 14328 15730 14331
rect 11388 14300 15730 14328
rect 11388 14288 11394 14300
rect 15718 14297 15730 14300
rect 15764 14297 15776 14331
rect 15718 14291 15776 14297
rect 18230 14220 18236 14272
rect 18288 14220 18294 14272
rect 1104 14170 18860 14192
rect 1104 14118 2610 14170
rect 2662 14118 2674 14170
rect 2726 14118 2738 14170
rect 2790 14118 2802 14170
rect 2854 14118 2866 14170
rect 2918 14118 7610 14170
rect 7662 14118 7674 14170
rect 7726 14118 7738 14170
rect 7790 14118 7802 14170
rect 7854 14118 7866 14170
rect 7918 14118 12610 14170
rect 12662 14118 12674 14170
rect 12726 14118 12738 14170
rect 12790 14118 12802 14170
rect 12854 14118 12866 14170
rect 12918 14118 17610 14170
rect 17662 14118 17674 14170
rect 17726 14118 17738 14170
rect 17790 14118 17802 14170
rect 17854 14118 17866 14170
rect 17918 14118 18860 14170
rect 1104 14096 18860 14118
rect 6549 14059 6607 14065
rect 6549 14025 6561 14059
rect 6595 14025 6607 14059
rect 6549 14019 6607 14025
rect 6564 13988 6592 14019
rect 11054 14016 11060 14068
rect 11112 14056 11118 14068
rect 16114 14056 16120 14068
rect 11112 14028 16120 14056
rect 11112 14016 11118 14028
rect 16114 14016 16120 14028
rect 16172 14016 16178 14068
rect 11146 13988 11152 14000
rect 6564 13960 11152 13988
rect 11146 13948 11152 13960
rect 11204 13948 11210 14000
rect 6733 13923 6791 13929
rect 6733 13889 6745 13923
rect 6779 13920 6791 13923
rect 11238 13920 11244 13932
rect 6779 13892 11244 13920
rect 6779 13889 6791 13892
rect 6733 13883 6791 13889
rect 11238 13880 11244 13892
rect 11296 13880 11302 13932
rect 10594 13744 10600 13796
rect 10652 13784 10658 13796
rect 10778 13784 10784 13796
rect 10652 13756 10784 13784
rect 10652 13744 10658 13756
rect 10778 13744 10784 13756
rect 10836 13784 10842 13796
rect 15470 13784 15476 13796
rect 10836 13756 15476 13784
rect 10836 13744 10842 13756
rect 15470 13744 15476 13756
rect 15528 13784 15534 13796
rect 16850 13784 16856 13796
rect 15528 13756 16856 13784
rect 15528 13744 15534 13756
rect 16850 13744 16856 13756
rect 16908 13744 16914 13796
rect 1104 13626 18860 13648
rect 1104 13574 1950 13626
rect 2002 13574 2014 13626
rect 2066 13574 2078 13626
rect 2130 13574 2142 13626
rect 2194 13574 2206 13626
rect 2258 13574 6950 13626
rect 7002 13574 7014 13626
rect 7066 13574 7078 13626
rect 7130 13574 7142 13626
rect 7194 13574 7206 13626
rect 7258 13574 11950 13626
rect 12002 13574 12014 13626
rect 12066 13574 12078 13626
rect 12130 13574 12142 13626
rect 12194 13574 12206 13626
rect 12258 13574 16950 13626
rect 17002 13574 17014 13626
rect 17066 13574 17078 13626
rect 17130 13574 17142 13626
rect 17194 13574 17206 13626
rect 17258 13574 18860 13626
rect 1104 13552 18860 13574
rect 8570 13472 8576 13524
rect 8628 13512 8634 13524
rect 16117 13515 16175 13521
rect 16117 13512 16129 13515
rect 8628 13484 16129 13512
rect 8628 13472 8634 13484
rect 16117 13481 16129 13484
rect 16163 13481 16175 13515
rect 16117 13475 16175 13481
rect 16390 13268 16396 13320
rect 16448 13268 16454 13320
rect 7282 13200 7288 13252
rect 7340 13240 7346 13252
rect 16669 13243 16727 13249
rect 16669 13240 16681 13243
rect 7340 13212 16681 13240
rect 7340 13200 7346 13212
rect 16669 13209 16681 13212
rect 16715 13209 16727 13243
rect 16669 13203 16727 13209
rect 16574 13132 16580 13184
rect 16632 13132 16638 13184
rect 1104 13082 18860 13104
rect 1104 13030 2610 13082
rect 2662 13030 2674 13082
rect 2726 13030 2738 13082
rect 2790 13030 2802 13082
rect 2854 13030 2866 13082
rect 2918 13030 7610 13082
rect 7662 13030 7674 13082
rect 7726 13030 7738 13082
rect 7790 13030 7802 13082
rect 7854 13030 7866 13082
rect 7918 13030 12610 13082
rect 12662 13030 12674 13082
rect 12726 13030 12738 13082
rect 12790 13030 12802 13082
rect 12854 13030 12866 13082
rect 12918 13030 17610 13082
rect 17662 13030 17674 13082
rect 17726 13030 17738 13082
rect 17790 13030 17802 13082
rect 17854 13030 17866 13082
rect 17918 13030 18860 13082
rect 1104 13008 18860 13030
rect 4525 12971 4583 12977
rect 4525 12937 4537 12971
rect 4571 12968 4583 12971
rect 11054 12968 11060 12980
rect 4571 12940 11060 12968
rect 4571 12937 4583 12940
rect 4525 12931 4583 12937
rect 11054 12928 11060 12940
rect 11112 12928 11118 12980
rect 11698 12928 11704 12980
rect 11756 12968 11762 12980
rect 18046 12968 18052 12980
rect 11756 12940 18052 12968
rect 11756 12928 11762 12940
rect 18046 12928 18052 12940
rect 18104 12968 18110 12980
rect 18233 12971 18291 12977
rect 18233 12968 18245 12971
rect 18104 12940 18245 12968
rect 18104 12928 18110 12940
rect 18233 12937 18245 12940
rect 18279 12937 18291 12971
rect 18233 12931 18291 12937
rect 2501 12903 2559 12909
rect 2501 12869 2513 12903
rect 2547 12900 2559 12903
rect 2869 12903 2927 12909
rect 2869 12900 2881 12903
rect 2547 12872 2881 12900
rect 2547 12869 2559 12872
rect 2501 12863 2559 12869
rect 2869 12869 2881 12872
rect 2915 12900 2927 12903
rect 3412 12903 3470 12909
rect 3412 12900 3424 12903
rect 2915 12872 3424 12900
rect 2915 12869 2927 12872
rect 2869 12863 2927 12869
rect 3412 12869 3424 12872
rect 3458 12900 3470 12903
rect 4985 12903 5043 12909
rect 4985 12900 4997 12903
rect 3458 12872 4997 12900
rect 3458 12869 3470 12872
rect 3412 12863 3470 12869
rect 4985 12869 4997 12872
rect 5031 12900 5043 12903
rect 5258 12900 5264 12912
rect 5031 12872 5264 12900
rect 5031 12869 5043 12872
rect 4985 12863 5043 12869
rect 5258 12860 5264 12872
rect 5316 12860 5322 12912
rect 17120 12903 17178 12909
rect 17120 12869 17132 12903
rect 17166 12900 17178 12903
rect 17310 12900 17316 12912
rect 17166 12872 17316 12900
rect 17166 12869 17178 12872
rect 17120 12863 17178 12869
rect 17310 12860 17316 12872
rect 17368 12860 17374 12912
rect 16850 12792 16856 12844
rect 16908 12792 16914 12844
rect 3145 12767 3203 12773
rect 3145 12733 3157 12767
rect 3191 12733 3203 12767
rect 3145 12727 3203 12733
rect 3160 12628 3188 12727
rect 3878 12628 3884 12640
rect 3160 12600 3884 12628
rect 3878 12588 3884 12600
rect 3936 12588 3942 12640
rect 1104 12538 18860 12560
rect 1104 12486 1950 12538
rect 2002 12486 2014 12538
rect 2066 12486 2078 12538
rect 2130 12486 2142 12538
rect 2194 12486 2206 12538
rect 2258 12486 6950 12538
rect 7002 12486 7014 12538
rect 7066 12486 7078 12538
rect 7130 12486 7142 12538
rect 7194 12486 7206 12538
rect 7258 12486 11950 12538
rect 12002 12486 12014 12538
rect 12066 12486 12078 12538
rect 12130 12486 12142 12538
rect 12194 12486 12206 12538
rect 12258 12486 16950 12538
rect 17002 12486 17014 12538
rect 17066 12486 17078 12538
rect 17130 12486 17142 12538
rect 17194 12486 17206 12538
rect 17258 12486 18860 12538
rect 1104 12464 18860 12486
rect 7374 12384 7380 12436
rect 7432 12384 7438 12436
rect 12158 12316 12164 12368
rect 12216 12316 12222 12368
rect 18230 12316 18236 12368
rect 18288 12316 18294 12368
rect 8573 12291 8631 12297
rect 8573 12257 8585 12291
rect 8619 12288 8631 12291
rect 9125 12291 9183 12297
rect 9125 12288 9137 12291
rect 8619 12260 9137 12288
rect 8619 12257 8631 12260
rect 8573 12251 8631 12257
rect 9125 12257 9137 12260
rect 9171 12288 9183 12291
rect 9171 12260 10364 12288
rect 9171 12257 9183 12260
rect 9125 12251 9183 12257
rect 3878 12180 3884 12232
rect 3936 12220 3942 12232
rect 5997 12223 6055 12229
rect 5997 12220 6009 12223
rect 3936 12192 6009 12220
rect 3936 12180 3942 12192
rect 5997 12189 6009 12192
rect 6043 12189 6055 12223
rect 8938 12220 8944 12232
rect 5997 12183 6055 12189
rect 6886 12192 8944 12220
rect 6264 12155 6322 12161
rect 6264 12121 6276 12155
rect 6310 12152 6322 12155
rect 6886 12152 6914 12192
rect 8938 12180 8944 12192
rect 8996 12180 9002 12232
rect 10336 12229 10364 12260
rect 9401 12223 9459 12229
rect 9401 12189 9413 12223
rect 9447 12189 9459 12223
rect 9401 12183 9459 12189
rect 10321 12223 10379 12229
rect 10321 12189 10333 12223
rect 10367 12220 10379 12223
rect 10686 12220 10692 12232
rect 10367 12192 10692 12220
rect 10367 12189 10379 12192
rect 10321 12183 10379 12189
rect 9416 12152 9444 12183
rect 10686 12180 10692 12192
rect 10744 12180 10750 12232
rect 10778 12180 10784 12232
rect 10836 12180 10842 12232
rect 11054 12229 11060 12232
rect 11048 12183 11060 12229
rect 11054 12180 11060 12183
rect 11112 12180 11118 12232
rect 18046 12180 18052 12232
rect 18104 12180 18110 12232
rect 6310 12124 6914 12152
rect 7300 12124 9444 12152
rect 6310 12121 6322 12124
rect 6264 12115 6322 12121
rect 1486 12044 1492 12096
rect 1544 12084 1550 12096
rect 7300 12084 7328 12124
rect 1544 12056 7328 12084
rect 1544 12044 1550 12056
rect 1104 11994 18860 12016
rect 1104 11942 2610 11994
rect 2662 11942 2674 11994
rect 2726 11942 2738 11994
rect 2790 11942 2802 11994
rect 2854 11942 2866 11994
rect 2918 11942 7610 11994
rect 7662 11942 7674 11994
rect 7726 11942 7738 11994
rect 7790 11942 7802 11994
rect 7854 11942 7866 11994
rect 7918 11942 12610 11994
rect 12662 11942 12674 11994
rect 12726 11942 12738 11994
rect 12790 11942 12802 11994
rect 12854 11942 12866 11994
rect 12918 11942 17610 11994
rect 17662 11942 17674 11994
rect 17726 11942 17738 11994
rect 17790 11942 17802 11994
rect 17854 11942 17866 11994
rect 17918 11942 18860 11994
rect 1104 11920 18860 11942
rect 4798 11772 4804 11824
rect 4856 11812 4862 11824
rect 6270 11812 6276 11824
rect 4856 11784 6276 11812
rect 4856 11772 4862 11784
rect 6270 11772 6276 11784
rect 6328 11772 6334 11824
rect 3142 11500 3148 11552
rect 3200 11540 3206 11552
rect 5718 11540 5724 11552
rect 3200 11512 5724 11540
rect 3200 11500 3206 11512
rect 5718 11500 5724 11512
rect 5776 11500 5782 11552
rect 1104 11450 18860 11472
rect 1104 11398 1950 11450
rect 2002 11398 2014 11450
rect 2066 11398 2078 11450
rect 2130 11398 2142 11450
rect 2194 11398 2206 11450
rect 2258 11398 6950 11450
rect 7002 11398 7014 11450
rect 7066 11398 7078 11450
rect 7130 11398 7142 11450
rect 7194 11398 7206 11450
rect 7258 11398 11950 11450
rect 12002 11398 12014 11450
rect 12066 11398 12078 11450
rect 12130 11398 12142 11450
rect 12194 11398 12206 11450
rect 12258 11398 16950 11450
rect 17002 11398 17014 11450
rect 17066 11398 17078 11450
rect 17130 11398 17142 11450
rect 17194 11398 17206 11450
rect 17258 11398 18860 11450
rect 1104 11376 18860 11398
rect 14553 11203 14611 11209
rect 14553 11200 14565 11203
rect 12406 11172 14565 11200
rect 6638 11092 6644 11144
rect 6696 11132 6702 11144
rect 12406 11132 12434 11172
rect 14553 11169 14565 11172
rect 14599 11200 14611 11203
rect 15194 11200 15200 11212
rect 14599 11172 15200 11200
rect 14599 11169 14611 11172
rect 14553 11163 14611 11169
rect 15194 11160 15200 11172
rect 15252 11160 15258 11212
rect 15286 11160 15292 11212
rect 15344 11160 15350 11212
rect 6696 11104 12434 11132
rect 14645 11135 14703 11141
rect 6696 11092 6702 11104
rect 14645 11101 14657 11135
rect 14691 11101 14703 11135
rect 14645 11095 14703 11101
rect 14660 11064 14688 11095
rect 14826 11092 14832 11144
rect 14884 11092 14890 11144
rect 16022 11064 16028 11076
rect 14660 11036 16028 11064
rect 16022 11024 16028 11036
rect 16080 11024 16086 11076
rect 1104 10906 18860 10928
rect 1104 10854 2610 10906
rect 2662 10854 2674 10906
rect 2726 10854 2738 10906
rect 2790 10854 2802 10906
rect 2854 10854 2866 10906
rect 2918 10854 7610 10906
rect 7662 10854 7674 10906
rect 7726 10854 7738 10906
rect 7790 10854 7802 10906
rect 7854 10854 7866 10906
rect 7918 10854 12610 10906
rect 12662 10854 12674 10906
rect 12726 10854 12738 10906
rect 12790 10854 12802 10906
rect 12854 10854 12866 10906
rect 12918 10854 17610 10906
rect 17662 10854 17674 10906
rect 17726 10854 17738 10906
rect 17790 10854 17802 10906
rect 17854 10854 17866 10906
rect 17918 10854 18860 10906
rect 1104 10832 18860 10854
rect 1854 10752 1860 10804
rect 1912 10792 1918 10804
rect 2685 10795 2743 10801
rect 2685 10792 2697 10795
rect 1912 10764 2697 10792
rect 1912 10752 1918 10764
rect 2685 10761 2697 10764
rect 2731 10792 2743 10795
rect 3142 10792 3148 10804
rect 2731 10764 3148 10792
rect 2731 10761 2743 10764
rect 2685 10755 2743 10761
rect 3142 10752 3148 10764
rect 3200 10752 3206 10804
rect 2225 10727 2283 10733
rect 2225 10693 2237 10727
rect 2271 10724 2283 10727
rect 2590 10724 2596 10736
rect 2271 10696 2596 10724
rect 2271 10693 2283 10696
rect 2225 10687 2283 10693
rect 2590 10684 2596 10696
rect 2648 10684 2654 10736
rect 15194 10616 15200 10668
rect 15252 10656 15258 10668
rect 18049 10659 18107 10665
rect 18049 10656 18061 10659
rect 15252 10628 18061 10656
rect 15252 10616 15258 10628
rect 18049 10625 18061 10628
rect 18095 10625 18107 10659
rect 18049 10619 18107 10625
rect 4890 10412 4896 10464
rect 4948 10452 4954 10464
rect 14366 10452 14372 10464
rect 4948 10424 14372 10452
rect 4948 10412 4954 10424
rect 14366 10412 14372 10424
rect 14424 10412 14430 10464
rect 18230 10412 18236 10464
rect 18288 10412 18294 10464
rect 1104 10362 18860 10384
rect 1104 10310 1950 10362
rect 2002 10310 2014 10362
rect 2066 10310 2078 10362
rect 2130 10310 2142 10362
rect 2194 10310 2206 10362
rect 2258 10310 6950 10362
rect 7002 10310 7014 10362
rect 7066 10310 7078 10362
rect 7130 10310 7142 10362
rect 7194 10310 7206 10362
rect 7258 10310 11950 10362
rect 12002 10310 12014 10362
rect 12066 10310 12078 10362
rect 12130 10310 12142 10362
rect 12194 10310 12206 10362
rect 12258 10310 16950 10362
rect 17002 10310 17014 10362
rect 17066 10310 17078 10362
rect 17130 10310 17142 10362
rect 17194 10310 17206 10362
rect 17258 10310 18860 10362
rect 1104 10288 18860 10310
rect 1854 10208 1860 10260
rect 1912 10208 1918 10260
rect 6914 10208 6920 10260
rect 6972 10248 6978 10260
rect 8202 10248 8208 10260
rect 6972 10220 8208 10248
rect 6972 10208 6978 10220
rect 8202 10208 8208 10220
rect 8260 10208 8266 10260
rect 10502 10180 10508 10192
rect 6886 10152 10508 10180
rect 6886 10112 6914 10152
rect 10502 10140 10508 10152
rect 10560 10140 10566 10192
rect 7374 10112 7380 10124
rect 5184 10084 6914 10112
rect 7024 10084 7380 10112
rect 5184 10053 5212 10084
rect 5169 10047 5227 10053
rect 5169 10013 5181 10047
rect 5215 10013 5227 10047
rect 5169 10007 5227 10013
rect 6914 10004 6920 10056
rect 6972 10004 6978 10056
rect 7024 10053 7052 10084
rect 7374 10072 7380 10084
rect 7432 10072 7438 10124
rect 7653 10115 7711 10121
rect 7653 10081 7665 10115
rect 7699 10112 7711 10115
rect 7926 10112 7932 10124
rect 7699 10084 7932 10112
rect 7699 10081 7711 10084
rect 7653 10075 7711 10081
rect 7926 10072 7932 10084
rect 7984 10072 7990 10124
rect 7009 10047 7067 10053
rect 7009 10013 7021 10047
rect 7055 10013 7067 10047
rect 7009 10007 7067 10013
rect 7193 10047 7251 10053
rect 7193 10013 7205 10047
rect 7239 10044 7251 10047
rect 7282 10044 7288 10056
rect 7239 10016 7288 10044
rect 7239 10013 7251 10016
rect 7193 10007 7251 10013
rect 7282 10004 7288 10016
rect 7340 10004 7346 10056
rect 15930 9976 15936 9988
rect 5000 9948 15936 9976
rect 5000 9917 5028 9948
rect 15930 9936 15936 9948
rect 15988 9936 15994 9988
rect 4985 9911 5043 9917
rect 4985 9877 4997 9911
rect 5031 9877 5043 9911
rect 4985 9871 5043 9877
rect 5997 9911 6055 9917
rect 5997 9877 6009 9911
rect 6043 9908 6055 9911
rect 6273 9911 6331 9917
rect 6273 9908 6285 9911
rect 6043 9880 6285 9908
rect 6043 9877 6055 9880
rect 5997 9871 6055 9877
rect 6273 9877 6285 9880
rect 6319 9908 6331 9911
rect 7926 9908 7932 9920
rect 6319 9880 7932 9908
rect 6319 9877 6331 9880
rect 6273 9871 6331 9877
rect 7926 9868 7932 9880
rect 7984 9868 7990 9920
rect 1104 9818 18860 9840
rect 1104 9766 2610 9818
rect 2662 9766 2674 9818
rect 2726 9766 2738 9818
rect 2790 9766 2802 9818
rect 2854 9766 2866 9818
rect 2918 9766 7610 9818
rect 7662 9766 7674 9818
rect 7726 9766 7738 9818
rect 7790 9766 7802 9818
rect 7854 9766 7866 9818
rect 7918 9766 12610 9818
rect 12662 9766 12674 9818
rect 12726 9766 12738 9818
rect 12790 9766 12802 9818
rect 12854 9766 12866 9818
rect 12918 9766 17610 9818
rect 17662 9766 17674 9818
rect 17726 9766 17738 9818
rect 17790 9766 17802 9818
rect 17854 9766 17866 9818
rect 17918 9766 18860 9818
rect 1104 9744 18860 9766
rect 2314 9596 2320 9648
rect 2372 9636 2378 9648
rect 3878 9636 3884 9648
rect 2372 9608 3884 9636
rect 2372 9596 2378 9608
rect 3878 9596 3884 9608
rect 3936 9636 3942 9648
rect 6181 9639 6239 9645
rect 3936 9608 4292 9636
rect 3936 9596 3942 9608
rect 4264 9580 4292 9608
rect 6181 9605 6193 9639
rect 6227 9636 6239 9639
rect 7469 9639 7527 9645
rect 7469 9636 7481 9639
rect 6227 9608 7481 9636
rect 6227 9605 6239 9608
rect 6181 9599 6239 9605
rect 7469 9605 7481 9608
rect 7515 9605 7527 9639
rect 7469 9599 7527 9605
rect 7561 9639 7619 9645
rect 7561 9605 7573 9639
rect 7607 9636 7619 9639
rect 13078 9636 13084 9648
rect 7607 9608 13084 9636
rect 7607 9605 7619 9608
rect 7561 9599 7619 9605
rect 1765 9571 1823 9577
rect 1765 9537 1777 9571
rect 1811 9568 1823 9571
rect 2133 9571 2191 9577
rect 2133 9568 2145 9571
rect 1811 9540 2145 9568
rect 1811 9537 1823 9540
rect 1765 9531 1823 9537
rect 2133 9537 2145 9540
rect 2179 9568 2191 9571
rect 2501 9571 2559 9577
rect 2501 9568 2513 9571
rect 2179 9540 2513 9568
rect 2179 9537 2191 9540
rect 2133 9531 2191 9537
rect 2501 9537 2513 9540
rect 2547 9568 2559 9571
rect 3993 9571 4051 9577
rect 3993 9568 4005 9571
rect 2547 9540 4005 9568
rect 2547 9537 2559 9540
rect 2501 9531 2559 9537
rect 3993 9537 4005 9540
rect 4039 9568 4051 9571
rect 4039 9540 4200 9568
rect 4039 9537 4051 9540
rect 3993 9531 4051 9537
rect 4172 9500 4200 9540
rect 4246 9528 4252 9580
rect 4304 9528 4310 9580
rect 4617 9571 4675 9577
rect 4617 9537 4629 9571
rect 4663 9568 4675 9571
rect 4985 9571 5043 9577
rect 4985 9568 4997 9571
rect 4663 9540 4997 9568
rect 4663 9537 4675 9540
rect 4617 9531 4675 9537
rect 4985 9537 4997 9540
rect 5031 9568 5043 9571
rect 5353 9571 5411 9577
rect 5353 9568 5365 9571
rect 5031 9540 5365 9568
rect 5031 9537 5043 9540
rect 4985 9531 5043 9537
rect 5353 9537 5365 9540
rect 5399 9568 5411 9571
rect 5534 9568 5540 9580
rect 5399 9540 5540 9568
rect 5399 9537 5411 9540
rect 5353 9531 5411 9537
rect 4632 9500 4660 9531
rect 5534 9528 5540 9540
rect 5592 9568 5598 9580
rect 5721 9571 5779 9577
rect 5721 9568 5733 9571
rect 5592 9540 5733 9568
rect 5592 9528 5598 9540
rect 5721 9537 5733 9540
rect 5767 9568 5779 9571
rect 6638 9568 6644 9580
rect 5767 9540 6644 9568
rect 5767 9537 5779 9540
rect 5721 9531 5779 9537
rect 6638 9528 6644 9540
rect 6696 9528 6702 9580
rect 7484 9568 7512 9599
rect 13078 9596 13084 9608
rect 13136 9596 13142 9648
rect 15378 9568 15384 9580
rect 7484 9540 15384 9568
rect 15378 9528 15384 9540
rect 15436 9528 15442 9580
rect 4172 9472 4660 9500
rect 7469 9503 7527 9509
rect 7469 9469 7481 9503
rect 7515 9469 7527 9503
rect 7469 9463 7527 9469
rect 7006 9392 7012 9444
rect 7064 9392 7070 9444
rect 7484 9432 7512 9463
rect 18138 9432 18144 9444
rect 7484 9404 18144 9432
rect 18138 9392 18144 9404
rect 18196 9392 18202 9444
rect 2869 9367 2927 9373
rect 2869 9333 2881 9367
rect 2915 9364 2927 9367
rect 3970 9364 3976 9376
rect 2915 9336 3976 9364
rect 2915 9333 2927 9336
rect 2869 9327 2927 9333
rect 3970 9324 3976 9336
rect 4028 9324 4034 9376
rect 7926 9324 7932 9376
rect 7984 9364 7990 9376
rect 9582 9364 9588 9376
rect 7984 9336 9588 9364
rect 7984 9324 7990 9336
rect 9582 9324 9588 9336
rect 9640 9324 9646 9376
rect 1104 9274 18860 9296
rect 1104 9222 1950 9274
rect 2002 9222 2014 9274
rect 2066 9222 2078 9274
rect 2130 9222 2142 9274
rect 2194 9222 2206 9274
rect 2258 9222 6950 9274
rect 7002 9222 7014 9274
rect 7066 9222 7078 9274
rect 7130 9222 7142 9274
rect 7194 9222 7206 9274
rect 7258 9222 11950 9274
rect 12002 9222 12014 9274
rect 12066 9222 12078 9274
rect 12130 9222 12142 9274
rect 12194 9222 12206 9274
rect 12258 9222 16950 9274
rect 17002 9222 17014 9274
rect 17066 9222 17078 9274
rect 17130 9222 17142 9274
rect 17194 9222 17206 9274
rect 17258 9222 18860 9274
rect 1104 9200 18860 9222
rect 4157 9163 4215 9169
rect 4157 9129 4169 9163
rect 4203 9160 4215 9163
rect 4525 9163 4583 9169
rect 4525 9160 4537 9163
rect 4203 9132 4537 9160
rect 4203 9129 4215 9132
rect 4157 9123 4215 9129
rect 4525 9129 4537 9132
rect 4571 9160 4583 9163
rect 4893 9163 4951 9169
rect 4893 9160 4905 9163
rect 4571 9132 4905 9160
rect 4571 9129 4583 9132
rect 4525 9123 4583 9129
rect 4893 9129 4905 9132
rect 4939 9160 4951 9163
rect 5534 9160 5540 9172
rect 4939 9132 5540 9160
rect 4939 9129 4951 9132
rect 4893 9123 4951 9129
rect 5534 9120 5540 9132
rect 5592 9120 5598 9172
rect 8021 9163 8079 9169
rect 8021 9129 8033 9163
rect 8067 9160 8079 9163
rect 8110 9160 8116 9172
rect 8067 9132 8116 9160
rect 8067 9129 8079 9132
rect 8021 9123 8079 9129
rect 8110 9120 8116 9132
rect 8168 9120 8174 9172
rect 17402 9120 17408 9172
rect 17460 9160 17466 9172
rect 17681 9163 17739 9169
rect 17681 9160 17693 9163
rect 17460 9132 17693 9160
rect 17460 9120 17466 9132
rect 17681 9129 17693 9132
rect 17727 9129 17739 9163
rect 17681 9123 17739 9129
rect 5721 9027 5779 9033
rect 5721 8993 5733 9027
rect 5767 9024 5779 9027
rect 7466 9024 7472 9036
rect 5767 8996 7472 9024
rect 5767 8993 5779 8996
rect 5721 8987 5779 8993
rect 7466 8984 7472 8996
rect 7524 9024 7530 9036
rect 7926 9024 7932 9036
rect 7524 8996 7932 9024
rect 7524 8984 7530 8996
rect 7926 8984 7932 8996
rect 7984 8984 7990 9036
rect 5169 8959 5227 8965
rect 5169 8925 5181 8959
rect 5215 8956 5227 8959
rect 8110 8956 8116 8968
rect 5215 8928 8116 8956
rect 5215 8925 5227 8928
rect 5169 8919 5227 8925
rect 8110 8916 8116 8928
rect 8168 8916 8174 8968
rect 8202 8916 8208 8968
rect 8260 8916 8266 8968
rect 17696 8956 17724 9123
rect 18049 8959 18107 8965
rect 18049 8956 18061 8959
rect 17696 8928 18061 8956
rect 18049 8925 18061 8928
rect 18095 8925 18107 8959
rect 18049 8919 18107 8925
rect 8018 8848 8024 8900
rect 8076 8888 8082 8900
rect 10137 8891 10195 8897
rect 10137 8888 10149 8891
rect 8076 8860 10149 8888
rect 8076 8848 8082 8860
rect 10137 8857 10149 8860
rect 10183 8857 10195 8891
rect 10137 8851 10195 8857
rect 5166 8780 5172 8832
rect 5224 8820 5230 8832
rect 8481 8823 8539 8829
rect 8481 8820 8493 8823
rect 5224 8792 8493 8820
rect 5224 8780 5230 8792
rect 8481 8789 8493 8792
rect 8527 8820 8539 8823
rect 9309 8823 9367 8829
rect 9309 8820 9321 8823
rect 8527 8792 9321 8820
rect 8527 8789 8539 8792
rect 8481 8783 8539 8789
rect 9309 8789 9321 8792
rect 9355 8820 9367 8823
rect 9677 8823 9735 8829
rect 9677 8820 9689 8823
rect 9355 8792 9689 8820
rect 9355 8789 9367 8792
rect 9309 8783 9367 8789
rect 9677 8789 9689 8792
rect 9723 8820 9735 8823
rect 10229 8823 10287 8829
rect 10229 8820 10241 8823
rect 9723 8792 10241 8820
rect 9723 8789 9735 8792
rect 9677 8783 9735 8789
rect 10229 8789 10241 8792
rect 10275 8820 10287 8823
rect 10597 8823 10655 8829
rect 10597 8820 10609 8823
rect 10275 8792 10609 8820
rect 10275 8789 10287 8792
rect 10229 8783 10287 8789
rect 10597 8789 10609 8792
rect 10643 8820 10655 8823
rect 10965 8823 11023 8829
rect 10965 8820 10977 8823
rect 10643 8792 10977 8820
rect 10643 8789 10655 8792
rect 10597 8783 10655 8789
rect 10965 8789 10977 8792
rect 11011 8789 11023 8823
rect 10965 8783 11023 8789
rect 18230 8780 18236 8832
rect 18288 8780 18294 8832
rect 1104 8730 18860 8752
rect 1104 8678 2610 8730
rect 2662 8678 2674 8730
rect 2726 8678 2738 8730
rect 2790 8678 2802 8730
rect 2854 8678 2866 8730
rect 2918 8678 7610 8730
rect 7662 8678 7674 8730
rect 7726 8678 7738 8730
rect 7790 8678 7802 8730
rect 7854 8678 7866 8730
rect 7918 8678 12610 8730
rect 12662 8678 12674 8730
rect 12726 8678 12738 8730
rect 12790 8678 12802 8730
rect 12854 8678 12866 8730
rect 12918 8678 17610 8730
rect 17662 8678 17674 8730
rect 17726 8678 17738 8730
rect 17790 8678 17802 8730
rect 17854 8678 17866 8730
rect 17918 8678 18860 8730
rect 1104 8656 18860 8678
rect 3694 8576 3700 8628
rect 3752 8576 3758 8628
rect 8110 8576 8116 8628
rect 8168 8616 8174 8628
rect 14642 8616 14648 8628
rect 8168 8588 14648 8616
rect 8168 8576 8174 8588
rect 14642 8576 14648 8588
rect 14700 8616 14706 8628
rect 17957 8619 18015 8625
rect 14700 8588 17908 8616
rect 14700 8576 14706 8588
rect 10778 8548 10784 8560
rect 9600 8520 10784 8548
rect 2041 8483 2099 8489
rect 2041 8449 2053 8483
rect 2087 8480 2099 8483
rect 2087 8452 2544 8480
rect 2087 8449 2099 8452
rect 2041 8443 2099 8449
rect 2516 8424 2544 8452
rect 4246 8440 4252 8492
rect 4304 8480 4310 8492
rect 9600 8489 9628 8520
rect 10778 8508 10784 8520
rect 10836 8548 10842 8560
rect 10962 8548 10968 8560
rect 10836 8520 10968 8548
rect 10836 8508 10842 8520
rect 10962 8508 10968 8520
rect 11020 8508 11026 8560
rect 14090 8548 14096 8560
rect 11440 8520 14096 8548
rect 9585 8483 9643 8489
rect 9585 8480 9597 8483
rect 4304 8452 9597 8480
rect 4304 8440 4310 8452
rect 9585 8449 9597 8452
rect 9631 8449 9643 8483
rect 9585 8443 9643 8449
rect 9852 8483 9910 8489
rect 9852 8449 9864 8483
rect 9898 8480 9910 8483
rect 11440 8480 11468 8520
rect 14090 8508 14096 8520
rect 14148 8508 14154 8560
rect 14550 8508 14556 8560
rect 14608 8548 14614 8560
rect 17880 8548 17908 8588
rect 17957 8585 17969 8619
rect 18003 8616 18015 8619
rect 19058 8616 19064 8628
rect 18003 8588 19064 8616
rect 18003 8585 18015 8588
rect 17957 8579 18015 8585
rect 19058 8576 19064 8588
rect 19116 8576 19122 8628
rect 18046 8548 18052 8560
rect 14608 8520 17816 8548
rect 17880 8520 18052 8548
rect 14608 8508 14614 8520
rect 9898 8452 11468 8480
rect 9898 8449 9910 8452
rect 9852 8443 9910 8449
rect 11514 8440 11520 8492
rect 11572 8480 11578 8492
rect 17788 8489 17816 8520
rect 18046 8508 18052 8520
rect 18104 8508 18110 8560
rect 14645 8483 14703 8489
rect 14645 8480 14657 8483
rect 11572 8452 14657 8480
rect 11572 8440 11578 8452
rect 14645 8449 14657 8452
rect 14691 8449 14703 8483
rect 14645 8443 14703 8449
rect 17773 8483 17831 8489
rect 17773 8449 17785 8483
rect 17819 8449 17831 8483
rect 17773 8443 17831 8449
rect 2314 8372 2320 8424
rect 2372 8372 2378 8424
rect 2498 8372 2504 8424
rect 2556 8412 2562 8424
rect 2593 8415 2651 8421
rect 2593 8412 2605 8415
rect 2556 8384 2605 8412
rect 2556 8372 2562 8384
rect 2593 8381 2605 8384
rect 2639 8381 2651 8415
rect 2593 8375 2651 8381
rect 14366 8372 14372 8424
rect 14424 8372 14430 8424
rect 10965 8347 11023 8353
rect 10965 8313 10977 8347
rect 11011 8344 11023 8347
rect 11606 8344 11612 8356
rect 11011 8316 11612 8344
rect 11011 8313 11023 8316
rect 10965 8307 11023 8313
rect 11606 8304 11612 8316
rect 11664 8304 11670 8356
rect 12434 8236 12440 8288
rect 12492 8276 12498 8288
rect 13262 8276 13268 8288
rect 12492 8248 13268 8276
rect 12492 8236 12498 8248
rect 13262 8236 13268 8248
rect 13320 8236 13326 8288
rect 1104 8186 18860 8208
rect 1104 8134 1950 8186
rect 2002 8134 2014 8186
rect 2066 8134 2078 8186
rect 2130 8134 2142 8186
rect 2194 8134 2206 8186
rect 2258 8134 6950 8186
rect 7002 8134 7014 8186
rect 7066 8134 7078 8186
rect 7130 8134 7142 8186
rect 7194 8134 7206 8186
rect 7258 8134 11950 8186
rect 12002 8134 12014 8186
rect 12066 8134 12078 8186
rect 12130 8134 12142 8186
rect 12194 8134 12206 8186
rect 12258 8134 16950 8186
rect 17002 8134 17014 8186
rect 17066 8134 17078 8186
rect 17130 8134 17142 8186
rect 17194 8134 17206 8186
rect 17258 8134 18860 8186
rect 1104 8112 18860 8134
rect 1302 8032 1308 8084
rect 1360 8072 1366 8084
rect 2961 8075 3019 8081
rect 2961 8072 2973 8075
rect 1360 8044 2973 8072
rect 1360 8032 1366 8044
rect 2961 8041 2973 8044
rect 3007 8072 3019 8075
rect 3329 8075 3387 8081
rect 3329 8072 3341 8075
rect 3007 8044 3341 8072
rect 3007 8041 3019 8044
rect 2961 8035 3019 8041
rect 3329 8041 3341 8044
rect 3375 8072 3387 8075
rect 4341 8075 4399 8081
rect 4341 8072 4353 8075
rect 3375 8044 4353 8072
rect 3375 8041 3387 8044
rect 3329 8035 3387 8041
rect 4341 8041 4353 8044
rect 4387 8072 4399 8075
rect 4709 8075 4767 8081
rect 4709 8072 4721 8075
rect 4387 8044 4721 8072
rect 4387 8041 4399 8044
rect 4341 8035 4399 8041
rect 4709 8041 4721 8044
rect 4755 8072 4767 8075
rect 5077 8075 5135 8081
rect 5077 8072 5089 8075
rect 4755 8044 5089 8072
rect 4755 8041 4767 8044
rect 4709 8035 4767 8041
rect 5077 8041 5089 8044
rect 5123 8072 5135 8075
rect 5445 8075 5503 8081
rect 5445 8072 5457 8075
rect 5123 8044 5457 8072
rect 5123 8041 5135 8044
rect 5077 8035 5135 8041
rect 5445 8041 5457 8044
rect 5491 8041 5503 8075
rect 5445 8035 5503 8041
rect 11514 8032 11520 8084
rect 11572 8072 11578 8084
rect 11885 8075 11943 8081
rect 11885 8072 11897 8075
rect 11572 8044 11897 8072
rect 11572 8032 11578 8044
rect 11885 8041 11897 8044
rect 11931 8072 11943 8075
rect 11931 8044 12572 8072
rect 11931 8041 11943 8044
rect 11885 8035 11943 8041
rect 8754 7896 8760 7948
rect 8812 7936 8818 7948
rect 9585 7939 9643 7945
rect 9585 7936 9597 7939
rect 8812 7908 9597 7936
rect 8812 7896 8818 7908
rect 9585 7905 9597 7908
rect 9631 7905 9643 7939
rect 9585 7899 9643 7905
rect 9769 7939 9827 7945
rect 9769 7905 9781 7939
rect 9815 7936 9827 7939
rect 12434 7936 12440 7948
rect 9815 7908 12440 7936
rect 9815 7905 9827 7908
rect 9769 7899 9827 7905
rect 12434 7896 12440 7908
rect 12492 7896 12498 7948
rect 2958 7828 2964 7880
rect 3016 7868 3022 7880
rect 4157 7871 4215 7877
rect 4157 7868 4169 7871
rect 3016 7840 4169 7868
rect 3016 7828 3022 7840
rect 4157 7837 4169 7840
rect 4203 7837 4215 7871
rect 4157 7831 4215 7837
rect 9493 7871 9551 7877
rect 9493 7837 9505 7871
rect 9539 7868 9551 7871
rect 10042 7868 10048 7880
rect 9539 7840 10048 7868
rect 9539 7837 9551 7840
rect 9493 7831 9551 7837
rect 10042 7828 10048 7840
rect 10100 7868 10106 7880
rect 10870 7868 10876 7880
rect 10100 7840 10876 7868
rect 10100 7828 10106 7840
rect 10870 7828 10876 7840
rect 10928 7828 10934 7880
rect 12250 7828 12256 7880
rect 12308 7828 12314 7880
rect 12544 7800 12572 8044
rect 12897 7803 12955 7809
rect 12897 7800 12909 7803
rect 12452 7772 12909 7800
rect 9122 7692 9128 7744
rect 9180 7692 9186 7744
rect 12452 7741 12480 7772
rect 12897 7769 12909 7772
rect 12943 7800 12955 7803
rect 13173 7803 13231 7809
rect 13173 7800 13185 7803
rect 12943 7772 13185 7800
rect 12943 7769 12955 7772
rect 12897 7763 12955 7769
rect 13173 7769 13185 7772
rect 13219 7769 13231 7803
rect 13173 7763 13231 7769
rect 12437 7735 12495 7741
rect 12437 7701 12449 7735
rect 12483 7701 12495 7735
rect 12437 7695 12495 7701
rect 1104 7642 18860 7664
rect 1104 7590 2610 7642
rect 2662 7590 2674 7642
rect 2726 7590 2738 7642
rect 2790 7590 2802 7642
rect 2854 7590 2866 7642
rect 2918 7590 7610 7642
rect 7662 7590 7674 7642
rect 7726 7590 7738 7642
rect 7790 7590 7802 7642
rect 7854 7590 7866 7642
rect 7918 7590 12610 7642
rect 12662 7590 12674 7642
rect 12726 7590 12738 7642
rect 12790 7590 12802 7642
rect 12854 7590 12866 7642
rect 12918 7590 17610 7642
rect 17662 7590 17674 7642
rect 17726 7590 17738 7642
rect 17790 7590 17802 7642
rect 17854 7590 17866 7642
rect 17918 7590 18860 7642
rect 1104 7568 18860 7590
rect 11977 7531 12035 7537
rect 11977 7497 11989 7531
rect 12023 7528 12035 7531
rect 12250 7528 12256 7540
rect 12023 7500 12256 7528
rect 12023 7497 12035 7500
rect 11977 7491 12035 7497
rect 12250 7488 12256 7500
rect 12308 7488 12314 7540
rect 14182 7420 14188 7472
rect 14240 7420 14246 7472
rect 13814 7216 13820 7268
rect 13872 7256 13878 7268
rect 14369 7259 14427 7265
rect 14369 7256 14381 7259
rect 13872 7228 14381 7256
rect 13872 7216 13878 7228
rect 14369 7225 14381 7228
rect 14415 7225 14427 7259
rect 14369 7219 14427 7225
rect 1104 7098 18860 7120
rect 1104 7046 1950 7098
rect 2002 7046 2014 7098
rect 2066 7046 2078 7098
rect 2130 7046 2142 7098
rect 2194 7046 2206 7098
rect 2258 7046 6950 7098
rect 7002 7046 7014 7098
rect 7066 7046 7078 7098
rect 7130 7046 7142 7098
rect 7194 7046 7206 7098
rect 7258 7046 11950 7098
rect 12002 7046 12014 7098
rect 12066 7046 12078 7098
rect 12130 7046 12142 7098
rect 12194 7046 12206 7098
rect 12258 7046 16950 7098
rect 17002 7046 17014 7098
rect 17066 7046 17078 7098
rect 17130 7046 17142 7098
rect 17194 7046 17206 7098
rect 17258 7046 18860 7098
rect 1104 7024 18860 7046
rect 6914 6876 6920 6928
rect 6972 6876 6978 6928
rect 9217 6919 9275 6925
rect 9217 6885 9229 6919
rect 9263 6914 9275 6919
rect 9263 6886 9297 6914
rect 9263 6885 9275 6886
rect 9217 6879 9275 6885
rect 7374 6808 7380 6860
rect 7432 6808 7438 6860
rect 7466 6808 7472 6860
rect 7524 6808 7530 6860
rect 9232 6848 9260 6879
rect 10318 6848 10324 6860
rect 9232 6820 10324 6848
rect 10318 6808 10324 6820
rect 10376 6808 10382 6860
rect 18049 6783 18107 6789
rect 18049 6780 18061 6783
rect 6886 6752 18061 6780
rect 6270 6672 6276 6724
rect 6328 6712 6334 6724
rect 6886 6712 6914 6752
rect 18049 6749 18061 6752
rect 18095 6749 18107 6783
rect 18049 6743 18107 6749
rect 6328 6684 6914 6712
rect 6328 6672 6334 6684
rect 9490 6672 9496 6724
rect 9548 6672 9554 6724
rect 9674 6672 9680 6724
rect 9732 6672 9738 6724
rect 9769 6715 9827 6721
rect 9769 6681 9781 6715
rect 9815 6712 9827 6715
rect 13538 6712 13544 6724
rect 9815 6684 13544 6712
rect 9815 6681 9827 6684
rect 9769 6675 9827 6681
rect 13538 6672 13544 6684
rect 13596 6672 13602 6724
rect 7377 6647 7435 6653
rect 7377 6613 7389 6647
rect 7423 6644 7435 6647
rect 12710 6644 12716 6656
rect 7423 6616 12716 6644
rect 7423 6613 7435 6616
rect 7377 6607 7435 6613
rect 12710 6604 12716 6616
rect 12768 6604 12774 6656
rect 18230 6604 18236 6656
rect 18288 6604 18294 6656
rect 1104 6554 18860 6576
rect 1104 6502 2610 6554
rect 2662 6502 2674 6554
rect 2726 6502 2738 6554
rect 2790 6502 2802 6554
rect 2854 6502 2866 6554
rect 2918 6502 7610 6554
rect 7662 6502 7674 6554
rect 7726 6502 7738 6554
rect 7790 6502 7802 6554
rect 7854 6502 7866 6554
rect 7918 6502 12610 6554
rect 12662 6502 12674 6554
rect 12726 6502 12738 6554
rect 12790 6502 12802 6554
rect 12854 6502 12866 6554
rect 12918 6502 17610 6554
rect 17662 6502 17674 6554
rect 17726 6502 17738 6554
rect 17790 6502 17802 6554
rect 17854 6502 17866 6554
rect 17918 6502 18860 6554
rect 1104 6480 18860 6502
rect 3602 6400 3608 6452
rect 3660 6440 3666 6452
rect 9490 6440 9496 6452
rect 3660 6412 9496 6440
rect 3660 6400 3666 6412
rect 9490 6400 9496 6412
rect 9548 6400 9554 6452
rect 5810 6332 5816 6384
rect 5868 6372 5874 6384
rect 8202 6372 8208 6384
rect 5868 6344 8208 6372
rect 5868 6332 5874 6344
rect 8202 6332 8208 6344
rect 8260 6332 8266 6384
rect 1104 6010 18860 6032
rect 1104 5958 1950 6010
rect 2002 5958 2014 6010
rect 2066 5958 2078 6010
rect 2130 5958 2142 6010
rect 2194 5958 2206 6010
rect 2258 5958 6950 6010
rect 7002 5958 7014 6010
rect 7066 5958 7078 6010
rect 7130 5958 7142 6010
rect 7194 5958 7206 6010
rect 7258 5958 11950 6010
rect 12002 5958 12014 6010
rect 12066 5958 12078 6010
rect 12130 5958 12142 6010
rect 12194 5958 12206 6010
rect 12258 5958 16950 6010
rect 17002 5958 17014 6010
rect 17066 5958 17078 6010
rect 17130 5958 17142 6010
rect 17194 5958 17206 6010
rect 17258 5958 18860 6010
rect 1104 5936 18860 5958
rect 2314 5652 2320 5704
rect 2372 5692 2378 5704
rect 5074 5692 5080 5704
rect 2372 5664 5080 5692
rect 2372 5652 2378 5664
rect 5074 5652 5080 5664
rect 5132 5652 5138 5704
rect 5344 5695 5402 5701
rect 5344 5661 5356 5695
rect 5390 5692 5402 5695
rect 6178 5692 6184 5704
rect 5390 5664 6184 5692
rect 5390 5661 5402 5664
rect 5344 5655 5402 5661
rect 6178 5652 6184 5664
rect 6236 5652 6242 5704
rect 6457 5559 6515 5565
rect 6457 5525 6469 5559
rect 6503 5556 6515 5559
rect 11422 5556 11428 5568
rect 6503 5528 11428 5556
rect 6503 5525 6515 5528
rect 6457 5519 6515 5525
rect 11422 5516 11428 5528
rect 11480 5516 11486 5568
rect 1104 5466 18860 5488
rect 1104 5414 2610 5466
rect 2662 5414 2674 5466
rect 2726 5414 2738 5466
rect 2790 5414 2802 5466
rect 2854 5414 2866 5466
rect 2918 5414 7610 5466
rect 7662 5414 7674 5466
rect 7726 5414 7738 5466
rect 7790 5414 7802 5466
rect 7854 5414 7866 5466
rect 7918 5414 12610 5466
rect 12662 5414 12674 5466
rect 12726 5414 12738 5466
rect 12790 5414 12802 5466
rect 12854 5414 12866 5466
rect 12918 5414 17610 5466
rect 17662 5414 17674 5466
rect 17726 5414 17738 5466
rect 17790 5414 17802 5466
rect 17854 5414 17866 5466
rect 17918 5414 18860 5466
rect 1104 5392 18860 5414
rect 1670 5312 1676 5364
rect 1728 5352 1734 5364
rect 1728 5324 16988 5352
rect 1728 5312 1734 5324
rect 13354 5244 13360 5296
rect 13412 5244 13418 5296
rect 16960 5293 16988 5324
rect 16945 5287 17003 5293
rect 16945 5253 16957 5287
rect 16991 5253 17003 5287
rect 16945 5247 17003 5253
rect 5905 5219 5963 5225
rect 5905 5185 5917 5219
rect 5951 5216 5963 5219
rect 9122 5216 9128 5228
rect 5951 5188 9128 5216
rect 5951 5185 5963 5188
rect 5905 5179 5963 5185
rect 9122 5176 9128 5188
rect 9180 5176 9186 5228
rect 11054 5176 11060 5228
rect 11112 5216 11118 5228
rect 11698 5216 11704 5228
rect 11112 5188 11704 5216
rect 11112 5176 11118 5188
rect 11698 5176 11704 5188
rect 11756 5176 11762 5228
rect 16206 5176 16212 5228
rect 16264 5216 16270 5228
rect 17129 5219 17187 5225
rect 17129 5216 17141 5219
rect 16264 5188 17141 5216
rect 16264 5176 16270 5188
rect 17129 5185 17141 5188
rect 17175 5216 17187 5219
rect 17405 5219 17463 5225
rect 17405 5216 17417 5219
rect 17175 5188 17417 5216
rect 17175 5185 17187 5188
rect 17129 5179 17187 5185
rect 17405 5185 17417 5188
rect 17451 5185 17463 5219
rect 17405 5179 17463 5185
rect 11977 5151 12035 5157
rect 11977 5148 11989 5151
rect 11072 5120 11989 5148
rect 6546 5040 6552 5092
rect 6604 5080 6610 5092
rect 11072 5089 11100 5120
rect 11977 5117 11989 5120
rect 12023 5148 12035 5151
rect 13633 5151 13691 5157
rect 13633 5148 13645 5151
rect 12023 5120 13645 5148
rect 12023 5117 12035 5120
rect 11977 5111 12035 5117
rect 13633 5117 13645 5120
rect 13679 5148 13691 5151
rect 14001 5151 14059 5157
rect 14001 5148 14013 5151
rect 13679 5120 14013 5148
rect 13679 5117 13691 5120
rect 13633 5111 13691 5117
rect 14001 5117 14013 5120
rect 14047 5148 14059 5151
rect 14369 5151 14427 5157
rect 14369 5148 14381 5151
rect 14047 5120 14381 5148
rect 14047 5117 14059 5120
rect 14001 5111 14059 5117
rect 14369 5117 14381 5120
rect 14415 5117 14427 5151
rect 17420 5148 17448 5179
rect 17494 5176 17500 5228
rect 17552 5216 17558 5228
rect 18049 5219 18107 5225
rect 18049 5216 18061 5219
rect 17552 5188 18061 5216
rect 17552 5176 17558 5188
rect 18049 5185 18061 5188
rect 18095 5185 18107 5219
rect 18049 5179 18107 5185
rect 17773 5151 17831 5157
rect 17773 5148 17785 5151
rect 17420 5120 17785 5148
rect 14369 5111 14427 5117
rect 17773 5117 17785 5120
rect 17819 5117 17831 5151
rect 17773 5111 17831 5117
rect 10689 5083 10747 5089
rect 10689 5080 10701 5083
rect 6604 5052 10701 5080
rect 6604 5040 6610 5052
rect 10689 5049 10701 5052
rect 10735 5080 10747 5083
rect 11057 5083 11115 5089
rect 11057 5080 11069 5083
rect 10735 5052 11069 5080
rect 10735 5049 10747 5052
rect 10689 5043 10747 5049
rect 11057 5049 11069 5052
rect 11103 5049 11115 5083
rect 11057 5043 11115 5049
rect 5721 5015 5779 5021
rect 5721 4981 5733 5015
rect 5767 5012 5779 5015
rect 8110 5012 8116 5024
rect 5767 4984 8116 5012
rect 5767 4981 5779 4984
rect 5721 4975 5779 4981
rect 8110 4972 8116 4984
rect 8168 4972 8174 5024
rect 18230 4972 18236 5024
rect 18288 4972 18294 5024
rect 1104 4922 18860 4944
rect 1104 4870 1950 4922
rect 2002 4870 2014 4922
rect 2066 4870 2078 4922
rect 2130 4870 2142 4922
rect 2194 4870 2206 4922
rect 2258 4870 6950 4922
rect 7002 4870 7014 4922
rect 7066 4870 7078 4922
rect 7130 4870 7142 4922
rect 7194 4870 7206 4922
rect 7258 4870 11950 4922
rect 12002 4870 12014 4922
rect 12066 4870 12078 4922
rect 12130 4870 12142 4922
rect 12194 4870 12206 4922
rect 12258 4870 16950 4922
rect 17002 4870 17014 4922
rect 17066 4870 17078 4922
rect 17130 4870 17142 4922
rect 17194 4870 17206 4922
rect 17258 4870 18860 4922
rect 1104 4848 18860 4870
rect 7282 4632 7288 4684
rect 7340 4672 7346 4684
rect 10321 4675 10379 4681
rect 10321 4672 10333 4675
rect 7340 4644 10333 4672
rect 7340 4632 7346 4644
rect 10321 4641 10333 4644
rect 10367 4641 10379 4675
rect 10321 4635 10379 4641
rect 10045 4607 10103 4613
rect 10045 4573 10057 4607
rect 10091 4604 10103 4607
rect 14458 4604 14464 4616
rect 10091 4576 14464 4604
rect 10091 4573 10103 4576
rect 10045 4567 10103 4573
rect 14458 4564 14464 4576
rect 14516 4564 14522 4616
rect 1104 4378 18860 4400
rect 1104 4326 2610 4378
rect 2662 4326 2674 4378
rect 2726 4326 2738 4378
rect 2790 4326 2802 4378
rect 2854 4326 2866 4378
rect 2918 4326 7610 4378
rect 7662 4326 7674 4378
rect 7726 4326 7738 4378
rect 7790 4326 7802 4378
rect 7854 4326 7866 4378
rect 7918 4326 12610 4378
rect 12662 4326 12674 4378
rect 12726 4326 12738 4378
rect 12790 4326 12802 4378
rect 12854 4326 12866 4378
rect 12918 4326 17610 4378
rect 17662 4326 17674 4378
rect 17726 4326 17738 4378
rect 17790 4326 17802 4378
rect 17854 4326 17866 4378
rect 17918 4326 18860 4378
rect 1104 4304 18860 4326
rect 5074 4088 5080 4140
rect 5132 4128 5138 4140
rect 6549 4131 6607 4137
rect 6549 4128 6561 4131
rect 5132 4100 6561 4128
rect 5132 4088 5138 4100
rect 6549 4097 6561 4100
rect 6595 4097 6607 4131
rect 6805 4131 6863 4137
rect 6805 4128 6817 4131
rect 6549 4091 6607 4097
rect 6656 4100 6817 4128
rect 1210 4020 1216 4072
rect 1268 4060 1274 4072
rect 6656 4060 6684 4100
rect 6805 4097 6817 4100
rect 6851 4097 6863 4131
rect 6805 4091 6863 4097
rect 9769 4131 9827 4137
rect 9769 4097 9781 4131
rect 9815 4128 9827 4131
rect 16666 4128 16672 4140
rect 9815 4100 16672 4128
rect 9815 4097 9827 4100
rect 9769 4091 9827 4097
rect 16666 4088 16672 4100
rect 16724 4088 16730 4140
rect 1268 4032 6684 4060
rect 1268 4020 1274 4032
rect 8202 4020 8208 4072
rect 8260 4060 8266 4072
rect 10045 4063 10103 4069
rect 10045 4060 10057 4063
rect 8260 4032 10057 4060
rect 8260 4020 8266 4032
rect 10045 4029 10057 4032
rect 10091 4029 10103 4063
rect 10045 4023 10103 4029
rect 7929 3995 7987 4001
rect 7929 3961 7941 3995
rect 7975 3992 7987 3995
rect 8294 3992 8300 4004
rect 7975 3964 8300 3992
rect 7975 3961 7987 3964
rect 7929 3955 7987 3961
rect 8294 3952 8300 3964
rect 8352 3952 8358 4004
rect 1104 3834 18860 3856
rect 1104 3782 1950 3834
rect 2002 3782 2014 3834
rect 2066 3782 2078 3834
rect 2130 3782 2142 3834
rect 2194 3782 2206 3834
rect 2258 3782 6950 3834
rect 7002 3782 7014 3834
rect 7066 3782 7078 3834
rect 7130 3782 7142 3834
rect 7194 3782 7206 3834
rect 7258 3782 11950 3834
rect 12002 3782 12014 3834
rect 12066 3782 12078 3834
rect 12130 3782 12142 3834
rect 12194 3782 12206 3834
rect 12258 3782 16950 3834
rect 17002 3782 17014 3834
rect 17066 3782 17078 3834
rect 17130 3782 17142 3834
rect 17194 3782 17206 3834
rect 17258 3782 18860 3834
rect 1104 3760 18860 3782
rect 10962 3680 10968 3732
rect 11020 3720 11026 3732
rect 13633 3723 13691 3729
rect 13633 3720 13645 3723
rect 11020 3692 13645 3720
rect 11020 3680 11026 3692
rect 13633 3689 13645 3692
rect 13679 3689 13691 3723
rect 13633 3683 13691 3689
rect 11698 3544 11704 3596
rect 11756 3584 11762 3596
rect 12253 3587 12311 3593
rect 12253 3584 12265 3587
rect 11756 3556 12265 3584
rect 11756 3544 11762 3556
rect 12253 3553 12265 3556
rect 12299 3553 12311 3587
rect 12253 3547 12311 3553
rect 8110 3476 8116 3528
rect 8168 3516 8174 3528
rect 12509 3519 12567 3525
rect 12509 3516 12521 3519
rect 8168 3488 12521 3516
rect 8168 3476 8174 3488
rect 12509 3485 12521 3488
rect 12555 3485 12567 3519
rect 12509 3479 12567 3485
rect 1104 3290 18860 3312
rect 1104 3238 2610 3290
rect 2662 3238 2674 3290
rect 2726 3238 2738 3290
rect 2790 3238 2802 3290
rect 2854 3238 2866 3290
rect 2918 3238 7610 3290
rect 7662 3238 7674 3290
rect 7726 3238 7738 3290
rect 7790 3238 7802 3290
rect 7854 3238 7866 3290
rect 7918 3238 12610 3290
rect 12662 3238 12674 3290
rect 12726 3238 12738 3290
rect 12790 3238 12802 3290
rect 12854 3238 12866 3290
rect 12918 3238 17610 3290
rect 17662 3238 17674 3290
rect 17726 3238 17738 3290
rect 17790 3238 17802 3290
rect 17854 3238 17866 3290
rect 17918 3238 18860 3290
rect 1104 3216 18860 3238
rect 3881 3179 3939 3185
rect 3881 3145 3893 3179
rect 3927 3176 3939 3179
rect 9306 3176 9312 3188
rect 3927 3148 9312 3176
rect 3927 3145 3939 3148
rect 3881 3139 3939 3145
rect 9306 3136 9312 3148
rect 9364 3136 9370 3188
rect 2768 3111 2826 3117
rect 2768 3077 2780 3111
rect 2814 3108 2826 3111
rect 5626 3108 5632 3120
rect 2814 3080 5632 3108
rect 2814 3077 2826 3080
rect 2768 3071 2826 3077
rect 5626 3068 5632 3080
rect 5684 3068 5690 3120
rect 18049 3043 18107 3049
rect 18049 3009 18061 3043
rect 18095 3040 18107 3043
rect 19702 3040 19708 3052
rect 18095 3012 19708 3040
rect 18095 3009 18107 3012
rect 18049 3003 18107 3009
rect 19702 3000 19708 3012
rect 19760 3000 19766 3052
rect 2314 2932 2320 2984
rect 2372 2972 2378 2984
rect 2501 2975 2559 2981
rect 2501 2972 2513 2975
rect 2372 2944 2513 2972
rect 2372 2932 2378 2944
rect 2501 2941 2513 2944
rect 2547 2941 2559 2975
rect 2501 2935 2559 2941
rect 18230 2796 18236 2848
rect 18288 2796 18294 2848
rect 1104 2746 18860 2768
rect 1104 2694 1950 2746
rect 2002 2694 2014 2746
rect 2066 2694 2078 2746
rect 2130 2694 2142 2746
rect 2194 2694 2206 2746
rect 2258 2694 6950 2746
rect 7002 2694 7014 2746
rect 7066 2694 7078 2746
rect 7130 2694 7142 2746
rect 7194 2694 7206 2746
rect 7258 2694 11950 2746
rect 12002 2694 12014 2746
rect 12066 2694 12078 2746
rect 12130 2694 12142 2746
rect 12194 2694 12206 2746
rect 12258 2694 16950 2746
rect 17002 2694 17014 2746
rect 17066 2694 17078 2746
rect 17130 2694 17142 2746
rect 17194 2694 17206 2746
rect 17258 2694 18860 2746
rect 1104 2672 18860 2694
rect 7193 2635 7251 2641
rect 7193 2601 7205 2635
rect 7239 2632 7251 2635
rect 7561 2635 7619 2641
rect 7561 2632 7573 2635
rect 7239 2604 7573 2632
rect 7239 2601 7251 2604
rect 7193 2595 7251 2601
rect 7561 2601 7573 2604
rect 7607 2632 7619 2635
rect 7929 2635 7987 2641
rect 7929 2632 7941 2635
rect 7607 2604 7941 2632
rect 7607 2601 7619 2604
rect 7561 2595 7619 2601
rect 7929 2601 7941 2604
rect 7975 2632 7987 2635
rect 9858 2632 9864 2644
rect 7975 2604 9864 2632
rect 7975 2601 7987 2604
rect 7929 2595 7987 2601
rect 5994 2388 6000 2440
rect 6052 2428 6058 2440
rect 6549 2431 6607 2437
rect 6549 2428 6561 2431
rect 6052 2400 6561 2428
rect 6052 2388 6058 2400
rect 6549 2397 6561 2400
rect 6595 2397 6607 2431
rect 6549 2391 6607 2397
rect 5629 2295 5687 2301
rect 5629 2261 5641 2295
rect 5675 2292 5687 2295
rect 5905 2295 5963 2301
rect 5905 2292 5917 2295
rect 5675 2264 5917 2292
rect 5675 2261 5687 2264
rect 5629 2255 5687 2261
rect 5905 2261 5917 2264
rect 5951 2292 5963 2295
rect 6733 2295 6791 2301
rect 6733 2292 6745 2295
rect 5951 2264 6745 2292
rect 5951 2261 5963 2264
rect 5905 2255 5963 2261
rect 6733 2261 6745 2264
rect 6779 2292 6791 2295
rect 7208 2292 7236 2595
rect 9858 2592 9864 2604
rect 9916 2592 9922 2644
rect 14458 2592 14464 2644
rect 14516 2592 14522 2644
rect 18046 2456 18052 2508
rect 18104 2456 18110 2508
rect 8846 2388 8852 2440
rect 8904 2428 8910 2440
rect 10045 2431 10103 2437
rect 10045 2428 10057 2431
rect 8904 2400 10057 2428
rect 8904 2388 8910 2400
rect 10045 2397 10057 2400
rect 10091 2397 10103 2431
rect 10045 2391 10103 2397
rect 17862 2388 17868 2440
rect 17920 2388 17926 2440
rect 13906 2320 13912 2372
rect 13964 2360 13970 2372
rect 14369 2363 14427 2369
rect 14369 2360 14381 2363
rect 13964 2332 14381 2360
rect 13964 2320 13970 2332
rect 14369 2329 14381 2332
rect 14415 2329 14427 2363
rect 14369 2323 14427 2329
rect 6779 2264 7236 2292
rect 6779 2261 6791 2264
rect 6733 2255 6791 2261
rect 9950 2252 9956 2304
rect 10008 2292 10014 2304
rect 10229 2295 10287 2301
rect 10229 2292 10241 2295
rect 10008 2264 10241 2292
rect 10008 2252 10014 2264
rect 10229 2261 10241 2264
rect 10275 2261 10287 2295
rect 10229 2255 10287 2261
rect 1104 2202 18860 2224
rect 1104 2150 2610 2202
rect 2662 2150 2674 2202
rect 2726 2150 2738 2202
rect 2790 2150 2802 2202
rect 2854 2150 2866 2202
rect 2918 2150 7610 2202
rect 7662 2150 7674 2202
rect 7726 2150 7738 2202
rect 7790 2150 7802 2202
rect 7854 2150 7866 2202
rect 7918 2150 12610 2202
rect 12662 2150 12674 2202
rect 12726 2150 12738 2202
rect 12790 2150 12802 2202
rect 12854 2150 12866 2202
rect 12918 2150 17610 2202
rect 17662 2150 17674 2202
rect 17726 2150 17738 2202
rect 17790 2150 17802 2202
rect 17854 2150 17866 2202
rect 17918 2150 18860 2202
rect 1104 2128 18860 2150
<< via1 >>
rect 1950 77766 2002 77818
rect 2014 77766 2066 77818
rect 2078 77766 2130 77818
rect 2142 77766 2194 77818
rect 2206 77766 2258 77818
rect 6950 77766 7002 77818
rect 7014 77766 7066 77818
rect 7078 77766 7130 77818
rect 7142 77766 7194 77818
rect 7206 77766 7258 77818
rect 11950 77766 12002 77818
rect 12014 77766 12066 77818
rect 12078 77766 12130 77818
rect 12142 77766 12194 77818
rect 12206 77766 12258 77818
rect 16950 77766 17002 77818
rect 17014 77766 17066 77818
rect 17078 77766 17130 77818
rect 17142 77766 17194 77818
rect 17206 77766 17258 77818
rect 18328 77460 18380 77512
rect 16856 77324 16908 77376
rect 18236 77367 18288 77376
rect 18236 77333 18245 77367
rect 18245 77333 18279 77367
rect 18279 77333 18288 77367
rect 18236 77324 18288 77333
rect 2610 77222 2662 77274
rect 2674 77222 2726 77274
rect 2738 77222 2790 77274
rect 2802 77222 2854 77274
rect 2866 77222 2918 77274
rect 7610 77222 7662 77274
rect 7674 77222 7726 77274
rect 7738 77222 7790 77274
rect 7802 77222 7854 77274
rect 7866 77222 7918 77274
rect 12610 77222 12662 77274
rect 12674 77222 12726 77274
rect 12738 77222 12790 77274
rect 12802 77222 12854 77274
rect 12866 77222 12918 77274
rect 17610 77222 17662 77274
rect 17674 77222 17726 77274
rect 17738 77222 17790 77274
rect 17802 77222 17854 77274
rect 17866 77222 17918 77274
rect 17500 76916 17552 76968
rect 14648 76823 14700 76832
rect 14648 76789 14657 76823
rect 14657 76789 14691 76823
rect 14691 76789 14700 76823
rect 14648 76780 14700 76789
rect 15936 76823 15988 76832
rect 15936 76789 15945 76823
rect 15945 76789 15979 76823
rect 15979 76789 15988 76823
rect 15936 76780 15988 76789
rect 16488 76780 16540 76832
rect 1950 76678 2002 76730
rect 2014 76678 2066 76730
rect 2078 76678 2130 76730
rect 2142 76678 2194 76730
rect 2206 76678 2258 76730
rect 6950 76678 7002 76730
rect 7014 76678 7066 76730
rect 7078 76678 7130 76730
rect 7142 76678 7194 76730
rect 7206 76678 7258 76730
rect 11950 76678 12002 76730
rect 12014 76678 12066 76730
rect 12078 76678 12130 76730
rect 12142 76678 12194 76730
rect 12206 76678 12258 76730
rect 16950 76678 17002 76730
rect 17014 76678 17066 76730
rect 17078 76678 17130 76730
rect 17142 76678 17194 76730
rect 17206 76678 17258 76730
rect 16488 76576 16540 76628
rect 7932 76440 7984 76492
rect 2964 76236 3016 76288
rect 7104 76236 7156 76288
rect 8208 76372 8260 76424
rect 14924 76415 14976 76424
rect 14924 76381 14933 76415
rect 14933 76381 14967 76415
rect 14967 76381 14976 76415
rect 14924 76372 14976 76381
rect 8484 76347 8536 76356
rect 8484 76313 8493 76347
rect 8493 76313 8527 76347
rect 8527 76313 8536 76347
rect 8484 76304 8536 76313
rect 8944 76236 8996 76288
rect 11244 76279 11296 76288
rect 11244 76245 11253 76279
rect 11253 76245 11287 76279
rect 11287 76245 11296 76279
rect 14648 76304 14700 76356
rect 16856 76304 16908 76356
rect 11244 76236 11296 76245
rect 11704 76279 11756 76288
rect 11704 76245 11713 76279
rect 11713 76245 11747 76279
rect 11747 76245 11756 76279
rect 11704 76236 11756 76245
rect 16304 76279 16356 76288
rect 16304 76245 16313 76279
rect 16313 76245 16347 76279
rect 16347 76245 16356 76279
rect 16304 76236 16356 76245
rect 2610 76134 2662 76186
rect 2674 76134 2726 76186
rect 2738 76134 2790 76186
rect 2802 76134 2854 76186
rect 2866 76134 2918 76186
rect 7610 76134 7662 76186
rect 7674 76134 7726 76186
rect 7738 76134 7790 76186
rect 7802 76134 7854 76186
rect 7866 76134 7918 76186
rect 12610 76134 12662 76186
rect 12674 76134 12726 76186
rect 12738 76134 12790 76186
rect 12802 76134 12854 76186
rect 12866 76134 12918 76186
rect 17610 76134 17662 76186
rect 17674 76134 17726 76186
rect 17738 76134 17790 76186
rect 17802 76134 17854 76186
rect 17866 76134 17918 76186
rect 5540 75964 5592 76016
rect 16672 76032 16724 76084
rect 6644 75828 6696 75880
rect 7104 75939 7156 75948
rect 7104 75905 7113 75939
rect 7113 75905 7147 75939
rect 7147 75905 7156 75939
rect 7104 75896 7156 75905
rect 7380 75896 7432 75948
rect 7564 76007 7616 76016
rect 7564 75973 7573 76007
rect 7573 75973 7607 76007
rect 7607 75973 7616 76007
rect 7564 75964 7616 75973
rect 8760 76007 8812 76016
rect 8760 75973 8769 76007
rect 8769 75973 8803 76007
rect 8803 75973 8812 76007
rect 8760 75964 8812 75973
rect 12440 75964 12492 76016
rect 14096 75939 14148 75948
rect 14096 75905 14105 75939
rect 14105 75905 14139 75939
rect 14139 75905 14148 75939
rect 14096 75896 14148 75905
rect 14188 75939 14240 75948
rect 14188 75905 14197 75939
rect 14197 75905 14231 75939
rect 14231 75905 14240 75939
rect 14188 75896 14240 75905
rect 14464 75828 14516 75880
rect 9220 75735 9272 75744
rect 9220 75701 9229 75735
rect 9229 75701 9263 75735
rect 9263 75701 9272 75735
rect 9220 75692 9272 75701
rect 13728 75735 13780 75744
rect 13728 75701 13737 75735
rect 13737 75701 13771 75735
rect 13771 75701 13780 75735
rect 13728 75692 13780 75701
rect 1950 75590 2002 75642
rect 2014 75590 2066 75642
rect 2078 75590 2130 75642
rect 2142 75590 2194 75642
rect 2206 75590 2258 75642
rect 6950 75590 7002 75642
rect 7014 75590 7066 75642
rect 7078 75590 7130 75642
rect 7142 75590 7194 75642
rect 7206 75590 7258 75642
rect 11950 75590 12002 75642
rect 12014 75590 12066 75642
rect 12078 75590 12130 75642
rect 12142 75590 12194 75642
rect 12206 75590 12258 75642
rect 16950 75590 17002 75642
rect 17014 75590 17066 75642
rect 17078 75590 17130 75642
rect 17142 75590 17194 75642
rect 17206 75590 17258 75642
rect 15200 75463 15252 75472
rect 15200 75429 15209 75463
rect 15209 75429 15243 75463
rect 15243 75429 15252 75463
rect 15200 75420 15252 75429
rect 11796 75352 11848 75404
rect 5448 75284 5500 75336
rect 7288 75284 7340 75336
rect 8116 75284 8168 75336
rect 5080 75191 5132 75200
rect 5080 75157 5089 75191
rect 5089 75157 5123 75191
rect 5123 75157 5132 75191
rect 5080 75148 5132 75157
rect 6552 75191 6604 75200
rect 6552 75157 6561 75191
rect 6561 75157 6595 75191
rect 6595 75157 6604 75191
rect 6552 75148 6604 75157
rect 14096 75216 14148 75268
rect 16028 75148 16080 75200
rect 18236 75191 18288 75200
rect 18236 75157 18245 75191
rect 18245 75157 18279 75191
rect 18279 75157 18288 75191
rect 18236 75148 18288 75157
rect 2610 75046 2662 75098
rect 2674 75046 2726 75098
rect 2738 75046 2790 75098
rect 2802 75046 2854 75098
rect 2866 75046 2918 75098
rect 7610 75046 7662 75098
rect 7674 75046 7726 75098
rect 7738 75046 7790 75098
rect 7802 75046 7854 75098
rect 7866 75046 7918 75098
rect 12610 75046 12662 75098
rect 12674 75046 12726 75098
rect 12738 75046 12790 75098
rect 12802 75046 12854 75098
rect 12866 75046 12918 75098
rect 17610 75046 17662 75098
rect 17674 75046 17726 75098
rect 17738 75046 17790 75098
rect 17802 75046 17854 75098
rect 17866 75046 17918 75098
rect 8116 74944 8168 74996
rect 15292 74944 15344 74996
rect 6552 74876 6604 74928
rect 6460 74808 6512 74860
rect 14924 74808 14976 74860
rect 15108 74851 15160 74860
rect 15108 74817 15142 74851
rect 15142 74817 15160 74851
rect 15108 74808 15160 74817
rect 16856 74851 16908 74860
rect 16856 74817 16865 74851
rect 16865 74817 16899 74851
rect 16899 74817 16908 74851
rect 16856 74808 16908 74817
rect 4620 74672 4672 74724
rect 9404 74740 9456 74792
rect 15844 74672 15896 74724
rect 17500 74672 17552 74724
rect 6736 74647 6788 74656
rect 6736 74613 6745 74647
rect 6745 74613 6779 74647
rect 6779 74613 6788 74647
rect 6736 74604 6788 74613
rect 18788 74604 18840 74656
rect 1950 74502 2002 74554
rect 2014 74502 2066 74554
rect 2078 74502 2130 74554
rect 2142 74502 2194 74554
rect 2206 74502 2258 74554
rect 6950 74502 7002 74554
rect 7014 74502 7066 74554
rect 7078 74502 7130 74554
rect 7142 74502 7194 74554
rect 7206 74502 7258 74554
rect 11950 74502 12002 74554
rect 12014 74502 12066 74554
rect 12078 74502 12130 74554
rect 12142 74502 12194 74554
rect 12206 74502 12258 74554
rect 16950 74502 17002 74554
rect 17014 74502 17066 74554
rect 17078 74502 17130 74554
rect 17142 74502 17194 74554
rect 17206 74502 17258 74554
rect 7380 74400 7432 74452
rect 10324 74400 10376 74452
rect 16856 74400 16908 74452
rect 13728 74264 13780 74316
rect 14280 74239 14332 74248
rect 14280 74205 14289 74239
rect 14289 74205 14323 74239
rect 14323 74205 14332 74239
rect 14280 74196 14332 74205
rect 14924 74196 14976 74248
rect 10508 74128 10560 74180
rect 12440 74103 12492 74112
rect 12440 74069 12449 74103
rect 12449 74069 12483 74103
rect 12483 74069 12492 74103
rect 12440 74060 12492 74069
rect 13452 74060 13504 74112
rect 15568 74060 15620 74112
rect 2610 73958 2662 74010
rect 2674 73958 2726 74010
rect 2738 73958 2790 74010
rect 2802 73958 2854 74010
rect 2866 73958 2918 74010
rect 7610 73958 7662 74010
rect 7674 73958 7726 74010
rect 7738 73958 7790 74010
rect 7802 73958 7854 74010
rect 7866 73958 7918 74010
rect 12610 73958 12662 74010
rect 12674 73958 12726 74010
rect 12738 73958 12790 74010
rect 12802 73958 12854 74010
rect 12866 73958 12918 74010
rect 17610 73958 17662 74010
rect 17674 73958 17726 74010
rect 17738 73958 17790 74010
rect 17802 73958 17854 74010
rect 17866 73958 17918 74010
rect 7288 73899 7340 73908
rect 7288 73865 7297 73899
rect 7297 73865 7331 73899
rect 7331 73865 7340 73899
rect 7288 73856 7340 73865
rect 15936 73788 15988 73840
rect 16304 73788 16356 73840
rect 7380 73720 7432 73772
rect 8208 73652 8260 73704
rect 17500 73652 17552 73704
rect 18236 73559 18288 73568
rect 18236 73525 18245 73559
rect 18245 73525 18279 73559
rect 18279 73525 18288 73559
rect 18236 73516 18288 73525
rect 1950 73414 2002 73466
rect 2014 73414 2066 73466
rect 2078 73414 2130 73466
rect 2142 73414 2194 73466
rect 2206 73414 2258 73466
rect 6950 73414 7002 73466
rect 7014 73414 7066 73466
rect 7078 73414 7130 73466
rect 7142 73414 7194 73466
rect 7206 73414 7258 73466
rect 11950 73414 12002 73466
rect 12014 73414 12066 73466
rect 12078 73414 12130 73466
rect 12142 73414 12194 73466
rect 12206 73414 12258 73466
rect 16950 73414 17002 73466
rect 17014 73414 17066 73466
rect 17078 73414 17130 73466
rect 17142 73414 17194 73466
rect 17206 73414 17258 73466
rect 5540 73176 5592 73228
rect 1308 72972 1360 73024
rect 8116 72972 8168 73024
rect 2610 72870 2662 72922
rect 2674 72870 2726 72922
rect 2738 72870 2790 72922
rect 2802 72870 2854 72922
rect 2866 72870 2918 72922
rect 7610 72870 7662 72922
rect 7674 72870 7726 72922
rect 7738 72870 7790 72922
rect 7802 72870 7854 72922
rect 7866 72870 7918 72922
rect 12610 72870 12662 72922
rect 12674 72870 12726 72922
rect 12738 72870 12790 72922
rect 12802 72870 12854 72922
rect 12866 72870 12918 72922
rect 17610 72870 17662 72922
rect 17674 72870 17726 72922
rect 17738 72870 17790 72922
rect 17802 72870 17854 72922
rect 17866 72870 17918 72922
rect 8208 72700 8260 72752
rect 12348 72632 12400 72684
rect 7380 72564 7432 72616
rect 16580 72564 16632 72616
rect 13268 72428 13320 72480
rect 1950 72326 2002 72378
rect 2014 72326 2066 72378
rect 2078 72326 2130 72378
rect 2142 72326 2194 72378
rect 2206 72326 2258 72378
rect 6950 72326 7002 72378
rect 7014 72326 7066 72378
rect 7078 72326 7130 72378
rect 7142 72326 7194 72378
rect 7206 72326 7258 72378
rect 11950 72326 12002 72378
rect 12014 72326 12066 72378
rect 12078 72326 12130 72378
rect 12142 72326 12194 72378
rect 12206 72326 12258 72378
rect 16950 72326 17002 72378
rect 17014 72326 17066 72378
rect 17078 72326 17130 72378
rect 17142 72326 17194 72378
rect 17206 72326 17258 72378
rect 16672 72224 16724 72276
rect 16856 72020 16908 72072
rect 16580 71884 16632 71936
rect 16856 71884 16908 71936
rect 2610 71782 2662 71834
rect 2674 71782 2726 71834
rect 2738 71782 2790 71834
rect 2802 71782 2854 71834
rect 2866 71782 2918 71834
rect 7610 71782 7662 71834
rect 7674 71782 7726 71834
rect 7738 71782 7790 71834
rect 7802 71782 7854 71834
rect 7866 71782 7918 71834
rect 12610 71782 12662 71834
rect 12674 71782 12726 71834
rect 12738 71782 12790 71834
rect 12802 71782 12854 71834
rect 12866 71782 12918 71834
rect 17610 71782 17662 71834
rect 17674 71782 17726 71834
rect 17738 71782 17790 71834
rect 17802 71782 17854 71834
rect 17866 71782 17918 71834
rect 12440 71680 12492 71732
rect 18972 71680 19024 71732
rect 5540 71612 5592 71664
rect 3332 71587 3384 71596
rect 3332 71553 3366 71587
rect 3366 71553 3384 71587
rect 3332 71544 3384 71553
rect 15660 71544 15712 71596
rect 8208 71340 8260 71392
rect 18236 71383 18288 71392
rect 18236 71349 18245 71383
rect 18245 71349 18279 71383
rect 18279 71349 18288 71383
rect 18236 71340 18288 71349
rect 1950 71238 2002 71290
rect 2014 71238 2066 71290
rect 2078 71238 2130 71290
rect 2142 71238 2194 71290
rect 2206 71238 2258 71290
rect 6950 71238 7002 71290
rect 7014 71238 7066 71290
rect 7078 71238 7130 71290
rect 7142 71238 7194 71290
rect 7206 71238 7258 71290
rect 11950 71238 12002 71290
rect 12014 71238 12066 71290
rect 12078 71238 12130 71290
rect 12142 71238 12194 71290
rect 12206 71238 12258 71290
rect 16950 71238 17002 71290
rect 17014 71238 17066 71290
rect 17078 71238 17130 71290
rect 17142 71238 17194 71290
rect 17206 71238 17258 71290
rect 6276 71136 6328 71188
rect 15200 71136 15252 71188
rect 10508 71111 10560 71120
rect 10508 71077 10517 71111
rect 10517 71077 10551 71111
rect 10551 71077 10560 71111
rect 10508 71068 10560 71077
rect 5540 71000 5592 71052
rect 6828 70932 6880 70984
rect 9128 70975 9180 70984
rect 9128 70941 9137 70975
rect 9137 70941 9171 70975
rect 9171 70941 9180 70975
rect 9128 70932 9180 70941
rect 9864 70932 9916 70984
rect 14280 70932 14332 70984
rect 6276 70907 6328 70916
rect 6276 70873 6310 70907
rect 6310 70873 6328 70907
rect 6276 70864 6328 70873
rect 1124 70796 1176 70848
rect 15752 70907 15804 70916
rect 15752 70873 15786 70907
rect 15786 70873 15804 70907
rect 15752 70864 15804 70873
rect 6552 70796 6604 70848
rect 9036 70796 9088 70848
rect 16672 70796 16724 70848
rect 2610 70694 2662 70746
rect 2674 70694 2726 70746
rect 2738 70694 2790 70746
rect 2802 70694 2854 70746
rect 2866 70694 2918 70746
rect 7610 70694 7662 70746
rect 7674 70694 7726 70746
rect 7738 70694 7790 70746
rect 7802 70694 7854 70746
rect 7866 70694 7918 70746
rect 12610 70694 12662 70746
rect 12674 70694 12726 70746
rect 12738 70694 12790 70746
rect 12802 70694 12854 70746
rect 12866 70694 12918 70746
rect 17610 70694 17662 70746
rect 17674 70694 17726 70746
rect 17738 70694 17790 70746
rect 17802 70694 17854 70746
rect 17866 70694 17918 70746
rect 1950 70150 2002 70202
rect 2014 70150 2066 70202
rect 2078 70150 2130 70202
rect 2142 70150 2194 70202
rect 2206 70150 2258 70202
rect 6950 70150 7002 70202
rect 7014 70150 7066 70202
rect 7078 70150 7130 70202
rect 7142 70150 7194 70202
rect 7206 70150 7258 70202
rect 11950 70150 12002 70202
rect 12014 70150 12066 70202
rect 12078 70150 12130 70202
rect 12142 70150 12194 70202
rect 12206 70150 12258 70202
rect 16950 70150 17002 70202
rect 17014 70150 17066 70202
rect 17078 70150 17130 70202
rect 17142 70150 17194 70202
rect 17206 70150 17258 70202
rect 2044 70023 2096 70032
rect 2044 69989 2053 70023
rect 2053 69989 2087 70023
rect 2087 69989 2096 70023
rect 2044 69980 2096 69989
rect 16672 70048 16724 70100
rect 12440 69912 12492 69964
rect 13728 69912 13780 69964
rect 2964 69844 3016 69896
rect 3976 69887 4028 69896
rect 3976 69853 3985 69887
rect 3985 69853 4019 69887
rect 4019 69853 4028 69887
rect 3976 69844 4028 69853
rect 7012 69844 7064 69896
rect 8300 69844 8352 69896
rect 9312 69844 9364 69896
rect 15016 69887 15068 69896
rect 15016 69853 15025 69887
rect 15025 69853 15059 69887
rect 15059 69853 15068 69887
rect 15016 69844 15068 69853
rect 15108 69844 15160 69896
rect 3792 69776 3844 69828
rect 6552 69776 6604 69828
rect 2504 69751 2556 69760
rect 2504 69717 2513 69751
rect 2513 69717 2547 69751
rect 2547 69717 2556 69751
rect 2504 69708 2556 69717
rect 5264 69708 5316 69760
rect 6644 69708 6696 69760
rect 6828 69708 6880 69760
rect 15476 69708 15528 69760
rect 18236 69751 18288 69760
rect 18236 69717 18245 69751
rect 18245 69717 18279 69751
rect 18279 69717 18288 69751
rect 18236 69708 18288 69717
rect 2610 69606 2662 69658
rect 2674 69606 2726 69658
rect 2738 69606 2790 69658
rect 2802 69606 2854 69658
rect 2866 69606 2918 69658
rect 7610 69606 7662 69658
rect 7674 69606 7726 69658
rect 7738 69606 7790 69658
rect 7802 69606 7854 69658
rect 7866 69606 7918 69658
rect 12610 69606 12662 69658
rect 12674 69606 12726 69658
rect 12738 69606 12790 69658
rect 12802 69606 12854 69658
rect 12866 69606 12918 69658
rect 17610 69606 17662 69658
rect 17674 69606 17726 69658
rect 17738 69606 17790 69658
rect 17802 69606 17854 69658
rect 17866 69606 17918 69658
rect 3976 69436 4028 69488
rect 13176 69504 13228 69556
rect 7472 69436 7524 69488
rect 9128 69368 9180 69420
rect 11060 69207 11112 69216
rect 11060 69173 11069 69207
rect 11069 69173 11103 69207
rect 11103 69173 11112 69207
rect 11060 69164 11112 69173
rect 1950 69062 2002 69114
rect 2014 69062 2066 69114
rect 2078 69062 2130 69114
rect 2142 69062 2194 69114
rect 2206 69062 2258 69114
rect 6950 69062 7002 69114
rect 7014 69062 7066 69114
rect 7078 69062 7130 69114
rect 7142 69062 7194 69114
rect 7206 69062 7258 69114
rect 11950 69062 12002 69114
rect 12014 69062 12066 69114
rect 12078 69062 12130 69114
rect 12142 69062 12194 69114
rect 12206 69062 12258 69114
rect 16950 69062 17002 69114
rect 17014 69062 17066 69114
rect 17078 69062 17130 69114
rect 17142 69062 17194 69114
rect 17206 69062 17258 69114
rect 9128 68867 9180 68876
rect 9128 68833 9137 68867
rect 9137 68833 9171 68867
rect 9171 68833 9180 68867
rect 9128 68824 9180 68833
rect 13820 68756 13872 68808
rect 14280 68799 14332 68808
rect 14280 68765 14289 68799
rect 14289 68765 14323 68799
rect 14323 68765 14332 68799
rect 14280 68756 14332 68765
rect 9588 68688 9640 68740
rect 14556 68731 14608 68740
rect 14556 68697 14590 68731
rect 14590 68697 14608 68731
rect 14556 68688 14608 68697
rect 10508 68663 10560 68672
rect 10508 68629 10517 68663
rect 10517 68629 10551 68663
rect 10551 68629 10560 68663
rect 10508 68620 10560 68629
rect 15660 68663 15712 68672
rect 15660 68629 15669 68663
rect 15669 68629 15703 68663
rect 15703 68629 15712 68663
rect 15660 68620 15712 68629
rect 2610 68518 2662 68570
rect 2674 68518 2726 68570
rect 2738 68518 2790 68570
rect 2802 68518 2854 68570
rect 2866 68518 2918 68570
rect 7610 68518 7662 68570
rect 7674 68518 7726 68570
rect 7738 68518 7790 68570
rect 7802 68518 7854 68570
rect 7866 68518 7918 68570
rect 12610 68518 12662 68570
rect 12674 68518 12726 68570
rect 12738 68518 12790 68570
rect 12802 68518 12854 68570
rect 12866 68518 12918 68570
rect 17610 68518 17662 68570
rect 17674 68518 17726 68570
rect 17738 68518 17790 68570
rect 17802 68518 17854 68570
rect 17866 68518 17918 68570
rect 6184 68280 6236 68332
rect 14924 68280 14976 68332
rect 1950 67974 2002 68026
rect 2014 67974 2066 68026
rect 2078 67974 2130 68026
rect 2142 67974 2194 68026
rect 2206 67974 2258 68026
rect 6950 67974 7002 68026
rect 7014 67974 7066 68026
rect 7078 67974 7130 68026
rect 7142 67974 7194 68026
rect 7206 67974 7258 68026
rect 11950 67974 12002 68026
rect 12014 67974 12066 68026
rect 12078 67974 12130 68026
rect 12142 67974 12194 68026
rect 12206 67974 12258 68026
rect 16950 67974 17002 68026
rect 17014 67974 17066 68026
rect 17078 67974 17130 68026
rect 17142 67974 17194 68026
rect 17206 67974 17258 68026
rect 10416 67804 10468 67856
rect 18236 67847 18288 67856
rect 18236 67813 18245 67847
rect 18245 67813 18279 67847
rect 18279 67813 18288 67847
rect 18236 67804 18288 67813
rect 17408 67668 17460 67720
rect 12072 67643 12124 67652
rect 12072 67609 12081 67643
rect 12081 67609 12115 67643
rect 12115 67609 12124 67643
rect 12072 67600 12124 67609
rect 2610 67430 2662 67482
rect 2674 67430 2726 67482
rect 2738 67430 2790 67482
rect 2802 67430 2854 67482
rect 2866 67430 2918 67482
rect 7610 67430 7662 67482
rect 7674 67430 7726 67482
rect 7738 67430 7790 67482
rect 7802 67430 7854 67482
rect 7866 67430 7918 67482
rect 12610 67430 12662 67482
rect 12674 67430 12726 67482
rect 12738 67430 12790 67482
rect 12802 67430 12854 67482
rect 12866 67430 12918 67482
rect 17610 67430 17662 67482
rect 17674 67430 17726 67482
rect 17738 67430 17790 67482
rect 17802 67430 17854 67482
rect 17866 67430 17918 67482
rect 11796 67260 11848 67312
rect 3700 67192 3752 67244
rect 14004 67192 14056 67244
rect 16028 67124 16080 67176
rect 16488 67124 16540 67176
rect 1216 66988 1268 67040
rect 17316 66988 17368 67040
rect 1950 66886 2002 66938
rect 2014 66886 2066 66938
rect 2078 66886 2130 66938
rect 2142 66886 2194 66938
rect 2206 66886 2258 66938
rect 6950 66886 7002 66938
rect 7014 66886 7066 66938
rect 7078 66886 7130 66938
rect 7142 66886 7194 66938
rect 7206 66886 7258 66938
rect 11950 66886 12002 66938
rect 12014 66886 12066 66938
rect 12078 66886 12130 66938
rect 12142 66886 12194 66938
rect 12206 66886 12258 66938
rect 16950 66886 17002 66938
rect 17014 66886 17066 66938
rect 17078 66886 17130 66938
rect 17142 66886 17194 66938
rect 17206 66886 17258 66938
rect 2610 66342 2662 66394
rect 2674 66342 2726 66394
rect 2738 66342 2790 66394
rect 2802 66342 2854 66394
rect 2866 66342 2918 66394
rect 7610 66342 7662 66394
rect 7674 66342 7726 66394
rect 7738 66342 7790 66394
rect 7802 66342 7854 66394
rect 7866 66342 7918 66394
rect 12610 66342 12662 66394
rect 12674 66342 12726 66394
rect 12738 66342 12790 66394
rect 12802 66342 12854 66394
rect 12866 66342 12918 66394
rect 17610 66342 17662 66394
rect 17674 66342 17726 66394
rect 17738 66342 17790 66394
rect 17802 66342 17854 66394
rect 17866 66342 17918 66394
rect 13912 66172 13964 66224
rect 16580 66172 16632 66224
rect 17500 66172 17552 66224
rect 13636 66104 13688 66156
rect 17408 66104 17460 66156
rect 14280 65900 14332 65952
rect 14832 65900 14884 65952
rect 17500 65943 17552 65952
rect 17500 65909 17509 65943
rect 17509 65909 17543 65943
rect 17543 65909 17552 65943
rect 17500 65900 17552 65909
rect 1950 65798 2002 65850
rect 2014 65798 2066 65850
rect 2078 65798 2130 65850
rect 2142 65798 2194 65850
rect 2206 65798 2258 65850
rect 6950 65798 7002 65850
rect 7014 65798 7066 65850
rect 7078 65798 7130 65850
rect 7142 65798 7194 65850
rect 7206 65798 7258 65850
rect 11950 65798 12002 65850
rect 12014 65798 12066 65850
rect 12078 65798 12130 65850
rect 12142 65798 12194 65850
rect 12206 65798 12258 65850
rect 16950 65798 17002 65850
rect 17014 65798 17066 65850
rect 17078 65798 17130 65850
rect 17142 65798 17194 65850
rect 17206 65798 17258 65850
rect 4068 65671 4120 65680
rect 4068 65637 4077 65671
rect 4077 65637 4111 65671
rect 4111 65637 4120 65671
rect 4068 65628 4120 65637
rect 11796 65628 11848 65680
rect 18236 65671 18288 65680
rect 18236 65637 18245 65671
rect 18245 65637 18279 65671
rect 18279 65637 18288 65671
rect 18236 65628 18288 65637
rect 4620 65603 4672 65612
rect 4620 65569 4629 65603
rect 4629 65569 4663 65603
rect 4663 65569 4672 65603
rect 4620 65560 4672 65569
rect 11520 65560 11572 65612
rect 11796 65535 11848 65544
rect 11796 65501 11805 65535
rect 11805 65501 11839 65535
rect 11839 65501 11848 65535
rect 11796 65492 11848 65501
rect 11888 65535 11940 65544
rect 11888 65501 11897 65535
rect 11897 65501 11931 65535
rect 11931 65501 11940 65535
rect 11888 65492 11940 65501
rect 15568 65492 15620 65544
rect 16212 65492 16264 65544
rect 9496 65424 9548 65476
rect 11428 65424 11480 65476
rect 3608 65356 3660 65408
rect 2610 65254 2662 65306
rect 2674 65254 2726 65306
rect 2738 65254 2790 65306
rect 2802 65254 2854 65306
rect 2866 65254 2918 65306
rect 7610 65254 7662 65306
rect 7674 65254 7726 65306
rect 7738 65254 7790 65306
rect 7802 65254 7854 65306
rect 7866 65254 7918 65306
rect 12610 65254 12662 65306
rect 12674 65254 12726 65306
rect 12738 65254 12790 65306
rect 12802 65254 12854 65306
rect 12866 65254 12918 65306
rect 17610 65254 17662 65306
rect 17674 65254 17726 65306
rect 17738 65254 17790 65306
rect 17802 65254 17854 65306
rect 17866 65254 17918 65306
rect 8300 65152 8352 65204
rect 14372 65195 14424 65204
rect 14372 65161 14381 65195
rect 14381 65161 14415 65195
rect 14415 65161 14424 65195
rect 14372 65152 14424 65161
rect 15108 65152 15160 65204
rect 17408 65152 17460 65204
rect 17592 65152 17644 65204
rect 19156 65084 19208 65136
rect 7932 65016 7984 65068
rect 8668 65016 8720 65068
rect 19340 65016 19392 65068
rect 8300 64880 8352 64932
rect 12440 64948 12492 65000
rect 11888 64880 11940 64932
rect 17040 64880 17092 64932
rect 17408 64880 17460 64932
rect 18420 64880 18472 64932
rect 13728 64812 13780 64864
rect 16488 64812 16540 64864
rect 16948 64812 17000 64864
rect 1950 64710 2002 64762
rect 2014 64710 2066 64762
rect 2078 64710 2130 64762
rect 2142 64710 2194 64762
rect 2206 64710 2258 64762
rect 6950 64710 7002 64762
rect 7014 64710 7066 64762
rect 7078 64710 7130 64762
rect 7142 64710 7194 64762
rect 7206 64710 7258 64762
rect 11950 64710 12002 64762
rect 12014 64710 12066 64762
rect 12078 64710 12130 64762
rect 12142 64710 12194 64762
rect 12206 64710 12258 64762
rect 16950 64710 17002 64762
rect 17014 64710 17066 64762
rect 17078 64710 17130 64762
rect 17142 64710 17194 64762
rect 17206 64710 17258 64762
rect 13268 64608 13320 64660
rect 8116 64472 8168 64524
rect 8392 64472 8444 64524
rect 7288 64404 7340 64456
rect 13728 64404 13780 64456
rect 11336 64336 11388 64388
rect 1768 64268 1820 64320
rect 7932 64268 7984 64320
rect 8116 64268 8168 64320
rect 13912 64268 13964 64320
rect 2610 64166 2662 64218
rect 2674 64166 2726 64218
rect 2738 64166 2790 64218
rect 2802 64166 2854 64218
rect 2866 64166 2918 64218
rect 7610 64166 7662 64218
rect 7674 64166 7726 64218
rect 7738 64166 7790 64218
rect 7802 64166 7854 64218
rect 7866 64166 7918 64218
rect 12610 64166 12662 64218
rect 12674 64166 12726 64218
rect 12738 64166 12790 64218
rect 12802 64166 12854 64218
rect 12866 64166 12918 64218
rect 17610 64166 17662 64218
rect 17674 64166 17726 64218
rect 17738 64166 17790 64218
rect 17802 64166 17854 64218
rect 17866 64166 17918 64218
rect 11244 63928 11296 63980
rect 18512 63928 18564 63980
rect 9680 63792 9732 63844
rect 9956 63724 10008 63776
rect 15384 63860 15436 63912
rect 18236 63767 18288 63776
rect 18236 63733 18245 63767
rect 18245 63733 18279 63767
rect 18279 63733 18288 63767
rect 18236 63724 18288 63733
rect 1950 63622 2002 63674
rect 2014 63622 2066 63674
rect 2078 63622 2130 63674
rect 2142 63622 2194 63674
rect 2206 63622 2258 63674
rect 6950 63622 7002 63674
rect 7014 63622 7066 63674
rect 7078 63622 7130 63674
rect 7142 63622 7194 63674
rect 7206 63622 7258 63674
rect 11950 63622 12002 63674
rect 12014 63622 12066 63674
rect 12078 63622 12130 63674
rect 12142 63622 12194 63674
rect 12206 63622 12258 63674
rect 16950 63622 17002 63674
rect 17014 63622 17066 63674
rect 17078 63622 17130 63674
rect 17142 63622 17194 63674
rect 17206 63622 17258 63674
rect 13912 63520 13964 63572
rect 14924 63520 14976 63572
rect 6552 63452 6604 63504
rect 7288 63452 7340 63504
rect 14556 63452 14608 63504
rect 15568 63316 15620 63368
rect 16488 63359 16540 63368
rect 16488 63325 16497 63359
rect 16497 63325 16531 63359
rect 16531 63325 16540 63359
rect 16488 63316 16540 63325
rect 9680 63248 9732 63300
rect 6368 63223 6420 63232
rect 6368 63189 6377 63223
rect 6377 63189 6411 63223
rect 6411 63189 6420 63223
rect 6368 63180 6420 63189
rect 14464 63223 14516 63232
rect 14464 63189 14473 63223
rect 14473 63189 14507 63223
rect 14507 63189 14516 63223
rect 14464 63180 14516 63189
rect 2610 63078 2662 63130
rect 2674 63078 2726 63130
rect 2738 63078 2790 63130
rect 2802 63078 2854 63130
rect 2866 63078 2918 63130
rect 7610 63078 7662 63130
rect 7674 63078 7726 63130
rect 7738 63078 7790 63130
rect 7802 63078 7854 63130
rect 7866 63078 7918 63130
rect 12610 63078 12662 63130
rect 12674 63078 12726 63130
rect 12738 63078 12790 63130
rect 12802 63078 12854 63130
rect 12866 63078 12918 63130
rect 17610 63078 17662 63130
rect 17674 63078 17726 63130
rect 17738 63078 17790 63130
rect 17802 63078 17854 63130
rect 17866 63078 17918 63130
rect 5448 62976 5500 63028
rect 11152 62976 11204 63028
rect 6552 62883 6604 62892
rect 6552 62849 6561 62883
rect 6561 62849 6595 62883
rect 6595 62849 6604 62883
rect 6552 62840 6604 62849
rect 9588 62772 9640 62824
rect 19064 62772 19116 62824
rect 8760 62679 8812 62688
rect 8760 62645 8769 62679
rect 8769 62645 8803 62679
rect 8803 62645 8812 62679
rect 8760 62636 8812 62645
rect 1950 62534 2002 62586
rect 2014 62534 2066 62586
rect 2078 62534 2130 62586
rect 2142 62534 2194 62586
rect 2206 62534 2258 62586
rect 6950 62534 7002 62586
rect 7014 62534 7066 62586
rect 7078 62534 7130 62586
rect 7142 62534 7194 62586
rect 7206 62534 7258 62586
rect 11950 62534 12002 62586
rect 12014 62534 12066 62586
rect 12078 62534 12130 62586
rect 12142 62534 12194 62586
rect 12206 62534 12258 62586
rect 16950 62534 17002 62586
rect 17014 62534 17066 62586
rect 17078 62534 17130 62586
rect 17142 62534 17194 62586
rect 17206 62534 17258 62586
rect 4160 62432 4212 62484
rect 13820 62432 13872 62484
rect 11152 62364 11204 62416
rect 11796 62364 11848 62416
rect 18604 62228 18656 62280
rect 4252 62203 4304 62212
rect 4252 62169 4261 62203
rect 4261 62169 4295 62203
rect 4295 62169 4304 62203
rect 4252 62160 4304 62169
rect 4344 62135 4396 62144
rect 4344 62101 4353 62135
rect 4353 62101 4387 62135
rect 4387 62101 4396 62135
rect 4344 62092 4396 62101
rect 18236 62135 18288 62144
rect 18236 62101 18245 62135
rect 18245 62101 18279 62135
rect 18279 62101 18288 62135
rect 18236 62092 18288 62101
rect 2610 61990 2662 62042
rect 2674 61990 2726 62042
rect 2738 61990 2790 62042
rect 2802 61990 2854 62042
rect 2866 61990 2918 62042
rect 7610 61990 7662 62042
rect 7674 61990 7726 62042
rect 7738 61990 7790 62042
rect 7802 61990 7854 62042
rect 7866 61990 7918 62042
rect 12610 61990 12662 62042
rect 12674 61990 12726 62042
rect 12738 61990 12790 62042
rect 12802 61990 12854 62042
rect 12866 61990 12918 62042
rect 17610 61990 17662 62042
rect 17674 61990 17726 62042
rect 17738 61990 17790 62042
rect 17802 61990 17854 62042
rect 17866 61990 17918 62042
rect 16488 61888 16540 61940
rect 15660 61820 15712 61872
rect 11612 61684 11664 61736
rect 12348 61752 12400 61804
rect 13544 61684 13596 61736
rect 14280 61684 14332 61736
rect 1950 61446 2002 61498
rect 2014 61446 2066 61498
rect 2078 61446 2130 61498
rect 2142 61446 2194 61498
rect 2206 61446 2258 61498
rect 6950 61446 7002 61498
rect 7014 61446 7066 61498
rect 7078 61446 7130 61498
rect 7142 61446 7194 61498
rect 7206 61446 7258 61498
rect 11950 61446 12002 61498
rect 12014 61446 12066 61498
rect 12078 61446 12130 61498
rect 12142 61446 12194 61498
rect 12206 61446 12258 61498
rect 16950 61446 17002 61498
rect 17014 61446 17066 61498
rect 17078 61446 17130 61498
rect 17142 61446 17194 61498
rect 17206 61446 17258 61498
rect 4804 61344 4856 61396
rect 16212 61344 16264 61396
rect 13820 61140 13872 61192
rect 14280 61140 14332 61192
rect 16212 61115 16264 61124
rect 16212 61081 16246 61115
rect 16246 61081 16264 61115
rect 16212 61072 16264 61081
rect 17960 61004 18012 61056
rect 2610 60902 2662 60954
rect 2674 60902 2726 60954
rect 2738 60902 2790 60954
rect 2802 60902 2854 60954
rect 2866 60902 2918 60954
rect 7610 60902 7662 60954
rect 7674 60902 7726 60954
rect 7738 60902 7790 60954
rect 7802 60902 7854 60954
rect 7866 60902 7918 60954
rect 12610 60902 12662 60954
rect 12674 60902 12726 60954
rect 12738 60902 12790 60954
rect 12802 60902 12854 60954
rect 12866 60902 12918 60954
rect 17610 60902 17662 60954
rect 17674 60902 17726 60954
rect 17738 60902 17790 60954
rect 17802 60902 17854 60954
rect 17866 60902 17918 60954
rect 8484 60732 8536 60784
rect 9496 60775 9548 60784
rect 9496 60741 9505 60775
rect 9505 60741 9539 60775
rect 9539 60741 9548 60775
rect 9496 60732 9548 60741
rect 6552 60707 6604 60716
rect 6552 60673 6561 60707
rect 6561 60673 6595 60707
rect 6595 60673 6604 60707
rect 6552 60664 6604 60673
rect 5908 60639 5960 60648
rect 5908 60605 5917 60639
rect 5917 60605 5951 60639
rect 5951 60605 5960 60639
rect 5908 60596 5960 60605
rect 9404 60639 9456 60648
rect 9404 60605 9413 60639
rect 9413 60605 9447 60639
rect 9447 60605 9456 60639
rect 9404 60596 9456 60605
rect 4620 60460 4672 60512
rect 10968 60528 11020 60580
rect 7932 60503 7984 60512
rect 7932 60469 7941 60503
rect 7941 60469 7975 60503
rect 7975 60469 7984 60503
rect 7932 60460 7984 60469
rect 8024 60460 8076 60512
rect 1950 60358 2002 60410
rect 2014 60358 2066 60410
rect 2078 60358 2130 60410
rect 2142 60358 2194 60410
rect 2206 60358 2258 60410
rect 6950 60358 7002 60410
rect 7014 60358 7066 60410
rect 7078 60358 7130 60410
rect 7142 60358 7194 60410
rect 7206 60358 7258 60410
rect 11950 60358 12002 60410
rect 12014 60358 12066 60410
rect 12078 60358 12130 60410
rect 12142 60358 12194 60410
rect 12206 60358 12258 60410
rect 16950 60358 17002 60410
rect 17014 60358 17066 60410
rect 17078 60358 17130 60410
rect 17142 60358 17194 60410
rect 17206 60358 17258 60410
rect 1032 60256 1084 60308
rect 8024 60256 8076 60308
rect 13176 60256 13228 60308
rect 10508 60188 10560 60240
rect 16488 60188 16540 60240
rect 7196 60120 7248 60172
rect 8116 60120 8168 60172
rect 10784 60120 10836 60172
rect 15476 60120 15528 60172
rect 16396 60120 16448 60172
rect 6276 59984 6328 60036
rect 6828 59984 6880 60036
rect 8116 59984 8168 60036
rect 13084 59984 13136 60036
rect 7288 59916 7340 59968
rect 9588 59959 9640 59968
rect 9588 59925 9597 59959
rect 9597 59925 9631 59959
rect 9631 59925 9640 59959
rect 9588 59916 9640 59925
rect 14280 60095 14332 60104
rect 14280 60061 14289 60095
rect 14289 60061 14323 60095
rect 14323 60061 14332 60095
rect 14280 60052 14332 60061
rect 15384 60052 15436 60104
rect 19248 60052 19300 60104
rect 14556 60027 14608 60036
rect 14556 59993 14590 60027
rect 14590 59993 14608 60027
rect 14556 59984 14608 59993
rect 16120 59916 16172 59968
rect 18236 59959 18288 59968
rect 18236 59925 18245 59959
rect 18245 59925 18279 59959
rect 18279 59925 18288 59959
rect 18236 59916 18288 59925
rect 2610 59814 2662 59866
rect 2674 59814 2726 59866
rect 2738 59814 2790 59866
rect 2802 59814 2854 59866
rect 2866 59814 2918 59866
rect 7610 59814 7662 59866
rect 7674 59814 7726 59866
rect 7738 59814 7790 59866
rect 7802 59814 7854 59866
rect 7866 59814 7918 59866
rect 12610 59814 12662 59866
rect 12674 59814 12726 59866
rect 12738 59814 12790 59866
rect 12802 59814 12854 59866
rect 12866 59814 12918 59866
rect 17610 59814 17662 59866
rect 17674 59814 17726 59866
rect 17738 59814 17790 59866
rect 17802 59814 17854 59866
rect 17866 59814 17918 59866
rect 6552 59644 6604 59696
rect 7196 59644 7248 59696
rect 8208 59644 8260 59696
rect 3240 59619 3292 59628
rect 3240 59585 3249 59619
rect 3249 59585 3283 59619
rect 3283 59585 3292 59619
rect 3240 59576 3292 59585
rect 5172 59372 5224 59424
rect 1950 59270 2002 59322
rect 2014 59270 2066 59322
rect 2078 59270 2130 59322
rect 2142 59270 2194 59322
rect 2206 59270 2258 59322
rect 6950 59270 7002 59322
rect 7014 59270 7066 59322
rect 7078 59270 7130 59322
rect 7142 59270 7194 59322
rect 7206 59270 7258 59322
rect 11950 59270 12002 59322
rect 12014 59270 12066 59322
rect 12078 59270 12130 59322
rect 12142 59270 12194 59322
rect 12206 59270 12258 59322
rect 16950 59270 17002 59322
rect 17014 59270 17066 59322
rect 17078 59270 17130 59322
rect 17142 59270 17194 59322
rect 17206 59270 17258 59322
rect 15200 59075 15252 59084
rect 15200 59041 15209 59075
rect 15209 59041 15243 59075
rect 15243 59041 15252 59075
rect 15200 59032 15252 59041
rect 15384 59075 15436 59084
rect 15384 59041 15393 59075
rect 15393 59041 15427 59075
rect 15427 59041 15436 59075
rect 15384 59032 15436 59041
rect 4068 58964 4120 59016
rect 18880 58964 18932 59016
rect 15292 58939 15344 58948
rect 15292 58905 15301 58939
rect 15301 58905 15335 58939
rect 15335 58905 15344 58939
rect 15292 58896 15344 58905
rect 15476 58896 15528 58948
rect 13728 58871 13780 58880
rect 13728 58837 13737 58871
rect 13737 58837 13771 58871
rect 13771 58837 13780 58871
rect 13728 58828 13780 58837
rect 2610 58726 2662 58778
rect 2674 58726 2726 58778
rect 2738 58726 2790 58778
rect 2802 58726 2854 58778
rect 2866 58726 2918 58778
rect 7610 58726 7662 58778
rect 7674 58726 7726 58778
rect 7738 58726 7790 58778
rect 7802 58726 7854 58778
rect 7866 58726 7918 58778
rect 12610 58726 12662 58778
rect 12674 58726 12726 58778
rect 12738 58726 12790 58778
rect 12802 58726 12854 58778
rect 12866 58726 12918 58778
rect 17610 58726 17662 58778
rect 17674 58726 17726 58778
rect 17738 58726 17790 58778
rect 17802 58726 17854 58778
rect 17866 58726 17918 58778
rect 16672 58488 16724 58540
rect 18236 58327 18288 58336
rect 18236 58293 18245 58327
rect 18245 58293 18279 58327
rect 18279 58293 18288 58327
rect 18236 58284 18288 58293
rect 1950 58182 2002 58234
rect 2014 58182 2066 58234
rect 2078 58182 2130 58234
rect 2142 58182 2194 58234
rect 2206 58182 2258 58234
rect 6950 58182 7002 58234
rect 7014 58182 7066 58234
rect 7078 58182 7130 58234
rect 7142 58182 7194 58234
rect 7206 58182 7258 58234
rect 11950 58182 12002 58234
rect 12014 58182 12066 58234
rect 12078 58182 12130 58234
rect 12142 58182 12194 58234
rect 12206 58182 12258 58234
rect 16950 58182 17002 58234
rect 17014 58182 17066 58234
rect 17078 58182 17130 58234
rect 17142 58182 17194 58234
rect 17206 58182 17258 58234
rect 2320 57740 2372 57792
rect 8116 57740 8168 57792
rect 10048 57740 10100 57792
rect 2610 57638 2662 57690
rect 2674 57638 2726 57690
rect 2738 57638 2790 57690
rect 2802 57638 2854 57690
rect 2866 57638 2918 57690
rect 7610 57638 7662 57690
rect 7674 57638 7726 57690
rect 7738 57638 7790 57690
rect 7802 57638 7854 57690
rect 7866 57638 7918 57690
rect 12610 57638 12662 57690
rect 12674 57638 12726 57690
rect 12738 57638 12790 57690
rect 12802 57638 12854 57690
rect 12866 57638 12918 57690
rect 17610 57638 17662 57690
rect 17674 57638 17726 57690
rect 17738 57638 17790 57690
rect 17802 57638 17854 57690
rect 17866 57638 17918 57690
rect 8116 57536 8168 57588
rect 8392 57536 8444 57588
rect 15568 57536 15620 57588
rect 3240 57468 3292 57520
rect 4988 57468 5040 57520
rect 16580 57468 16632 57520
rect 3056 57443 3108 57452
rect 3056 57409 3090 57443
rect 3090 57409 3108 57443
rect 3056 57400 3108 57409
rect 16856 57400 16908 57452
rect 15292 57332 15344 57384
rect 17408 57264 17460 57316
rect 4160 57239 4212 57248
rect 4160 57205 4169 57239
rect 4169 57205 4203 57239
rect 4203 57205 4212 57239
rect 4160 57196 4212 57205
rect 8300 57196 8352 57248
rect 1950 57094 2002 57146
rect 2014 57094 2066 57146
rect 2078 57094 2130 57146
rect 2142 57094 2194 57146
rect 2206 57094 2258 57146
rect 6950 57094 7002 57146
rect 7014 57094 7066 57146
rect 7078 57094 7130 57146
rect 7142 57094 7194 57146
rect 7206 57094 7258 57146
rect 11950 57094 12002 57146
rect 12014 57094 12066 57146
rect 12078 57094 12130 57146
rect 12142 57094 12194 57146
rect 12206 57094 12258 57146
rect 16950 57094 17002 57146
rect 17014 57094 17066 57146
rect 17078 57094 17130 57146
rect 17142 57094 17194 57146
rect 17206 57094 17258 57146
rect 4160 56992 4212 57044
rect 13176 56992 13228 57044
rect 3516 56924 3568 56976
rect 1492 56856 1544 56908
rect 2320 56856 2372 56908
rect 2412 56652 2464 56704
rect 17960 56652 18012 56704
rect 2610 56550 2662 56602
rect 2674 56550 2726 56602
rect 2738 56550 2790 56602
rect 2802 56550 2854 56602
rect 2866 56550 2918 56602
rect 7610 56550 7662 56602
rect 7674 56550 7726 56602
rect 7738 56550 7790 56602
rect 7802 56550 7854 56602
rect 7866 56550 7918 56602
rect 12610 56550 12662 56602
rect 12674 56550 12726 56602
rect 12738 56550 12790 56602
rect 12802 56550 12854 56602
rect 12866 56550 12918 56602
rect 17610 56550 17662 56602
rect 17674 56550 17726 56602
rect 17738 56550 17790 56602
rect 17802 56550 17854 56602
rect 17866 56550 17918 56602
rect 1676 56312 1728 56364
rect 940 56176 992 56228
rect 2964 56312 3016 56364
rect 3240 56312 3292 56364
rect 8116 56312 8168 56364
rect 12440 56287 12492 56296
rect 12440 56253 12449 56287
rect 12449 56253 12483 56287
rect 12483 56253 12492 56287
rect 12440 56244 12492 56253
rect 12992 56244 13044 56296
rect 2320 56151 2372 56160
rect 2320 56117 2329 56151
rect 2329 56117 2363 56151
rect 2363 56117 2372 56151
rect 2320 56108 2372 56117
rect 4528 56151 4580 56160
rect 4528 56117 4537 56151
rect 4537 56117 4571 56151
rect 4571 56117 4580 56151
rect 4528 56108 4580 56117
rect 18236 56151 18288 56160
rect 18236 56117 18245 56151
rect 18245 56117 18279 56151
rect 18279 56117 18288 56151
rect 18236 56108 18288 56117
rect 1950 56006 2002 56058
rect 2014 56006 2066 56058
rect 2078 56006 2130 56058
rect 2142 56006 2194 56058
rect 2206 56006 2258 56058
rect 6950 56006 7002 56058
rect 7014 56006 7066 56058
rect 7078 56006 7130 56058
rect 7142 56006 7194 56058
rect 7206 56006 7258 56058
rect 11950 56006 12002 56058
rect 12014 56006 12066 56058
rect 12078 56006 12130 56058
rect 12142 56006 12194 56058
rect 12206 56006 12258 56058
rect 16950 56006 17002 56058
rect 17014 56006 17066 56058
rect 17078 56006 17130 56058
rect 17142 56006 17194 56058
rect 17206 56006 17258 56058
rect 4896 55836 4948 55888
rect 11704 55836 11756 55888
rect 10968 55768 11020 55820
rect 2964 55700 3016 55752
rect 11704 55700 11756 55752
rect 848 55632 900 55684
rect 17132 55632 17184 55684
rect 10232 55564 10284 55616
rect 2610 55462 2662 55514
rect 2674 55462 2726 55514
rect 2738 55462 2790 55514
rect 2802 55462 2854 55514
rect 2866 55462 2918 55514
rect 7610 55462 7662 55514
rect 7674 55462 7726 55514
rect 7738 55462 7790 55514
rect 7802 55462 7854 55514
rect 7866 55462 7918 55514
rect 12610 55462 12662 55514
rect 12674 55462 12726 55514
rect 12738 55462 12790 55514
rect 12802 55462 12854 55514
rect 12866 55462 12918 55514
rect 17610 55462 17662 55514
rect 17674 55462 17726 55514
rect 17738 55462 17790 55514
rect 17802 55462 17854 55514
rect 17866 55462 17918 55514
rect 3608 55403 3660 55412
rect 3608 55369 3617 55403
rect 3617 55369 3651 55403
rect 3651 55369 3660 55403
rect 3608 55360 3660 55369
rect 5724 55360 5776 55412
rect 16856 55403 16908 55412
rect 16856 55369 16865 55403
rect 16865 55369 16899 55403
rect 16899 55369 16908 55403
rect 16856 55360 16908 55369
rect 2964 55292 3016 55344
rect 10416 55292 10468 55344
rect 16580 55292 16632 55344
rect 5540 55267 5592 55276
rect 5540 55233 5549 55267
rect 5549 55233 5583 55267
rect 5583 55233 5592 55267
rect 5540 55224 5592 55233
rect 5724 55267 5776 55276
rect 5724 55233 5733 55267
rect 5733 55233 5767 55267
rect 5767 55233 5776 55267
rect 6552 55267 6604 55276
rect 5724 55224 5776 55233
rect 6552 55233 6561 55267
rect 6561 55233 6595 55267
rect 6595 55233 6604 55267
rect 6552 55224 6604 55233
rect 16856 55224 16908 55276
rect 17132 55156 17184 55208
rect 1950 54918 2002 54970
rect 2014 54918 2066 54970
rect 2078 54918 2130 54970
rect 2142 54918 2194 54970
rect 2206 54918 2258 54970
rect 6950 54918 7002 54970
rect 7014 54918 7066 54970
rect 7078 54918 7130 54970
rect 7142 54918 7194 54970
rect 7206 54918 7258 54970
rect 11950 54918 12002 54970
rect 12014 54918 12066 54970
rect 12078 54918 12130 54970
rect 12142 54918 12194 54970
rect 12206 54918 12258 54970
rect 16950 54918 17002 54970
rect 17014 54918 17066 54970
rect 17078 54918 17130 54970
rect 17142 54918 17194 54970
rect 17206 54918 17258 54970
rect 18144 54612 18196 54664
rect 18236 54519 18288 54528
rect 18236 54485 18245 54519
rect 18245 54485 18279 54519
rect 18279 54485 18288 54519
rect 18236 54476 18288 54485
rect 2610 54374 2662 54426
rect 2674 54374 2726 54426
rect 2738 54374 2790 54426
rect 2802 54374 2854 54426
rect 2866 54374 2918 54426
rect 7610 54374 7662 54426
rect 7674 54374 7726 54426
rect 7738 54374 7790 54426
rect 7802 54374 7854 54426
rect 7866 54374 7918 54426
rect 12610 54374 12662 54426
rect 12674 54374 12726 54426
rect 12738 54374 12790 54426
rect 12802 54374 12854 54426
rect 12866 54374 12918 54426
rect 17610 54374 17662 54426
rect 17674 54374 17726 54426
rect 17738 54374 17790 54426
rect 17802 54374 17854 54426
rect 17866 54374 17918 54426
rect 8116 54272 8168 54324
rect 8392 54272 8444 54324
rect 11060 54272 11112 54324
rect 11428 54272 11480 54324
rect 7380 54136 7432 54188
rect 8116 54136 8168 54188
rect 10600 54179 10652 54188
rect 10600 54145 10609 54179
rect 10609 54145 10643 54179
rect 10643 54145 10652 54179
rect 10600 54136 10652 54145
rect 11060 54136 11112 54188
rect 11244 54136 11296 54188
rect 12440 54136 12492 54188
rect 10784 54068 10836 54120
rect 10968 54068 11020 54120
rect 7380 54000 7432 54052
rect 12532 53932 12584 53984
rect 1950 53830 2002 53882
rect 2014 53830 2066 53882
rect 2078 53830 2130 53882
rect 2142 53830 2194 53882
rect 2206 53830 2258 53882
rect 6950 53830 7002 53882
rect 7014 53830 7066 53882
rect 7078 53830 7130 53882
rect 7142 53830 7194 53882
rect 7206 53830 7258 53882
rect 11950 53830 12002 53882
rect 12014 53830 12066 53882
rect 12078 53830 12130 53882
rect 12142 53830 12194 53882
rect 12206 53830 12258 53882
rect 16950 53830 17002 53882
rect 17014 53830 17066 53882
rect 17078 53830 17130 53882
rect 17142 53830 17194 53882
rect 17206 53830 17258 53882
rect 1952 53388 2004 53440
rect 15936 53388 15988 53440
rect 2610 53286 2662 53338
rect 2674 53286 2726 53338
rect 2738 53286 2790 53338
rect 2802 53286 2854 53338
rect 2866 53286 2918 53338
rect 7610 53286 7662 53338
rect 7674 53286 7726 53338
rect 7738 53286 7790 53338
rect 7802 53286 7854 53338
rect 7866 53286 7918 53338
rect 12610 53286 12662 53338
rect 12674 53286 12726 53338
rect 12738 53286 12790 53338
rect 12802 53286 12854 53338
rect 12866 53286 12918 53338
rect 17610 53286 17662 53338
rect 17674 53286 17726 53338
rect 17738 53286 17790 53338
rect 17802 53286 17854 53338
rect 17866 53286 17918 53338
rect 7840 53184 7892 53236
rect 15292 53184 15344 53236
rect 1952 53159 2004 53168
rect 1952 53125 1961 53159
rect 1961 53125 1995 53159
rect 1995 53125 2004 53159
rect 1952 53116 2004 53125
rect 9128 53048 9180 53100
rect 10140 53116 10192 53168
rect 11428 53048 11480 53100
rect 3332 52980 3384 53032
rect 9864 53023 9916 53032
rect 9864 52989 9873 53023
rect 9873 52989 9907 53023
rect 9907 52989 9916 53023
rect 9864 52980 9916 52989
rect 756 52912 808 52964
rect 1768 52844 1820 52896
rect 8024 52844 8076 52896
rect 8576 52844 8628 52896
rect 9496 52887 9548 52896
rect 9496 52853 9505 52887
rect 9505 52853 9539 52887
rect 9539 52853 9548 52887
rect 9496 52844 9548 52853
rect 10416 52980 10468 53032
rect 14280 53116 14332 53168
rect 15844 53048 15896 53100
rect 10876 52844 10928 52896
rect 13268 52844 13320 52896
rect 1950 52742 2002 52794
rect 2014 52742 2066 52794
rect 2078 52742 2130 52794
rect 2142 52742 2194 52794
rect 2206 52742 2258 52794
rect 6950 52742 7002 52794
rect 7014 52742 7066 52794
rect 7078 52742 7130 52794
rect 7142 52742 7194 52794
rect 7206 52742 7258 52794
rect 11950 52742 12002 52794
rect 12014 52742 12066 52794
rect 12078 52742 12130 52794
rect 12142 52742 12194 52794
rect 12206 52742 12258 52794
rect 16950 52742 17002 52794
rect 17014 52742 17066 52794
rect 17078 52742 17130 52794
rect 17142 52742 17194 52794
rect 17206 52742 17258 52794
rect 6920 52640 6972 52692
rect 7840 52640 7892 52692
rect 18236 52615 18288 52624
rect 18236 52581 18245 52615
rect 18245 52581 18279 52615
rect 18279 52581 18288 52615
rect 18236 52572 18288 52581
rect 14280 52547 14332 52556
rect 14280 52513 14289 52547
rect 14289 52513 14323 52547
rect 14323 52513 14332 52547
rect 14280 52504 14332 52513
rect 8760 52436 8812 52488
rect 9312 52436 9364 52488
rect 15568 52436 15620 52488
rect 17960 52436 18012 52488
rect 15660 52343 15712 52352
rect 15660 52309 15669 52343
rect 15669 52309 15703 52343
rect 15703 52309 15712 52343
rect 15660 52300 15712 52309
rect 2610 52198 2662 52250
rect 2674 52198 2726 52250
rect 2738 52198 2790 52250
rect 2802 52198 2854 52250
rect 2866 52198 2918 52250
rect 7610 52198 7662 52250
rect 7674 52198 7726 52250
rect 7738 52198 7790 52250
rect 7802 52198 7854 52250
rect 7866 52198 7918 52250
rect 12610 52198 12662 52250
rect 12674 52198 12726 52250
rect 12738 52198 12790 52250
rect 12802 52198 12854 52250
rect 12866 52198 12918 52250
rect 17610 52198 17662 52250
rect 17674 52198 17726 52250
rect 17738 52198 17790 52250
rect 17802 52198 17854 52250
rect 17866 52198 17918 52250
rect 14556 52096 14608 52148
rect 18696 51960 18748 52012
rect 1950 51654 2002 51706
rect 2014 51654 2066 51706
rect 2078 51654 2130 51706
rect 2142 51654 2194 51706
rect 2206 51654 2258 51706
rect 6950 51654 7002 51706
rect 7014 51654 7066 51706
rect 7078 51654 7130 51706
rect 7142 51654 7194 51706
rect 7206 51654 7258 51706
rect 11950 51654 12002 51706
rect 12014 51654 12066 51706
rect 12078 51654 12130 51706
rect 12142 51654 12194 51706
rect 12206 51654 12258 51706
rect 16950 51654 17002 51706
rect 17014 51654 17066 51706
rect 17078 51654 17130 51706
rect 17142 51654 17194 51706
rect 17206 51654 17258 51706
rect 7840 51552 7892 51604
rect 2964 51416 3016 51468
rect 10416 51459 10468 51468
rect 10416 51425 10425 51459
rect 10425 51425 10459 51459
rect 10459 51425 10468 51459
rect 10416 51416 10468 51425
rect 13360 51416 13412 51468
rect 1400 51348 1452 51400
rect 14096 51348 14148 51400
rect 14280 51391 14332 51400
rect 14280 51357 14289 51391
rect 14289 51357 14323 51391
rect 14323 51357 14332 51391
rect 14280 51348 14332 51357
rect 4160 51212 4212 51264
rect 10600 51212 10652 51264
rect 11244 51212 11296 51264
rect 2610 51110 2662 51162
rect 2674 51110 2726 51162
rect 2738 51110 2790 51162
rect 2802 51110 2854 51162
rect 2866 51110 2918 51162
rect 7610 51110 7662 51162
rect 7674 51110 7726 51162
rect 7738 51110 7790 51162
rect 7802 51110 7854 51162
rect 7866 51110 7918 51162
rect 12610 51110 12662 51162
rect 12674 51110 12726 51162
rect 12738 51110 12790 51162
rect 12802 51110 12854 51162
rect 12866 51110 12918 51162
rect 17610 51110 17662 51162
rect 17674 51110 17726 51162
rect 17738 51110 17790 51162
rect 17802 51110 17854 51162
rect 17866 51110 17918 51162
rect 6092 50940 6144 50992
rect 8024 50940 8076 50992
rect 10692 50872 10744 50924
rect 13176 50872 13228 50924
rect 8024 50804 8076 50856
rect 8116 50736 8168 50788
rect 8760 50736 8812 50788
rect 2320 50668 2372 50720
rect 2596 50668 2648 50720
rect 9312 50668 9364 50720
rect 10692 50711 10744 50720
rect 10692 50677 10701 50711
rect 10701 50677 10735 50711
rect 10735 50677 10744 50711
rect 10692 50668 10744 50677
rect 18236 50711 18288 50720
rect 18236 50677 18245 50711
rect 18245 50677 18279 50711
rect 18279 50677 18288 50711
rect 18236 50668 18288 50677
rect 1950 50566 2002 50618
rect 2014 50566 2066 50618
rect 2078 50566 2130 50618
rect 2142 50566 2194 50618
rect 2206 50566 2258 50618
rect 6950 50566 7002 50618
rect 7014 50566 7066 50618
rect 7078 50566 7130 50618
rect 7142 50566 7194 50618
rect 7206 50566 7258 50618
rect 11950 50566 12002 50618
rect 12014 50566 12066 50618
rect 12078 50566 12130 50618
rect 12142 50566 12194 50618
rect 12206 50566 12258 50618
rect 16950 50566 17002 50618
rect 17014 50566 17066 50618
rect 17078 50566 17130 50618
rect 17142 50566 17194 50618
rect 17206 50566 17258 50618
rect 3148 50396 3200 50448
rect 4804 50328 4856 50380
rect 3332 50303 3384 50312
rect 3332 50269 3341 50303
rect 3341 50269 3375 50303
rect 3375 50269 3384 50303
rect 3332 50260 3384 50269
rect 5080 50260 5132 50312
rect 7564 50124 7616 50176
rect 14556 50124 14608 50176
rect 2610 50022 2662 50074
rect 2674 50022 2726 50074
rect 2738 50022 2790 50074
rect 2802 50022 2854 50074
rect 2866 50022 2918 50074
rect 7610 50022 7662 50074
rect 7674 50022 7726 50074
rect 7738 50022 7790 50074
rect 7802 50022 7854 50074
rect 7866 50022 7918 50074
rect 12610 50022 12662 50074
rect 12674 50022 12726 50074
rect 12738 50022 12790 50074
rect 12802 50022 12854 50074
rect 12866 50022 12918 50074
rect 17610 50022 17662 50074
rect 17674 50022 17726 50074
rect 17738 50022 17790 50074
rect 17802 50022 17854 50074
rect 17866 50022 17918 50074
rect 1860 49920 1912 49972
rect 3700 49920 3752 49972
rect 4436 49963 4488 49972
rect 4436 49929 4445 49963
rect 4445 49929 4479 49963
rect 4479 49929 4488 49963
rect 4436 49920 4488 49929
rect 4160 49852 4212 49904
rect 8300 49895 8352 49904
rect 8300 49861 8334 49895
rect 8334 49861 8352 49895
rect 8300 49852 8352 49861
rect 2964 49716 3016 49768
rect 8024 49759 8076 49768
rect 8024 49725 8033 49759
rect 8033 49725 8067 49759
rect 8067 49725 8076 49759
rect 8024 49716 8076 49725
rect 9588 49716 9640 49768
rect 16856 49716 16908 49768
rect 3424 49580 3476 49632
rect 1950 49478 2002 49530
rect 2014 49478 2066 49530
rect 2078 49478 2130 49530
rect 2142 49478 2194 49530
rect 2206 49478 2258 49530
rect 6950 49478 7002 49530
rect 7014 49478 7066 49530
rect 7078 49478 7130 49530
rect 7142 49478 7194 49530
rect 7206 49478 7258 49530
rect 11950 49478 12002 49530
rect 12014 49478 12066 49530
rect 12078 49478 12130 49530
rect 12142 49478 12194 49530
rect 12206 49478 12258 49530
rect 16950 49478 17002 49530
rect 17014 49478 17066 49530
rect 17078 49478 17130 49530
rect 17142 49478 17194 49530
rect 17206 49478 17258 49530
rect 14004 49308 14056 49360
rect 3424 49172 3476 49224
rect 8024 49172 8076 49224
rect 16396 49104 16448 49156
rect 8024 49036 8076 49088
rect 8576 49036 8628 49088
rect 2610 48934 2662 48986
rect 2674 48934 2726 48986
rect 2738 48934 2790 48986
rect 2802 48934 2854 48986
rect 2866 48934 2918 48986
rect 7610 48934 7662 48986
rect 7674 48934 7726 48986
rect 7738 48934 7790 48986
rect 7802 48934 7854 48986
rect 7866 48934 7918 48986
rect 12610 48934 12662 48986
rect 12674 48934 12726 48986
rect 12738 48934 12790 48986
rect 12802 48934 12854 48986
rect 12866 48934 12918 48986
rect 17610 48934 17662 48986
rect 17674 48934 17726 48986
rect 17738 48934 17790 48986
rect 17802 48934 17854 48986
rect 17866 48934 17918 48986
rect 7472 48875 7524 48884
rect 7472 48841 7481 48875
rect 7481 48841 7515 48875
rect 7515 48841 7524 48875
rect 7472 48832 7524 48841
rect 14096 48832 14148 48884
rect 10232 48764 10284 48816
rect 10784 48764 10836 48816
rect 3700 48739 3752 48748
rect 3700 48705 3734 48739
rect 3734 48705 3752 48739
rect 3700 48696 3752 48705
rect 8576 48696 8628 48748
rect 3424 48671 3476 48680
rect 3424 48637 3433 48671
rect 3433 48637 3467 48671
rect 3467 48637 3476 48671
rect 3424 48628 3476 48637
rect 6276 48560 6328 48612
rect 14648 48739 14700 48748
rect 14648 48705 14657 48739
rect 14657 48705 14691 48739
rect 14691 48705 14700 48739
rect 14648 48696 14700 48705
rect 16028 48739 16080 48748
rect 16028 48705 16037 48739
rect 16037 48705 16071 48739
rect 16071 48705 16080 48739
rect 16028 48696 16080 48705
rect 10692 48628 10744 48680
rect 10048 48560 10100 48612
rect 10232 48560 10284 48612
rect 11060 48628 11112 48680
rect 14740 48671 14792 48680
rect 14740 48637 14749 48671
rect 14749 48637 14783 48671
rect 14783 48637 14792 48671
rect 14740 48628 14792 48637
rect 15016 48628 15068 48680
rect 15384 48628 15436 48680
rect 16672 48560 16724 48612
rect 6644 48492 6696 48544
rect 10692 48492 10744 48544
rect 15660 48492 15712 48544
rect 18236 48535 18288 48544
rect 18236 48501 18245 48535
rect 18245 48501 18279 48535
rect 18279 48501 18288 48535
rect 18236 48492 18288 48501
rect 1950 48390 2002 48442
rect 2014 48390 2066 48442
rect 2078 48390 2130 48442
rect 2142 48390 2194 48442
rect 2206 48390 2258 48442
rect 6950 48390 7002 48442
rect 7014 48390 7066 48442
rect 7078 48390 7130 48442
rect 7142 48390 7194 48442
rect 7206 48390 7258 48442
rect 11950 48390 12002 48442
rect 12014 48390 12066 48442
rect 12078 48390 12130 48442
rect 12142 48390 12194 48442
rect 12206 48390 12258 48442
rect 16950 48390 17002 48442
rect 17014 48390 17066 48442
rect 17078 48390 17130 48442
rect 17142 48390 17194 48442
rect 17206 48390 17258 48442
rect 1584 48288 1636 48340
rect 6644 48288 6696 48340
rect 10048 48288 10100 48340
rect 10692 48288 10744 48340
rect 2610 47846 2662 47898
rect 2674 47846 2726 47898
rect 2738 47846 2790 47898
rect 2802 47846 2854 47898
rect 2866 47846 2918 47898
rect 7610 47846 7662 47898
rect 7674 47846 7726 47898
rect 7738 47846 7790 47898
rect 7802 47846 7854 47898
rect 7866 47846 7918 47898
rect 12610 47846 12662 47898
rect 12674 47846 12726 47898
rect 12738 47846 12790 47898
rect 12802 47846 12854 47898
rect 12866 47846 12918 47898
rect 17610 47846 17662 47898
rect 17674 47846 17726 47898
rect 17738 47846 17790 47898
rect 17802 47846 17854 47898
rect 17866 47846 17918 47898
rect 6184 47744 6236 47796
rect 6460 47744 6512 47796
rect 7656 47744 7708 47796
rect 8392 47744 8444 47796
rect 8852 47676 8904 47728
rect 2964 47608 3016 47660
rect 3056 47651 3108 47660
rect 3056 47617 3065 47651
rect 3065 47617 3099 47651
rect 3099 47617 3108 47651
rect 3056 47608 3108 47617
rect 3976 47472 4028 47524
rect 7380 47608 7432 47660
rect 7472 47608 7524 47660
rect 7748 47608 7800 47660
rect 10508 47608 10560 47660
rect 11520 47540 11572 47592
rect 12440 47540 12492 47592
rect 7564 47472 7616 47524
rect 4804 47447 4856 47456
rect 4804 47413 4813 47447
rect 4813 47413 4847 47447
rect 4847 47413 4856 47447
rect 4804 47404 4856 47413
rect 13084 47404 13136 47456
rect 19248 47404 19300 47456
rect 1950 47302 2002 47354
rect 2014 47302 2066 47354
rect 2078 47302 2130 47354
rect 2142 47302 2194 47354
rect 2206 47302 2258 47354
rect 6950 47302 7002 47354
rect 7014 47302 7066 47354
rect 7078 47302 7130 47354
rect 7142 47302 7194 47354
rect 7206 47302 7258 47354
rect 11950 47302 12002 47354
rect 12014 47302 12066 47354
rect 12078 47302 12130 47354
rect 12142 47302 12194 47354
rect 12206 47302 12258 47354
rect 16950 47302 17002 47354
rect 17014 47302 17066 47354
rect 17078 47302 17130 47354
rect 17142 47302 17194 47354
rect 17206 47302 17258 47354
rect 3056 47132 3108 47184
rect 11428 47132 11480 47184
rect 2964 47064 3016 47116
rect 15108 47064 15160 47116
rect 3240 46971 3292 46980
rect 3240 46937 3249 46971
rect 3249 46937 3283 46971
rect 3283 46937 3292 46971
rect 3240 46928 3292 46937
rect 3792 46928 3844 46980
rect 7748 46996 7800 47048
rect 15844 46996 15896 47048
rect 16488 46996 16540 47048
rect 7656 46928 7708 46980
rect 18236 46903 18288 46912
rect 18236 46869 18245 46903
rect 18245 46869 18279 46903
rect 18279 46869 18288 46903
rect 18236 46860 18288 46869
rect 2610 46758 2662 46810
rect 2674 46758 2726 46810
rect 2738 46758 2790 46810
rect 2802 46758 2854 46810
rect 2866 46758 2918 46810
rect 7610 46758 7662 46810
rect 7674 46758 7726 46810
rect 7738 46758 7790 46810
rect 7802 46758 7854 46810
rect 7866 46758 7918 46810
rect 12610 46758 12662 46810
rect 12674 46758 12726 46810
rect 12738 46758 12790 46810
rect 12802 46758 12854 46810
rect 12866 46758 12918 46810
rect 17610 46758 17662 46810
rect 17674 46758 17726 46810
rect 17738 46758 17790 46810
rect 17802 46758 17854 46810
rect 17866 46758 17918 46810
rect 3976 46656 4028 46708
rect 12532 46631 12584 46640
rect 12532 46597 12566 46631
rect 12566 46597 12584 46631
rect 12532 46588 12584 46597
rect 16856 46520 16908 46572
rect 6460 46316 6512 46368
rect 8024 46316 8076 46368
rect 12440 46316 12492 46368
rect 13636 46359 13688 46368
rect 13636 46325 13645 46359
rect 13645 46325 13679 46359
rect 13679 46325 13688 46359
rect 13636 46316 13688 46325
rect 1950 46214 2002 46266
rect 2014 46214 2066 46266
rect 2078 46214 2130 46266
rect 2142 46214 2194 46266
rect 2206 46214 2258 46266
rect 6950 46214 7002 46266
rect 7014 46214 7066 46266
rect 7078 46214 7130 46266
rect 7142 46214 7194 46266
rect 7206 46214 7258 46266
rect 11950 46214 12002 46266
rect 12014 46214 12066 46266
rect 12078 46214 12130 46266
rect 12142 46214 12194 46266
rect 12206 46214 12258 46266
rect 16950 46214 17002 46266
rect 17014 46214 17066 46266
rect 17078 46214 17130 46266
rect 17142 46214 17194 46266
rect 17206 46214 17258 46266
rect 7288 46112 7340 46164
rect 8024 46112 8076 46164
rect 2610 45670 2662 45722
rect 2674 45670 2726 45722
rect 2738 45670 2790 45722
rect 2802 45670 2854 45722
rect 2866 45670 2918 45722
rect 7610 45670 7662 45722
rect 7674 45670 7726 45722
rect 7738 45670 7790 45722
rect 7802 45670 7854 45722
rect 7866 45670 7918 45722
rect 12610 45670 12662 45722
rect 12674 45670 12726 45722
rect 12738 45670 12790 45722
rect 12802 45670 12854 45722
rect 12866 45670 12918 45722
rect 17610 45670 17662 45722
rect 17674 45670 17726 45722
rect 17738 45670 17790 45722
rect 17802 45670 17854 45722
rect 17866 45670 17918 45722
rect 7288 45568 7340 45620
rect 12440 45568 12492 45620
rect 1950 45126 2002 45178
rect 2014 45126 2066 45178
rect 2078 45126 2130 45178
rect 2142 45126 2194 45178
rect 2206 45126 2258 45178
rect 6950 45126 7002 45178
rect 7014 45126 7066 45178
rect 7078 45126 7130 45178
rect 7142 45126 7194 45178
rect 7206 45126 7258 45178
rect 11950 45126 12002 45178
rect 12014 45126 12066 45178
rect 12078 45126 12130 45178
rect 12142 45126 12194 45178
rect 12206 45126 12258 45178
rect 16950 45126 17002 45178
rect 17014 45126 17066 45178
rect 17078 45126 17130 45178
rect 17142 45126 17194 45178
rect 17206 45126 17258 45178
rect 13544 45024 13596 45076
rect 13820 45024 13872 45076
rect 16396 45067 16448 45076
rect 16396 45033 16405 45067
rect 16405 45033 16439 45067
rect 16439 45033 16448 45067
rect 16396 45024 16448 45033
rect 12440 44888 12492 44940
rect 14556 44931 14608 44940
rect 14556 44897 14565 44931
rect 14565 44897 14599 44931
rect 14599 44897 14608 44931
rect 14556 44888 14608 44897
rect 11704 44820 11756 44872
rect 2504 44752 2556 44804
rect 4436 44752 4488 44804
rect 11520 44752 11572 44804
rect 13452 44795 13504 44804
rect 13452 44761 13461 44795
rect 13461 44761 13495 44795
rect 13495 44761 13504 44795
rect 13452 44752 13504 44761
rect 13728 44820 13780 44872
rect 19524 44820 19576 44872
rect 14004 44752 14056 44804
rect 2136 44684 2188 44736
rect 3884 44684 3936 44736
rect 6092 44684 6144 44736
rect 15292 44684 15344 44736
rect 16764 44684 16816 44736
rect 18236 44727 18288 44736
rect 18236 44693 18245 44727
rect 18245 44693 18279 44727
rect 18279 44693 18288 44727
rect 18236 44684 18288 44693
rect 2610 44582 2662 44634
rect 2674 44582 2726 44634
rect 2738 44582 2790 44634
rect 2802 44582 2854 44634
rect 2866 44582 2918 44634
rect 7610 44582 7662 44634
rect 7674 44582 7726 44634
rect 7738 44582 7790 44634
rect 7802 44582 7854 44634
rect 7866 44582 7918 44634
rect 12610 44582 12662 44634
rect 12674 44582 12726 44634
rect 12738 44582 12790 44634
rect 12802 44582 12854 44634
rect 12866 44582 12918 44634
rect 17610 44582 17662 44634
rect 17674 44582 17726 44634
rect 17738 44582 17790 44634
rect 17802 44582 17854 44634
rect 17866 44582 17918 44634
rect 14372 44480 14424 44532
rect 2136 44455 2188 44464
rect 2136 44421 2145 44455
rect 2145 44421 2179 44455
rect 2179 44421 2188 44455
rect 2136 44412 2188 44421
rect 3332 44412 3384 44464
rect 7288 44412 7340 44464
rect 2320 44276 2372 44328
rect 3424 44276 3476 44328
rect 4436 44344 4488 44396
rect 18328 44344 18380 44396
rect 2228 44208 2280 44260
rect 2504 44208 2556 44260
rect 5724 44183 5776 44192
rect 5724 44149 5733 44183
rect 5733 44149 5767 44183
rect 5767 44149 5776 44183
rect 5724 44140 5776 44149
rect 8392 44140 8444 44192
rect 10600 44140 10652 44192
rect 18144 44140 18196 44192
rect 1950 44038 2002 44090
rect 2014 44038 2066 44090
rect 2078 44038 2130 44090
rect 2142 44038 2194 44090
rect 2206 44038 2258 44090
rect 6950 44038 7002 44090
rect 7014 44038 7066 44090
rect 7078 44038 7130 44090
rect 7142 44038 7194 44090
rect 7206 44038 7258 44090
rect 11950 44038 12002 44090
rect 12014 44038 12066 44090
rect 12078 44038 12130 44090
rect 12142 44038 12194 44090
rect 12206 44038 12258 44090
rect 16950 44038 17002 44090
rect 17014 44038 17066 44090
rect 17078 44038 17130 44090
rect 17142 44038 17194 44090
rect 17206 44038 17258 44090
rect 19432 44072 19484 44124
rect 3332 43800 3384 43852
rect 9772 43800 9824 43852
rect 8760 43732 8812 43784
rect 14832 43732 14884 43784
rect 19432 43664 19484 43716
rect 6736 43639 6788 43648
rect 6736 43605 6745 43639
rect 6745 43605 6779 43639
rect 6779 43605 6788 43639
rect 6736 43596 6788 43605
rect 2610 43494 2662 43546
rect 2674 43494 2726 43546
rect 2738 43494 2790 43546
rect 2802 43494 2854 43546
rect 2866 43494 2918 43546
rect 7610 43494 7662 43546
rect 7674 43494 7726 43546
rect 7738 43494 7790 43546
rect 7802 43494 7854 43546
rect 7866 43494 7918 43546
rect 12610 43494 12662 43546
rect 12674 43494 12726 43546
rect 12738 43494 12790 43546
rect 12802 43494 12854 43546
rect 12866 43494 12918 43546
rect 17610 43494 17662 43546
rect 17674 43494 17726 43546
rect 17738 43494 17790 43546
rect 17802 43494 17854 43546
rect 17866 43494 17918 43546
rect 13728 43392 13780 43444
rect 18512 43392 18564 43444
rect 18512 43256 18564 43308
rect 8944 43188 8996 43240
rect 12532 43188 12584 43240
rect 18236 43095 18288 43104
rect 18236 43061 18245 43095
rect 18245 43061 18279 43095
rect 18279 43061 18288 43095
rect 18236 43052 18288 43061
rect 1950 42950 2002 43002
rect 2014 42950 2066 43002
rect 2078 42950 2130 43002
rect 2142 42950 2194 43002
rect 2206 42950 2258 43002
rect 6950 42950 7002 43002
rect 7014 42950 7066 43002
rect 7078 42950 7130 43002
rect 7142 42950 7194 43002
rect 7206 42950 7258 43002
rect 11950 42950 12002 43002
rect 12014 42950 12066 43002
rect 12078 42950 12130 43002
rect 12142 42950 12194 43002
rect 12206 42950 12258 43002
rect 16950 42950 17002 43002
rect 17014 42950 17066 43002
rect 17078 42950 17130 43002
rect 17142 42950 17194 43002
rect 17206 42950 17258 43002
rect 6460 42780 6512 42832
rect 6736 42780 6788 42832
rect 10968 42780 11020 42832
rect 1676 42712 1728 42764
rect 1952 42712 2004 42764
rect 1492 42644 1544 42696
rect 5448 42644 5500 42696
rect 3608 42576 3660 42628
rect 1676 42551 1728 42560
rect 1676 42517 1709 42551
rect 1709 42517 1728 42551
rect 1676 42508 1728 42517
rect 3332 42508 3384 42560
rect 7472 42712 7524 42764
rect 6460 42644 6512 42696
rect 13360 42780 13412 42832
rect 13912 42780 13964 42832
rect 13820 42712 13872 42764
rect 9312 42508 9364 42560
rect 10416 42576 10468 42628
rect 11704 42576 11756 42628
rect 9680 42508 9732 42560
rect 10508 42551 10560 42560
rect 10508 42517 10517 42551
rect 10517 42517 10551 42551
rect 10551 42517 10560 42551
rect 10508 42508 10560 42517
rect 10692 42508 10744 42560
rect 15200 42644 15252 42696
rect 13728 42576 13780 42628
rect 13176 42508 13228 42560
rect 16764 42508 16816 42560
rect 17316 42508 17368 42560
rect 17408 42508 17460 42560
rect 17592 42508 17644 42560
rect 2610 42406 2662 42458
rect 2674 42406 2726 42458
rect 2738 42406 2790 42458
rect 2802 42406 2854 42458
rect 2866 42406 2918 42458
rect 7610 42406 7662 42458
rect 7674 42406 7726 42458
rect 7738 42406 7790 42458
rect 7802 42406 7854 42458
rect 7866 42406 7918 42458
rect 12610 42406 12662 42458
rect 12674 42406 12726 42458
rect 12738 42406 12790 42458
rect 12802 42406 12854 42458
rect 12866 42406 12918 42458
rect 17610 42406 17662 42458
rect 17674 42406 17726 42458
rect 17738 42406 17790 42458
rect 17802 42406 17854 42458
rect 17866 42406 17918 42458
rect 1952 42236 2004 42288
rect 8116 42236 8168 42288
rect 2228 42168 2280 42220
rect 7288 42211 7340 42220
rect 7288 42177 7297 42211
rect 7297 42177 7331 42211
rect 7331 42177 7340 42211
rect 7288 42168 7340 42177
rect 8668 42347 8720 42356
rect 8668 42313 8677 42347
rect 8677 42313 8711 42347
rect 8711 42313 8720 42347
rect 8668 42304 8720 42313
rect 9128 42347 9180 42356
rect 9128 42313 9137 42347
rect 9137 42313 9171 42347
rect 9171 42313 9180 42347
rect 9128 42304 9180 42313
rect 8300 42236 8352 42288
rect 13176 42304 13228 42356
rect 9312 42236 9364 42288
rect 10508 42236 10560 42288
rect 17316 42236 17368 42288
rect 9772 42143 9824 42152
rect 9772 42109 9781 42143
rect 9781 42109 9815 42143
rect 9815 42109 9824 42143
rect 9772 42100 9824 42109
rect 13820 42100 13872 42152
rect 9496 42032 9548 42084
rect 18604 42100 18656 42152
rect 11612 41964 11664 42016
rect 1950 41862 2002 41914
rect 2014 41862 2066 41914
rect 2078 41862 2130 41914
rect 2142 41862 2194 41914
rect 2206 41862 2258 41914
rect 6950 41862 7002 41914
rect 7014 41862 7066 41914
rect 7078 41862 7130 41914
rect 7142 41862 7194 41914
rect 7206 41862 7258 41914
rect 11950 41862 12002 41914
rect 12014 41862 12066 41914
rect 12078 41862 12130 41914
rect 12142 41862 12194 41914
rect 12206 41862 12258 41914
rect 16950 41862 17002 41914
rect 17014 41862 17066 41914
rect 17078 41862 17130 41914
rect 17142 41862 17194 41914
rect 17206 41862 17258 41914
rect 7196 41760 7248 41812
rect 7380 41760 7432 41812
rect 8116 41760 8168 41812
rect 8392 41760 8444 41812
rect 6276 41624 6328 41676
rect 10968 41624 11020 41676
rect 664 41556 716 41608
rect 6460 41556 6512 41608
rect 6736 41556 6788 41608
rect 7472 41556 7524 41608
rect 9312 41556 9364 41608
rect 15200 41488 15252 41540
rect 6092 41463 6144 41472
rect 6092 41429 6101 41463
rect 6101 41429 6135 41463
rect 6135 41429 6144 41463
rect 6092 41420 6144 41429
rect 6184 41463 6236 41472
rect 6184 41429 6193 41463
rect 6193 41429 6227 41463
rect 6227 41429 6236 41463
rect 6184 41420 6236 41429
rect 2610 41318 2662 41370
rect 2674 41318 2726 41370
rect 2738 41318 2790 41370
rect 2802 41318 2854 41370
rect 2866 41318 2918 41370
rect 7610 41318 7662 41370
rect 7674 41318 7726 41370
rect 7738 41318 7790 41370
rect 7802 41318 7854 41370
rect 7866 41318 7918 41370
rect 12610 41318 12662 41370
rect 12674 41318 12726 41370
rect 12738 41318 12790 41370
rect 12802 41318 12854 41370
rect 12866 41318 12918 41370
rect 17610 41318 17662 41370
rect 17674 41318 17726 41370
rect 17738 41318 17790 41370
rect 17802 41318 17854 41370
rect 17866 41318 17918 41370
rect 19800 41080 19852 41132
rect 7196 40876 7248 40928
rect 7656 40876 7708 40928
rect 18236 40919 18288 40928
rect 18236 40885 18245 40919
rect 18245 40885 18279 40919
rect 18279 40885 18288 40919
rect 18236 40876 18288 40885
rect 1950 40774 2002 40826
rect 2014 40774 2066 40826
rect 2078 40774 2130 40826
rect 2142 40774 2194 40826
rect 2206 40774 2258 40826
rect 6950 40774 7002 40826
rect 7014 40774 7066 40826
rect 7078 40774 7130 40826
rect 7142 40774 7194 40826
rect 7206 40774 7258 40826
rect 11950 40774 12002 40826
rect 12014 40774 12066 40826
rect 12078 40774 12130 40826
rect 12142 40774 12194 40826
rect 12206 40774 12258 40826
rect 16950 40774 17002 40826
rect 17014 40774 17066 40826
rect 17078 40774 17130 40826
rect 17142 40774 17194 40826
rect 17206 40774 17258 40826
rect 8668 40468 8720 40520
rect 8944 40468 8996 40520
rect 6644 40332 6696 40384
rect 7656 40332 7708 40384
rect 10968 40332 11020 40384
rect 2610 40230 2662 40282
rect 2674 40230 2726 40282
rect 2738 40230 2790 40282
rect 2802 40230 2854 40282
rect 2866 40230 2918 40282
rect 7610 40230 7662 40282
rect 7674 40230 7726 40282
rect 7738 40230 7790 40282
rect 7802 40230 7854 40282
rect 7866 40230 7918 40282
rect 12610 40230 12662 40282
rect 12674 40230 12726 40282
rect 12738 40230 12790 40282
rect 12802 40230 12854 40282
rect 12866 40230 12918 40282
rect 17610 40230 17662 40282
rect 17674 40230 17726 40282
rect 17738 40230 17790 40282
rect 17802 40230 17854 40282
rect 17866 40230 17918 40282
rect 5080 40128 5132 40180
rect 8484 40128 8536 40180
rect 9312 40128 9364 40180
rect 10968 40171 11020 40180
rect 10968 40137 10977 40171
rect 10977 40137 11011 40171
rect 11011 40137 11020 40171
rect 10968 40128 11020 40137
rect 8852 40060 8904 40112
rect 6828 39992 6880 40044
rect 11336 39992 11388 40044
rect 8392 39924 8444 39976
rect 8484 39967 8536 39976
rect 8484 39933 8493 39967
rect 8493 39933 8527 39967
rect 8527 39933 8536 39967
rect 8484 39924 8536 39933
rect 8760 39924 8812 39976
rect 16764 39924 16816 39976
rect 7288 39856 7340 39908
rect 8484 39788 8536 39840
rect 8668 39788 8720 39840
rect 15016 39788 15068 39840
rect 16764 39788 16816 39840
rect 16948 39788 17000 39840
rect 1950 39686 2002 39738
rect 2014 39686 2066 39738
rect 2078 39686 2130 39738
rect 2142 39686 2194 39738
rect 2206 39686 2258 39738
rect 6950 39686 7002 39738
rect 7014 39686 7066 39738
rect 7078 39686 7130 39738
rect 7142 39686 7194 39738
rect 7206 39686 7258 39738
rect 11950 39686 12002 39738
rect 12014 39686 12066 39738
rect 12078 39686 12130 39738
rect 12142 39686 12194 39738
rect 12206 39686 12258 39738
rect 16950 39686 17002 39738
rect 17014 39686 17066 39738
rect 17078 39686 17130 39738
rect 17142 39686 17194 39738
rect 17206 39686 17258 39738
rect 2504 39584 2556 39636
rect 8392 39584 8444 39636
rect 11796 39584 11848 39636
rect 14188 39584 14240 39636
rect 8944 39516 8996 39568
rect 12532 39448 12584 39500
rect 13452 39448 13504 39500
rect 8484 39380 8536 39432
rect 9128 39312 9180 39364
rect 10508 39312 10560 39364
rect 12348 39287 12400 39296
rect 12348 39253 12357 39287
rect 12357 39253 12391 39287
rect 12391 39253 12400 39287
rect 12348 39244 12400 39253
rect 18236 39287 18288 39296
rect 18236 39253 18245 39287
rect 18245 39253 18279 39287
rect 18279 39253 18288 39287
rect 18236 39244 18288 39253
rect 2610 39142 2662 39194
rect 2674 39142 2726 39194
rect 2738 39142 2790 39194
rect 2802 39142 2854 39194
rect 2866 39142 2918 39194
rect 7610 39142 7662 39194
rect 7674 39142 7726 39194
rect 7738 39142 7790 39194
rect 7802 39142 7854 39194
rect 7866 39142 7918 39194
rect 12610 39142 12662 39194
rect 12674 39142 12726 39194
rect 12738 39142 12790 39194
rect 12802 39142 12854 39194
rect 12866 39142 12918 39194
rect 17610 39142 17662 39194
rect 17674 39142 17726 39194
rect 17738 39142 17790 39194
rect 17802 39142 17854 39194
rect 17866 39142 17918 39194
rect 4896 38972 4948 39024
rect 2320 38904 2372 38956
rect 17316 38904 17368 38956
rect 2964 38700 3016 38752
rect 7288 38768 7340 38820
rect 15016 38768 15068 38820
rect 19616 38836 19668 38888
rect 6828 38700 6880 38752
rect 14004 38700 14056 38752
rect 14464 38700 14516 38752
rect 17316 38700 17368 38752
rect 1950 38598 2002 38650
rect 2014 38598 2066 38650
rect 2078 38598 2130 38650
rect 2142 38598 2194 38650
rect 2206 38598 2258 38650
rect 6950 38598 7002 38650
rect 7014 38598 7066 38650
rect 7078 38598 7130 38650
rect 7142 38598 7194 38650
rect 7206 38598 7258 38650
rect 11950 38598 12002 38650
rect 12014 38598 12066 38650
rect 12078 38598 12130 38650
rect 12142 38598 12194 38650
rect 12206 38598 12258 38650
rect 16950 38598 17002 38650
rect 17014 38598 17066 38650
rect 17078 38598 17130 38650
rect 17142 38598 17194 38650
rect 17206 38598 17258 38650
rect 6644 38496 6696 38548
rect 7288 38496 7340 38548
rect 15200 38292 15252 38344
rect 13544 38224 13596 38276
rect 19892 38224 19944 38276
rect 11336 38156 11388 38208
rect 2610 38054 2662 38106
rect 2674 38054 2726 38106
rect 2738 38054 2790 38106
rect 2802 38054 2854 38106
rect 2866 38054 2918 38106
rect 7610 38054 7662 38106
rect 7674 38054 7726 38106
rect 7738 38054 7790 38106
rect 7802 38054 7854 38106
rect 7866 38054 7918 38106
rect 12610 38054 12662 38106
rect 12674 38054 12726 38106
rect 12738 38054 12790 38106
rect 12802 38054 12854 38106
rect 12866 38054 12918 38106
rect 17610 38054 17662 38106
rect 17674 38054 17726 38106
rect 17738 38054 17790 38106
rect 17802 38054 17854 38106
rect 17866 38054 17918 38106
rect 15936 37995 15988 38004
rect 15936 37961 15945 37995
rect 15945 37961 15979 37995
rect 15979 37961 15988 37995
rect 15936 37952 15988 37961
rect 18328 37952 18380 38004
rect 5540 37884 5592 37936
rect 15384 37884 15436 37936
rect 16488 37816 16540 37868
rect 13544 37748 13596 37800
rect 15200 37612 15252 37664
rect 1950 37510 2002 37562
rect 2014 37510 2066 37562
rect 2078 37510 2130 37562
rect 2142 37510 2194 37562
rect 2206 37510 2258 37562
rect 6950 37510 7002 37562
rect 7014 37510 7066 37562
rect 7078 37510 7130 37562
rect 7142 37510 7194 37562
rect 7206 37510 7258 37562
rect 11950 37510 12002 37562
rect 12014 37510 12066 37562
rect 12078 37510 12130 37562
rect 12142 37510 12194 37562
rect 12206 37510 12258 37562
rect 16950 37510 17002 37562
rect 17014 37510 17066 37562
rect 17078 37510 17130 37562
rect 17142 37510 17194 37562
rect 17206 37510 17258 37562
rect 9588 37408 9640 37460
rect 9772 37408 9824 37460
rect 12624 37451 12676 37460
rect 12624 37417 12633 37451
rect 12633 37417 12667 37451
rect 12667 37417 12676 37451
rect 12624 37408 12676 37417
rect 12440 37340 12492 37392
rect 15016 37340 15068 37392
rect 13544 37272 13596 37324
rect 14832 37272 14884 37324
rect 15752 37272 15804 37324
rect 2964 37204 3016 37256
rect 13084 37204 13136 37256
rect 18052 37247 18104 37256
rect 18052 37213 18061 37247
rect 18061 37213 18095 37247
rect 18095 37213 18104 37247
rect 18052 37204 18104 37213
rect 1860 37136 1912 37188
rect 12624 37136 12676 37188
rect 13452 37136 13504 37188
rect 8392 37068 8444 37120
rect 9036 37068 9088 37120
rect 13176 37068 13228 37120
rect 18236 37111 18288 37120
rect 18236 37077 18245 37111
rect 18245 37077 18279 37111
rect 18279 37077 18288 37111
rect 18236 37068 18288 37077
rect 2610 36966 2662 37018
rect 2674 36966 2726 37018
rect 2738 36966 2790 37018
rect 2802 36966 2854 37018
rect 2866 36966 2918 37018
rect 7610 36966 7662 37018
rect 7674 36966 7726 37018
rect 7738 36966 7790 37018
rect 7802 36966 7854 37018
rect 7866 36966 7918 37018
rect 12610 36966 12662 37018
rect 12674 36966 12726 37018
rect 12738 36966 12790 37018
rect 12802 36966 12854 37018
rect 12866 36966 12918 37018
rect 17610 36966 17662 37018
rect 17674 36966 17726 37018
rect 17738 36966 17790 37018
rect 17802 36966 17854 37018
rect 17866 36966 17918 37018
rect 4068 36864 4120 36916
rect 8392 36864 8444 36916
rect 10692 36864 10744 36916
rect 11612 36864 11664 36916
rect 9128 36728 9180 36780
rect 12992 36864 13044 36916
rect 13360 36864 13412 36916
rect 17500 36864 17552 36916
rect 15936 36728 15988 36780
rect 8668 36703 8720 36712
rect 8668 36669 8677 36703
rect 8677 36669 8711 36703
rect 8711 36669 8720 36703
rect 8668 36660 8720 36669
rect 9772 36660 9824 36712
rect 10416 36660 10468 36712
rect 13268 36660 13320 36712
rect 17408 36660 17460 36712
rect 6644 36592 6696 36644
rect 14004 36592 14056 36644
rect 15108 36524 15160 36576
rect 15660 36524 15712 36576
rect 18328 36524 18380 36576
rect 19432 36524 19484 36576
rect 1950 36422 2002 36474
rect 2014 36422 2066 36474
rect 2078 36422 2130 36474
rect 2142 36422 2194 36474
rect 2206 36422 2258 36474
rect 6950 36422 7002 36474
rect 7014 36422 7066 36474
rect 7078 36422 7130 36474
rect 7142 36422 7194 36474
rect 7206 36422 7258 36474
rect 11950 36422 12002 36474
rect 12014 36422 12066 36474
rect 12078 36422 12130 36474
rect 12142 36422 12194 36474
rect 12206 36422 12258 36474
rect 16950 36422 17002 36474
rect 17014 36422 17066 36474
rect 17078 36422 17130 36474
rect 17142 36422 17194 36474
rect 17206 36422 17258 36474
rect 6644 36320 6696 36372
rect 10232 36320 10284 36372
rect 10600 36320 10652 36372
rect 4528 36252 4580 36304
rect 9772 36184 9824 36236
rect 9864 36116 9916 36168
rect 9312 36048 9364 36100
rect 18052 36048 18104 36100
rect 10048 35980 10100 36032
rect 11520 35980 11572 36032
rect 2610 35878 2662 35930
rect 2674 35878 2726 35930
rect 2738 35878 2790 35930
rect 2802 35878 2854 35930
rect 2866 35878 2918 35930
rect 7610 35878 7662 35930
rect 7674 35878 7726 35930
rect 7738 35878 7790 35930
rect 7802 35878 7854 35930
rect 7866 35878 7918 35930
rect 12610 35878 12662 35930
rect 12674 35878 12726 35930
rect 12738 35878 12790 35930
rect 12802 35878 12854 35930
rect 12866 35878 12918 35930
rect 17610 35878 17662 35930
rect 17674 35878 17726 35930
rect 17738 35878 17790 35930
rect 17802 35878 17854 35930
rect 17866 35878 17918 35930
rect 3700 35776 3752 35828
rect 4988 35776 5040 35828
rect 6828 35776 6880 35828
rect 9772 35776 9824 35828
rect 11888 35776 11940 35828
rect 11428 35708 11480 35760
rect 8024 35640 8076 35692
rect 11428 35572 11480 35624
rect 11796 35572 11848 35624
rect 11888 35572 11940 35624
rect 5724 35504 5776 35556
rect 12992 35504 13044 35556
rect 12440 35479 12492 35488
rect 12440 35445 12449 35479
rect 12449 35445 12483 35479
rect 12483 35445 12492 35479
rect 12440 35436 12492 35445
rect 14096 35504 14148 35556
rect 19708 35504 19760 35556
rect 13820 35436 13872 35488
rect 18236 35479 18288 35488
rect 18236 35445 18245 35479
rect 18245 35445 18279 35479
rect 18279 35445 18288 35479
rect 18236 35436 18288 35445
rect 1950 35334 2002 35386
rect 2014 35334 2066 35386
rect 2078 35334 2130 35386
rect 2142 35334 2194 35386
rect 2206 35334 2258 35386
rect 6950 35334 7002 35386
rect 7014 35334 7066 35386
rect 7078 35334 7130 35386
rect 7142 35334 7194 35386
rect 7206 35334 7258 35386
rect 11950 35334 12002 35386
rect 12014 35334 12066 35386
rect 12078 35334 12130 35386
rect 12142 35334 12194 35386
rect 12206 35334 12258 35386
rect 16950 35334 17002 35386
rect 17014 35334 17066 35386
rect 17078 35334 17130 35386
rect 17142 35334 17194 35386
rect 17206 35334 17258 35386
rect 13728 35232 13780 35284
rect 18696 35164 18748 35216
rect 8392 35096 8444 35148
rect 8208 35071 8260 35080
rect 8208 35037 8217 35071
rect 8217 35037 8251 35071
rect 8251 35037 8260 35071
rect 8208 35028 8260 35037
rect 8760 35028 8812 35080
rect 13544 35096 13596 35148
rect 13728 35096 13780 35148
rect 12532 35028 12584 35080
rect 12992 35028 13044 35080
rect 15844 35028 15896 35080
rect 4804 34960 4856 35012
rect 10324 34960 10376 35012
rect 12440 34960 12492 35012
rect 13084 34960 13136 35012
rect 8208 34892 8260 34944
rect 9680 34892 9732 34944
rect 13268 34892 13320 34944
rect 13544 34892 13596 34944
rect 15016 34892 15068 34944
rect 2610 34790 2662 34842
rect 2674 34790 2726 34842
rect 2738 34790 2790 34842
rect 2802 34790 2854 34842
rect 2866 34790 2918 34842
rect 7610 34790 7662 34842
rect 7674 34790 7726 34842
rect 7738 34790 7790 34842
rect 7802 34790 7854 34842
rect 7866 34790 7918 34842
rect 12610 34790 12662 34842
rect 12674 34790 12726 34842
rect 12738 34790 12790 34842
rect 12802 34790 12854 34842
rect 12866 34790 12918 34842
rect 17610 34790 17662 34842
rect 17674 34790 17726 34842
rect 17738 34790 17790 34842
rect 17802 34790 17854 34842
rect 17866 34790 17918 34842
rect 2412 34620 2464 34672
rect 5356 34688 5408 34740
rect 3240 34663 3292 34672
rect 3240 34629 3249 34663
rect 3249 34629 3283 34663
rect 3283 34629 3292 34663
rect 3240 34620 3292 34629
rect 4896 34552 4948 34604
rect 8024 34552 8076 34604
rect 10140 34731 10192 34740
rect 10140 34697 10149 34731
rect 10149 34697 10183 34731
rect 10183 34697 10192 34731
rect 10140 34688 10192 34697
rect 9496 34620 9548 34672
rect 13176 34552 13228 34604
rect 13268 34552 13320 34604
rect 13820 34620 13872 34672
rect 15108 34688 15160 34740
rect 15384 34731 15436 34740
rect 15384 34697 15393 34731
rect 15393 34697 15427 34731
rect 15427 34697 15436 34731
rect 15384 34688 15436 34697
rect 7288 34484 7340 34536
rect 8760 34527 8812 34536
rect 8760 34493 8769 34527
rect 8769 34493 8803 34527
rect 8803 34493 8812 34527
rect 8760 34484 8812 34493
rect 12440 34484 12492 34536
rect 15016 34595 15068 34604
rect 15016 34561 15025 34595
rect 15025 34561 15059 34595
rect 15059 34561 15068 34595
rect 15016 34552 15068 34561
rect 12992 34416 13044 34468
rect 13268 34416 13320 34468
rect 7288 34348 7340 34400
rect 17408 34416 17460 34468
rect 1950 34246 2002 34298
rect 2014 34246 2066 34298
rect 2078 34246 2130 34298
rect 2142 34246 2194 34298
rect 2206 34246 2258 34298
rect 6950 34246 7002 34298
rect 7014 34246 7066 34298
rect 7078 34246 7130 34298
rect 7142 34246 7194 34298
rect 7206 34246 7258 34298
rect 11950 34246 12002 34298
rect 12014 34246 12066 34298
rect 12078 34246 12130 34298
rect 12142 34246 12194 34298
rect 12206 34246 12258 34298
rect 16950 34246 17002 34298
rect 17014 34246 17066 34298
rect 17078 34246 17130 34298
rect 17142 34246 17194 34298
rect 17206 34246 17258 34298
rect 16764 34076 16816 34128
rect 17408 34051 17460 34060
rect 17408 34017 17417 34051
rect 17417 34017 17451 34051
rect 17451 34017 17460 34051
rect 17408 34008 17460 34017
rect 16304 33983 16356 33992
rect 16304 33949 16313 33983
rect 16313 33949 16347 33983
rect 16347 33949 16356 33983
rect 16304 33940 16356 33949
rect 7012 33872 7064 33924
rect 16120 33847 16172 33856
rect 16120 33813 16129 33847
rect 16129 33813 16163 33847
rect 16163 33813 16172 33847
rect 16120 33804 16172 33813
rect 16488 33804 16540 33856
rect 2610 33702 2662 33754
rect 2674 33702 2726 33754
rect 2738 33702 2790 33754
rect 2802 33702 2854 33754
rect 2866 33702 2918 33754
rect 7610 33702 7662 33754
rect 7674 33702 7726 33754
rect 7738 33702 7790 33754
rect 7802 33702 7854 33754
rect 7866 33702 7918 33754
rect 12610 33702 12662 33754
rect 12674 33702 12726 33754
rect 12738 33702 12790 33754
rect 12802 33702 12854 33754
rect 12866 33702 12918 33754
rect 17610 33702 17662 33754
rect 17674 33702 17726 33754
rect 17738 33702 17790 33754
rect 17802 33702 17854 33754
rect 17866 33702 17918 33754
rect 15568 33643 15620 33652
rect 15568 33609 15577 33643
rect 15577 33609 15611 33643
rect 15611 33609 15620 33643
rect 15568 33600 15620 33609
rect 15752 33600 15804 33652
rect 16488 33600 16540 33652
rect 14004 33464 14056 33516
rect 9036 33396 9088 33448
rect 3240 33260 3292 33312
rect 6644 33260 6696 33312
rect 7012 33260 7064 33312
rect 18236 33303 18288 33312
rect 18236 33269 18245 33303
rect 18245 33269 18279 33303
rect 18279 33269 18288 33303
rect 18236 33260 18288 33269
rect 1950 33158 2002 33210
rect 2014 33158 2066 33210
rect 2078 33158 2130 33210
rect 2142 33158 2194 33210
rect 2206 33158 2258 33210
rect 6950 33158 7002 33210
rect 7014 33158 7066 33210
rect 7078 33158 7130 33210
rect 7142 33158 7194 33210
rect 7206 33158 7258 33210
rect 11950 33158 12002 33210
rect 12014 33158 12066 33210
rect 12078 33158 12130 33210
rect 12142 33158 12194 33210
rect 12206 33158 12258 33210
rect 16950 33158 17002 33210
rect 17014 33158 17066 33210
rect 17078 33158 17130 33210
rect 17142 33158 17194 33210
rect 17206 33158 17258 33210
rect 4620 33056 4672 33108
rect 6736 33056 6788 33108
rect 16488 33056 16540 33108
rect 19524 33056 19576 33108
rect 13820 32920 13872 32972
rect 16856 32852 16908 32904
rect 16120 32784 16172 32836
rect 2610 32614 2662 32666
rect 2674 32614 2726 32666
rect 2738 32614 2790 32666
rect 2802 32614 2854 32666
rect 2866 32614 2918 32666
rect 7610 32614 7662 32666
rect 7674 32614 7726 32666
rect 7738 32614 7790 32666
rect 7802 32614 7854 32666
rect 7866 32614 7918 32666
rect 12610 32614 12662 32666
rect 12674 32614 12726 32666
rect 12738 32614 12790 32666
rect 12802 32614 12854 32666
rect 12866 32614 12918 32666
rect 17610 32614 17662 32666
rect 17674 32614 17726 32666
rect 17738 32614 17790 32666
rect 17802 32614 17854 32666
rect 17866 32614 17918 32666
rect 7472 32512 7524 32564
rect 13360 32512 13412 32564
rect 7472 32376 7524 32428
rect 8300 32376 8352 32428
rect 13820 32444 13872 32496
rect 16856 32419 16908 32428
rect 16856 32385 16865 32419
rect 16865 32385 16899 32419
rect 16899 32385 16908 32419
rect 16856 32376 16908 32385
rect 18420 32376 18472 32428
rect 7288 32308 7340 32360
rect 8392 32308 8444 32360
rect 2412 32240 2464 32292
rect 11520 32240 11572 32292
rect 6736 32172 6788 32224
rect 6920 32172 6972 32224
rect 7288 32172 7340 32224
rect 11796 32172 11848 32224
rect 17960 32172 18012 32224
rect 18420 32172 18472 32224
rect 1950 32070 2002 32122
rect 2014 32070 2066 32122
rect 2078 32070 2130 32122
rect 2142 32070 2194 32122
rect 2206 32070 2258 32122
rect 6950 32070 7002 32122
rect 7014 32070 7066 32122
rect 7078 32070 7130 32122
rect 7142 32070 7194 32122
rect 7206 32070 7258 32122
rect 11950 32070 12002 32122
rect 12014 32070 12066 32122
rect 12078 32070 12130 32122
rect 12142 32070 12194 32122
rect 12206 32070 12258 32122
rect 16950 32070 17002 32122
rect 17014 32070 17066 32122
rect 17078 32070 17130 32122
rect 17142 32070 17194 32122
rect 17206 32070 17258 32122
rect 11336 31968 11388 32020
rect 11520 31968 11572 32020
rect 16488 31968 16540 32020
rect 6460 31832 6512 31884
rect 9496 31832 9548 31884
rect 16764 31832 16816 31884
rect 16488 31764 16540 31816
rect 16580 31764 16632 31816
rect 18052 31807 18104 31816
rect 18052 31773 18061 31807
rect 18061 31773 18095 31807
rect 18095 31773 18104 31807
rect 18052 31764 18104 31773
rect 8024 31696 8076 31748
rect 6920 31628 6972 31680
rect 8116 31628 8168 31680
rect 8300 31628 8352 31680
rect 18236 31671 18288 31680
rect 18236 31637 18245 31671
rect 18245 31637 18279 31671
rect 18279 31637 18288 31671
rect 18236 31628 18288 31637
rect 2610 31526 2662 31578
rect 2674 31526 2726 31578
rect 2738 31526 2790 31578
rect 2802 31526 2854 31578
rect 2866 31526 2918 31578
rect 7610 31526 7662 31578
rect 7674 31526 7726 31578
rect 7738 31526 7790 31578
rect 7802 31526 7854 31578
rect 7866 31526 7918 31578
rect 12610 31526 12662 31578
rect 12674 31526 12726 31578
rect 12738 31526 12790 31578
rect 12802 31526 12854 31578
rect 12866 31526 12918 31578
rect 17610 31526 17662 31578
rect 17674 31526 17726 31578
rect 17738 31526 17790 31578
rect 17802 31526 17854 31578
rect 17866 31526 17918 31578
rect 6920 31424 6972 31476
rect 14740 31424 14792 31476
rect 6368 31356 6420 31408
rect 1768 31331 1820 31340
rect 1768 31297 1777 31331
rect 1777 31297 1811 31331
rect 1811 31297 1820 31331
rect 1768 31288 1820 31297
rect 7288 31288 7340 31340
rect 7380 31288 7432 31340
rect 8208 31288 8260 31340
rect 16856 31331 16908 31340
rect 16856 31297 16865 31331
rect 16865 31297 16899 31331
rect 16899 31297 16908 31331
rect 16856 31288 16908 31297
rect 7288 31084 7340 31136
rect 1950 30982 2002 31034
rect 2014 30982 2066 31034
rect 2078 30982 2130 31034
rect 2142 30982 2194 31034
rect 2206 30982 2258 31034
rect 6950 30982 7002 31034
rect 7014 30982 7066 31034
rect 7078 30982 7130 31034
rect 7142 30982 7194 31034
rect 7206 30982 7258 31034
rect 11950 30982 12002 31034
rect 12014 30982 12066 31034
rect 12078 30982 12130 31034
rect 12142 30982 12194 31034
rect 12206 30982 12258 31034
rect 16950 30982 17002 31034
rect 17014 30982 17066 31034
rect 17078 30982 17130 31034
rect 17142 30982 17194 31034
rect 17206 30982 17258 31034
rect 6368 30787 6420 30796
rect 6368 30753 6377 30787
rect 6377 30753 6411 30787
rect 6411 30753 6420 30787
rect 6368 30744 6420 30753
rect 11244 30608 11296 30660
rect 5724 30583 5776 30592
rect 5724 30549 5733 30583
rect 5733 30549 5767 30583
rect 5767 30549 5776 30583
rect 5724 30540 5776 30549
rect 9128 30540 9180 30592
rect 13268 30608 13320 30660
rect 13728 30608 13780 30660
rect 19524 30540 19576 30592
rect 2610 30438 2662 30490
rect 2674 30438 2726 30490
rect 2738 30438 2790 30490
rect 2802 30438 2854 30490
rect 2866 30438 2918 30490
rect 7610 30438 7662 30490
rect 7674 30438 7726 30490
rect 7738 30438 7790 30490
rect 7802 30438 7854 30490
rect 7866 30438 7918 30490
rect 12610 30438 12662 30490
rect 12674 30438 12726 30490
rect 12738 30438 12790 30490
rect 12802 30438 12854 30490
rect 12866 30438 12918 30490
rect 17610 30438 17662 30490
rect 17674 30438 17726 30490
rect 17738 30438 17790 30490
rect 17802 30438 17854 30490
rect 17866 30438 17918 30490
rect 7288 30268 7340 30320
rect 7564 30268 7616 30320
rect 8024 30311 8076 30320
rect 8024 30277 8047 30311
rect 8047 30277 8076 30311
rect 8024 30268 8076 30277
rect 3240 30243 3292 30252
rect 3240 30209 3249 30243
rect 3249 30209 3283 30243
rect 3283 30209 3292 30243
rect 3240 30200 3292 30209
rect 3792 30243 3844 30252
rect 3792 30209 3801 30243
rect 3801 30209 3835 30243
rect 3835 30209 3844 30243
rect 3792 30200 3844 30209
rect 7748 30243 7800 30252
rect 7748 30209 7757 30243
rect 7757 30209 7791 30243
rect 7791 30209 7800 30243
rect 7748 30200 7800 30209
rect 13268 30268 13320 30320
rect 13636 30268 13688 30320
rect 18880 30268 18932 30320
rect 13820 30200 13872 30252
rect 6644 30039 6696 30048
rect 6644 30005 6653 30039
rect 6653 30005 6687 30039
rect 6687 30005 6696 30039
rect 6644 29996 6696 30005
rect 11796 30132 11848 30184
rect 17500 30200 17552 30252
rect 10048 29996 10100 30048
rect 16396 30064 16448 30116
rect 15936 30039 15988 30048
rect 15936 30005 15945 30039
rect 15945 30005 15979 30039
rect 15979 30005 15988 30039
rect 15936 29996 15988 30005
rect 1950 29894 2002 29946
rect 2014 29894 2066 29946
rect 2078 29894 2130 29946
rect 2142 29894 2194 29946
rect 2206 29894 2258 29946
rect 6950 29894 7002 29946
rect 7014 29894 7066 29946
rect 7078 29894 7130 29946
rect 7142 29894 7194 29946
rect 7206 29894 7258 29946
rect 11950 29894 12002 29946
rect 12014 29894 12066 29946
rect 12078 29894 12130 29946
rect 12142 29894 12194 29946
rect 12206 29894 12258 29946
rect 16950 29894 17002 29946
rect 17014 29894 17066 29946
rect 17078 29894 17130 29946
rect 17142 29894 17194 29946
rect 17206 29894 17258 29946
rect 3240 29792 3292 29844
rect 14188 29792 14240 29844
rect 15660 29835 15712 29844
rect 15660 29801 15669 29835
rect 15669 29801 15703 29835
rect 15703 29801 15712 29835
rect 15660 29792 15712 29801
rect 6644 29724 6696 29776
rect 19340 29724 19392 29776
rect 7288 29656 7340 29708
rect 7748 29656 7800 29708
rect 8760 29656 8812 29708
rect 9128 29656 9180 29708
rect 15936 29656 15988 29708
rect 17960 29656 18012 29708
rect 19616 29656 19668 29708
rect 18604 29588 18656 29640
rect 7564 29452 7616 29504
rect 9404 29452 9456 29504
rect 15476 29452 15528 29504
rect 16028 29495 16080 29504
rect 16028 29461 16037 29495
rect 16037 29461 16071 29495
rect 16071 29461 16080 29495
rect 16028 29452 16080 29461
rect 16120 29495 16172 29504
rect 16120 29461 16129 29495
rect 16129 29461 16163 29495
rect 16163 29461 16172 29495
rect 16120 29452 16172 29461
rect 18236 29495 18288 29504
rect 18236 29461 18245 29495
rect 18245 29461 18279 29495
rect 18279 29461 18288 29495
rect 18236 29452 18288 29461
rect 2610 29350 2662 29402
rect 2674 29350 2726 29402
rect 2738 29350 2790 29402
rect 2802 29350 2854 29402
rect 2866 29350 2918 29402
rect 7610 29350 7662 29402
rect 7674 29350 7726 29402
rect 7738 29350 7790 29402
rect 7802 29350 7854 29402
rect 7866 29350 7918 29402
rect 12610 29350 12662 29402
rect 12674 29350 12726 29402
rect 12738 29350 12790 29402
rect 12802 29350 12854 29402
rect 12866 29350 12918 29402
rect 17610 29350 17662 29402
rect 17674 29350 17726 29402
rect 17738 29350 17790 29402
rect 17802 29350 17854 29402
rect 17866 29350 17918 29402
rect 5448 29248 5500 29300
rect 4620 29223 4672 29232
rect 4620 29189 4629 29223
rect 4629 29189 4663 29223
rect 4663 29189 4672 29223
rect 4620 29180 4672 29189
rect 7932 29180 7984 29232
rect 8392 29180 8444 29232
rect 4436 29155 4488 29164
rect 4436 29121 4445 29155
rect 4445 29121 4479 29155
rect 4479 29121 4488 29155
rect 4436 29112 4488 29121
rect 10968 29112 11020 29164
rect 8760 29044 8812 29096
rect 9128 29044 9180 29096
rect 10048 29087 10100 29096
rect 10048 29053 10057 29087
rect 10057 29053 10091 29087
rect 10091 29053 10100 29087
rect 10048 29044 10100 29053
rect 6368 28976 6420 29028
rect 10692 29044 10744 29096
rect 1950 28806 2002 28858
rect 2014 28806 2066 28858
rect 2078 28806 2130 28858
rect 2142 28806 2194 28858
rect 2206 28806 2258 28858
rect 6950 28806 7002 28858
rect 7014 28806 7066 28858
rect 7078 28806 7130 28858
rect 7142 28806 7194 28858
rect 7206 28806 7258 28858
rect 11950 28806 12002 28858
rect 12014 28806 12066 28858
rect 12078 28806 12130 28858
rect 12142 28806 12194 28858
rect 12206 28806 12258 28858
rect 16950 28806 17002 28858
rect 17014 28806 17066 28858
rect 17078 28806 17130 28858
rect 17142 28806 17194 28858
rect 17206 28806 17258 28858
rect 11060 28704 11112 28756
rect 9128 28568 9180 28620
rect 9772 28611 9824 28620
rect 9772 28577 9781 28611
rect 9781 28577 9815 28611
rect 9815 28577 9824 28611
rect 9772 28568 9824 28577
rect 5632 28543 5684 28552
rect 5632 28509 5641 28543
rect 5641 28509 5675 28543
rect 5675 28509 5684 28543
rect 5632 28500 5684 28509
rect 9864 28475 9916 28484
rect 9864 28441 9873 28475
rect 9873 28441 9907 28475
rect 9907 28441 9916 28475
rect 9864 28432 9916 28441
rect 10600 28432 10652 28484
rect 10508 28364 10560 28416
rect 2610 28262 2662 28314
rect 2674 28262 2726 28314
rect 2738 28262 2790 28314
rect 2802 28262 2854 28314
rect 2866 28262 2918 28314
rect 7610 28262 7662 28314
rect 7674 28262 7726 28314
rect 7738 28262 7790 28314
rect 7802 28262 7854 28314
rect 7866 28262 7918 28314
rect 12610 28262 12662 28314
rect 12674 28262 12726 28314
rect 12738 28262 12790 28314
rect 12802 28262 12854 28314
rect 12866 28262 12918 28314
rect 17610 28262 17662 28314
rect 17674 28262 17726 28314
rect 17738 28262 17790 28314
rect 17802 28262 17854 28314
rect 17866 28262 17918 28314
rect 3332 28092 3384 28144
rect 10784 28024 10836 28076
rect 4068 27999 4120 28008
rect 4068 27965 4077 27999
rect 4077 27965 4111 27999
rect 4111 27965 4120 27999
rect 4068 27956 4120 27965
rect 10968 27820 11020 27872
rect 17868 27820 17920 27872
rect 1950 27718 2002 27770
rect 2014 27718 2066 27770
rect 2078 27718 2130 27770
rect 2142 27718 2194 27770
rect 2206 27718 2258 27770
rect 6950 27718 7002 27770
rect 7014 27718 7066 27770
rect 7078 27718 7130 27770
rect 7142 27718 7194 27770
rect 7206 27718 7258 27770
rect 11950 27718 12002 27770
rect 12014 27718 12066 27770
rect 12078 27718 12130 27770
rect 12142 27718 12194 27770
rect 12206 27718 12258 27770
rect 16950 27718 17002 27770
rect 17014 27718 17066 27770
rect 17078 27718 17130 27770
rect 17142 27718 17194 27770
rect 17206 27718 17258 27770
rect 4068 27548 4120 27600
rect 7288 27548 7340 27600
rect 10876 27548 10928 27600
rect 13912 27548 13964 27600
rect 19156 27548 19208 27600
rect 4160 27480 4212 27532
rect 5080 27412 5132 27464
rect 18144 27412 18196 27464
rect 2610 27174 2662 27226
rect 2674 27174 2726 27226
rect 2738 27174 2790 27226
rect 2802 27174 2854 27226
rect 2866 27174 2918 27226
rect 7610 27174 7662 27226
rect 7674 27174 7726 27226
rect 7738 27174 7790 27226
rect 7802 27174 7854 27226
rect 7866 27174 7918 27226
rect 12610 27174 12662 27226
rect 12674 27174 12726 27226
rect 12738 27174 12790 27226
rect 12802 27174 12854 27226
rect 12866 27174 12918 27226
rect 17610 27174 17662 27226
rect 17674 27174 17726 27226
rect 17738 27174 17790 27226
rect 17802 27174 17854 27226
rect 17866 27174 17918 27226
rect 8392 27072 8444 27124
rect 9496 27072 9548 27124
rect 13820 27004 13872 27056
rect 1584 26936 1636 26988
rect 13268 26979 13320 26988
rect 13268 26945 13277 26979
rect 13277 26945 13311 26979
rect 13311 26945 13320 26979
rect 13268 26936 13320 26945
rect 1492 26732 1544 26784
rect 8668 26868 8720 26920
rect 9036 26868 9088 26920
rect 11796 26868 11848 26920
rect 1950 26630 2002 26682
rect 2014 26630 2066 26682
rect 2078 26630 2130 26682
rect 2142 26630 2194 26682
rect 2206 26630 2258 26682
rect 6950 26630 7002 26682
rect 7014 26630 7066 26682
rect 7078 26630 7130 26682
rect 7142 26630 7194 26682
rect 7206 26630 7258 26682
rect 11950 26630 12002 26682
rect 12014 26630 12066 26682
rect 12078 26630 12130 26682
rect 12142 26630 12194 26682
rect 12206 26630 12258 26682
rect 16950 26630 17002 26682
rect 17014 26630 17066 26682
rect 17078 26630 17130 26682
rect 17142 26630 17194 26682
rect 17206 26630 17258 26682
rect 6184 26528 6236 26580
rect 7380 26528 7432 26580
rect 4068 26392 4120 26444
rect 11520 26324 11572 26376
rect 5816 26299 5868 26308
rect 5816 26265 5850 26299
rect 5850 26265 5868 26299
rect 5816 26256 5868 26265
rect 7288 26256 7340 26308
rect 13268 26256 13320 26308
rect 7380 26188 7432 26240
rect 8300 26188 8352 26240
rect 2610 26086 2662 26138
rect 2674 26086 2726 26138
rect 2738 26086 2790 26138
rect 2802 26086 2854 26138
rect 2866 26086 2918 26138
rect 7610 26086 7662 26138
rect 7674 26086 7726 26138
rect 7738 26086 7790 26138
rect 7802 26086 7854 26138
rect 7866 26086 7918 26138
rect 12610 26086 12662 26138
rect 12674 26086 12726 26138
rect 12738 26086 12790 26138
rect 12802 26086 12854 26138
rect 12866 26086 12918 26138
rect 17610 26086 17662 26138
rect 17674 26086 17726 26138
rect 17738 26086 17790 26138
rect 17802 26086 17854 26138
rect 17866 26086 17918 26138
rect 10140 26027 10192 26036
rect 10140 25993 10149 26027
rect 10149 25993 10183 26027
rect 10183 25993 10192 26027
rect 10140 25984 10192 25993
rect 13728 25984 13780 26036
rect 17500 25984 17552 26036
rect 9680 25780 9732 25832
rect 14648 25848 14700 25900
rect 18972 25848 19024 25900
rect 10784 25823 10836 25832
rect 10784 25789 10793 25823
rect 10793 25789 10827 25823
rect 10827 25789 10836 25823
rect 10784 25780 10836 25789
rect 18236 25687 18288 25696
rect 18236 25653 18245 25687
rect 18245 25653 18279 25687
rect 18279 25653 18288 25687
rect 18236 25644 18288 25653
rect 1950 25542 2002 25594
rect 2014 25542 2066 25594
rect 2078 25542 2130 25594
rect 2142 25542 2194 25594
rect 2206 25542 2258 25594
rect 6950 25542 7002 25594
rect 7014 25542 7066 25594
rect 7078 25542 7130 25594
rect 7142 25542 7194 25594
rect 7206 25542 7258 25594
rect 11950 25542 12002 25594
rect 12014 25542 12066 25594
rect 12078 25542 12130 25594
rect 12142 25542 12194 25594
rect 12206 25542 12258 25594
rect 16950 25542 17002 25594
rect 17014 25542 17066 25594
rect 17078 25542 17130 25594
rect 17142 25542 17194 25594
rect 17206 25542 17258 25594
rect 1768 25440 1820 25492
rect 5356 25483 5408 25492
rect 5356 25449 5365 25483
rect 5365 25449 5399 25483
rect 5399 25449 5408 25483
rect 5356 25440 5408 25449
rect 1492 25304 1544 25356
rect 1768 25304 1820 25356
rect 5724 25304 5776 25356
rect 7380 25304 7432 25356
rect 10324 25347 10376 25356
rect 10324 25313 10333 25347
rect 10333 25313 10367 25347
rect 10367 25313 10376 25347
rect 10324 25304 10376 25313
rect 10416 25347 10468 25356
rect 10416 25313 10425 25347
rect 10425 25313 10459 25347
rect 10459 25313 10468 25347
rect 10416 25304 10468 25313
rect 12532 25304 12584 25356
rect 13360 25304 13412 25356
rect 4068 25236 4120 25288
rect 10232 25279 10284 25288
rect 10232 25245 10241 25279
rect 10241 25245 10275 25279
rect 10275 25245 10284 25279
rect 10232 25236 10284 25245
rect 12440 25236 12492 25288
rect 12992 25236 13044 25288
rect 1492 25168 1544 25220
rect 2320 25168 2372 25220
rect 11520 25168 11572 25220
rect 13084 25168 13136 25220
rect 15844 25168 15896 25220
rect 10508 25100 10560 25152
rect 2610 24998 2662 25050
rect 2674 24998 2726 25050
rect 2738 24998 2790 25050
rect 2802 24998 2854 25050
rect 2866 24998 2918 25050
rect 7610 24998 7662 25050
rect 7674 24998 7726 25050
rect 7738 24998 7790 25050
rect 7802 24998 7854 25050
rect 7866 24998 7918 25050
rect 12610 24998 12662 25050
rect 12674 24998 12726 25050
rect 12738 24998 12790 25050
rect 12802 24998 12854 25050
rect 12866 24998 12918 25050
rect 17610 24998 17662 25050
rect 17674 24998 17726 25050
rect 17738 24998 17790 25050
rect 17802 24998 17854 25050
rect 17866 24998 17918 25050
rect 11428 24896 11480 24948
rect 13820 24896 13872 24948
rect 6736 24760 6788 24812
rect 9772 24803 9824 24812
rect 9772 24769 9781 24803
rect 9781 24769 9815 24803
rect 9815 24769 9824 24803
rect 9772 24760 9824 24769
rect 14832 24760 14884 24812
rect 17960 24760 18012 24812
rect 14740 24692 14792 24744
rect 15108 24692 15160 24744
rect 16396 24692 16448 24744
rect 18144 24735 18196 24744
rect 18144 24701 18153 24735
rect 18153 24701 18187 24735
rect 18187 24701 18196 24735
rect 18144 24692 18196 24701
rect 14280 24624 14332 24676
rect 8944 24556 8996 24608
rect 1950 24454 2002 24506
rect 2014 24454 2066 24506
rect 2078 24454 2130 24506
rect 2142 24454 2194 24506
rect 2206 24454 2258 24506
rect 6950 24454 7002 24506
rect 7014 24454 7066 24506
rect 7078 24454 7130 24506
rect 7142 24454 7194 24506
rect 7206 24454 7258 24506
rect 11950 24454 12002 24506
rect 12014 24454 12066 24506
rect 12078 24454 12130 24506
rect 12142 24454 12194 24506
rect 12206 24454 12258 24506
rect 16950 24454 17002 24506
rect 17014 24454 17066 24506
rect 17078 24454 17130 24506
rect 17142 24454 17194 24506
rect 17206 24454 17258 24506
rect 14740 24148 14792 24200
rect 6276 24080 6328 24132
rect 13084 24080 13136 24132
rect 13728 24080 13780 24132
rect 18236 24055 18288 24064
rect 18236 24021 18245 24055
rect 18245 24021 18279 24055
rect 18279 24021 18288 24055
rect 18236 24012 18288 24021
rect 2610 23910 2662 23962
rect 2674 23910 2726 23962
rect 2738 23910 2790 23962
rect 2802 23910 2854 23962
rect 2866 23910 2918 23962
rect 7610 23910 7662 23962
rect 7674 23910 7726 23962
rect 7738 23910 7790 23962
rect 7802 23910 7854 23962
rect 7866 23910 7918 23962
rect 12610 23910 12662 23962
rect 12674 23910 12726 23962
rect 12738 23910 12790 23962
rect 12802 23910 12854 23962
rect 12866 23910 12918 23962
rect 17610 23910 17662 23962
rect 17674 23910 17726 23962
rect 17738 23910 17790 23962
rect 17802 23910 17854 23962
rect 17866 23910 17918 23962
rect 9312 23851 9364 23860
rect 9312 23817 9321 23851
rect 9321 23817 9355 23851
rect 9355 23817 9364 23851
rect 9312 23808 9364 23817
rect 16672 23808 16724 23860
rect 7380 23740 7432 23792
rect 13728 23740 13780 23792
rect 6460 23672 6512 23724
rect 7288 23672 7340 23724
rect 12532 23672 12584 23724
rect 16580 23604 16632 23656
rect 11336 23468 11388 23520
rect 16948 23579 17000 23588
rect 16948 23545 16957 23579
rect 16957 23545 16991 23579
rect 16991 23545 17000 23579
rect 16948 23536 17000 23545
rect 16764 23468 16816 23520
rect 1950 23366 2002 23418
rect 2014 23366 2066 23418
rect 2078 23366 2130 23418
rect 2142 23366 2194 23418
rect 2206 23366 2258 23418
rect 6950 23366 7002 23418
rect 7014 23366 7066 23418
rect 7078 23366 7130 23418
rect 7142 23366 7194 23418
rect 7206 23366 7258 23418
rect 11950 23366 12002 23418
rect 12014 23366 12066 23418
rect 12078 23366 12130 23418
rect 12142 23366 12194 23418
rect 12206 23366 12258 23418
rect 16950 23366 17002 23418
rect 17014 23366 17066 23418
rect 17078 23366 17130 23418
rect 17142 23366 17194 23418
rect 17206 23366 17258 23418
rect 18052 23264 18104 23316
rect 18420 23264 18472 23316
rect 2610 22822 2662 22874
rect 2674 22822 2726 22874
rect 2738 22822 2790 22874
rect 2802 22822 2854 22874
rect 2866 22822 2918 22874
rect 7610 22822 7662 22874
rect 7674 22822 7726 22874
rect 7738 22822 7790 22874
rect 7802 22822 7854 22874
rect 7866 22822 7918 22874
rect 12610 22822 12662 22874
rect 12674 22822 12726 22874
rect 12738 22822 12790 22874
rect 12802 22822 12854 22874
rect 12866 22822 12918 22874
rect 17610 22822 17662 22874
rect 17674 22822 17726 22874
rect 17738 22822 17790 22874
rect 17802 22822 17854 22874
rect 17866 22822 17918 22874
rect 7932 22720 7984 22772
rect 8208 22720 8260 22772
rect 10324 22720 10376 22772
rect 13360 22720 13412 22772
rect 5540 22584 5592 22636
rect 9864 22584 9916 22636
rect 18052 22516 18104 22568
rect 17224 22491 17276 22500
rect 17224 22457 17233 22491
rect 17233 22457 17267 22491
rect 17267 22457 17276 22491
rect 17224 22448 17276 22457
rect 1950 22278 2002 22330
rect 2014 22278 2066 22330
rect 2078 22278 2130 22330
rect 2142 22278 2194 22330
rect 2206 22278 2258 22330
rect 6950 22278 7002 22330
rect 7014 22278 7066 22330
rect 7078 22278 7130 22330
rect 7142 22278 7194 22330
rect 7206 22278 7258 22330
rect 11950 22278 12002 22330
rect 12014 22278 12066 22330
rect 12078 22278 12130 22330
rect 12142 22278 12194 22330
rect 12206 22278 12258 22330
rect 16950 22278 17002 22330
rect 17014 22278 17066 22330
rect 17078 22278 17130 22330
rect 17142 22278 17194 22330
rect 17206 22278 17258 22330
rect 1400 22040 1452 22092
rect 4160 22040 4212 22092
rect 6184 22040 6236 22092
rect 9220 22108 9272 22160
rect 9772 22108 9824 22160
rect 16212 22108 16264 22160
rect 7104 22040 7156 22092
rect 6920 21972 6972 22024
rect 9496 21972 9548 22024
rect 15200 21972 15252 22024
rect 18052 22015 18104 22024
rect 18052 21981 18061 22015
rect 18061 21981 18095 22015
rect 18095 21981 18104 22015
rect 18052 21972 18104 21981
rect 3332 21904 3384 21956
rect 6460 21836 6512 21888
rect 6644 21836 6696 21888
rect 7288 21904 7340 21956
rect 7104 21836 7156 21888
rect 7932 21836 7984 21888
rect 8208 21836 8260 21888
rect 11244 21836 11296 21888
rect 12348 21836 12400 21888
rect 14096 21836 14148 21888
rect 18236 21879 18288 21888
rect 18236 21845 18245 21879
rect 18245 21845 18279 21879
rect 18279 21845 18288 21879
rect 18236 21836 18288 21845
rect 2610 21734 2662 21786
rect 2674 21734 2726 21786
rect 2738 21734 2790 21786
rect 2802 21734 2854 21786
rect 2866 21734 2918 21786
rect 7610 21734 7662 21786
rect 7674 21734 7726 21786
rect 7738 21734 7790 21786
rect 7802 21734 7854 21786
rect 7866 21734 7918 21786
rect 12610 21734 12662 21786
rect 12674 21734 12726 21786
rect 12738 21734 12790 21786
rect 12802 21734 12854 21786
rect 12866 21734 12918 21786
rect 17610 21734 17662 21786
rect 17674 21734 17726 21786
rect 17738 21734 17790 21786
rect 17802 21734 17854 21786
rect 17866 21734 17918 21786
rect 3332 21632 3384 21684
rect 10784 21632 10836 21684
rect 19892 21632 19944 21684
rect 3148 21496 3200 21548
rect 6460 21428 6512 21480
rect 11428 21428 11480 21480
rect 12348 21292 12400 21344
rect 18788 21292 18840 21344
rect 1950 21190 2002 21242
rect 2014 21190 2066 21242
rect 2078 21190 2130 21242
rect 2142 21190 2194 21242
rect 2206 21190 2258 21242
rect 6950 21190 7002 21242
rect 7014 21190 7066 21242
rect 7078 21190 7130 21242
rect 7142 21190 7194 21242
rect 7206 21190 7258 21242
rect 11950 21190 12002 21242
rect 12014 21190 12066 21242
rect 12078 21190 12130 21242
rect 12142 21190 12194 21242
rect 12206 21190 12258 21242
rect 16950 21190 17002 21242
rect 17014 21190 17066 21242
rect 17078 21190 17130 21242
rect 17142 21190 17194 21242
rect 17206 21190 17258 21242
rect 9128 21131 9180 21140
rect 9128 21097 9137 21131
rect 9137 21097 9171 21131
rect 9171 21097 9180 21131
rect 9128 21088 9180 21097
rect 12992 21088 13044 21140
rect 9680 21020 9732 21072
rect 6828 20952 6880 21004
rect 9404 20952 9456 21004
rect 13268 21020 13320 21072
rect 15016 21020 15068 21072
rect 13728 20952 13780 21004
rect 12348 20884 12400 20936
rect 14188 20884 14240 20936
rect 14648 20927 14700 20936
rect 14648 20893 14657 20927
rect 14657 20893 14691 20927
rect 14691 20893 14700 20927
rect 14648 20884 14700 20893
rect 10784 20816 10836 20868
rect 14832 20816 14884 20868
rect 9312 20748 9364 20800
rect 15660 20748 15712 20800
rect 15936 20748 15988 20800
rect 2610 20646 2662 20698
rect 2674 20646 2726 20698
rect 2738 20646 2790 20698
rect 2802 20646 2854 20698
rect 2866 20646 2918 20698
rect 7610 20646 7662 20698
rect 7674 20646 7726 20698
rect 7738 20646 7790 20698
rect 7802 20646 7854 20698
rect 7866 20646 7918 20698
rect 12610 20646 12662 20698
rect 12674 20646 12726 20698
rect 12738 20646 12790 20698
rect 12802 20646 12854 20698
rect 12866 20646 12918 20698
rect 17610 20646 17662 20698
rect 17674 20646 17726 20698
rect 17738 20646 17790 20698
rect 17802 20646 17854 20698
rect 17866 20646 17918 20698
rect 4344 20544 4396 20596
rect 8392 20476 8444 20528
rect 5540 20408 5592 20460
rect 11980 20544 12032 20596
rect 17224 20544 17276 20596
rect 14924 20519 14976 20528
rect 14924 20485 14933 20519
rect 14933 20485 14967 20519
rect 14967 20485 14976 20519
rect 14924 20476 14976 20485
rect 16488 20408 16540 20460
rect 1860 20272 1912 20324
rect 11428 20340 11480 20392
rect 13544 20340 13596 20392
rect 8668 20272 8720 20324
rect 13084 20315 13136 20324
rect 13084 20281 13093 20315
rect 13093 20281 13127 20315
rect 13127 20281 13136 20315
rect 13084 20272 13136 20281
rect 16304 20272 16356 20324
rect 16856 20272 16908 20324
rect 4436 20204 4488 20256
rect 11980 20204 12032 20256
rect 13268 20204 13320 20256
rect 18144 20340 18196 20392
rect 1950 20102 2002 20154
rect 2014 20102 2066 20154
rect 2078 20102 2130 20154
rect 2142 20102 2194 20154
rect 2206 20102 2258 20154
rect 6950 20102 7002 20154
rect 7014 20102 7066 20154
rect 7078 20102 7130 20154
rect 7142 20102 7194 20154
rect 7206 20102 7258 20154
rect 11950 20102 12002 20154
rect 12014 20102 12066 20154
rect 12078 20102 12130 20154
rect 12142 20102 12194 20154
rect 12206 20102 12258 20154
rect 16950 20102 17002 20154
rect 17014 20102 17066 20154
rect 17078 20102 17130 20154
rect 17142 20102 17194 20154
rect 17206 20102 17258 20154
rect 10600 20000 10652 20052
rect 11428 20000 11480 20052
rect 13728 20000 13780 20052
rect 14556 20000 14608 20052
rect 16856 20000 16908 20052
rect 18236 19975 18288 19984
rect 18236 19941 18245 19975
rect 18245 19941 18279 19975
rect 18279 19941 18288 19975
rect 18236 19932 18288 19941
rect 6000 19796 6052 19848
rect 2610 19558 2662 19610
rect 2674 19558 2726 19610
rect 2738 19558 2790 19610
rect 2802 19558 2854 19610
rect 2866 19558 2918 19610
rect 7610 19558 7662 19610
rect 7674 19558 7726 19610
rect 7738 19558 7790 19610
rect 7802 19558 7854 19610
rect 7866 19558 7918 19610
rect 12610 19558 12662 19610
rect 12674 19558 12726 19610
rect 12738 19558 12790 19610
rect 12802 19558 12854 19610
rect 12866 19558 12918 19610
rect 17610 19558 17662 19610
rect 17674 19558 17726 19610
rect 17738 19558 17790 19610
rect 17802 19558 17854 19610
rect 17866 19558 17918 19610
rect 14188 19456 14240 19508
rect 12164 19363 12216 19372
rect 12164 19329 12173 19363
rect 12173 19329 12207 19363
rect 12207 19329 12216 19363
rect 12164 19320 12216 19329
rect 1950 19014 2002 19066
rect 2014 19014 2066 19066
rect 2078 19014 2130 19066
rect 2142 19014 2194 19066
rect 2206 19014 2258 19066
rect 6950 19014 7002 19066
rect 7014 19014 7066 19066
rect 7078 19014 7130 19066
rect 7142 19014 7194 19066
rect 7206 19014 7258 19066
rect 11950 19014 12002 19066
rect 12014 19014 12066 19066
rect 12078 19014 12130 19066
rect 12142 19014 12194 19066
rect 12206 19014 12258 19066
rect 16950 19014 17002 19066
rect 17014 19014 17066 19066
rect 17078 19014 17130 19066
rect 17142 19014 17194 19066
rect 17206 19014 17258 19066
rect 2610 18470 2662 18522
rect 2674 18470 2726 18522
rect 2738 18470 2790 18522
rect 2802 18470 2854 18522
rect 2866 18470 2918 18522
rect 7610 18470 7662 18522
rect 7674 18470 7726 18522
rect 7738 18470 7790 18522
rect 7802 18470 7854 18522
rect 7866 18470 7918 18522
rect 12610 18470 12662 18522
rect 12674 18470 12726 18522
rect 12738 18470 12790 18522
rect 12802 18470 12854 18522
rect 12866 18470 12918 18522
rect 17610 18470 17662 18522
rect 17674 18470 17726 18522
rect 17738 18470 17790 18522
rect 17802 18470 17854 18522
rect 17866 18470 17918 18522
rect 18328 18368 18380 18420
rect 14188 18343 14240 18352
rect 14188 18309 14222 18343
rect 14222 18309 14240 18343
rect 14188 18300 14240 18309
rect 13728 18232 13780 18284
rect 19248 18232 19300 18284
rect 10324 18028 10376 18080
rect 11060 18028 11112 18080
rect 18236 18071 18288 18080
rect 18236 18037 18245 18071
rect 18245 18037 18279 18071
rect 18279 18037 18288 18071
rect 18236 18028 18288 18037
rect 1950 17926 2002 17978
rect 2014 17926 2066 17978
rect 2078 17926 2130 17978
rect 2142 17926 2194 17978
rect 2206 17926 2258 17978
rect 6950 17926 7002 17978
rect 7014 17926 7066 17978
rect 7078 17926 7130 17978
rect 7142 17926 7194 17978
rect 7206 17926 7258 17978
rect 11950 17926 12002 17978
rect 12014 17926 12066 17978
rect 12078 17926 12130 17978
rect 12142 17926 12194 17978
rect 12206 17926 12258 17978
rect 16950 17926 17002 17978
rect 17014 17926 17066 17978
rect 17078 17926 17130 17978
rect 17142 17926 17194 17978
rect 17206 17926 17258 17978
rect 13820 17824 13872 17876
rect 14556 17756 14608 17808
rect 7288 17688 7340 17740
rect 10600 17731 10652 17740
rect 10600 17697 10609 17731
rect 10609 17697 10643 17731
rect 10643 17697 10652 17731
rect 10600 17688 10652 17697
rect 13084 17688 13136 17740
rect 10876 17663 10928 17672
rect 10876 17629 10910 17663
rect 10910 17629 10928 17663
rect 10876 17620 10928 17629
rect 13360 17663 13412 17672
rect 13360 17629 13369 17663
rect 13369 17629 13403 17663
rect 13403 17629 13412 17663
rect 13360 17620 13412 17629
rect 12532 17552 12584 17604
rect 13544 17552 13596 17604
rect 2610 17382 2662 17434
rect 2674 17382 2726 17434
rect 2738 17382 2790 17434
rect 2802 17382 2854 17434
rect 2866 17382 2918 17434
rect 7610 17382 7662 17434
rect 7674 17382 7726 17434
rect 7738 17382 7790 17434
rect 7802 17382 7854 17434
rect 7866 17382 7918 17434
rect 12610 17382 12662 17434
rect 12674 17382 12726 17434
rect 12738 17382 12790 17434
rect 12802 17382 12854 17434
rect 12866 17382 12918 17434
rect 17610 17382 17662 17434
rect 17674 17382 17726 17434
rect 17738 17382 17790 17434
rect 17802 17382 17854 17434
rect 17866 17382 17918 17434
rect 5724 17280 5776 17332
rect 5908 17280 5960 17332
rect 1584 17212 1636 17264
rect 5908 17008 5960 17060
rect 10232 17008 10284 17060
rect 848 16940 900 16992
rect 1950 16838 2002 16890
rect 2014 16838 2066 16890
rect 2078 16838 2130 16890
rect 2142 16838 2194 16890
rect 2206 16838 2258 16890
rect 6950 16838 7002 16890
rect 7014 16838 7066 16890
rect 7078 16838 7130 16890
rect 7142 16838 7194 16890
rect 7206 16838 7258 16890
rect 11950 16838 12002 16890
rect 12014 16838 12066 16890
rect 12078 16838 12130 16890
rect 12142 16838 12194 16890
rect 12206 16838 12258 16890
rect 16950 16838 17002 16890
rect 17014 16838 17066 16890
rect 17078 16838 17130 16890
rect 17142 16838 17194 16890
rect 17206 16838 17258 16890
rect 5540 16600 5592 16652
rect 7288 16736 7340 16788
rect 17960 16779 18012 16788
rect 17960 16745 17969 16779
rect 17969 16745 18003 16779
rect 18003 16745 18012 16779
rect 17960 16736 18012 16745
rect 756 16464 808 16516
rect 13452 16532 13504 16584
rect 14740 16464 14792 16516
rect 664 16396 716 16448
rect 5908 16439 5960 16448
rect 5908 16405 5917 16439
rect 5917 16405 5951 16439
rect 5951 16405 5960 16439
rect 5908 16396 5960 16405
rect 8484 16439 8536 16448
rect 8484 16405 8493 16439
rect 8493 16405 8527 16439
rect 8527 16405 8536 16439
rect 8484 16396 8536 16405
rect 2610 16294 2662 16346
rect 2674 16294 2726 16346
rect 2738 16294 2790 16346
rect 2802 16294 2854 16346
rect 2866 16294 2918 16346
rect 7610 16294 7662 16346
rect 7674 16294 7726 16346
rect 7738 16294 7790 16346
rect 7802 16294 7854 16346
rect 7866 16294 7918 16346
rect 12610 16294 12662 16346
rect 12674 16294 12726 16346
rect 12738 16294 12790 16346
rect 12802 16294 12854 16346
rect 12866 16294 12918 16346
rect 17610 16294 17662 16346
rect 17674 16294 17726 16346
rect 17738 16294 17790 16346
rect 17802 16294 17854 16346
rect 17866 16294 17918 16346
rect 9036 16235 9088 16244
rect 9036 16201 9045 16235
rect 9045 16201 9079 16235
rect 9079 16201 9088 16235
rect 9036 16192 9088 16201
rect 9772 16235 9824 16244
rect 9772 16201 9781 16235
rect 9781 16201 9815 16235
rect 9815 16201 9824 16235
rect 9772 16192 9824 16201
rect 18236 16235 18288 16244
rect 18236 16201 18245 16235
rect 18245 16201 18279 16235
rect 18279 16201 18288 16235
rect 18236 16192 18288 16201
rect 3516 16124 3568 16176
rect 1768 16056 1820 16108
rect 10968 16056 11020 16108
rect 7288 15988 7340 16040
rect 8300 15988 8352 16040
rect 1950 15750 2002 15802
rect 2014 15750 2066 15802
rect 2078 15750 2130 15802
rect 2142 15750 2194 15802
rect 2206 15750 2258 15802
rect 6950 15750 7002 15802
rect 7014 15750 7066 15802
rect 7078 15750 7130 15802
rect 7142 15750 7194 15802
rect 7206 15750 7258 15802
rect 11950 15750 12002 15802
rect 12014 15750 12066 15802
rect 12078 15750 12130 15802
rect 12142 15750 12194 15802
rect 12206 15750 12258 15802
rect 16950 15750 17002 15802
rect 17014 15750 17066 15802
rect 17078 15750 17130 15802
rect 17142 15750 17194 15802
rect 17206 15750 17258 15802
rect 9772 15648 9824 15700
rect 11796 15648 11848 15700
rect 9496 15580 9548 15632
rect 12992 15555 13044 15564
rect 12992 15521 13001 15555
rect 13001 15521 13035 15555
rect 13035 15521 13044 15555
rect 12992 15512 13044 15521
rect 13084 15555 13136 15564
rect 13084 15521 13093 15555
rect 13093 15521 13127 15555
rect 13127 15521 13136 15555
rect 13084 15512 13136 15521
rect 13636 15512 13688 15564
rect 1032 15444 1084 15496
rect 16856 15487 16908 15496
rect 16856 15453 16865 15487
rect 16865 15453 16899 15487
rect 16899 15453 16908 15487
rect 16856 15444 16908 15453
rect 16580 15376 16632 15428
rect 11428 15308 11480 15360
rect 19800 15376 19852 15428
rect 18236 15351 18288 15360
rect 18236 15317 18245 15351
rect 18245 15317 18279 15351
rect 18279 15317 18288 15351
rect 18236 15308 18288 15317
rect 18512 15308 18564 15360
rect 2610 15206 2662 15258
rect 2674 15206 2726 15258
rect 2738 15206 2790 15258
rect 2802 15206 2854 15258
rect 2866 15206 2918 15258
rect 7610 15206 7662 15258
rect 7674 15206 7726 15258
rect 7738 15206 7790 15258
rect 7802 15206 7854 15258
rect 7866 15206 7918 15258
rect 12610 15206 12662 15258
rect 12674 15206 12726 15258
rect 12738 15206 12790 15258
rect 12802 15206 12854 15258
rect 12866 15206 12918 15258
rect 17610 15206 17662 15258
rect 17674 15206 17726 15258
rect 17738 15206 17790 15258
rect 17802 15206 17854 15258
rect 17866 15206 17918 15258
rect 940 15104 992 15156
rect 14924 15104 14976 15156
rect 2320 15079 2372 15088
rect 2320 15045 2329 15079
rect 2329 15045 2363 15079
rect 2363 15045 2372 15079
rect 2320 15036 2372 15045
rect 15844 15036 15896 15088
rect 15016 14968 15068 15020
rect 17684 14875 17736 14884
rect 17684 14841 17693 14875
rect 17693 14841 17727 14875
rect 17727 14841 17736 14875
rect 17684 14832 17736 14841
rect 1950 14662 2002 14714
rect 2014 14662 2066 14714
rect 2078 14662 2130 14714
rect 2142 14662 2194 14714
rect 2206 14662 2258 14714
rect 6950 14662 7002 14714
rect 7014 14662 7066 14714
rect 7078 14662 7130 14714
rect 7142 14662 7194 14714
rect 7206 14662 7258 14714
rect 11950 14662 12002 14714
rect 12014 14662 12066 14714
rect 12078 14662 12130 14714
rect 12142 14662 12194 14714
rect 12206 14662 12258 14714
rect 16950 14662 17002 14714
rect 17014 14662 17066 14714
rect 17078 14662 17130 14714
rect 17142 14662 17194 14714
rect 17206 14662 17258 14714
rect 7380 14560 7432 14612
rect 13176 14560 13228 14612
rect 1124 14492 1176 14544
rect 7840 14399 7892 14408
rect 7840 14365 7849 14399
rect 7849 14365 7883 14399
rect 7883 14365 7892 14399
rect 7840 14356 7892 14365
rect 8392 14399 8444 14408
rect 8392 14365 8401 14399
rect 8401 14365 8435 14399
rect 8435 14365 8444 14399
rect 8392 14356 8444 14365
rect 15476 14399 15528 14408
rect 15476 14365 15485 14399
rect 15485 14365 15519 14399
rect 15519 14365 15528 14399
rect 15476 14356 15528 14365
rect 19524 14356 19576 14408
rect 11336 14288 11388 14340
rect 18236 14263 18288 14272
rect 18236 14229 18245 14263
rect 18245 14229 18279 14263
rect 18279 14229 18288 14263
rect 18236 14220 18288 14229
rect 2610 14118 2662 14170
rect 2674 14118 2726 14170
rect 2738 14118 2790 14170
rect 2802 14118 2854 14170
rect 2866 14118 2918 14170
rect 7610 14118 7662 14170
rect 7674 14118 7726 14170
rect 7738 14118 7790 14170
rect 7802 14118 7854 14170
rect 7866 14118 7918 14170
rect 12610 14118 12662 14170
rect 12674 14118 12726 14170
rect 12738 14118 12790 14170
rect 12802 14118 12854 14170
rect 12866 14118 12918 14170
rect 17610 14118 17662 14170
rect 17674 14118 17726 14170
rect 17738 14118 17790 14170
rect 17802 14118 17854 14170
rect 17866 14118 17918 14170
rect 11060 14016 11112 14068
rect 16120 14016 16172 14068
rect 11152 13948 11204 14000
rect 11244 13880 11296 13932
rect 10600 13744 10652 13796
rect 10784 13744 10836 13796
rect 15476 13744 15528 13796
rect 16856 13744 16908 13796
rect 1950 13574 2002 13626
rect 2014 13574 2066 13626
rect 2078 13574 2130 13626
rect 2142 13574 2194 13626
rect 2206 13574 2258 13626
rect 6950 13574 7002 13626
rect 7014 13574 7066 13626
rect 7078 13574 7130 13626
rect 7142 13574 7194 13626
rect 7206 13574 7258 13626
rect 11950 13574 12002 13626
rect 12014 13574 12066 13626
rect 12078 13574 12130 13626
rect 12142 13574 12194 13626
rect 12206 13574 12258 13626
rect 16950 13574 17002 13626
rect 17014 13574 17066 13626
rect 17078 13574 17130 13626
rect 17142 13574 17194 13626
rect 17206 13574 17258 13626
rect 8576 13472 8628 13524
rect 16396 13311 16448 13320
rect 16396 13277 16405 13311
rect 16405 13277 16439 13311
rect 16439 13277 16448 13311
rect 16396 13268 16448 13277
rect 7288 13200 7340 13252
rect 16580 13175 16632 13184
rect 16580 13141 16589 13175
rect 16589 13141 16623 13175
rect 16623 13141 16632 13175
rect 16580 13132 16632 13141
rect 2610 13030 2662 13082
rect 2674 13030 2726 13082
rect 2738 13030 2790 13082
rect 2802 13030 2854 13082
rect 2866 13030 2918 13082
rect 7610 13030 7662 13082
rect 7674 13030 7726 13082
rect 7738 13030 7790 13082
rect 7802 13030 7854 13082
rect 7866 13030 7918 13082
rect 12610 13030 12662 13082
rect 12674 13030 12726 13082
rect 12738 13030 12790 13082
rect 12802 13030 12854 13082
rect 12866 13030 12918 13082
rect 17610 13030 17662 13082
rect 17674 13030 17726 13082
rect 17738 13030 17790 13082
rect 17802 13030 17854 13082
rect 17866 13030 17918 13082
rect 11060 12928 11112 12980
rect 11704 12928 11756 12980
rect 18052 12928 18104 12980
rect 5264 12903 5316 12912
rect 5264 12869 5273 12903
rect 5273 12869 5307 12903
rect 5307 12869 5316 12903
rect 5264 12860 5316 12869
rect 17316 12860 17368 12912
rect 16856 12835 16908 12844
rect 16856 12801 16865 12835
rect 16865 12801 16899 12835
rect 16899 12801 16908 12835
rect 16856 12792 16908 12801
rect 3884 12588 3936 12640
rect 1950 12486 2002 12538
rect 2014 12486 2066 12538
rect 2078 12486 2130 12538
rect 2142 12486 2194 12538
rect 2206 12486 2258 12538
rect 6950 12486 7002 12538
rect 7014 12486 7066 12538
rect 7078 12486 7130 12538
rect 7142 12486 7194 12538
rect 7206 12486 7258 12538
rect 11950 12486 12002 12538
rect 12014 12486 12066 12538
rect 12078 12486 12130 12538
rect 12142 12486 12194 12538
rect 12206 12486 12258 12538
rect 16950 12486 17002 12538
rect 17014 12486 17066 12538
rect 17078 12486 17130 12538
rect 17142 12486 17194 12538
rect 17206 12486 17258 12538
rect 7380 12427 7432 12436
rect 7380 12393 7389 12427
rect 7389 12393 7423 12427
rect 7423 12393 7432 12427
rect 7380 12384 7432 12393
rect 12164 12359 12216 12368
rect 12164 12325 12173 12359
rect 12173 12325 12207 12359
rect 12207 12325 12216 12359
rect 12164 12316 12216 12325
rect 18236 12359 18288 12368
rect 18236 12325 18245 12359
rect 18245 12325 18279 12359
rect 18279 12325 18288 12359
rect 18236 12316 18288 12325
rect 3884 12180 3936 12232
rect 8944 12180 8996 12232
rect 10692 12223 10744 12232
rect 10692 12189 10701 12223
rect 10701 12189 10735 12223
rect 10735 12189 10744 12223
rect 10692 12180 10744 12189
rect 10784 12223 10836 12232
rect 10784 12189 10793 12223
rect 10793 12189 10827 12223
rect 10827 12189 10836 12223
rect 10784 12180 10836 12189
rect 11060 12223 11112 12232
rect 11060 12189 11094 12223
rect 11094 12189 11112 12223
rect 11060 12180 11112 12189
rect 18052 12223 18104 12232
rect 18052 12189 18061 12223
rect 18061 12189 18095 12223
rect 18095 12189 18104 12223
rect 18052 12180 18104 12189
rect 1492 12044 1544 12096
rect 2610 11942 2662 11994
rect 2674 11942 2726 11994
rect 2738 11942 2790 11994
rect 2802 11942 2854 11994
rect 2866 11942 2918 11994
rect 7610 11942 7662 11994
rect 7674 11942 7726 11994
rect 7738 11942 7790 11994
rect 7802 11942 7854 11994
rect 7866 11942 7918 11994
rect 12610 11942 12662 11994
rect 12674 11942 12726 11994
rect 12738 11942 12790 11994
rect 12802 11942 12854 11994
rect 12866 11942 12918 11994
rect 17610 11942 17662 11994
rect 17674 11942 17726 11994
rect 17738 11942 17790 11994
rect 17802 11942 17854 11994
rect 17866 11942 17918 11994
rect 4804 11772 4856 11824
rect 6276 11772 6328 11824
rect 3148 11500 3200 11552
rect 5724 11500 5776 11552
rect 1950 11398 2002 11450
rect 2014 11398 2066 11450
rect 2078 11398 2130 11450
rect 2142 11398 2194 11450
rect 2206 11398 2258 11450
rect 6950 11398 7002 11450
rect 7014 11398 7066 11450
rect 7078 11398 7130 11450
rect 7142 11398 7194 11450
rect 7206 11398 7258 11450
rect 11950 11398 12002 11450
rect 12014 11398 12066 11450
rect 12078 11398 12130 11450
rect 12142 11398 12194 11450
rect 12206 11398 12258 11450
rect 16950 11398 17002 11450
rect 17014 11398 17066 11450
rect 17078 11398 17130 11450
rect 17142 11398 17194 11450
rect 17206 11398 17258 11450
rect 6644 11092 6696 11144
rect 15200 11160 15252 11212
rect 15292 11203 15344 11212
rect 15292 11169 15301 11203
rect 15301 11169 15335 11203
rect 15335 11169 15344 11203
rect 15292 11160 15344 11169
rect 14832 11135 14884 11144
rect 14832 11101 14841 11135
rect 14841 11101 14875 11135
rect 14875 11101 14884 11135
rect 14832 11092 14884 11101
rect 16028 11024 16080 11076
rect 2610 10854 2662 10906
rect 2674 10854 2726 10906
rect 2738 10854 2790 10906
rect 2802 10854 2854 10906
rect 2866 10854 2918 10906
rect 7610 10854 7662 10906
rect 7674 10854 7726 10906
rect 7738 10854 7790 10906
rect 7802 10854 7854 10906
rect 7866 10854 7918 10906
rect 12610 10854 12662 10906
rect 12674 10854 12726 10906
rect 12738 10854 12790 10906
rect 12802 10854 12854 10906
rect 12866 10854 12918 10906
rect 17610 10854 17662 10906
rect 17674 10854 17726 10906
rect 17738 10854 17790 10906
rect 17802 10854 17854 10906
rect 17866 10854 17918 10906
rect 1860 10795 1912 10804
rect 1860 10761 1869 10795
rect 1869 10761 1903 10795
rect 1903 10761 1912 10795
rect 1860 10752 1912 10761
rect 3148 10795 3200 10804
rect 3148 10761 3157 10795
rect 3157 10761 3191 10795
rect 3191 10761 3200 10795
rect 3148 10752 3200 10761
rect 2596 10727 2648 10736
rect 2596 10693 2605 10727
rect 2605 10693 2639 10727
rect 2639 10693 2648 10727
rect 2596 10684 2648 10693
rect 15200 10616 15252 10668
rect 4896 10412 4948 10464
rect 14372 10412 14424 10464
rect 18236 10455 18288 10464
rect 18236 10421 18245 10455
rect 18245 10421 18279 10455
rect 18279 10421 18288 10455
rect 18236 10412 18288 10421
rect 1950 10310 2002 10362
rect 2014 10310 2066 10362
rect 2078 10310 2130 10362
rect 2142 10310 2194 10362
rect 2206 10310 2258 10362
rect 6950 10310 7002 10362
rect 7014 10310 7066 10362
rect 7078 10310 7130 10362
rect 7142 10310 7194 10362
rect 7206 10310 7258 10362
rect 11950 10310 12002 10362
rect 12014 10310 12066 10362
rect 12078 10310 12130 10362
rect 12142 10310 12194 10362
rect 12206 10310 12258 10362
rect 16950 10310 17002 10362
rect 17014 10310 17066 10362
rect 17078 10310 17130 10362
rect 17142 10310 17194 10362
rect 17206 10310 17258 10362
rect 1860 10251 1912 10260
rect 1860 10217 1869 10251
rect 1869 10217 1903 10251
rect 1903 10217 1912 10251
rect 1860 10208 1912 10217
rect 6920 10208 6972 10260
rect 8208 10208 8260 10260
rect 10508 10140 10560 10192
rect 6920 10047 6972 10056
rect 6920 10013 6929 10047
rect 6929 10013 6963 10047
rect 6963 10013 6972 10047
rect 6920 10004 6972 10013
rect 7380 10072 7432 10124
rect 7932 10115 7984 10124
rect 7932 10081 7941 10115
rect 7941 10081 7975 10115
rect 7975 10081 7984 10115
rect 7932 10072 7984 10081
rect 7288 10004 7340 10056
rect 15936 9936 15988 9988
rect 7932 9868 7984 9920
rect 2610 9766 2662 9818
rect 2674 9766 2726 9818
rect 2738 9766 2790 9818
rect 2802 9766 2854 9818
rect 2866 9766 2918 9818
rect 7610 9766 7662 9818
rect 7674 9766 7726 9818
rect 7738 9766 7790 9818
rect 7802 9766 7854 9818
rect 7866 9766 7918 9818
rect 12610 9766 12662 9818
rect 12674 9766 12726 9818
rect 12738 9766 12790 9818
rect 12802 9766 12854 9818
rect 12866 9766 12918 9818
rect 17610 9766 17662 9818
rect 17674 9766 17726 9818
rect 17738 9766 17790 9818
rect 17802 9766 17854 9818
rect 17866 9766 17918 9818
rect 2320 9596 2372 9648
rect 3884 9596 3936 9648
rect 4252 9571 4304 9580
rect 4252 9537 4261 9571
rect 4261 9537 4295 9571
rect 4295 9537 4304 9571
rect 4252 9528 4304 9537
rect 5540 9528 5592 9580
rect 6644 9571 6696 9580
rect 6644 9537 6653 9571
rect 6653 9537 6687 9571
rect 6687 9537 6696 9571
rect 6644 9528 6696 9537
rect 13084 9596 13136 9648
rect 15384 9528 15436 9580
rect 7012 9435 7064 9444
rect 7012 9401 7021 9435
rect 7021 9401 7055 9435
rect 7055 9401 7064 9435
rect 7012 9392 7064 9401
rect 18144 9392 18196 9444
rect 3976 9324 4028 9376
rect 7932 9324 7984 9376
rect 9588 9324 9640 9376
rect 1950 9222 2002 9274
rect 2014 9222 2066 9274
rect 2078 9222 2130 9274
rect 2142 9222 2194 9274
rect 2206 9222 2258 9274
rect 6950 9222 7002 9274
rect 7014 9222 7066 9274
rect 7078 9222 7130 9274
rect 7142 9222 7194 9274
rect 7206 9222 7258 9274
rect 11950 9222 12002 9274
rect 12014 9222 12066 9274
rect 12078 9222 12130 9274
rect 12142 9222 12194 9274
rect 12206 9222 12258 9274
rect 16950 9222 17002 9274
rect 17014 9222 17066 9274
rect 17078 9222 17130 9274
rect 17142 9222 17194 9274
rect 17206 9222 17258 9274
rect 5540 9120 5592 9172
rect 8116 9120 8168 9172
rect 17408 9120 17460 9172
rect 7472 8984 7524 9036
rect 7932 8984 7984 9036
rect 8116 8916 8168 8968
rect 8208 8959 8260 8968
rect 8208 8925 8217 8959
rect 8217 8925 8251 8959
rect 8251 8925 8260 8959
rect 8208 8916 8260 8925
rect 8024 8848 8076 8900
rect 5172 8780 5224 8832
rect 18236 8823 18288 8832
rect 18236 8789 18245 8823
rect 18245 8789 18279 8823
rect 18279 8789 18288 8823
rect 18236 8780 18288 8789
rect 2610 8678 2662 8730
rect 2674 8678 2726 8730
rect 2738 8678 2790 8730
rect 2802 8678 2854 8730
rect 2866 8678 2918 8730
rect 7610 8678 7662 8730
rect 7674 8678 7726 8730
rect 7738 8678 7790 8730
rect 7802 8678 7854 8730
rect 7866 8678 7918 8730
rect 12610 8678 12662 8730
rect 12674 8678 12726 8730
rect 12738 8678 12790 8730
rect 12802 8678 12854 8730
rect 12866 8678 12918 8730
rect 17610 8678 17662 8730
rect 17674 8678 17726 8730
rect 17738 8678 17790 8730
rect 17802 8678 17854 8730
rect 17866 8678 17918 8730
rect 3700 8619 3752 8628
rect 3700 8585 3709 8619
rect 3709 8585 3743 8619
rect 3743 8585 3752 8619
rect 3700 8576 3752 8585
rect 8116 8576 8168 8628
rect 14648 8576 14700 8628
rect 4252 8440 4304 8492
rect 10784 8508 10836 8560
rect 10968 8508 11020 8560
rect 14096 8508 14148 8560
rect 14556 8508 14608 8560
rect 19064 8576 19116 8628
rect 11520 8440 11572 8492
rect 18052 8508 18104 8560
rect 2320 8415 2372 8424
rect 2320 8381 2329 8415
rect 2329 8381 2363 8415
rect 2363 8381 2372 8415
rect 2320 8372 2372 8381
rect 2504 8372 2556 8424
rect 14372 8415 14424 8424
rect 14372 8381 14381 8415
rect 14381 8381 14415 8415
rect 14415 8381 14424 8415
rect 14372 8372 14424 8381
rect 11612 8304 11664 8356
rect 12440 8236 12492 8288
rect 13268 8236 13320 8288
rect 1950 8134 2002 8186
rect 2014 8134 2066 8186
rect 2078 8134 2130 8186
rect 2142 8134 2194 8186
rect 2206 8134 2258 8186
rect 6950 8134 7002 8186
rect 7014 8134 7066 8186
rect 7078 8134 7130 8186
rect 7142 8134 7194 8186
rect 7206 8134 7258 8186
rect 11950 8134 12002 8186
rect 12014 8134 12066 8186
rect 12078 8134 12130 8186
rect 12142 8134 12194 8186
rect 12206 8134 12258 8186
rect 16950 8134 17002 8186
rect 17014 8134 17066 8186
rect 17078 8134 17130 8186
rect 17142 8134 17194 8186
rect 17206 8134 17258 8186
rect 1308 8032 1360 8084
rect 11520 8075 11572 8084
rect 11520 8041 11529 8075
rect 11529 8041 11563 8075
rect 11563 8041 11572 8075
rect 11520 8032 11572 8041
rect 8760 7896 8812 7948
rect 12440 7896 12492 7948
rect 2964 7828 3016 7880
rect 10048 7828 10100 7880
rect 10876 7828 10928 7880
rect 12256 7871 12308 7880
rect 12256 7837 12265 7871
rect 12265 7837 12299 7871
rect 12299 7837 12308 7871
rect 12256 7828 12308 7837
rect 9128 7735 9180 7744
rect 9128 7701 9137 7735
rect 9137 7701 9171 7735
rect 9171 7701 9180 7735
rect 9128 7692 9180 7701
rect 2610 7590 2662 7642
rect 2674 7590 2726 7642
rect 2738 7590 2790 7642
rect 2802 7590 2854 7642
rect 2866 7590 2918 7642
rect 7610 7590 7662 7642
rect 7674 7590 7726 7642
rect 7738 7590 7790 7642
rect 7802 7590 7854 7642
rect 7866 7590 7918 7642
rect 12610 7590 12662 7642
rect 12674 7590 12726 7642
rect 12738 7590 12790 7642
rect 12802 7590 12854 7642
rect 12866 7590 12918 7642
rect 17610 7590 17662 7642
rect 17674 7590 17726 7642
rect 17738 7590 17790 7642
rect 17802 7590 17854 7642
rect 17866 7590 17918 7642
rect 12256 7488 12308 7540
rect 14188 7463 14240 7472
rect 14188 7429 14197 7463
rect 14197 7429 14231 7463
rect 14231 7429 14240 7463
rect 14188 7420 14240 7429
rect 13820 7259 13872 7268
rect 13820 7225 13829 7259
rect 13829 7225 13863 7259
rect 13863 7225 13872 7259
rect 13820 7216 13872 7225
rect 1950 7046 2002 7098
rect 2014 7046 2066 7098
rect 2078 7046 2130 7098
rect 2142 7046 2194 7098
rect 2206 7046 2258 7098
rect 6950 7046 7002 7098
rect 7014 7046 7066 7098
rect 7078 7046 7130 7098
rect 7142 7046 7194 7098
rect 7206 7046 7258 7098
rect 11950 7046 12002 7098
rect 12014 7046 12066 7098
rect 12078 7046 12130 7098
rect 12142 7046 12194 7098
rect 12206 7046 12258 7098
rect 16950 7046 17002 7098
rect 17014 7046 17066 7098
rect 17078 7046 17130 7098
rect 17142 7046 17194 7098
rect 17206 7046 17258 7098
rect 6920 6919 6972 6928
rect 6920 6885 6929 6919
rect 6929 6885 6963 6919
rect 6963 6885 6972 6919
rect 6920 6876 6972 6885
rect 7380 6851 7432 6860
rect 7380 6817 7389 6851
rect 7389 6817 7423 6851
rect 7423 6817 7432 6851
rect 7380 6808 7432 6817
rect 7472 6851 7524 6860
rect 7472 6817 7481 6851
rect 7481 6817 7515 6851
rect 7515 6817 7524 6851
rect 7472 6808 7524 6817
rect 10324 6808 10376 6860
rect 6276 6672 6328 6724
rect 9496 6715 9548 6724
rect 9496 6681 9505 6715
rect 9505 6681 9539 6715
rect 9539 6681 9548 6715
rect 9496 6672 9548 6681
rect 9680 6715 9732 6724
rect 9680 6681 9689 6715
rect 9689 6681 9723 6715
rect 9723 6681 9732 6715
rect 9680 6672 9732 6681
rect 13544 6672 13596 6724
rect 12716 6604 12768 6656
rect 18236 6647 18288 6656
rect 18236 6613 18245 6647
rect 18245 6613 18279 6647
rect 18279 6613 18288 6647
rect 18236 6604 18288 6613
rect 2610 6502 2662 6554
rect 2674 6502 2726 6554
rect 2738 6502 2790 6554
rect 2802 6502 2854 6554
rect 2866 6502 2918 6554
rect 7610 6502 7662 6554
rect 7674 6502 7726 6554
rect 7738 6502 7790 6554
rect 7802 6502 7854 6554
rect 7866 6502 7918 6554
rect 12610 6502 12662 6554
rect 12674 6502 12726 6554
rect 12738 6502 12790 6554
rect 12802 6502 12854 6554
rect 12866 6502 12918 6554
rect 17610 6502 17662 6554
rect 17674 6502 17726 6554
rect 17738 6502 17790 6554
rect 17802 6502 17854 6554
rect 17866 6502 17918 6554
rect 3608 6400 3660 6452
rect 9496 6400 9548 6452
rect 5816 6332 5868 6384
rect 8208 6332 8260 6384
rect 1950 5958 2002 6010
rect 2014 5958 2066 6010
rect 2078 5958 2130 6010
rect 2142 5958 2194 6010
rect 2206 5958 2258 6010
rect 6950 5958 7002 6010
rect 7014 5958 7066 6010
rect 7078 5958 7130 6010
rect 7142 5958 7194 6010
rect 7206 5958 7258 6010
rect 11950 5958 12002 6010
rect 12014 5958 12066 6010
rect 12078 5958 12130 6010
rect 12142 5958 12194 6010
rect 12206 5958 12258 6010
rect 16950 5958 17002 6010
rect 17014 5958 17066 6010
rect 17078 5958 17130 6010
rect 17142 5958 17194 6010
rect 17206 5958 17258 6010
rect 2320 5652 2372 5704
rect 5080 5695 5132 5704
rect 5080 5661 5089 5695
rect 5089 5661 5123 5695
rect 5123 5661 5132 5695
rect 5080 5652 5132 5661
rect 6184 5652 6236 5704
rect 11428 5516 11480 5568
rect 2610 5414 2662 5466
rect 2674 5414 2726 5466
rect 2738 5414 2790 5466
rect 2802 5414 2854 5466
rect 2866 5414 2918 5466
rect 7610 5414 7662 5466
rect 7674 5414 7726 5466
rect 7738 5414 7790 5466
rect 7802 5414 7854 5466
rect 7866 5414 7918 5466
rect 12610 5414 12662 5466
rect 12674 5414 12726 5466
rect 12738 5414 12790 5466
rect 12802 5414 12854 5466
rect 12866 5414 12918 5466
rect 17610 5414 17662 5466
rect 17674 5414 17726 5466
rect 17738 5414 17790 5466
rect 17802 5414 17854 5466
rect 17866 5414 17918 5466
rect 1676 5312 1728 5364
rect 13360 5287 13412 5296
rect 13360 5253 13369 5287
rect 13369 5253 13403 5287
rect 13403 5253 13412 5287
rect 13360 5244 13412 5253
rect 9128 5176 9180 5228
rect 11060 5176 11112 5228
rect 11704 5219 11756 5228
rect 11704 5185 11713 5219
rect 11713 5185 11747 5219
rect 11747 5185 11756 5219
rect 11704 5176 11756 5185
rect 16212 5219 16264 5228
rect 16212 5185 16221 5219
rect 16221 5185 16255 5219
rect 16255 5185 16264 5219
rect 16212 5176 16264 5185
rect 6552 5040 6604 5092
rect 17500 5176 17552 5228
rect 8116 4972 8168 5024
rect 18236 5015 18288 5024
rect 18236 4981 18245 5015
rect 18245 4981 18279 5015
rect 18279 4981 18288 5015
rect 18236 4972 18288 4981
rect 1950 4870 2002 4922
rect 2014 4870 2066 4922
rect 2078 4870 2130 4922
rect 2142 4870 2194 4922
rect 2206 4870 2258 4922
rect 6950 4870 7002 4922
rect 7014 4870 7066 4922
rect 7078 4870 7130 4922
rect 7142 4870 7194 4922
rect 7206 4870 7258 4922
rect 11950 4870 12002 4922
rect 12014 4870 12066 4922
rect 12078 4870 12130 4922
rect 12142 4870 12194 4922
rect 12206 4870 12258 4922
rect 16950 4870 17002 4922
rect 17014 4870 17066 4922
rect 17078 4870 17130 4922
rect 17142 4870 17194 4922
rect 17206 4870 17258 4922
rect 7288 4632 7340 4684
rect 14464 4564 14516 4616
rect 2610 4326 2662 4378
rect 2674 4326 2726 4378
rect 2738 4326 2790 4378
rect 2802 4326 2854 4378
rect 2866 4326 2918 4378
rect 7610 4326 7662 4378
rect 7674 4326 7726 4378
rect 7738 4326 7790 4378
rect 7802 4326 7854 4378
rect 7866 4326 7918 4378
rect 12610 4326 12662 4378
rect 12674 4326 12726 4378
rect 12738 4326 12790 4378
rect 12802 4326 12854 4378
rect 12866 4326 12918 4378
rect 17610 4326 17662 4378
rect 17674 4326 17726 4378
rect 17738 4326 17790 4378
rect 17802 4326 17854 4378
rect 17866 4326 17918 4378
rect 5080 4088 5132 4140
rect 1216 4020 1268 4072
rect 16672 4088 16724 4140
rect 8208 4020 8260 4072
rect 8300 3952 8352 4004
rect 1950 3782 2002 3834
rect 2014 3782 2066 3834
rect 2078 3782 2130 3834
rect 2142 3782 2194 3834
rect 2206 3782 2258 3834
rect 6950 3782 7002 3834
rect 7014 3782 7066 3834
rect 7078 3782 7130 3834
rect 7142 3782 7194 3834
rect 7206 3782 7258 3834
rect 11950 3782 12002 3834
rect 12014 3782 12066 3834
rect 12078 3782 12130 3834
rect 12142 3782 12194 3834
rect 12206 3782 12258 3834
rect 16950 3782 17002 3834
rect 17014 3782 17066 3834
rect 17078 3782 17130 3834
rect 17142 3782 17194 3834
rect 17206 3782 17258 3834
rect 10968 3680 11020 3732
rect 11704 3544 11756 3596
rect 8116 3476 8168 3528
rect 2610 3238 2662 3290
rect 2674 3238 2726 3290
rect 2738 3238 2790 3290
rect 2802 3238 2854 3290
rect 2866 3238 2918 3290
rect 7610 3238 7662 3290
rect 7674 3238 7726 3290
rect 7738 3238 7790 3290
rect 7802 3238 7854 3290
rect 7866 3238 7918 3290
rect 12610 3238 12662 3290
rect 12674 3238 12726 3290
rect 12738 3238 12790 3290
rect 12802 3238 12854 3290
rect 12866 3238 12918 3290
rect 17610 3238 17662 3290
rect 17674 3238 17726 3290
rect 17738 3238 17790 3290
rect 17802 3238 17854 3290
rect 17866 3238 17918 3290
rect 9312 3136 9364 3188
rect 5632 3068 5684 3120
rect 19708 3000 19760 3052
rect 2320 2932 2372 2984
rect 18236 2839 18288 2848
rect 18236 2805 18245 2839
rect 18245 2805 18279 2839
rect 18279 2805 18288 2839
rect 18236 2796 18288 2805
rect 1950 2694 2002 2746
rect 2014 2694 2066 2746
rect 2078 2694 2130 2746
rect 2142 2694 2194 2746
rect 2206 2694 2258 2746
rect 6950 2694 7002 2746
rect 7014 2694 7066 2746
rect 7078 2694 7130 2746
rect 7142 2694 7194 2746
rect 7206 2694 7258 2746
rect 11950 2694 12002 2746
rect 12014 2694 12066 2746
rect 12078 2694 12130 2746
rect 12142 2694 12194 2746
rect 12206 2694 12258 2746
rect 16950 2694 17002 2746
rect 17014 2694 17066 2746
rect 17078 2694 17130 2746
rect 17142 2694 17194 2746
rect 17206 2694 17258 2746
rect 6000 2388 6052 2440
rect 9864 2592 9916 2644
rect 14464 2635 14516 2644
rect 14464 2601 14473 2635
rect 14473 2601 14507 2635
rect 14507 2601 14516 2635
rect 14464 2592 14516 2601
rect 18052 2499 18104 2508
rect 18052 2465 18061 2499
rect 18061 2465 18095 2499
rect 18095 2465 18104 2499
rect 18052 2456 18104 2465
rect 8852 2388 8904 2440
rect 17868 2431 17920 2440
rect 17868 2397 17877 2431
rect 17877 2397 17911 2431
rect 17911 2397 17920 2431
rect 17868 2388 17920 2397
rect 13912 2320 13964 2372
rect 9956 2252 10008 2304
rect 2610 2150 2662 2202
rect 2674 2150 2726 2202
rect 2738 2150 2790 2202
rect 2802 2150 2854 2202
rect 2866 2150 2918 2202
rect 7610 2150 7662 2202
rect 7674 2150 7726 2202
rect 7738 2150 7790 2202
rect 7802 2150 7854 2202
rect 7866 2150 7918 2202
rect 12610 2150 12662 2202
rect 12674 2150 12726 2202
rect 12738 2150 12790 2202
rect 12802 2150 12854 2202
rect 12866 2150 12918 2202
rect 17610 2150 17662 2202
rect 17674 2150 17726 2202
rect 17738 2150 17790 2202
rect 17802 2150 17854 2202
rect 17866 2150 17918 2202
<< metal2 >>
rect 1950 77820 2258 77829
rect 1950 77818 1956 77820
rect 2012 77818 2036 77820
rect 2092 77818 2116 77820
rect 2172 77818 2196 77820
rect 2252 77818 2258 77820
rect 2012 77766 2014 77818
rect 2194 77766 2196 77818
rect 1950 77764 1956 77766
rect 2012 77764 2036 77766
rect 2092 77764 2116 77766
rect 2172 77764 2196 77766
rect 2252 77764 2258 77766
rect 1950 77755 2258 77764
rect 6950 77820 7258 77829
rect 6950 77818 6956 77820
rect 7012 77818 7036 77820
rect 7092 77818 7116 77820
rect 7172 77818 7196 77820
rect 7252 77818 7258 77820
rect 7012 77766 7014 77818
rect 7194 77766 7196 77818
rect 6950 77764 6956 77766
rect 7012 77764 7036 77766
rect 7092 77764 7116 77766
rect 7172 77764 7196 77766
rect 7252 77764 7258 77766
rect 6950 77755 7258 77764
rect 11950 77820 12258 77829
rect 11950 77818 11956 77820
rect 12012 77818 12036 77820
rect 12092 77818 12116 77820
rect 12172 77818 12196 77820
rect 12252 77818 12258 77820
rect 12012 77766 12014 77818
rect 12194 77766 12196 77818
rect 11950 77764 11956 77766
rect 12012 77764 12036 77766
rect 12092 77764 12116 77766
rect 12172 77764 12196 77766
rect 12252 77764 12258 77766
rect 11950 77755 12258 77764
rect 16950 77820 17258 77829
rect 16950 77818 16956 77820
rect 17012 77818 17036 77820
rect 17092 77818 17116 77820
rect 17172 77818 17196 77820
rect 17252 77818 17258 77820
rect 17012 77766 17014 77818
rect 17194 77766 17196 77818
rect 16950 77764 16956 77766
rect 17012 77764 17036 77766
rect 17092 77764 17116 77766
rect 17172 77764 17196 77766
rect 17252 77764 17258 77766
rect 16950 77755 17258 77764
rect 18328 77512 18380 77518
rect 18328 77454 18380 77460
rect 16856 77376 16908 77382
rect 16856 77318 16908 77324
rect 18236 77376 18288 77382
rect 18236 77318 18288 77324
rect 2610 77276 2918 77285
rect 2610 77274 2616 77276
rect 2672 77274 2696 77276
rect 2752 77274 2776 77276
rect 2832 77274 2856 77276
rect 2912 77274 2918 77276
rect 2672 77222 2674 77274
rect 2854 77222 2856 77274
rect 2610 77220 2616 77222
rect 2672 77220 2696 77222
rect 2752 77220 2776 77222
rect 2832 77220 2856 77222
rect 2912 77220 2918 77222
rect 2610 77211 2918 77220
rect 7610 77276 7918 77285
rect 7610 77274 7616 77276
rect 7672 77274 7696 77276
rect 7752 77274 7776 77276
rect 7832 77274 7856 77276
rect 7912 77274 7918 77276
rect 7672 77222 7674 77274
rect 7854 77222 7856 77274
rect 7610 77220 7616 77222
rect 7672 77220 7696 77222
rect 7752 77220 7776 77222
rect 7832 77220 7856 77222
rect 7912 77220 7918 77222
rect 7610 77211 7918 77220
rect 12610 77276 12918 77285
rect 12610 77274 12616 77276
rect 12672 77274 12696 77276
rect 12752 77274 12776 77276
rect 12832 77274 12856 77276
rect 12912 77274 12918 77276
rect 12672 77222 12674 77274
rect 12854 77222 12856 77274
rect 12610 77220 12616 77222
rect 12672 77220 12696 77222
rect 12752 77220 12776 77222
rect 12832 77220 12856 77222
rect 12912 77220 12918 77222
rect 12610 77211 12918 77220
rect 14648 76832 14700 76838
rect 14646 76800 14648 76809
rect 15936 76832 15988 76838
rect 14700 76800 14702 76809
rect 1950 76732 2258 76741
rect 1950 76730 1956 76732
rect 2012 76730 2036 76732
rect 2092 76730 2116 76732
rect 2172 76730 2196 76732
rect 2252 76730 2258 76732
rect 2012 76678 2014 76730
rect 2194 76678 2196 76730
rect 1950 76676 1956 76678
rect 2012 76676 2036 76678
rect 2092 76676 2116 76678
rect 2172 76676 2196 76678
rect 2252 76676 2258 76678
rect 1950 76667 2258 76676
rect 6950 76732 7258 76741
rect 6950 76730 6956 76732
rect 7012 76730 7036 76732
rect 7092 76730 7116 76732
rect 7172 76730 7196 76732
rect 7252 76730 7258 76732
rect 7012 76678 7014 76730
rect 7194 76678 7196 76730
rect 6950 76676 6956 76678
rect 7012 76676 7036 76678
rect 7092 76676 7116 76678
rect 7172 76676 7196 76678
rect 7252 76676 7258 76678
rect 6950 76667 7258 76676
rect 11950 76732 12258 76741
rect 14646 76735 14702 76744
rect 15934 76800 15936 76809
rect 16488 76832 16540 76838
rect 15988 76800 15990 76809
rect 16488 76774 16540 76780
rect 15934 76735 15990 76744
rect 11950 76730 11956 76732
rect 12012 76730 12036 76732
rect 12092 76730 12116 76732
rect 12172 76730 12196 76732
rect 12252 76730 12258 76732
rect 12012 76678 12014 76730
rect 12194 76678 12196 76730
rect 11950 76676 11956 76678
rect 12012 76676 12036 76678
rect 12092 76676 12116 76678
rect 12172 76676 12196 76678
rect 12252 76676 12258 76678
rect 11950 76667 12258 76676
rect 7932 76492 7984 76498
rect 7932 76434 7984 76440
rect 2964 76288 3016 76294
rect 2964 76230 3016 76236
rect 7104 76288 7156 76294
rect 7104 76230 7156 76236
rect 7944 76242 7972 76434
rect 8208 76424 8260 76430
rect 8208 76366 8260 76372
rect 8482 76392 8538 76401
rect 2610 76188 2918 76197
rect 2610 76186 2616 76188
rect 2672 76186 2696 76188
rect 2752 76186 2776 76188
rect 2832 76186 2856 76188
rect 2912 76186 2918 76188
rect 2672 76134 2674 76186
rect 2854 76134 2856 76186
rect 2610 76132 2616 76134
rect 2672 76132 2696 76134
rect 2752 76132 2776 76134
rect 2832 76132 2856 76134
rect 2912 76132 2918 76134
rect 2610 76123 2918 76132
rect 1950 75644 2258 75653
rect 1950 75642 1956 75644
rect 2012 75642 2036 75644
rect 2092 75642 2116 75644
rect 2172 75642 2196 75644
rect 2252 75642 2258 75644
rect 2012 75590 2014 75642
rect 2194 75590 2196 75642
rect 1950 75588 1956 75590
rect 2012 75588 2036 75590
rect 2092 75588 2116 75590
rect 2172 75588 2196 75590
rect 2252 75588 2258 75590
rect 1950 75579 2258 75588
rect 2610 75100 2918 75109
rect 2610 75098 2616 75100
rect 2672 75098 2696 75100
rect 2752 75098 2776 75100
rect 2832 75098 2856 75100
rect 2912 75098 2918 75100
rect 2672 75046 2674 75098
rect 2854 75046 2856 75098
rect 2610 75044 2616 75046
rect 2672 75044 2696 75046
rect 2752 75044 2776 75046
rect 2832 75044 2856 75046
rect 2912 75044 2918 75046
rect 2610 75035 2918 75044
rect 1950 74556 2258 74565
rect 1950 74554 1956 74556
rect 2012 74554 2036 74556
rect 2092 74554 2116 74556
rect 2172 74554 2196 74556
rect 2252 74554 2258 74556
rect 2012 74502 2014 74554
rect 2194 74502 2196 74554
rect 1950 74500 1956 74502
rect 2012 74500 2036 74502
rect 2092 74500 2116 74502
rect 2172 74500 2196 74502
rect 2252 74500 2258 74502
rect 1950 74491 2258 74500
rect 2610 74012 2918 74021
rect 2610 74010 2616 74012
rect 2672 74010 2696 74012
rect 2752 74010 2776 74012
rect 2832 74010 2856 74012
rect 2912 74010 2918 74012
rect 2672 73958 2674 74010
rect 2854 73958 2856 74010
rect 2610 73956 2616 73958
rect 2672 73956 2696 73958
rect 2752 73956 2776 73958
rect 2832 73956 2856 73958
rect 2912 73956 2918 73958
rect 2610 73947 2918 73956
rect 1950 73468 2258 73477
rect 1950 73466 1956 73468
rect 2012 73466 2036 73468
rect 2092 73466 2116 73468
rect 2172 73466 2196 73468
rect 2252 73466 2258 73468
rect 2012 73414 2014 73466
rect 2194 73414 2196 73466
rect 1950 73412 1956 73414
rect 2012 73412 2036 73414
rect 2092 73412 2116 73414
rect 2172 73412 2196 73414
rect 2252 73412 2258 73414
rect 1950 73403 2258 73412
rect 1308 73024 1360 73030
rect 1308 72966 1360 72972
rect 1124 70848 1176 70854
rect 1124 70790 1176 70796
rect 1032 60308 1084 60314
rect 1032 60250 1084 60256
rect 940 56228 992 56234
rect 940 56170 992 56176
rect 848 55684 900 55690
rect 848 55626 900 55632
rect 756 52964 808 52970
rect 756 52906 808 52912
rect 664 41608 716 41614
rect 664 41550 716 41556
rect 676 16454 704 41550
rect 768 16522 796 52906
rect 860 16998 888 55626
rect 848 16992 900 16998
rect 848 16934 900 16940
rect 756 16516 808 16522
rect 756 16458 808 16464
rect 664 16448 716 16454
rect 664 16390 716 16396
rect 952 15162 980 56170
rect 1044 15502 1072 60250
rect 1032 15496 1084 15502
rect 1032 15438 1084 15444
rect 940 15156 992 15162
rect 940 15098 992 15104
rect 1136 14550 1164 70790
rect 1216 67040 1268 67046
rect 1216 66982 1268 66988
rect 1124 14544 1176 14550
rect 1124 14486 1176 14492
rect 1228 4078 1256 66982
rect 1320 8090 1348 72966
rect 2610 72924 2918 72933
rect 2610 72922 2616 72924
rect 2672 72922 2696 72924
rect 2752 72922 2776 72924
rect 2832 72922 2856 72924
rect 2912 72922 2918 72924
rect 2672 72870 2674 72922
rect 2854 72870 2856 72922
rect 2610 72868 2616 72870
rect 2672 72868 2696 72870
rect 2752 72868 2776 72870
rect 2832 72868 2856 72870
rect 2912 72868 2918 72870
rect 2610 72859 2918 72868
rect 1950 72380 2258 72389
rect 1950 72378 1956 72380
rect 2012 72378 2036 72380
rect 2092 72378 2116 72380
rect 2172 72378 2196 72380
rect 2252 72378 2258 72380
rect 2012 72326 2014 72378
rect 2194 72326 2196 72378
rect 1950 72324 1956 72326
rect 2012 72324 2036 72326
rect 2092 72324 2116 72326
rect 2172 72324 2196 72326
rect 2252 72324 2258 72326
rect 1950 72315 2258 72324
rect 2610 71836 2918 71845
rect 2610 71834 2616 71836
rect 2672 71834 2696 71836
rect 2752 71834 2776 71836
rect 2832 71834 2856 71836
rect 2912 71834 2918 71836
rect 2672 71782 2674 71834
rect 2854 71782 2856 71834
rect 2610 71780 2616 71782
rect 2672 71780 2696 71782
rect 2752 71780 2776 71782
rect 2832 71780 2856 71782
rect 2912 71780 2918 71782
rect 2610 71771 2918 71780
rect 1950 71292 2258 71301
rect 1950 71290 1956 71292
rect 2012 71290 2036 71292
rect 2092 71290 2116 71292
rect 2172 71290 2196 71292
rect 2252 71290 2258 71292
rect 2012 71238 2014 71290
rect 2194 71238 2196 71290
rect 1950 71236 1956 71238
rect 2012 71236 2036 71238
rect 2092 71236 2116 71238
rect 2172 71236 2196 71238
rect 2252 71236 2258 71238
rect 1950 71227 2258 71236
rect 2610 70748 2918 70757
rect 2610 70746 2616 70748
rect 2672 70746 2696 70748
rect 2752 70746 2776 70748
rect 2832 70746 2856 70748
rect 2912 70746 2918 70748
rect 2672 70694 2674 70746
rect 2854 70694 2856 70746
rect 2610 70692 2616 70694
rect 2672 70692 2696 70694
rect 2752 70692 2776 70694
rect 2832 70692 2856 70694
rect 2912 70692 2918 70694
rect 2610 70683 2918 70692
rect 1950 70204 2258 70213
rect 1950 70202 1956 70204
rect 2012 70202 2036 70204
rect 2092 70202 2116 70204
rect 2172 70202 2196 70204
rect 2252 70202 2258 70204
rect 2012 70150 2014 70202
rect 2194 70150 2196 70202
rect 1950 70148 1956 70150
rect 2012 70148 2036 70150
rect 2092 70148 2116 70150
rect 2172 70148 2196 70150
rect 2252 70148 2258 70150
rect 1950 70139 2258 70148
rect 2044 70032 2096 70038
rect 2044 69974 2096 69980
rect 2056 69329 2084 69974
rect 2976 69902 3004 76230
rect 5540 76016 5592 76022
rect 5540 75958 5592 75964
rect 5448 75336 5500 75342
rect 5448 75278 5500 75284
rect 5080 75200 5132 75206
rect 5080 75142 5132 75148
rect 4620 74724 4672 74730
rect 4620 74666 4672 74672
rect 3332 71596 3384 71602
rect 3332 71538 3384 71544
rect 3344 70961 3372 71538
rect 3330 70952 3386 70961
rect 3330 70887 3386 70896
rect 2964 69896 3016 69902
rect 2964 69838 3016 69844
rect 3976 69896 4028 69902
rect 3976 69838 4028 69844
rect 3792 69828 3844 69834
rect 3792 69770 3844 69776
rect 2504 69760 2556 69766
rect 2504 69702 2556 69708
rect 2042 69320 2098 69329
rect 2042 69255 2098 69264
rect 1950 69116 2258 69125
rect 1950 69114 1956 69116
rect 2012 69114 2036 69116
rect 2092 69114 2116 69116
rect 2172 69114 2196 69116
rect 2252 69114 2258 69116
rect 2012 69062 2014 69114
rect 2194 69062 2196 69114
rect 1950 69060 1956 69062
rect 2012 69060 2036 69062
rect 2092 69060 2116 69062
rect 2172 69060 2196 69062
rect 2252 69060 2258 69062
rect 1950 69051 2258 69060
rect 1950 68028 2258 68037
rect 1950 68026 1956 68028
rect 2012 68026 2036 68028
rect 2092 68026 2116 68028
rect 2172 68026 2196 68028
rect 2252 68026 2258 68028
rect 2012 67974 2014 68026
rect 2194 67974 2196 68026
rect 1950 67972 1956 67974
rect 2012 67972 2036 67974
rect 2092 67972 2116 67974
rect 2172 67972 2196 67974
rect 2252 67972 2258 67974
rect 1950 67963 2258 67972
rect 1950 66940 2258 66949
rect 1950 66938 1956 66940
rect 2012 66938 2036 66940
rect 2092 66938 2116 66940
rect 2172 66938 2196 66940
rect 2252 66938 2258 66940
rect 2012 66886 2014 66938
rect 2194 66886 2196 66938
rect 1950 66884 1956 66886
rect 2012 66884 2036 66886
rect 2092 66884 2116 66886
rect 2172 66884 2196 66886
rect 2252 66884 2258 66886
rect 1950 66875 2258 66884
rect 1950 65852 2258 65861
rect 1950 65850 1956 65852
rect 2012 65850 2036 65852
rect 2092 65850 2116 65852
rect 2172 65850 2196 65852
rect 2252 65850 2258 65852
rect 2012 65798 2014 65850
rect 2194 65798 2196 65850
rect 1950 65796 1956 65798
rect 2012 65796 2036 65798
rect 2092 65796 2116 65798
rect 2172 65796 2196 65798
rect 2252 65796 2258 65798
rect 1950 65787 2258 65796
rect 1950 64764 2258 64773
rect 1950 64762 1956 64764
rect 2012 64762 2036 64764
rect 2092 64762 2116 64764
rect 2172 64762 2196 64764
rect 2252 64762 2258 64764
rect 2012 64710 2014 64762
rect 2194 64710 2196 64762
rect 1950 64708 1956 64710
rect 2012 64708 2036 64710
rect 2092 64708 2116 64710
rect 2172 64708 2196 64710
rect 2252 64708 2258 64710
rect 1950 64699 2258 64708
rect 1768 64320 1820 64326
rect 1768 64262 1820 64268
rect 1492 56908 1544 56914
rect 1492 56850 1544 56856
rect 1400 51400 1452 51406
rect 1400 51342 1452 51348
rect 1412 22098 1440 51342
rect 1504 42702 1532 56850
rect 1676 56364 1728 56370
rect 1676 56306 1728 56312
rect 1688 55729 1716 56306
rect 1674 55720 1730 55729
rect 1674 55655 1730 55664
rect 1780 55214 1808 64262
rect 1950 63676 2258 63685
rect 1950 63674 1956 63676
rect 2012 63674 2036 63676
rect 2092 63674 2116 63676
rect 2172 63674 2196 63676
rect 2252 63674 2258 63676
rect 2012 63622 2014 63674
rect 2194 63622 2196 63674
rect 1950 63620 1956 63622
rect 2012 63620 2036 63622
rect 2092 63620 2116 63622
rect 2172 63620 2196 63622
rect 2252 63620 2258 63622
rect 1950 63611 2258 63620
rect 1950 62588 2258 62597
rect 1950 62586 1956 62588
rect 2012 62586 2036 62588
rect 2092 62586 2116 62588
rect 2172 62586 2196 62588
rect 2252 62586 2258 62588
rect 2012 62534 2014 62586
rect 2194 62534 2196 62586
rect 1950 62532 1956 62534
rect 2012 62532 2036 62534
rect 2092 62532 2116 62534
rect 2172 62532 2196 62534
rect 2252 62532 2258 62534
rect 1950 62523 2258 62532
rect 1950 61500 2258 61509
rect 1950 61498 1956 61500
rect 2012 61498 2036 61500
rect 2092 61498 2116 61500
rect 2172 61498 2196 61500
rect 2252 61498 2258 61500
rect 2012 61446 2014 61498
rect 2194 61446 2196 61498
rect 1950 61444 1956 61446
rect 2012 61444 2036 61446
rect 2092 61444 2116 61446
rect 2172 61444 2196 61446
rect 2252 61444 2258 61446
rect 1950 61435 2258 61444
rect 1950 60412 2258 60421
rect 1950 60410 1956 60412
rect 2012 60410 2036 60412
rect 2092 60410 2116 60412
rect 2172 60410 2196 60412
rect 2252 60410 2258 60412
rect 2012 60358 2014 60410
rect 2194 60358 2196 60410
rect 1950 60356 1956 60358
rect 2012 60356 2036 60358
rect 2092 60356 2116 60358
rect 2172 60356 2196 60358
rect 2252 60356 2258 60358
rect 1950 60347 2258 60356
rect 1950 59324 2258 59333
rect 1950 59322 1956 59324
rect 2012 59322 2036 59324
rect 2092 59322 2116 59324
rect 2172 59322 2196 59324
rect 2252 59322 2258 59324
rect 2012 59270 2014 59322
rect 2194 59270 2196 59322
rect 1950 59268 1956 59270
rect 2012 59268 2036 59270
rect 2092 59268 2116 59270
rect 2172 59268 2196 59270
rect 2252 59268 2258 59270
rect 1950 59259 2258 59268
rect 1950 58236 2258 58245
rect 1950 58234 1956 58236
rect 2012 58234 2036 58236
rect 2092 58234 2116 58236
rect 2172 58234 2196 58236
rect 2252 58234 2258 58236
rect 2012 58182 2014 58234
rect 2194 58182 2196 58234
rect 1950 58180 1956 58182
rect 2012 58180 2036 58182
rect 2092 58180 2116 58182
rect 2172 58180 2196 58182
rect 2252 58180 2258 58182
rect 1950 58171 2258 58180
rect 2320 57792 2372 57798
rect 2320 57734 2372 57740
rect 1950 57148 2258 57157
rect 1950 57146 1956 57148
rect 2012 57146 2036 57148
rect 2092 57146 2116 57148
rect 2172 57146 2196 57148
rect 2252 57146 2258 57148
rect 2012 57094 2014 57146
rect 2194 57094 2196 57146
rect 1950 57092 1956 57094
rect 2012 57092 2036 57094
rect 2092 57092 2116 57094
rect 2172 57092 2196 57094
rect 2252 57092 2258 57094
rect 1950 57083 2258 57092
rect 2332 56914 2360 57734
rect 2320 56908 2372 56914
rect 2320 56850 2372 56856
rect 2412 56704 2464 56710
rect 2412 56646 2464 56652
rect 2320 56160 2372 56166
rect 2320 56102 2372 56108
rect 1950 56060 2258 56069
rect 1950 56058 1956 56060
rect 2012 56058 2036 56060
rect 2092 56058 2116 56060
rect 2172 56058 2196 56060
rect 2252 56058 2258 56060
rect 2012 56006 2014 56058
rect 2194 56006 2196 56058
rect 1950 56004 1956 56006
rect 2012 56004 2036 56006
rect 2092 56004 2116 56006
rect 2172 56004 2196 56006
rect 2252 56004 2258 56006
rect 1950 55995 2258 56004
rect 1688 55186 1808 55214
rect 1584 48340 1636 48346
rect 1584 48282 1636 48288
rect 1492 42696 1544 42702
rect 1492 42638 1544 42644
rect 1596 40746 1624 48282
rect 1688 42770 1716 55186
rect 1950 54972 2258 54981
rect 1950 54970 1956 54972
rect 2012 54970 2036 54972
rect 2092 54970 2116 54972
rect 2172 54970 2196 54972
rect 2252 54970 2258 54972
rect 2012 54918 2014 54970
rect 2194 54918 2196 54970
rect 1950 54916 1956 54918
rect 2012 54916 2036 54918
rect 2092 54916 2116 54918
rect 2172 54916 2196 54918
rect 2252 54916 2258 54918
rect 1950 54907 2258 54916
rect 1950 53884 2258 53893
rect 1950 53882 1956 53884
rect 2012 53882 2036 53884
rect 2092 53882 2116 53884
rect 2172 53882 2196 53884
rect 2252 53882 2258 53884
rect 2012 53830 2014 53882
rect 2194 53830 2196 53882
rect 1950 53828 1956 53830
rect 2012 53828 2036 53830
rect 2092 53828 2116 53830
rect 2172 53828 2196 53830
rect 2252 53828 2258 53830
rect 1950 53819 2258 53828
rect 1952 53440 2004 53446
rect 1952 53382 2004 53388
rect 1964 53174 1992 53382
rect 1952 53168 2004 53174
rect 1952 53110 2004 53116
rect 1768 52896 1820 52902
rect 1768 52838 1820 52844
rect 1676 42764 1728 42770
rect 1676 42706 1728 42712
rect 1676 42560 1728 42566
rect 1676 42502 1728 42508
rect 1504 40718 1624 40746
rect 1504 26874 1532 40718
rect 1582 40624 1638 40633
rect 1582 40559 1638 40568
rect 1596 26994 1624 40559
rect 1584 26988 1636 26994
rect 1584 26930 1636 26936
rect 1504 26846 1624 26874
rect 1492 26784 1544 26790
rect 1492 26726 1544 26732
rect 1504 25362 1532 26726
rect 1492 25356 1544 25362
rect 1492 25298 1544 25304
rect 1492 25220 1544 25226
rect 1492 25162 1544 25168
rect 1400 22092 1452 22098
rect 1400 22034 1452 22040
rect 1504 12102 1532 25162
rect 1596 17270 1624 26846
rect 1584 17264 1636 17270
rect 1584 17206 1636 17212
rect 1492 12096 1544 12102
rect 1492 12038 1544 12044
rect 1308 8084 1360 8090
rect 1308 8026 1360 8032
rect 1688 5370 1716 42502
rect 1780 40905 1808 52838
rect 1950 52796 2258 52805
rect 1950 52794 1956 52796
rect 2012 52794 2036 52796
rect 2092 52794 2116 52796
rect 2172 52794 2196 52796
rect 2252 52794 2258 52796
rect 2012 52742 2014 52794
rect 2194 52742 2196 52794
rect 1950 52740 1956 52742
rect 2012 52740 2036 52742
rect 2092 52740 2116 52742
rect 2172 52740 2196 52742
rect 2252 52740 2258 52742
rect 1950 52731 2258 52740
rect 1950 51708 2258 51717
rect 1950 51706 1956 51708
rect 2012 51706 2036 51708
rect 2092 51706 2116 51708
rect 2172 51706 2196 51708
rect 2252 51706 2258 51708
rect 2012 51654 2014 51706
rect 2194 51654 2196 51706
rect 1950 51652 1956 51654
rect 2012 51652 2036 51654
rect 2092 51652 2116 51654
rect 2172 51652 2196 51654
rect 2252 51652 2258 51654
rect 1950 51643 2258 51652
rect 2332 50726 2360 56102
rect 2320 50720 2372 50726
rect 2320 50662 2372 50668
rect 1950 50620 2258 50629
rect 1950 50618 1956 50620
rect 2012 50618 2036 50620
rect 2092 50618 2116 50620
rect 2172 50618 2196 50620
rect 2252 50618 2258 50620
rect 2012 50566 2014 50618
rect 2194 50566 2196 50618
rect 1950 50564 1956 50566
rect 2012 50564 2036 50566
rect 2092 50564 2116 50566
rect 2172 50564 2196 50566
rect 2252 50564 2258 50566
rect 1950 50555 2258 50564
rect 2424 50538 2452 56646
rect 2332 50510 2452 50538
rect 1860 49972 1912 49978
rect 1860 49914 1912 49920
rect 1766 40896 1822 40905
rect 1766 40831 1822 40840
rect 1872 40746 1900 49914
rect 1950 49532 2258 49541
rect 1950 49530 1956 49532
rect 2012 49530 2036 49532
rect 2092 49530 2116 49532
rect 2172 49530 2196 49532
rect 2252 49530 2258 49532
rect 2012 49478 2014 49530
rect 2194 49478 2196 49530
rect 1950 49476 1956 49478
rect 2012 49476 2036 49478
rect 2092 49476 2116 49478
rect 2172 49476 2196 49478
rect 2252 49476 2258 49478
rect 1950 49467 2258 49476
rect 1950 48444 2258 48453
rect 1950 48442 1956 48444
rect 2012 48442 2036 48444
rect 2092 48442 2116 48444
rect 2172 48442 2196 48444
rect 2252 48442 2258 48444
rect 2012 48390 2014 48442
rect 2194 48390 2196 48442
rect 1950 48388 1956 48390
rect 2012 48388 2036 48390
rect 2092 48388 2116 48390
rect 2172 48388 2196 48390
rect 2252 48388 2258 48390
rect 1950 48379 2258 48388
rect 1950 47356 2258 47365
rect 1950 47354 1956 47356
rect 2012 47354 2036 47356
rect 2092 47354 2116 47356
rect 2172 47354 2196 47356
rect 2252 47354 2258 47356
rect 2012 47302 2014 47354
rect 2194 47302 2196 47354
rect 1950 47300 1956 47302
rect 2012 47300 2036 47302
rect 2092 47300 2116 47302
rect 2172 47300 2196 47302
rect 2252 47300 2258 47302
rect 1950 47291 2258 47300
rect 1950 46268 2258 46277
rect 1950 46266 1956 46268
rect 2012 46266 2036 46268
rect 2092 46266 2116 46268
rect 2172 46266 2196 46268
rect 2252 46266 2258 46268
rect 2012 46214 2014 46266
rect 2194 46214 2196 46266
rect 1950 46212 1956 46214
rect 2012 46212 2036 46214
rect 2092 46212 2116 46214
rect 2172 46212 2196 46214
rect 2252 46212 2258 46214
rect 1950 46203 2258 46212
rect 1950 45180 2258 45189
rect 1950 45178 1956 45180
rect 2012 45178 2036 45180
rect 2092 45178 2116 45180
rect 2172 45178 2196 45180
rect 2252 45178 2258 45180
rect 2012 45126 2014 45178
rect 2194 45126 2196 45178
rect 1950 45124 1956 45126
rect 2012 45124 2036 45126
rect 2092 45124 2116 45126
rect 2172 45124 2196 45126
rect 2252 45124 2258 45126
rect 1950 45115 2258 45124
rect 2136 44736 2188 44742
rect 2136 44678 2188 44684
rect 2148 44470 2176 44678
rect 2136 44464 2188 44470
rect 2332 44418 2360 50510
rect 2516 50402 2544 69702
rect 2610 69660 2918 69669
rect 2610 69658 2616 69660
rect 2672 69658 2696 69660
rect 2752 69658 2776 69660
rect 2832 69658 2856 69660
rect 2912 69658 2918 69660
rect 2672 69606 2674 69658
rect 2854 69606 2856 69658
rect 2610 69604 2616 69606
rect 2672 69604 2696 69606
rect 2752 69604 2776 69606
rect 2832 69604 2856 69606
rect 2912 69604 2918 69606
rect 2610 69595 2918 69604
rect 2610 68572 2918 68581
rect 2610 68570 2616 68572
rect 2672 68570 2696 68572
rect 2752 68570 2776 68572
rect 2832 68570 2856 68572
rect 2912 68570 2918 68572
rect 2672 68518 2674 68570
rect 2854 68518 2856 68570
rect 2610 68516 2616 68518
rect 2672 68516 2696 68518
rect 2752 68516 2776 68518
rect 2832 68516 2856 68518
rect 2912 68516 2918 68518
rect 2610 68507 2918 68516
rect 2610 67484 2918 67493
rect 2610 67482 2616 67484
rect 2672 67482 2696 67484
rect 2752 67482 2776 67484
rect 2832 67482 2856 67484
rect 2912 67482 2918 67484
rect 2672 67430 2674 67482
rect 2854 67430 2856 67482
rect 2610 67428 2616 67430
rect 2672 67428 2696 67430
rect 2752 67428 2776 67430
rect 2832 67428 2856 67430
rect 2912 67428 2918 67430
rect 2610 67419 2918 67428
rect 3700 67244 3752 67250
rect 3700 67186 3752 67192
rect 2610 66396 2918 66405
rect 2610 66394 2616 66396
rect 2672 66394 2696 66396
rect 2752 66394 2776 66396
rect 2832 66394 2856 66396
rect 2912 66394 2918 66396
rect 2672 66342 2674 66394
rect 2854 66342 2856 66394
rect 2610 66340 2616 66342
rect 2672 66340 2696 66342
rect 2752 66340 2776 66342
rect 2832 66340 2856 66342
rect 2912 66340 2918 66342
rect 2610 66331 2918 66340
rect 3608 65408 3660 65414
rect 3608 65350 3660 65356
rect 2610 65308 2918 65317
rect 2610 65306 2616 65308
rect 2672 65306 2696 65308
rect 2752 65306 2776 65308
rect 2832 65306 2856 65308
rect 2912 65306 2918 65308
rect 2672 65254 2674 65306
rect 2854 65254 2856 65306
rect 2610 65252 2616 65254
rect 2672 65252 2696 65254
rect 2752 65252 2776 65254
rect 2832 65252 2856 65254
rect 2912 65252 2918 65254
rect 2610 65243 2918 65252
rect 2610 64220 2918 64229
rect 2610 64218 2616 64220
rect 2672 64218 2696 64220
rect 2752 64218 2776 64220
rect 2832 64218 2856 64220
rect 2912 64218 2918 64220
rect 2672 64166 2674 64218
rect 2854 64166 2856 64218
rect 2610 64164 2616 64166
rect 2672 64164 2696 64166
rect 2752 64164 2776 64166
rect 2832 64164 2856 64166
rect 2912 64164 2918 64166
rect 2610 64155 2918 64164
rect 2610 63132 2918 63141
rect 2610 63130 2616 63132
rect 2672 63130 2696 63132
rect 2752 63130 2776 63132
rect 2832 63130 2856 63132
rect 2912 63130 2918 63132
rect 2672 63078 2674 63130
rect 2854 63078 2856 63130
rect 2610 63076 2616 63078
rect 2672 63076 2696 63078
rect 2752 63076 2776 63078
rect 2832 63076 2856 63078
rect 2912 63076 2918 63078
rect 2610 63067 2918 63076
rect 2610 62044 2918 62053
rect 2610 62042 2616 62044
rect 2672 62042 2696 62044
rect 2752 62042 2776 62044
rect 2832 62042 2856 62044
rect 2912 62042 2918 62044
rect 2672 61990 2674 62042
rect 2854 61990 2856 62042
rect 2610 61988 2616 61990
rect 2672 61988 2696 61990
rect 2752 61988 2776 61990
rect 2832 61988 2856 61990
rect 2912 61988 2918 61990
rect 2610 61979 2918 61988
rect 2610 60956 2918 60965
rect 2610 60954 2616 60956
rect 2672 60954 2696 60956
rect 2752 60954 2776 60956
rect 2832 60954 2856 60956
rect 2912 60954 2918 60956
rect 2672 60902 2674 60954
rect 2854 60902 2856 60954
rect 2610 60900 2616 60902
rect 2672 60900 2696 60902
rect 2752 60900 2776 60902
rect 2832 60900 2856 60902
rect 2912 60900 2918 60902
rect 2610 60891 2918 60900
rect 2610 59868 2918 59877
rect 2610 59866 2616 59868
rect 2672 59866 2696 59868
rect 2752 59866 2776 59868
rect 2832 59866 2856 59868
rect 2912 59866 2918 59868
rect 2672 59814 2674 59866
rect 2854 59814 2856 59866
rect 2610 59812 2616 59814
rect 2672 59812 2696 59814
rect 2752 59812 2776 59814
rect 2832 59812 2856 59814
rect 2912 59812 2918 59814
rect 2610 59803 2918 59812
rect 3240 59628 3292 59634
rect 3240 59570 3292 59576
rect 2610 58780 2918 58789
rect 2610 58778 2616 58780
rect 2672 58778 2696 58780
rect 2752 58778 2776 58780
rect 2832 58778 2856 58780
rect 2912 58778 2918 58780
rect 2672 58726 2674 58778
rect 2854 58726 2856 58778
rect 2610 58724 2616 58726
rect 2672 58724 2696 58726
rect 2752 58724 2776 58726
rect 2832 58724 2856 58726
rect 2912 58724 2918 58726
rect 2610 58715 2918 58724
rect 2610 57692 2918 57701
rect 2610 57690 2616 57692
rect 2672 57690 2696 57692
rect 2752 57690 2776 57692
rect 2832 57690 2856 57692
rect 2912 57690 2918 57692
rect 2672 57638 2674 57690
rect 2854 57638 2856 57690
rect 2610 57636 2616 57638
rect 2672 57636 2696 57638
rect 2752 57636 2776 57638
rect 2832 57636 2856 57638
rect 2912 57636 2918 57638
rect 2610 57627 2918 57636
rect 3252 57526 3280 59570
rect 3240 57520 3292 57526
rect 3240 57462 3292 57468
rect 3056 57452 3108 57458
rect 3056 57394 3108 57400
rect 3068 56681 3096 57394
rect 3054 56672 3110 56681
rect 2610 56604 2918 56613
rect 3054 56607 3110 56616
rect 2610 56602 2616 56604
rect 2672 56602 2696 56604
rect 2752 56602 2776 56604
rect 2832 56602 2856 56604
rect 2912 56602 2918 56604
rect 2672 56550 2674 56602
rect 2854 56550 2856 56602
rect 2610 56548 2616 56550
rect 2672 56548 2696 56550
rect 2752 56548 2776 56550
rect 2832 56548 2856 56550
rect 2912 56548 2918 56550
rect 2610 56539 2918 56548
rect 3252 56370 3280 57462
rect 3516 56976 3568 56982
rect 3516 56918 3568 56924
rect 2964 56364 3016 56370
rect 2964 56306 3016 56312
rect 3240 56364 3292 56370
rect 3240 56306 3292 56312
rect 2976 55758 3004 56306
rect 2964 55752 3016 55758
rect 2964 55694 3016 55700
rect 2610 55516 2918 55525
rect 2610 55514 2616 55516
rect 2672 55514 2696 55516
rect 2752 55514 2776 55516
rect 2832 55514 2856 55516
rect 2912 55514 2918 55516
rect 2672 55462 2674 55514
rect 2854 55462 2856 55514
rect 2610 55460 2616 55462
rect 2672 55460 2696 55462
rect 2752 55460 2776 55462
rect 2832 55460 2856 55462
rect 2912 55460 2918 55462
rect 2610 55451 2918 55460
rect 2976 55350 3004 55694
rect 2964 55344 3016 55350
rect 2964 55286 3016 55292
rect 2610 54428 2918 54437
rect 2610 54426 2616 54428
rect 2672 54426 2696 54428
rect 2752 54426 2776 54428
rect 2832 54426 2856 54428
rect 2912 54426 2918 54428
rect 2672 54374 2674 54426
rect 2854 54374 2856 54426
rect 2610 54372 2616 54374
rect 2672 54372 2696 54374
rect 2752 54372 2776 54374
rect 2832 54372 2856 54374
rect 2912 54372 2918 54374
rect 2610 54363 2918 54372
rect 2610 53340 2918 53349
rect 2610 53338 2616 53340
rect 2672 53338 2696 53340
rect 2752 53338 2776 53340
rect 2832 53338 2856 53340
rect 2912 53338 2918 53340
rect 2672 53286 2674 53338
rect 2854 53286 2856 53338
rect 2610 53284 2616 53286
rect 2672 53284 2696 53286
rect 2752 53284 2776 53286
rect 2832 53284 2856 53286
rect 2912 53284 2918 53286
rect 2610 53275 2918 53284
rect 2610 52252 2918 52261
rect 2610 52250 2616 52252
rect 2672 52250 2696 52252
rect 2752 52250 2776 52252
rect 2832 52250 2856 52252
rect 2912 52250 2918 52252
rect 2672 52198 2674 52250
rect 2854 52198 2856 52250
rect 2610 52196 2616 52198
rect 2672 52196 2696 52198
rect 2752 52196 2776 52198
rect 2832 52196 2856 52198
rect 2912 52196 2918 52198
rect 2610 52187 2918 52196
rect 2976 51474 3004 55286
rect 3332 53032 3384 53038
rect 3332 52974 3384 52980
rect 2964 51468 3016 51474
rect 2964 51410 3016 51416
rect 2610 51164 2918 51173
rect 2610 51162 2616 51164
rect 2672 51162 2696 51164
rect 2752 51162 2776 51164
rect 2832 51162 2856 51164
rect 2912 51162 2918 51164
rect 2672 51110 2674 51162
rect 2854 51110 2856 51162
rect 2610 51108 2616 51110
rect 2672 51108 2696 51110
rect 2752 51108 2776 51110
rect 2832 51108 2856 51110
rect 2912 51108 2918 51110
rect 2610 51099 2918 51108
rect 2596 50720 2648 50726
rect 2596 50662 2648 50668
rect 2136 44406 2188 44412
rect 2240 44390 2360 44418
rect 2424 50374 2544 50402
rect 2240 44266 2268 44390
rect 2320 44328 2372 44334
rect 2320 44270 2372 44276
rect 2228 44260 2280 44266
rect 2228 44202 2280 44208
rect 1950 44092 2258 44101
rect 1950 44090 1956 44092
rect 2012 44090 2036 44092
rect 2092 44090 2116 44092
rect 2172 44090 2196 44092
rect 2252 44090 2258 44092
rect 2012 44038 2014 44090
rect 2194 44038 2196 44090
rect 1950 44036 1956 44038
rect 2012 44036 2036 44038
rect 2092 44036 2116 44038
rect 2172 44036 2196 44038
rect 2252 44036 2258 44038
rect 1950 44027 2258 44036
rect 1950 43004 2258 43013
rect 1950 43002 1956 43004
rect 2012 43002 2036 43004
rect 2092 43002 2116 43004
rect 2172 43002 2196 43004
rect 2252 43002 2258 43004
rect 2012 42950 2014 43002
rect 2194 42950 2196 43002
rect 1950 42948 1956 42950
rect 2012 42948 2036 42950
rect 2092 42948 2116 42950
rect 2172 42948 2196 42950
rect 2252 42948 2258 42950
rect 1950 42939 2258 42948
rect 1952 42764 2004 42770
rect 1952 42706 2004 42712
rect 1964 42294 1992 42706
rect 1952 42288 2004 42294
rect 1952 42230 2004 42236
rect 2228 42220 2280 42226
rect 2332 42208 2360 44270
rect 2280 42180 2360 42208
rect 2228 42162 2280 42168
rect 1950 41916 2258 41925
rect 1950 41914 1956 41916
rect 2012 41914 2036 41916
rect 2092 41914 2116 41916
rect 2172 41914 2196 41916
rect 2252 41914 2258 41916
rect 2012 41862 2014 41914
rect 2194 41862 2196 41914
rect 1950 41860 1956 41862
rect 2012 41860 2036 41862
rect 2092 41860 2116 41862
rect 2172 41860 2196 41862
rect 2252 41860 2258 41862
rect 1950 41851 2258 41860
rect 1950 40828 2258 40837
rect 1950 40826 1956 40828
rect 2012 40826 2036 40828
rect 2092 40826 2116 40828
rect 2172 40826 2196 40828
rect 2252 40826 2258 40828
rect 2012 40774 2014 40826
rect 2194 40774 2196 40826
rect 1950 40772 1956 40774
rect 2012 40772 2036 40774
rect 2092 40772 2116 40774
rect 2172 40772 2196 40774
rect 2252 40772 2258 40774
rect 1950 40763 2258 40772
rect 1780 40718 1900 40746
rect 1780 31754 1808 40718
rect 1950 39740 2258 39749
rect 1950 39738 1956 39740
rect 2012 39738 2036 39740
rect 2092 39738 2116 39740
rect 2172 39738 2196 39740
rect 2252 39738 2258 39740
rect 2012 39686 2014 39738
rect 2194 39686 2196 39738
rect 1950 39684 1956 39686
rect 2012 39684 2036 39686
rect 2092 39684 2116 39686
rect 2172 39684 2196 39686
rect 2252 39684 2258 39686
rect 1950 39675 2258 39684
rect 2332 38962 2360 42180
rect 2320 38956 2372 38962
rect 2320 38898 2372 38904
rect 1950 38652 2258 38661
rect 1950 38650 1956 38652
rect 2012 38650 2036 38652
rect 2092 38650 2116 38652
rect 2172 38650 2196 38652
rect 2252 38650 2258 38652
rect 2012 38598 2014 38650
rect 2194 38598 2196 38650
rect 1950 38596 1956 38598
rect 2012 38596 2036 38598
rect 2092 38596 2116 38598
rect 2172 38596 2196 38598
rect 2252 38596 2258 38598
rect 1950 38587 2258 38596
rect 1950 37564 2258 37573
rect 1950 37562 1956 37564
rect 2012 37562 2036 37564
rect 2092 37562 2116 37564
rect 2172 37562 2196 37564
rect 2252 37562 2258 37564
rect 2012 37510 2014 37562
rect 2194 37510 2196 37562
rect 1950 37508 1956 37510
rect 2012 37508 2036 37510
rect 2092 37508 2116 37510
rect 2172 37508 2196 37510
rect 2252 37508 2258 37510
rect 1950 37499 2258 37508
rect 1860 37188 1912 37194
rect 1860 37130 1912 37136
rect 1872 35894 1900 37130
rect 1950 36476 2258 36485
rect 1950 36474 1956 36476
rect 2012 36474 2036 36476
rect 2092 36474 2116 36476
rect 2172 36474 2196 36476
rect 2252 36474 2258 36476
rect 2012 36422 2014 36474
rect 2194 36422 2196 36474
rect 1950 36420 1956 36422
rect 2012 36420 2036 36422
rect 2092 36420 2116 36422
rect 2172 36420 2196 36422
rect 2252 36420 2258 36422
rect 1950 36411 2258 36420
rect 1872 35866 2360 35894
rect 1950 35388 2258 35397
rect 1950 35386 1956 35388
rect 2012 35386 2036 35388
rect 2092 35386 2116 35388
rect 2172 35386 2196 35388
rect 2252 35386 2258 35388
rect 2012 35334 2014 35386
rect 2194 35334 2196 35386
rect 1950 35332 1956 35334
rect 2012 35332 2036 35334
rect 2092 35332 2116 35334
rect 2172 35332 2196 35334
rect 2252 35332 2258 35334
rect 1950 35323 2258 35332
rect 1950 34300 2258 34309
rect 1950 34298 1956 34300
rect 2012 34298 2036 34300
rect 2092 34298 2116 34300
rect 2172 34298 2196 34300
rect 2252 34298 2258 34300
rect 2012 34246 2014 34298
rect 2194 34246 2196 34298
rect 1950 34244 1956 34246
rect 2012 34244 2036 34246
rect 2092 34244 2116 34246
rect 2172 34244 2196 34246
rect 2252 34244 2258 34246
rect 1950 34235 2258 34244
rect 1950 33212 2258 33221
rect 1950 33210 1956 33212
rect 2012 33210 2036 33212
rect 2092 33210 2116 33212
rect 2172 33210 2196 33212
rect 2252 33210 2258 33212
rect 2012 33158 2014 33210
rect 2194 33158 2196 33210
rect 1950 33156 1956 33158
rect 2012 33156 2036 33158
rect 2092 33156 2116 33158
rect 2172 33156 2196 33158
rect 2252 33156 2258 33158
rect 1950 33147 2258 33156
rect 1950 32124 2258 32133
rect 1950 32122 1956 32124
rect 2012 32122 2036 32124
rect 2092 32122 2116 32124
rect 2172 32122 2196 32124
rect 2252 32122 2258 32124
rect 2012 32070 2014 32122
rect 2194 32070 2196 32122
rect 1950 32068 1956 32070
rect 2012 32068 2036 32070
rect 2092 32068 2116 32070
rect 2172 32068 2196 32070
rect 2252 32068 2258 32070
rect 1950 32059 2258 32068
rect 1780 31726 1900 31754
rect 1768 31340 1820 31346
rect 1768 31282 1820 31288
rect 1780 25498 1808 31282
rect 1768 25492 1820 25498
rect 1768 25434 1820 25440
rect 1768 25356 1820 25362
rect 1768 25298 1820 25304
rect 1780 16114 1808 25298
rect 1872 20330 1900 31726
rect 1950 31036 2258 31045
rect 1950 31034 1956 31036
rect 2012 31034 2036 31036
rect 2092 31034 2116 31036
rect 2172 31034 2196 31036
rect 2252 31034 2258 31036
rect 2012 30982 2014 31034
rect 2194 30982 2196 31034
rect 1950 30980 1956 30982
rect 2012 30980 2036 30982
rect 2092 30980 2116 30982
rect 2172 30980 2196 30982
rect 2252 30980 2258 30982
rect 1950 30971 2258 30980
rect 1950 29948 2258 29957
rect 1950 29946 1956 29948
rect 2012 29946 2036 29948
rect 2092 29946 2116 29948
rect 2172 29946 2196 29948
rect 2252 29946 2258 29948
rect 2012 29894 2014 29946
rect 2194 29894 2196 29946
rect 1950 29892 1956 29894
rect 2012 29892 2036 29894
rect 2092 29892 2116 29894
rect 2172 29892 2196 29894
rect 2252 29892 2258 29894
rect 1950 29883 2258 29892
rect 1950 28860 2258 28869
rect 1950 28858 1956 28860
rect 2012 28858 2036 28860
rect 2092 28858 2116 28860
rect 2172 28858 2196 28860
rect 2252 28858 2258 28860
rect 2012 28806 2014 28858
rect 2194 28806 2196 28858
rect 1950 28804 1956 28806
rect 2012 28804 2036 28806
rect 2092 28804 2116 28806
rect 2172 28804 2196 28806
rect 2252 28804 2258 28806
rect 1950 28795 2258 28804
rect 1950 27772 2258 27781
rect 1950 27770 1956 27772
rect 2012 27770 2036 27772
rect 2092 27770 2116 27772
rect 2172 27770 2196 27772
rect 2252 27770 2258 27772
rect 2012 27718 2014 27770
rect 2194 27718 2196 27770
rect 1950 27716 1956 27718
rect 2012 27716 2036 27718
rect 2092 27716 2116 27718
rect 2172 27716 2196 27718
rect 2252 27716 2258 27718
rect 1950 27707 2258 27716
rect 1950 26684 2258 26693
rect 1950 26682 1956 26684
rect 2012 26682 2036 26684
rect 2092 26682 2116 26684
rect 2172 26682 2196 26684
rect 2252 26682 2258 26684
rect 2012 26630 2014 26682
rect 2194 26630 2196 26682
rect 1950 26628 1956 26630
rect 2012 26628 2036 26630
rect 2092 26628 2116 26630
rect 2172 26628 2196 26630
rect 2252 26628 2258 26630
rect 1950 26619 2258 26628
rect 1950 25596 2258 25605
rect 1950 25594 1956 25596
rect 2012 25594 2036 25596
rect 2092 25594 2116 25596
rect 2172 25594 2196 25596
rect 2252 25594 2258 25596
rect 2012 25542 2014 25594
rect 2194 25542 2196 25594
rect 1950 25540 1956 25542
rect 2012 25540 2036 25542
rect 2092 25540 2116 25542
rect 2172 25540 2196 25542
rect 2252 25540 2258 25542
rect 1950 25531 2258 25540
rect 2332 25226 2360 35866
rect 2424 34678 2452 50374
rect 2608 50266 2636 50662
rect 2516 50238 2636 50266
rect 2516 44810 2544 50238
rect 2610 50076 2918 50085
rect 2610 50074 2616 50076
rect 2672 50074 2696 50076
rect 2752 50074 2776 50076
rect 2832 50074 2856 50076
rect 2912 50074 2918 50076
rect 2672 50022 2674 50074
rect 2854 50022 2856 50074
rect 2610 50020 2616 50022
rect 2672 50020 2696 50022
rect 2752 50020 2776 50022
rect 2832 50020 2856 50022
rect 2912 50020 2918 50022
rect 2610 50011 2918 50020
rect 2976 49774 3004 51410
rect 3148 50448 3200 50454
rect 3148 50390 3200 50396
rect 2964 49768 3016 49774
rect 2964 49710 3016 49716
rect 2610 48988 2918 48997
rect 2610 48986 2616 48988
rect 2672 48986 2696 48988
rect 2752 48986 2776 48988
rect 2832 48986 2856 48988
rect 2912 48986 2918 48988
rect 2672 48934 2674 48986
rect 2854 48934 2856 48986
rect 2610 48932 2616 48934
rect 2672 48932 2696 48934
rect 2752 48932 2776 48934
rect 2832 48932 2856 48934
rect 2912 48932 2918 48934
rect 2610 48923 2918 48932
rect 2610 47900 2918 47909
rect 2610 47898 2616 47900
rect 2672 47898 2696 47900
rect 2752 47898 2776 47900
rect 2832 47898 2856 47900
rect 2912 47898 2918 47900
rect 2672 47846 2674 47898
rect 2854 47846 2856 47898
rect 2610 47844 2616 47846
rect 2672 47844 2696 47846
rect 2752 47844 2776 47846
rect 2832 47844 2856 47846
rect 2912 47844 2918 47846
rect 2610 47835 2918 47844
rect 2964 47660 3016 47666
rect 2964 47602 3016 47608
rect 3056 47660 3108 47666
rect 3056 47602 3108 47608
rect 2976 47122 3004 47602
rect 3068 47297 3096 47602
rect 3054 47288 3110 47297
rect 3054 47223 3110 47232
rect 3056 47184 3108 47190
rect 3056 47126 3108 47132
rect 2964 47116 3016 47122
rect 2964 47058 3016 47064
rect 2610 46812 2918 46821
rect 2610 46810 2616 46812
rect 2672 46810 2696 46812
rect 2752 46810 2776 46812
rect 2832 46810 2856 46812
rect 2912 46810 2918 46812
rect 2672 46758 2674 46810
rect 2854 46758 2856 46810
rect 2610 46756 2616 46758
rect 2672 46756 2696 46758
rect 2752 46756 2776 46758
rect 2832 46756 2856 46758
rect 2912 46756 2918 46758
rect 2610 46747 2918 46756
rect 2610 45724 2918 45733
rect 2610 45722 2616 45724
rect 2672 45722 2696 45724
rect 2752 45722 2776 45724
rect 2832 45722 2856 45724
rect 2912 45722 2918 45724
rect 2672 45670 2674 45722
rect 2854 45670 2856 45722
rect 2610 45668 2616 45670
rect 2672 45668 2696 45670
rect 2752 45668 2776 45670
rect 2832 45668 2856 45670
rect 2912 45668 2918 45670
rect 2610 45659 2918 45668
rect 2504 44804 2556 44810
rect 2504 44746 2556 44752
rect 2610 44636 2918 44645
rect 2610 44634 2616 44636
rect 2672 44634 2696 44636
rect 2752 44634 2776 44636
rect 2832 44634 2856 44636
rect 2912 44634 2918 44636
rect 2672 44582 2674 44634
rect 2854 44582 2856 44634
rect 2610 44580 2616 44582
rect 2672 44580 2696 44582
rect 2752 44580 2776 44582
rect 2832 44580 2856 44582
rect 2912 44580 2918 44582
rect 2610 44571 2918 44580
rect 2504 44260 2556 44266
rect 2504 44202 2556 44208
rect 2516 39642 2544 44202
rect 2610 43548 2918 43557
rect 2610 43546 2616 43548
rect 2672 43546 2696 43548
rect 2752 43546 2776 43548
rect 2832 43546 2856 43548
rect 2912 43546 2918 43548
rect 2672 43494 2674 43546
rect 2854 43494 2856 43546
rect 2610 43492 2616 43494
rect 2672 43492 2696 43494
rect 2752 43492 2776 43494
rect 2832 43492 2856 43494
rect 2912 43492 2918 43494
rect 2610 43483 2918 43492
rect 2610 42460 2918 42469
rect 2610 42458 2616 42460
rect 2672 42458 2696 42460
rect 2752 42458 2776 42460
rect 2832 42458 2856 42460
rect 2912 42458 2918 42460
rect 2672 42406 2674 42458
rect 2854 42406 2856 42458
rect 2610 42404 2616 42406
rect 2672 42404 2696 42406
rect 2752 42404 2776 42406
rect 2832 42404 2856 42406
rect 2912 42404 2918 42406
rect 2610 42395 2918 42404
rect 2610 41372 2918 41381
rect 2610 41370 2616 41372
rect 2672 41370 2696 41372
rect 2752 41370 2776 41372
rect 2832 41370 2856 41372
rect 2912 41370 2918 41372
rect 2672 41318 2674 41370
rect 2854 41318 2856 41370
rect 2610 41316 2616 41318
rect 2672 41316 2696 41318
rect 2752 41316 2776 41318
rect 2832 41316 2856 41318
rect 2912 41316 2918 41318
rect 2610 41307 2918 41316
rect 2610 40284 2918 40293
rect 2610 40282 2616 40284
rect 2672 40282 2696 40284
rect 2752 40282 2776 40284
rect 2832 40282 2856 40284
rect 2912 40282 2918 40284
rect 2672 40230 2674 40282
rect 2854 40230 2856 40282
rect 2610 40228 2616 40230
rect 2672 40228 2696 40230
rect 2752 40228 2776 40230
rect 2832 40228 2856 40230
rect 2912 40228 2918 40230
rect 2610 40219 2918 40228
rect 2504 39636 2556 39642
rect 2504 39578 2556 39584
rect 2610 39196 2918 39205
rect 2610 39194 2616 39196
rect 2672 39194 2696 39196
rect 2752 39194 2776 39196
rect 2832 39194 2856 39196
rect 2912 39194 2918 39196
rect 2672 39142 2674 39194
rect 2854 39142 2856 39194
rect 2610 39140 2616 39142
rect 2672 39140 2696 39142
rect 2752 39140 2776 39142
rect 2832 39140 2856 39142
rect 2912 39140 2918 39142
rect 2610 39131 2918 39140
rect 2964 38752 3016 38758
rect 2964 38694 3016 38700
rect 2610 38108 2918 38117
rect 2610 38106 2616 38108
rect 2672 38106 2696 38108
rect 2752 38106 2776 38108
rect 2832 38106 2856 38108
rect 2912 38106 2918 38108
rect 2672 38054 2674 38106
rect 2854 38054 2856 38106
rect 2610 38052 2616 38054
rect 2672 38052 2696 38054
rect 2752 38052 2776 38054
rect 2832 38052 2856 38054
rect 2912 38052 2918 38054
rect 2610 38043 2918 38052
rect 2976 37262 3004 38694
rect 2964 37256 3016 37262
rect 2964 37198 3016 37204
rect 2610 37020 2918 37029
rect 2610 37018 2616 37020
rect 2672 37018 2696 37020
rect 2752 37018 2776 37020
rect 2832 37018 2856 37020
rect 2912 37018 2918 37020
rect 2672 36966 2674 37018
rect 2854 36966 2856 37018
rect 2610 36964 2616 36966
rect 2672 36964 2696 36966
rect 2752 36964 2776 36966
rect 2832 36964 2856 36966
rect 2912 36964 2918 36966
rect 2610 36955 2918 36964
rect 2610 35932 2918 35941
rect 2610 35930 2616 35932
rect 2672 35930 2696 35932
rect 2752 35930 2776 35932
rect 2832 35930 2856 35932
rect 2912 35930 2918 35932
rect 2672 35878 2674 35930
rect 2854 35878 2856 35930
rect 2610 35876 2616 35878
rect 2672 35876 2696 35878
rect 2752 35876 2776 35878
rect 2832 35876 2856 35878
rect 2912 35876 2918 35878
rect 2610 35867 2918 35876
rect 2610 34844 2918 34853
rect 2610 34842 2616 34844
rect 2672 34842 2696 34844
rect 2752 34842 2776 34844
rect 2832 34842 2856 34844
rect 2912 34842 2918 34844
rect 2672 34790 2674 34842
rect 2854 34790 2856 34842
rect 2610 34788 2616 34790
rect 2672 34788 2696 34790
rect 2752 34788 2776 34790
rect 2832 34788 2856 34790
rect 2912 34788 2918 34790
rect 2610 34779 2918 34788
rect 2412 34672 2464 34678
rect 2412 34614 2464 34620
rect 2610 33756 2918 33765
rect 2610 33754 2616 33756
rect 2672 33754 2696 33756
rect 2752 33754 2776 33756
rect 2832 33754 2856 33756
rect 2912 33754 2918 33756
rect 2672 33702 2674 33754
rect 2854 33702 2856 33754
rect 2610 33700 2616 33702
rect 2672 33700 2696 33702
rect 2752 33700 2776 33702
rect 2832 33700 2856 33702
rect 2912 33700 2918 33702
rect 2610 33691 2918 33700
rect 2610 32668 2918 32677
rect 2610 32666 2616 32668
rect 2672 32666 2696 32668
rect 2752 32666 2776 32668
rect 2832 32666 2856 32668
rect 2912 32666 2918 32668
rect 2672 32614 2674 32666
rect 2854 32614 2856 32666
rect 2610 32612 2616 32614
rect 2672 32612 2696 32614
rect 2752 32612 2776 32614
rect 2832 32612 2856 32614
rect 2912 32612 2918 32614
rect 2610 32603 2918 32612
rect 2412 32292 2464 32298
rect 2412 32234 2464 32240
rect 2320 25220 2372 25226
rect 2320 25162 2372 25168
rect 1950 24508 2258 24517
rect 1950 24506 1956 24508
rect 2012 24506 2036 24508
rect 2092 24506 2116 24508
rect 2172 24506 2196 24508
rect 2252 24506 2258 24508
rect 2012 24454 2014 24506
rect 2194 24454 2196 24506
rect 1950 24452 1956 24454
rect 2012 24452 2036 24454
rect 2092 24452 2116 24454
rect 2172 24452 2196 24454
rect 2252 24452 2258 24454
rect 1950 24443 2258 24452
rect 1950 23420 2258 23429
rect 1950 23418 1956 23420
rect 2012 23418 2036 23420
rect 2092 23418 2116 23420
rect 2172 23418 2196 23420
rect 2252 23418 2258 23420
rect 2012 23366 2014 23418
rect 2194 23366 2196 23418
rect 1950 23364 1956 23366
rect 2012 23364 2036 23366
rect 2092 23364 2116 23366
rect 2172 23364 2196 23366
rect 2252 23364 2258 23366
rect 1950 23355 2258 23364
rect 1950 22332 2258 22341
rect 1950 22330 1956 22332
rect 2012 22330 2036 22332
rect 2092 22330 2116 22332
rect 2172 22330 2196 22332
rect 2252 22330 2258 22332
rect 2012 22278 2014 22330
rect 2194 22278 2196 22330
rect 1950 22276 1956 22278
rect 2012 22276 2036 22278
rect 2092 22276 2116 22278
rect 2172 22276 2196 22278
rect 2252 22276 2258 22278
rect 1950 22267 2258 22276
rect 2424 22094 2452 32234
rect 2502 31784 2558 31793
rect 2502 31719 2558 31728
rect 2332 22066 2452 22094
rect 1950 21244 2258 21253
rect 1950 21242 1956 21244
rect 2012 21242 2036 21244
rect 2092 21242 2116 21244
rect 2172 21242 2196 21244
rect 2252 21242 2258 21244
rect 2012 21190 2014 21242
rect 2194 21190 2196 21242
rect 1950 21188 1956 21190
rect 2012 21188 2036 21190
rect 2092 21188 2116 21190
rect 2172 21188 2196 21190
rect 2252 21188 2258 21190
rect 1950 21179 2258 21188
rect 1860 20324 1912 20330
rect 1860 20266 1912 20272
rect 1950 20156 2258 20165
rect 1950 20154 1956 20156
rect 2012 20154 2036 20156
rect 2092 20154 2116 20156
rect 2172 20154 2196 20156
rect 2252 20154 2258 20156
rect 2012 20102 2014 20154
rect 2194 20102 2196 20154
rect 1950 20100 1956 20102
rect 2012 20100 2036 20102
rect 2092 20100 2116 20102
rect 2172 20100 2196 20102
rect 2252 20100 2258 20102
rect 1950 20091 2258 20100
rect 1950 19068 2258 19077
rect 1950 19066 1956 19068
rect 2012 19066 2036 19068
rect 2092 19066 2116 19068
rect 2172 19066 2196 19068
rect 2252 19066 2258 19068
rect 2012 19014 2014 19066
rect 2194 19014 2196 19066
rect 1950 19012 1956 19014
rect 2012 19012 2036 19014
rect 2092 19012 2116 19014
rect 2172 19012 2196 19014
rect 2252 19012 2258 19014
rect 1950 19003 2258 19012
rect 1950 17980 2258 17989
rect 1950 17978 1956 17980
rect 2012 17978 2036 17980
rect 2092 17978 2116 17980
rect 2172 17978 2196 17980
rect 2252 17978 2258 17980
rect 2012 17926 2014 17978
rect 2194 17926 2196 17978
rect 1950 17924 1956 17926
rect 2012 17924 2036 17926
rect 2092 17924 2116 17926
rect 2172 17924 2196 17926
rect 2252 17924 2258 17926
rect 1950 17915 2258 17924
rect 1950 16892 2258 16901
rect 1950 16890 1956 16892
rect 2012 16890 2036 16892
rect 2092 16890 2116 16892
rect 2172 16890 2196 16892
rect 2252 16890 2258 16892
rect 2012 16838 2014 16890
rect 2194 16838 2196 16890
rect 1950 16836 1956 16838
rect 2012 16836 2036 16838
rect 2092 16836 2116 16838
rect 2172 16836 2196 16838
rect 2252 16836 2258 16838
rect 1950 16827 2258 16836
rect 1768 16108 1820 16114
rect 1768 16050 1820 16056
rect 1950 15804 2258 15813
rect 1950 15802 1956 15804
rect 2012 15802 2036 15804
rect 2092 15802 2116 15804
rect 2172 15802 2196 15804
rect 2252 15802 2258 15804
rect 2012 15750 2014 15802
rect 2194 15750 2196 15802
rect 1950 15748 1956 15750
rect 2012 15748 2036 15750
rect 2092 15748 2116 15750
rect 2172 15748 2196 15750
rect 2252 15748 2258 15750
rect 1950 15739 2258 15748
rect 2332 15094 2360 22066
rect 2320 15088 2372 15094
rect 2320 15030 2372 15036
rect 1950 14716 2258 14725
rect 1950 14714 1956 14716
rect 2012 14714 2036 14716
rect 2092 14714 2116 14716
rect 2172 14714 2196 14716
rect 2252 14714 2258 14716
rect 2012 14662 2014 14714
rect 2194 14662 2196 14714
rect 1950 14660 1956 14662
rect 2012 14660 2036 14662
rect 2092 14660 2116 14662
rect 2172 14660 2196 14662
rect 2252 14660 2258 14662
rect 1950 14651 2258 14660
rect 1950 13628 2258 13637
rect 1950 13626 1956 13628
rect 2012 13626 2036 13628
rect 2092 13626 2116 13628
rect 2172 13626 2196 13628
rect 2252 13626 2258 13628
rect 2012 13574 2014 13626
rect 2194 13574 2196 13626
rect 1950 13572 1956 13574
rect 2012 13572 2036 13574
rect 2092 13572 2116 13574
rect 2172 13572 2196 13574
rect 2252 13572 2258 13574
rect 1950 13563 2258 13572
rect 1950 12540 2258 12549
rect 1950 12538 1956 12540
rect 2012 12538 2036 12540
rect 2092 12538 2116 12540
rect 2172 12538 2196 12540
rect 2252 12538 2258 12540
rect 2012 12486 2014 12538
rect 2194 12486 2196 12538
rect 1950 12484 1956 12486
rect 2012 12484 2036 12486
rect 2092 12484 2116 12486
rect 2172 12484 2196 12486
rect 2252 12484 2258 12486
rect 1950 12475 2258 12484
rect 1950 11452 2258 11461
rect 1950 11450 1956 11452
rect 2012 11450 2036 11452
rect 2092 11450 2116 11452
rect 2172 11450 2196 11452
rect 2252 11450 2258 11452
rect 2012 11398 2014 11450
rect 2194 11398 2196 11450
rect 1950 11396 1956 11398
rect 2012 11396 2036 11398
rect 2092 11396 2116 11398
rect 2172 11396 2196 11398
rect 2252 11396 2258 11398
rect 1950 11387 2258 11396
rect 1860 10804 1912 10810
rect 1860 10746 1912 10752
rect 1872 10266 1900 10746
rect 1950 10364 2258 10373
rect 1950 10362 1956 10364
rect 2012 10362 2036 10364
rect 2092 10362 2116 10364
rect 2172 10362 2196 10364
rect 2252 10362 2258 10364
rect 2012 10310 2014 10362
rect 2194 10310 2196 10362
rect 1950 10308 1956 10310
rect 2012 10308 2036 10310
rect 2092 10308 2116 10310
rect 2172 10308 2196 10310
rect 2252 10308 2258 10310
rect 1950 10299 2258 10308
rect 1860 10260 1912 10266
rect 1860 10202 1912 10208
rect 2320 9648 2372 9654
rect 2320 9590 2372 9596
rect 1950 9276 2258 9285
rect 1950 9274 1956 9276
rect 2012 9274 2036 9276
rect 2092 9274 2116 9276
rect 2172 9274 2196 9276
rect 2252 9274 2258 9276
rect 2012 9222 2014 9274
rect 2194 9222 2196 9274
rect 1950 9220 1956 9222
rect 2012 9220 2036 9222
rect 2092 9220 2116 9222
rect 2172 9220 2196 9222
rect 2252 9220 2258 9222
rect 1950 9211 2258 9220
rect 2332 8430 2360 9590
rect 2516 8430 2544 31719
rect 2610 31580 2918 31589
rect 2610 31578 2616 31580
rect 2672 31578 2696 31580
rect 2752 31578 2776 31580
rect 2832 31578 2856 31580
rect 2912 31578 2918 31580
rect 2672 31526 2674 31578
rect 2854 31526 2856 31578
rect 2610 31524 2616 31526
rect 2672 31524 2696 31526
rect 2752 31524 2776 31526
rect 2832 31524 2856 31526
rect 2912 31524 2918 31526
rect 2610 31515 2918 31524
rect 2610 30492 2918 30501
rect 2610 30490 2616 30492
rect 2672 30490 2696 30492
rect 2752 30490 2776 30492
rect 2832 30490 2856 30492
rect 2912 30490 2918 30492
rect 2672 30438 2674 30490
rect 2854 30438 2856 30490
rect 2610 30436 2616 30438
rect 2672 30436 2696 30438
rect 2752 30436 2776 30438
rect 2832 30436 2856 30438
rect 2912 30436 2918 30438
rect 2610 30427 2918 30436
rect 2610 29404 2918 29413
rect 2610 29402 2616 29404
rect 2672 29402 2696 29404
rect 2752 29402 2776 29404
rect 2832 29402 2856 29404
rect 2912 29402 2918 29404
rect 2672 29350 2674 29402
rect 2854 29350 2856 29402
rect 2610 29348 2616 29350
rect 2672 29348 2696 29350
rect 2752 29348 2776 29350
rect 2832 29348 2856 29350
rect 2912 29348 2918 29350
rect 2610 29339 2918 29348
rect 2610 28316 2918 28325
rect 2610 28314 2616 28316
rect 2672 28314 2696 28316
rect 2752 28314 2776 28316
rect 2832 28314 2856 28316
rect 2912 28314 2918 28316
rect 2672 28262 2674 28314
rect 2854 28262 2856 28314
rect 2610 28260 2616 28262
rect 2672 28260 2696 28262
rect 2752 28260 2776 28262
rect 2832 28260 2856 28262
rect 2912 28260 2918 28262
rect 2610 28251 2918 28260
rect 2610 27228 2918 27237
rect 2610 27226 2616 27228
rect 2672 27226 2696 27228
rect 2752 27226 2776 27228
rect 2832 27226 2856 27228
rect 2912 27226 2918 27228
rect 2672 27174 2674 27226
rect 2854 27174 2856 27226
rect 2610 27172 2616 27174
rect 2672 27172 2696 27174
rect 2752 27172 2776 27174
rect 2832 27172 2856 27174
rect 2912 27172 2918 27174
rect 2610 27163 2918 27172
rect 2610 26140 2918 26149
rect 2610 26138 2616 26140
rect 2672 26138 2696 26140
rect 2752 26138 2776 26140
rect 2832 26138 2856 26140
rect 2912 26138 2918 26140
rect 2672 26086 2674 26138
rect 2854 26086 2856 26138
rect 2610 26084 2616 26086
rect 2672 26084 2696 26086
rect 2752 26084 2776 26086
rect 2832 26084 2856 26086
rect 2912 26084 2918 26086
rect 2610 26075 2918 26084
rect 2610 25052 2918 25061
rect 2610 25050 2616 25052
rect 2672 25050 2696 25052
rect 2752 25050 2776 25052
rect 2832 25050 2856 25052
rect 2912 25050 2918 25052
rect 2672 24998 2674 25050
rect 2854 24998 2856 25050
rect 2610 24996 2616 24998
rect 2672 24996 2696 24998
rect 2752 24996 2776 24998
rect 2832 24996 2856 24998
rect 2912 24996 2918 24998
rect 2610 24987 2918 24996
rect 2610 23964 2918 23973
rect 2610 23962 2616 23964
rect 2672 23962 2696 23964
rect 2752 23962 2776 23964
rect 2832 23962 2856 23964
rect 2912 23962 2918 23964
rect 2672 23910 2674 23962
rect 2854 23910 2856 23962
rect 2610 23908 2616 23910
rect 2672 23908 2696 23910
rect 2752 23908 2776 23910
rect 2832 23908 2856 23910
rect 2912 23908 2918 23910
rect 2610 23899 2918 23908
rect 2610 22876 2918 22885
rect 2610 22874 2616 22876
rect 2672 22874 2696 22876
rect 2752 22874 2776 22876
rect 2832 22874 2856 22876
rect 2912 22874 2918 22876
rect 2672 22822 2674 22874
rect 2854 22822 2856 22874
rect 2610 22820 2616 22822
rect 2672 22820 2696 22822
rect 2752 22820 2776 22822
rect 2832 22820 2856 22822
rect 2912 22820 2918 22822
rect 2610 22811 2918 22820
rect 3068 22094 3096 47126
rect 2976 22066 3096 22094
rect 2610 21788 2918 21797
rect 2610 21786 2616 21788
rect 2672 21786 2696 21788
rect 2752 21786 2776 21788
rect 2832 21786 2856 21788
rect 2912 21786 2918 21788
rect 2672 21734 2674 21786
rect 2854 21734 2856 21786
rect 2610 21732 2616 21734
rect 2672 21732 2696 21734
rect 2752 21732 2776 21734
rect 2832 21732 2856 21734
rect 2912 21732 2918 21734
rect 2610 21723 2918 21732
rect 2610 20700 2918 20709
rect 2610 20698 2616 20700
rect 2672 20698 2696 20700
rect 2752 20698 2776 20700
rect 2832 20698 2856 20700
rect 2912 20698 2918 20700
rect 2672 20646 2674 20698
rect 2854 20646 2856 20698
rect 2610 20644 2616 20646
rect 2672 20644 2696 20646
rect 2752 20644 2776 20646
rect 2832 20644 2856 20646
rect 2912 20644 2918 20646
rect 2610 20635 2918 20644
rect 2610 19612 2918 19621
rect 2610 19610 2616 19612
rect 2672 19610 2696 19612
rect 2752 19610 2776 19612
rect 2832 19610 2856 19612
rect 2912 19610 2918 19612
rect 2672 19558 2674 19610
rect 2854 19558 2856 19610
rect 2610 19556 2616 19558
rect 2672 19556 2696 19558
rect 2752 19556 2776 19558
rect 2832 19556 2856 19558
rect 2912 19556 2918 19558
rect 2610 19547 2918 19556
rect 2610 18524 2918 18533
rect 2610 18522 2616 18524
rect 2672 18522 2696 18524
rect 2752 18522 2776 18524
rect 2832 18522 2856 18524
rect 2912 18522 2918 18524
rect 2672 18470 2674 18522
rect 2854 18470 2856 18522
rect 2610 18468 2616 18470
rect 2672 18468 2696 18470
rect 2752 18468 2776 18470
rect 2832 18468 2856 18470
rect 2912 18468 2918 18470
rect 2610 18459 2918 18468
rect 2610 17436 2918 17445
rect 2610 17434 2616 17436
rect 2672 17434 2696 17436
rect 2752 17434 2776 17436
rect 2832 17434 2856 17436
rect 2912 17434 2918 17436
rect 2672 17382 2674 17434
rect 2854 17382 2856 17434
rect 2610 17380 2616 17382
rect 2672 17380 2696 17382
rect 2752 17380 2776 17382
rect 2832 17380 2856 17382
rect 2912 17380 2918 17382
rect 2610 17371 2918 17380
rect 2610 16348 2918 16357
rect 2610 16346 2616 16348
rect 2672 16346 2696 16348
rect 2752 16346 2776 16348
rect 2832 16346 2856 16348
rect 2912 16346 2918 16348
rect 2672 16294 2674 16346
rect 2854 16294 2856 16346
rect 2610 16292 2616 16294
rect 2672 16292 2696 16294
rect 2752 16292 2776 16294
rect 2832 16292 2856 16294
rect 2912 16292 2918 16294
rect 2610 16283 2918 16292
rect 2610 15260 2918 15269
rect 2610 15258 2616 15260
rect 2672 15258 2696 15260
rect 2752 15258 2776 15260
rect 2832 15258 2856 15260
rect 2912 15258 2918 15260
rect 2672 15206 2674 15258
rect 2854 15206 2856 15258
rect 2610 15204 2616 15206
rect 2672 15204 2696 15206
rect 2752 15204 2776 15206
rect 2832 15204 2856 15206
rect 2912 15204 2918 15206
rect 2610 15195 2918 15204
rect 2610 14172 2918 14181
rect 2610 14170 2616 14172
rect 2672 14170 2696 14172
rect 2752 14170 2776 14172
rect 2832 14170 2856 14172
rect 2912 14170 2918 14172
rect 2672 14118 2674 14170
rect 2854 14118 2856 14170
rect 2610 14116 2616 14118
rect 2672 14116 2696 14118
rect 2752 14116 2776 14118
rect 2832 14116 2856 14118
rect 2912 14116 2918 14118
rect 2610 14107 2918 14116
rect 2610 13084 2918 13093
rect 2610 13082 2616 13084
rect 2672 13082 2696 13084
rect 2752 13082 2776 13084
rect 2832 13082 2856 13084
rect 2912 13082 2918 13084
rect 2672 13030 2674 13082
rect 2854 13030 2856 13082
rect 2610 13028 2616 13030
rect 2672 13028 2696 13030
rect 2752 13028 2776 13030
rect 2832 13028 2856 13030
rect 2912 13028 2918 13030
rect 2610 13019 2918 13028
rect 2610 11996 2918 12005
rect 2610 11994 2616 11996
rect 2672 11994 2696 11996
rect 2752 11994 2776 11996
rect 2832 11994 2856 11996
rect 2912 11994 2918 11996
rect 2672 11942 2674 11994
rect 2854 11942 2856 11994
rect 2610 11940 2616 11942
rect 2672 11940 2696 11942
rect 2752 11940 2776 11942
rect 2832 11940 2856 11942
rect 2912 11940 2918 11942
rect 2610 11931 2918 11940
rect 2610 10908 2918 10917
rect 2610 10906 2616 10908
rect 2672 10906 2696 10908
rect 2752 10906 2776 10908
rect 2832 10906 2856 10908
rect 2912 10906 2918 10908
rect 2672 10854 2674 10906
rect 2854 10854 2856 10906
rect 2610 10852 2616 10854
rect 2672 10852 2696 10854
rect 2752 10852 2776 10854
rect 2832 10852 2856 10854
rect 2912 10852 2918 10854
rect 2610 10843 2918 10852
rect 2596 10736 2648 10742
rect 2594 10704 2596 10713
rect 2648 10704 2650 10713
rect 2594 10639 2650 10648
rect 2610 9820 2918 9829
rect 2610 9818 2616 9820
rect 2672 9818 2696 9820
rect 2752 9818 2776 9820
rect 2832 9818 2856 9820
rect 2912 9818 2918 9820
rect 2672 9766 2674 9818
rect 2854 9766 2856 9818
rect 2610 9764 2616 9766
rect 2672 9764 2696 9766
rect 2752 9764 2776 9766
rect 2832 9764 2856 9766
rect 2912 9764 2918 9766
rect 2610 9755 2918 9764
rect 2610 8732 2918 8741
rect 2610 8730 2616 8732
rect 2672 8730 2696 8732
rect 2752 8730 2776 8732
rect 2832 8730 2856 8732
rect 2912 8730 2918 8732
rect 2672 8678 2674 8730
rect 2854 8678 2856 8730
rect 2610 8676 2616 8678
rect 2672 8676 2696 8678
rect 2752 8676 2776 8678
rect 2832 8676 2856 8678
rect 2912 8676 2918 8678
rect 2610 8667 2918 8676
rect 2320 8424 2372 8430
rect 2320 8366 2372 8372
rect 2504 8424 2556 8430
rect 2504 8366 2556 8372
rect 1950 8188 2258 8197
rect 1950 8186 1956 8188
rect 2012 8186 2036 8188
rect 2092 8186 2116 8188
rect 2172 8186 2196 8188
rect 2252 8186 2258 8188
rect 2012 8134 2014 8186
rect 2194 8134 2196 8186
rect 1950 8132 1956 8134
rect 2012 8132 2036 8134
rect 2092 8132 2116 8134
rect 2172 8132 2196 8134
rect 2252 8132 2258 8134
rect 1950 8123 2258 8132
rect 1950 7100 2258 7109
rect 1950 7098 1956 7100
rect 2012 7098 2036 7100
rect 2092 7098 2116 7100
rect 2172 7098 2196 7100
rect 2252 7098 2258 7100
rect 2012 7046 2014 7098
rect 2194 7046 2196 7098
rect 1950 7044 1956 7046
rect 2012 7044 2036 7046
rect 2092 7044 2116 7046
rect 2172 7044 2196 7046
rect 2252 7044 2258 7046
rect 1950 7035 2258 7044
rect 1950 6012 2258 6021
rect 1950 6010 1956 6012
rect 2012 6010 2036 6012
rect 2092 6010 2116 6012
rect 2172 6010 2196 6012
rect 2252 6010 2258 6012
rect 2012 5958 2014 6010
rect 2194 5958 2196 6010
rect 1950 5956 1956 5958
rect 2012 5956 2036 5958
rect 2092 5956 2116 5958
rect 2172 5956 2196 5958
rect 2252 5956 2258 5958
rect 1950 5947 2258 5956
rect 2332 5710 2360 8366
rect 2976 7886 3004 22066
rect 3160 21554 3188 50390
rect 3344 50318 3372 52974
rect 3332 50312 3384 50318
rect 3332 50254 3384 50260
rect 3240 46980 3292 46986
rect 3240 46922 3292 46928
rect 3252 34678 3280 46922
rect 3344 44470 3372 50254
rect 3424 49632 3476 49638
rect 3424 49574 3476 49580
rect 3436 49230 3464 49574
rect 3424 49224 3476 49230
rect 3424 49166 3476 49172
rect 3436 48686 3464 49166
rect 3424 48680 3476 48686
rect 3424 48622 3476 48628
rect 3332 44464 3384 44470
rect 3332 44406 3384 44412
rect 3344 43858 3372 44406
rect 3436 44334 3464 48622
rect 3424 44328 3476 44334
rect 3424 44270 3476 44276
rect 3332 43852 3384 43858
rect 3332 43794 3384 43800
rect 3332 42560 3384 42566
rect 3332 42502 3384 42508
rect 3240 34672 3292 34678
rect 3240 34614 3292 34620
rect 3252 33318 3280 34614
rect 3240 33312 3292 33318
rect 3240 33254 3292 33260
rect 3240 30252 3292 30258
rect 3240 30194 3292 30200
rect 3252 29850 3280 30194
rect 3240 29844 3292 29850
rect 3240 29786 3292 29792
rect 3344 28150 3372 42502
rect 3332 28144 3384 28150
rect 3332 28086 3384 28092
rect 3332 21956 3384 21962
rect 3332 21898 3384 21904
rect 3344 21690 3372 21898
rect 3332 21684 3384 21690
rect 3332 21626 3384 21632
rect 3148 21548 3200 21554
rect 3148 21490 3200 21496
rect 3528 16182 3556 56918
rect 3620 55418 3648 65350
rect 3608 55412 3660 55418
rect 3608 55354 3660 55360
rect 3620 42634 3648 55354
rect 3712 49978 3740 67186
rect 3700 49972 3752 49978
rect 3700 49914 3752 49920
rect 3700 48748 3752 48754
rect 3700 48690 3752 48696
rect 3712 48249 3740 48690
rect 3698 48240 3754 48249
rect 3698 48175 3754 48184
rect 3804 46986 3832 69770
rect 3988 69494 4016 69838
rect 3976 69488 4028 69494
rect 3976 69430 4028 69436
rect 4068 65680 4120 65686
rect 4068 65622 4120 65628
rect 4080 65249 4108 65622
rect 4632 65618 4660 74666
rect 4620 65612 4672 65618
rect 4620 65554 4672 65560
rect 4066 65240 4122 65249
rect 4066 65175 4122 65184
rect 4160 62484 4212 62490
rect 4160 62426 4212 62432
rect 4068 59016 4120 59022
rect 4068 58958 4120 58964
rect 3976 47524 4028 47530
rect 3976 47466 4028 47472
rect 3792 46980 3844 46986
rect 3792 46922 3844 46928
rect 3608 42628 3660 42634
rect 3608 42570 3660 42576
rect 3516 16176 3568 16182
rect 3516 16118 3568 16124
rect 3148 11552 3200 11558
rect 3148 11494 3200 11500
rect 3160 10810 3188 11494
rect 3148 10804 3200 10810
rect 3148 10746 3200 10752
rect 2964 7880 3016 7886
rect 2964 7822 3016 7828
rect 2610 7644 2918 7653
rect 2610 7642 2616 7644
rect 2672 7642 2696 7644
rect 2752 7642 2776 7644
rect 2832 7642 2856 7644
rect 2912 7642 2918 7644
rect 2672 7590 2674 7642
rect 2854 7590 2856 7642
rect 2610 7588 2616 7590
rect 2672 7588 2696 7590
rect 2752 7588 2776 7590
rect 2832 7588 2856 7590
rect 2912 7588 2918 7590
rect 2610 7579 2918 7588
rect 2610 6556 2918 6565
rect 2610 6554 2616 6556
rect 2672 6554 2696 6556
rect 2752 6554 2776 6556
rect 2832 6554 2856 6556
rect 2912 6554 2918 6556
rect 2672 6502 2674 6554
rect 2854 6502 2856 6554
rect 2610 6500 2616 6502
rect 2672 6500 2696 6502
rect 2752 6500 2776 6502
rect 2832 6500 2856 6502
rect 2912 6500 2918 6502
rect 2610 6491 2918 6500
rect 3620 6458 3648 42570
rect 3700 35828 3752 35834
rect 3700 35770 3752 35776
rect 3712 8634 3740 35770
rect 3804 30258 3832 46922
rect 3988 46714 4016 47466
rect 3976 46708 4028 46714
rect 3976 46650 4028 46656
rect 3884 44736 3936 44742
rect 3884 44678 3936 44684
rect 3896 31754 3924 44678
rect 4080 36922 4108 58958
rect 4172 57338 4200 62426
rect 4250 62248 4306 62257
rect 4250 62183 4252 62192
rect 4304 62183 4306 62192
rect 4252 62154 4304 62160
rect 4344 62144 4396 62150
rect 4344 62086 4396 62092
rect 4172 57310 4292 57338
rect 4160 57248 4212 57254
rect 4160 57190 4212 57196
rect 4172 57050 4200 57190
rect 4160 57044 4212 57050
rect 4160 56986 4212 56992
rect 4160 51264 4212 51270
rect 4160 51206 4212 51212
rect 4172 49910 4200 51206
rect 4160 49904 4212 49910
rect 4160 49846 4212 49852
rect 4264 41414 4292 57310
rect 4172 41386 4292 41414
rect 4068 36916 4120 36922
rect 4068 36858 4120 36864
rect 3896 31726 4016 31754
rect 3792 30252 3844 30258
rect 3792 30194 3844 30200
rect 3884 12640 3936 12646
rect 3884 12582 3936 12588
rect 3896 12238 3924 12582
rect 3884 12232 3936 12238
rect 3884 12174 3936 12180
rect 3896 9654 3924 12174
rect 3884 9648 3936 9654
rect 3884 9590 3936 9596
rect 3988 9382 4016 31726
rect 4068 28008 4120 28014
rect 4068 27950 4120 27956
rect 4080 27606 4108 27950
rect 4068 27600 4120 27606
rect 4068 27542 4120 27548
rect 4080 26450 4108 27542
rect 4172 27538 4200 41386
rect 4160 27532 4212 27538
rect 4160 27474 4212 27480
rect 4068 26444 4120 26450
rect 4068 26386 4120 26392
rect 4080 25294 4108 26386
rect 4068 25288 4120 25294
rect 4068 25230 4120 25236
rect 4160 22092 4212 22098
rect 4160 22034 4212 22040
rect 4172 22001 4200 22034
rect 4158 21992 4214 22001
rect 4158 21927 4214 21936
rect 4356 20602 4384 62086
rect 4632 60518 4660 65554
rect 4804 61396 4856 61402
rect 4804 61338 4856 61344
rect 4620 60512 4672 60518
rect 4620 60454 4672 60460
rect 4528 56160 4580 56166
rect 4528 56102 4580 56108
rect 4436 49972 4488 49978
rect 4436 49914 4488 49920
rect 4448 49745 4476 49914
rect 4434 49736 4490 49745
rect 4434 49671 4490 49680
rect 4436 44804 4488 44810
rect 4436 44746 4488 44752
rect 4448 44402 4476 44746
rect 4436 44396 4488 44402
rect 4436 44338 4488 44344
rect 4540 36310 4568 56102
rect 4816 50386 4844 61338
rect 4988 57520 5040 57526
rect 4988 57462 5040 57468
rect 4896 55888 4948 55894
rect 4896 55830 4948 55836
rect 4804 50380 4856 50386
rect 4804 50322 4856 50328
rect 4804 47456 4856 47462
rect 4804 47398 4856 47404
rect 4528 36304 4580 36310
rect 4528 36246 4580 36252
rect 4816 35018 4844 47398
rect 4908 39030 4936 55830
rect 4896 39024 4948 39030
rect 4896 38966 4948 38972
rect 5000 35834 5028 57462
rect 5092 50318 5120 75142
rect 5264 69760 5316 69766
rect 5264 69702 5316 69708
rect 5172 59424 5224 59430
rect 5172 59366 5224 59372
rect 5080 50312 5132 50318
rect 5080 50254 5132 50260
rect 5080 40180 5132 40186
rect 5080 40122 5132 40128
rect 4988 35828 5040 35834
rect 4988 35770 5040 35776
rect 4804 35012 4856 35018
rect 4804 34954 4856 34960
rect 4896 34604 4948 34610
rect 4896 34546 4948 34552
rect 4620 33108 4672 33114
rect 4620 33050 4672 33056
rect 4632 29238 4660 33050
rect 4620 29232 4672 29238
rect 4620 29174 4672 29180
rect 4436 29164 4488 29170
rect 4436 29106 4488 29112
rect 4344 20596 4396 20602
rect 4344 20538 4396 20544
rect 4448 20262 4476 29106
rect 4802 20768 4858 20777
rect 4802 20703 4858 20712
rect 4436 20256 4488 20262
rect 4436 20198 4488 20204
rect 4816 11830 4844 20703
rect 4804 11824 4856 11830
rect 4804 11766 4856 11772
rect 4908 10470 4936 34546
rect 5092 27470 5120 40122
rect 5080 27464 5132 27470
rect 5080 27406 5132 27412
rect 4896 10464 4948 10470
rect 4896 10406 4948 10412
rect 4252 9580 4304 9586
rect 4252 9522 4304 9528
rect 3976 9376 4028 9382
rect 3976 9318 4028 9324
rect 3700 8628 3752 8634
rect 3700 8570 3752 8576
rect 4264 8498 4292 9522
rect 5184 8838 5212 59366
rect 5276 12918 5304 69702
rect 5460 63034 5488 75278
rect 5552 73234 5580 75958
rect 7116 75954 7144 76230
rect 7944 76214 8064 76242
rect 7610 76188 7918 76197
rect 7610 76186 7616 76188
rect 7672 76186 7696 76188
rect 7752 76186 7776 76188
rect 7832 76186 7856 76188
rect 7912 76186 7918 76188
rect 7672 76134 7674 76186
rect 7854 76134 7856 76186
rect 7610 76132 7616 76134
rect 7672 76132 7696 76134
rect 7752 76132 7776 76134
rect 7832 76132 7856 76134
rect 7912 76132 7918 76134
rect 7610 76123 7918 76132
rect 7564 76016 7616 76022
rect 7562 75984 7564 75993
rect 7616 75984 7618 75993
rect 7104 75948 7156 75954
rect 7104 75890 7156 75896
rect 7380 75948 7432 75954
rect 7562 75919 7618 75928
rect 7380 75890 7432 75896
rect 6644 75880 6696 75886
rect 6644 75822 6696 75828
rect 6552 75200 6604 75206
rect 6550 75168 6552 75177
rect 6604 75168 6606 75177
rect 6550 75103 6606 75112
rect 6552 74928 6604 74934
rect 6552 74870 6604 74876
rect 6460 74860 6512 74866
rect 6460 74802 6512 74808
rect 5540 73228 5592 73234
rect 5540 73170 5592 73176
rect 5552 71670 5580 73170
rect 5540 71664 5592 71670
rect 5540 71606 5592 71612
rect 5552 71058 5580 71606
rect 6276 71188 6328 71194
rect 6276 71130 6328 71136
rect 5540 71052 5592 71058
rect 5540 70994 5592 71000
rect 6288 70922 6316 71130
rect 6276 70916 6328 70922
rect 6276 70858 6328 70864
rect 6184 68332 6236 68338
rect 6184 68274 6236 68280
rect 5448 63028 5500 63034
rect 5448 62970 5500 62976
rect 5908 60648 5960 60654
rect 5908 60590 5960 60596
rect 5724 55412 5776 55418
rect 5724 55354 5776 55360
rect 5736 55282 5764 55354
rect 5540 55276 5592 55282
rect 5540 55218 5592 55224
rect 5724 55276 5776 55282
rect 5724 55218 5776 55224
rect 5448 42696 5500 42702
rect 5448 42638 5500 42644
rect 5356 34740 5408 34746
rect 5356 34682 5408 34688
rect 5368 25498 5396 34682
rect 5460 29306 5488 42638
rect 5552 37942 5580 55218
rect 5724 44192 5776 44198
rect 5724 44134 5776 44140
rect 5540 37936 5592 37942
rect 5540 37878 5592 37884
rect 5736 35562 5764 44134
rect 5724 35556 5776 35562
rect 5724 35498 5776 35504
rect 5724 30592 5776 30598
rect 5724 30534 5776 30540
rect 5448 29300 5500 29306
rect 5448 29242 5500 29248
rect 5632 28552 5684 28558
rect 5632 28494 5684 28500
rect 5356 25492 5408 25498
rect 5356 25434 5408 25440
rect 5540 22636 5592 22642
rect 5540 22578 5592 22584
rect 5552 20466 5580 22578
rect 5540 20460 5592 20466
rect 5540 20402 5592 20408
rect 5552 16658 5580 20402
rect 5540 16652 5592 16658
rect 5540 16594 5592 16600
rect 5264 12912 5316 12918
rect 5264 12854 5316 12860
rect 5540 9580 5592 9586
rect 5540 9522 5592 9528
rect 5552 9178 5580 9522
rect 5540 9172 5592 9178
rect 5540 9114 5592 9120
rect 5172 8832 5224 8838
rect 5172 8774 5224 8780
rect 4252 8492 4304 8498
rect 4252 8434 4304 8440
rect 3608 6452 3660 6458
rect 3608 6394 3660 6400
rect 2320 5704 2372 5710
rect 2320 5646 2372 5652
rect 5080 5704 5132 5710
rect 5080 5646 5132 5652
rect 1676 5364 1728 5370
rect 1676 5306 1728 5312
rect 1950 4924 2258 4933
rect 1950 4922 1956 4924
rect 2012 4922 2036 4924
rect 2092 4922 2116 4924
rect 2172 4922 2196 4924
rect 2252 4922 2258 4924
rect 2012 4870 2014 4922
rect 2194 4870 2196 4922
rect 1950 4868 1956 4870
rect 2012 4868 2036 4870
rect 2092 4868 2116 4870
rect 2172 4868 2196 4870
rect 2252 4868 2258 4870
rect 1950 4859 2258 4868
rect 1216 4072 1268 4078
rect 1216 4014 1268 4020
rect 1950 3836 2258 3845
rect 1950 3834 1956 3836
rect 2012 3834 2036 3836
rect 2092 3834 2116 3836
rect 2172 3834 2196 3836
rect 2252 3834 2258 3836
rect 2012 3782 2014 3834
rect 2194 3782 2196 3834
rect 1950 3780 1956 3782
rect 2012 3780 2036 3782
rect 2092 3780 2116 3782
rect 2172 3780 2196 3782
rect 2252 3780 2258 3782
rect 1950 3771 2258 3780
rect 2332 2990 2360 5646
rect 2610 5468 2918 5477
rect 2610 5466 2616 5468
rect 2672 5466 2696 5468
rect 2752 5466 2776 5468
rect 2832 5466 2856 5468
rect 2912 5466 2918 5468
rect 2672 5414 2674 5466
rect 2854 5414 2856 5466
rect 2610 5412 2616 5414
rect 2672 5412 2696 5414
rect 2752 5412 2776 5414
rect 2832 5412 2856 5414
rect 2912 5412 2918 5414
rect 2610 5403 2918 5412
rect 2610 4380 2918 4389
rect 2610 4378 2616 4380
rect 2672 4378 2696 4380
rect 2752 4378 2776 4380
rect 2832 4378 2856 4380
rect 2912 4378 2918 4380
rect 2672 4326 2674 4378
rect 2854 4326 2856 4378
rect 2610 4324 2616 4326
rect 2672 4324 2696 4326
rect 2752 4324 2776 4326
rect 2832 4324 2856 4326
rect 2912 4324 2918 4326
rect 2610 4315 2918 4324
rect 5092 4146 5120 5646
rect 5080 4140 5132 4146
rect 5080 4082 5132 4088
rect 2610 3292 2918 3301
rect 2610 3290 2616 3292
rect 2672 3290 2696 3292
rect 2752 3290 2776 3292
rect 2832 3290 2856 3292
rect 2912 3290 2918 3292
rect 2672 3238 2674 3290
rect 2854 3238 2856 3290
rect 2610 3236 2616 3238
rect 2672 3236 2696 3238
rect 2752 3236 2776 3238
rect 2832 3236 2856 3238
rect 2912 3236 2918 3238
rect 2610 3227 2918 3236
rect 5644 3126 5672 28494
rect 5736 25362 5764 30534
rect 5816 26308 5868 26314
rect 5816 26250 5868 26256
rect 5724 25356 5776 25362
rect 5724 25298 5776 25304
rect 5724 17332 5776 17338
rect 5724 17274 5776 17280
rect 5736 11558 5764 17274
rect 5724 11552 5776 11558
rect 5724 11494 5776 11500
rect 5828 6390 5856 26250
rect 5920 17338 5948 60590
rect 6092 50992 6144 50998
rect 6092 50934 6144 50940
rect 6104 44742 6132 50934
rect 6196 47802 6224 68274
rect 6368 63232 6420 63238
rect 6368 63174 6420 63180
rect 6276 60036 6328 60042
rect 6276 59978 6328 59984
rect 6288 48618 6316 59978
rect 6276 48612 6328 48618
rect 6276 48554 6328 48560
rect 6184 47796 6236 47802
rect 6184 47738 6236 47744
rect 6092 44736 6144 44742
rect 6092 44678 6144 44684
rect 6276 41676 6328 41682
rect 6276 41618 6328 41624
rect 6092 41472 6144 41478
rect 6092 41414 6144 41420
rect 6184 41472 6236 41478
rect 6184 41414 6236 41420
rect 6104 26602 6132 41414
rect 6196 27962 6224 41414
rect 6288 30818 6316 41618
rect 6380 31414 6408 63174
rect 6472 47802 6500 74802
rect 6564 70854 6592 74870
rect 6552 70848 6604 70854
rect 6552 70790 6604 70796
rect 6552 69828 6604 69834
rect 6552 69770 6604 69776
rect 6564 64874 6592 69770
rect 6656 69766 6684 75822
rect 6950 75644 7258 75653
rect 6950 75642 6956 75644
rect 7012 75642 7036 75644
rect 7092 75642 7116 75644
rect 7172 75642 7196 75644
rect 7252 75642 7258 75644
rect 7012 75590 7014 75642
rect 7194 75590 7196 75642
rect 6950 75588 6956 75590
rect 7012 75588 7036 75590
rect 7092 75588 7116 75590
rect 7172 75588 7196 75590
rect 7252 75588 7258 75590
rect 6950 75579 7258 75588
rect 7288 75336 7340 75342
rect 7288 75278 7340 75284
rect 6736 74656 6788 74662
rect 6736 74598 6788 74604
rect 6644 69760 6696 69766
rect 6644 69702 6696 69708
rect 6564 64846 6684 64874
rect 6552 63504 6604 63510
rect 6552 63446 6604 63452
rect 6564 62898 6592 63446
rect 6552 62892 6604 62898
rect 6552 62834 6604 62840
rect 6564 60722 6592 62834
rect 6552 60716 6604 60722
rect 6552 60658 6604 60664
rect 6564 59702 6592 60658
rect 6552 59696 6604 59702
rect 6552 59638 6604 59644
rect 6552 55276 6604 55282
rect 6552 55218 6604 55224
rect 6460 47796 6512 47802
rect 6460 47738 6512 47744
rect 6460 46368 6512 46374
rect 6460 46310 6512 46316
rect 6472 42838 6500 46310
rect 6460 42832 6512 42838
rect 6460 42774 6512 42780
rect 6460 42696 6512 42702
rect 6460 42638 6512 42644
rect 6472 41614 6500 42638
rect 6460 41608 6512 41614
rect 6460 41550 6512 41556
rect 6460 31884 6512 31890
rect 6460 31826 6512 31832
rect 6368 31408 6420 31414
rect 6368 31350 6420 31356
rect 6288 30802 6408 30818
rect 6288 30796 6420 30802
rect 6288 30790 6368 30796
rect 6368 30738 6420 30744
rect 6380 29034 6408 30738
rect 6368 29028 6420 29034
rect 6368 28970 6420 28976
rect 6196 27934 6316 27962
rect 6104 26586 6224 26602
rect 6104 26580 6236 26586
rect 6104 26574 6184 26580
rect 6104 22094 6132 26574
rect 6184 26522 6236 26528
rect 6288 24138 6316 27934
rect 6276 24132 6328 24138
rect 6276 24074 6328 24080
rect 6472 23730 6500 31826
rect 6460 23724 6512 23730
rect 6460 23666 6512 23672
rect 6012 22066 6132 22094
rect 6184 22092 6236 22098
rect 6012 19854 6040 22066
rect 6184 22034 6236 22040
rect 6000 19848 6052 19854
rect 6000 19790 6052 19796
rect 5908 17332 5960 17338
rect 5908 17274 5960 17280
rect 5908 17060 5960 17066
rect 5908 17002 5960 17008
rect 5920 16454 5948 17002
rect 5908 16448 5960 16454
rect 5908 16390 5960 16396
rect 5816 6384 5868 6390
rect 5816 6326 5868 6332
rect 6196 5710 6224 22034
rect 6460 21888 6512 21894
rect 6460 21830 6512 21836
rect 6472 21486 6500 21830
rect 6460 21480 6512 21486
rect 6460 21422 6512 21428
rect 6276 11824 6328 11830
rect 6276 11766 6328 11772
rect 6288 6730 6316 11766
rect 6276 6724 6328 6730
rect 6276 6666 6328 6672
rect 6184 5704 6236 5710
rect 6184 5646 6236 5652
rect 6564 5098 6592 55218
rect 6656 48634 6684 64846
rect 6748 51074 6776 74598
rect 6950 74556 7258 74565
rect 6950 74554 6956 74556
rect 7012 74554 7036 74556
rect 7092 74554 7116 74556
rect 7172 74554 7196 74556
rect 7252 74554 7258 74556
rect 7012 74502 7014 74554
rect 7194 74502 7196 74554
rect 6950 74500 6956 74502
rect 7012 74500 7036 74502
rect 7092 74500 7116 74502
rect 7172 74500 7196 74502
rect 7252 74500 7258 74502
rect 6950 74491 7258 74500
rect 7300 73914 7328 75278
rect 7392 74458 7420 75890
rect 7610 75100 7918 75109
rect 7610 75098 7616 75100
rect 7672 75098 7696 75100
rect 7752 75098 7776 75100
rect 7832 75098 7856 75100
rect 7912 75098 7918 75100
rect 7672 75046 7674 75098
rect 7854 75046 7856 75098
rect 7610 75044 7616 75046
rect 7672 75044 7696 75046
rect 7752 75044 7776 75046
rect 7832 75044 7856 75046
rect 7912 75044 7918 75046
rect 7610 75035 7918 75044
rect 7380 74452 7432 74458
rect 7380 74394 7432 74400
rect 7610 74012 7918 74021
rect 7610 74010 7616 74012
rect 7672 74010 7696 74012
rect 7752 74010 7776 74012
rect 7832 74010 7856 74012
rect 7912 74010 7918 74012
rect 7672 73958 7674 74010
rect 7854 73958 7856 74010
rect 7610 73956 7616 73958
rect 7672 73956 7696 73958
rect 7752 73956 7776 73958
rect 7832 73956 7856 73958
rect 7912 73956 7918 73958
rect 7610 73947 7918 73956
rect 7288 73908 7340 73914
rect 7288 73850 7340 73856
rect 7380 73772 7432 73778
rect 7380 73714 7432 73720
rect 6950 73468 7258 73477
rect 6950 73466 6956 73468
rect 7012 73466 7036 73468
rect 7092 73466 7116 73468
rect 7172 73466 7196 73468
rect 7252 73466 7258 73468
rect 7012 73414 7014 73466
rect 7194 73414 7196 73466
rect 6950 73412 6956 73414
rect 7012 73412 7036 73414
rect 7092 73412 7116 73414
rect 7172 73412 7196 73414
rect 7252 73412 7258 73414
rect 6950 73403 7258 73412
rect 7392 72622 7420 73714
rect 7610 72924 7918 72933
rect 7610 72922 7616 72924
rect 7672 72922 7696 72924
rect 7752 72922 7776 72924
rect 7832 72922 7856 72924
rect 7912 72922 7918 72924
rect 7672 72870 7674 72922
rect 7854 72870 7856 72922
rect 7610 72868 7616 72870
rect 7672 72868 7696 72870
rect 7752 72868 7776 72870
rect 7832 72868 7856 72870
rect 7912 72868 7918 72870
rect 7610 72859 7918 72868
rect 7380 72616 7432 72622
rect 7380 72558 7432 72564
rect 6950 72380 7258 72389
rect 6950 72378 6956 72380
rect 7012 72378 7036 72380
rect 7092 72378 7116 72380
rect 7172 72378 7196 72380
rect 7252 72378 7258 72380
rect 7012 72326 7014 72378
rect 7194 72326 7196 72378
rect 6950 72324 6956 72326
rect 7012 72324 7036 72326
rect 7092 72324 7116 72326
rect 7172 72324 7196 72326
rect 7252 72324 7258 72326
rect 6950 72315 7258 72324
rect 6950 71292 7258 71301
rect 6950 71290 6956 71292
rect 7012 71290 7036 71292
rect 7092 71290 7116 71292
rect 7172 71290 7196 71292
rect 7252 71290 7258 71292
rect 7012 71238 7014 71290
rect 7194 71238 7196 71290
rect 6950 71236 6956 71238
rect 7012 71236 7036 71238
rect 7092 71236 7116 71238
rect 7172 71236 7196 71238
rect 7252 71236 7258 71238
rect 6950 71227 7258 71236
rect 6828 70984 6880 70990
rect 6828 70926 6880 70932
rect 6840 69986 6868 70926
rect 6950 70204 7258 70213
rect 6950 70202 6956 70204
rect 7012 70202 7036 70204
rect 7092 70202 7116 70204
rect 7172 70202 7196 70204
rect 7252 70202 7258 70204
rect 7012 70150 7014 70202
rect 7194 70150 7196 70202
rect 6950 70148 6956 70150
rect 7012 70148 7036 70150
rect 7092 70148 7116 70150
rect 7172 70148 7196 70150
rect 7252 70148 7258 70150
rect 6950 70139 7258 70148
rect 6840 69958 7052 69986
rect 7024 69902 7052 69958
rect 7012 69896 7064 69902
rect 7012 69838 7064 69844
rect 6828 69760 6880 69766
rect 7024 69748 7052 69838
rect 7024 69720 7328 69748
rect 6828 69702 6880 69708
rect 6840 60042 6868 69702
rect 6950 69116 7258 69125
rect 6950 69114 6956 69116
rect 7012 69114 7036 69116
rect 7092 69114 7116 69116
rect 7172 69114 7196 69116
rect 7252 69114 7258 69116
rect 7012 69062 7014 69114
rect 7194 69062 7196 69114
rect 6950 69060 6956 69062
rect 7012 69060 7036 69062
rect 7092 69060 7116 69062
rect 7172 69060 7196 69062
rect 7252 69060 7258 69062
rect 6950 69051 7258 69060
rect 6950 68028 7258 68037
rect 6950 68026 6956 68028
rect 7012 68026 7036 68028
rect 7092 68026 7116 68028
rect 7172 68026 7196 68028
rect 7252 68026 7258 68028
rect 7012 67974 7014 68026
rect 7194 67974 7196 68026
rect 6950 67972 6956 67974
rect 7012 67972 7036 67974
rect 7092 67972 7116 67974
rect 7172 67972 7196 67974
rect 7252 67972 7258 67974
rect 6950 67963 7258 67972
rect 6950 66940 7258 66949
rect 6950 66938 6956 66940
rect 7012 66938 7036 66940
rect 7092 66938 7116 66940
rect 7172 66938 7196 66940
rect 7252 66938 7258 66940
rect 7012 66886 7014 66938
rect 7194 66886 7196 66938
rect 6950 66884 6956 66886
rect 7012 66884 7036 66886
rect 7092 66884 7116 66886
rect 7172 66884 7196 66886
rect 7252 66884 7258 66886
rect 6950 66875 7258 66884
rect 6950 65852 7258 65861
rect 6950 65850 6956 65852
rect 7012 65850 7036 65852
rect 7092 65850 7116 65852
rect 7172 65850 7196 65852
rect 7252 65850 7258 65852
rect 7012 65798 7014 65850
rect 7194 65798 7196 65850
rect 6950 65796 6956 65798
rect 7012 65796 7036 65798
rect 7092 65796 7116 65798
rect 7172 65796 7196 65798
rect 7252 65796 7258 65798
rect 6950 65787 7258 65796
rect 6950 64764 7258 64773
rect 6950 64762 6956 64764
rect 7012 64762 7036 64764
rect 7092 64762 7116 64764
rect 7172 64762 7196 64764
rect 7252 64762 7258 64764
rect 7012 64710 7014 64762
rect 7194 64710 7196 64762
rect 6950 64708 6956 64710
rect 7012 64708 7036 64710
rect 7092 64708 7116 64710
rect 7172 64708 7196 64710
rect 7252 64708 7258 64710
rect 6950 64699 7258 64708
rect 7300 64462 7328 69720
rect 7288 64456 7340 64462
rect 7288 64398 7340 64404
rect 6950 63676 7258 63685
rect 6950 63674 6956 63676
rect 7012 63674 7036 63676
rect 7092 63674 7116 63676
rect 7172 63674 7196 63676
rect 7252 63674 7258 63676
rect 7012 63622 7014 63674
rect 7194 63622 7196 63674
rect 6950 63620 6956 63622
rect 7012 63620 7036 63622
rect 7092 63620 7116 63622
rect 7172 63620 7196 63622
rect 7252 63620 7258 63622
rect 6950 63611 7258 63620
rect 7300 63510 7328 64398
rect 7288 63504 7340 63510
rect 7288 63446 7340 63452
rect 6950 62588 7258 62597
rect 6950 62586 6956 62588
rect 7012 62586 7036 62588
rect 7092 62586 7116 62588
rect 7172 62586 7196 62588
rect 7252 62586 7258 62588
rect 7012 62534 7014 62586
rect 7194 62534 7196 62586
rect 6950 62532 6956 62534
rect 7012 62532 7036 62534
rect 7092 62532 7116 62534
rect 7172 62532 7196 62534
rect 7252 62532 7258 62534
rect 6950 62523 7258 62532
rect 6950 61500 7258 61509
rect 6950 61498 6956 61500
rect 7012 61498 7036 61500
rect 7092 61498 7116 61500
rect 7172 61498 7196 61500
rect 7252 61498 7258 61500
rect 7012 61446 7014 61498
rect 7194 61446 7196 61498
rect 6950 61444 6956 61446
rect 7012 61444 7036 61446
rect 7092 61444 7116 61446
rect 7172 61444 7196 61446
rect 7252 61444 7258 61446
rect 6950 61435 7258 61444
rect 6950 60412 7258 60421
rect 6950 60410 6956 60412
rect 7012 60410 7036 60412
rect 7092 60410 7116 60412
rect 7172 60410 7196 60412
rect 7252 60410 7258 60412
rect 7012 60358 7014 60410
rect 7194 60358 7196 60410
rect 6950 60356 6956 60358
rect 7012 60356 7036 60358
rect 7092 60356 7116 60358
rect 7172 60356 7196 60358
rect 7252 60356 7258 60358
rect 6950 60347 7258 60356
rect 7196 60172 7248 60178
rect 7196 60114 7248 60120
rect 6828 60036 6880 60042
rect 6828 59978 6880 59984
rect 7208 59702 7236 60114
rect 7288 59968 7340 59974
rect 7288 59910 7340 59916
rect 7196 59696 7248 59702
rect 7196 59638 7248 59644
rect 6950 59324 7258 59333
rect 6950 59322 6956 59324
rect 7012 59322 7036 59324
rect 7092 59322 7116 59324
rect 7172 59322 7196 59324
rect 7252 59322 7258 59324
rect 7012 59270 7014 59322
rect 7194 59270 7196 59322
rect 6950 59268 6956 59270
rect 7012 59268 7036 59270
rect 7092 59268 7116 59270
rect 7172 59268 7196 59270
rect 7252 59268 7258 59270
rect 6950 59259 7258 59268
rect 6950 58236 7258 58245
rect 6950 58234 6956 58236
rect 7012 58234 7036 58236
rect 7092 58234 7116 58236
rect 7172 58234 7196 58236
rect 7252 58234 7258 58236
rect 7012 58182 7014 58234
rect 7194 58182 7196 58234
rect 6950 58180 6956 58182
rect 7012 58180 7036 58182
rect 7092 58180 7116 58182
rect 7172 58180 7196 58182
rect 7252 58180 7258 58182
rect 6950 58171 7258 58180
rect 6950 57148 7258 57157
rect 6950 57146 6956 57148
rect 7012 57146 7036 57148
rect 7092 57146 7116 57148
rect 7172 57146 7196 57148
rect 7252 57146 7258 57148
rect 7012 57094 7014 57146
rect 7194 57094 7196 57146
rect 6950 57092 6956 57094
rect 7012 57092 7036 57094
rect 7092 57092 7116 57094
rect 7172 57092 7196 57094
rect 7252 57092 7258 57094
rect 6950 57083 7258 57092
rect 6950 56060 7258 56069
rect 6950 56058 6956 56060
rect 7012 56058 7036 56060
rect 7092 56058 7116 56060
rect 7172 56058 7196 56060
rect 7252 56058 7258 56060
rect 7012 56006 7014 56058
rect 7194 56006 7196 56058
rect 6950 56004 6956 56006
rect 7012 56004 7036 56006
rect 7092 56004 7116 56006
rect 7172 56004 7196 56006
rect 7252 56004 7258 56006
rect 6950 55995 7258 56004
rect 6950 54972 7258 54981
rect 6950 54970 6956 54972
rect 7012 54970 7036 54972
rect 7092 54970 7116 54972
rect 7172 54970 7196 54972
rect 7252 54970 7258 54972
rect 7012 54918 7014 54970
rect 7194 54918 7196 54970
rect 6950 54916 6956 54918
rect 7012 54916 7036 54918
rect 7092 54916 7116 54918
rect 7172 54916 7196 54918
rect 7252 54916 7258 54918
rect 6950 54907 7258 54916
rect 6950 53884 7258 53893
rect 6950 53882 6956 53884
rect 7012 53882 7036 53884
rect 7092 53882 7116 53884
rect 7172 53882 7196 53884
rect 7252 53882 7258 53884
rect 7012 53830 7014 53882
rect 7194 53830 7196 53882
rect 6950 53828 6956 53830
rect 7012 53828 7036 53830
rect 7092 53828 7116 53830
rect 7172 53828 7196 53830
rect 7252 53828 7258 53830
rect 6950 53819 7258 53828
rect 6950 52796 7258 52805
rect 6950 52794 6956 52796
rect 7012 52794 7036 52796
rect 7092 52794 7116 52796
rect 7172 52794 7196 52796
rect 7252 52794 7258 52796
rect 7012 52742 7014 52794
rect 7194 52742 7196 52794
rect 6950 52740 6956 52742
rect 7012 52740 7036 52742
rect 7092 52740 7116 52742
rect 7172 52740 7196 52742
rect 7252 52740 7258 52742
rect 6950 52731 7258 52740
rect 6920 52692 6972 52698
rect 6920 52634 6972 52640
rect 6932 51898 6960 52634
rect 6840 51870 6960 51898
rect 6840 51490 6868 51870
rect 6950 51708 7258 51717
rect 6950 51706 6956 51708
rect 7012 51706 7036 51708
rect 7092 51706 7116 51708
rect 7172 51706 7196 51708
rect 7252 51706 7258 51708
rect 7012 51654 7014 51706
rect 7194 51654 7196 51706
rect 6950 51652 6956 51654
rect 7012 51652 7036 51654
rect 7092 51652 7116 51654
rect 7172 51652 7196 51654
rect 7252 51652 7258 51654
rect 6950 51643 7258 51652
rect 6840 51462 6960 51490
rect 6748 51046 6868 51074
rect 6656 48606 6776 48634
rect 6644 48544 6696 48550
rect 6644 48486 6696 48492
rect 6656 48346 6684 48486
rect 6644 48340 6696 48346
rect 6644 48282 6696 48288
rect 6748 48226 6776 48606
rect 6656 48198 6776 48226
rect 6656 41414 6684 48198
rect 6736 43648 6788 43654
rect 6736 43590 6788 43596
rect 6748 42945 6776 43590
rect 6734 42936 6790 42945
rect 6734 42871 6790 42880
rect 6736 42832 6788 42838
rect 6736 42774 6788 42780
rect 6748 41614 6776 42774
rect 6736 41608 6788 41614
rect 6736 41550 6788 41556
rect 6656 41386 6776 41414
rect 6644 40384 6696 40390
rect 6644 40326 6696 40332
rect 6656 38554 6684 40326
rect 6644 38548 6696 38554
rect 6644 38490 6696 38496
rect 6644 36644 6696 36650
rect 6644 36586 6696 36592
rect 6656 36378 6684 36586
rect 6644 36372 6696 36378
rect 6644 36314 6696 36320
rect 6644 33312 6696 33318
rect 6644 33254 6696 33260
rect 6656 32314 6684 33254
rect 6748 33114 6776 41386
rect 6840 40050 6868 51046
rect 6932 50833 6960 51462
rect 6918 50824 6974 50833
rect 6918 50759 6974 50768
rect 6950 50620 7258 50629
rect 6950 50618 6956 50620
rect 7012 50618 7036 50620
rect 7092 50618 7116 50620
rect 7172 50618 7196 50620
rect 7252 50618 7258 50620
rect 7012 50566 7014 50618
rect 7194 50566 7196 50618
rect 6950 50564 6956 50566
rect 7012 50564 7036 50566
rect 7092 50564 7116 50566
rect 7172 50564 7196 50566
rect 7252 50564 7258 50566
rect 6950 50555 7258 50564
rect 6950 49532 7258 49541
rect 6950 49530 6956 49532
rect 7012 49530 7036 49532
rect 7092 49530 7116 49532
rect 7172 49530 7196 49532
rect 7252 49530 7258 49532
rect 7012 49478 7014 49530
rect 7194 49478 7196 49530
rect 6950 49476 6956 49478
rect 7012 49476 7036 49478
rect 7092 49476 7116 49478
rect 7172 49476 7196 49478
rect 7252 49476 7258 49478
rect 6950 49467 7258 49476
rect 6950 48444 7258 48453
rect 6950 48442 6956 48444
rect 7012 48442 7036 48444
rect 7092 48442 7116 48444
rect 7172 48442 7196 48444
rect 7252 48442 7258 48444
rect 7012 48390 7014 48442
rect 7194 48390 7196 48442
rect 6950 48388 6956 48390
rect 7012 48388 7036 48390
rect 7092 48388 7116 48390
rect 7172 48388 7196 48390
rect 7252 48388 7258 48390
rect 6950 48379 7258 48388
rect 6950 47356 7258 47365
rect 6950 47354 6956 47356
rect 7012 47354 7036 47356
rect 7092 47354 7116 47356
rect 7172 47354 7196 47356
rect 7252 47354 7258 47356
rect 7012 47302 7014 47354
rect 7194 47302 7196 47354
rect 6950 47300 6956 47302
rect 7012 47300 7036 47302
rect 7092 47300 7116 47302
rect 7172 47300 7196 47302
rect 7252 47300 7258 47302
rect 6950 47291 7258 47300
rect 6950 46268 7258 46277
rect 6950 46266 6956 46268
rect 7012 46266 7036 46268
rect 7092 46266 7116 46268
rect 7172 46266 7196 46268
rect 7252 46266 7258 46268
rect 7012 46214 7014 46266
rect 7194 46214 7196 46266
rect 6950 46212 6956 46214
rect 7012 46212 7036 46214
rect 7092 46212 7116 46214
rect 7172 46212 7196 46214
rect 7252 46212 7258 46214
rect 6950 46203 7258 46212
rect 7300 46170 7328 59910
rect 7392 54194 7420 72558
rect 7610 71836 7918 71845
rect 7610 71834 7616 71836
rect 7672 71834 7696 71836
rect 7752 71834 7776 71836
rect 7832 71834 7856 71836
rect 7912 71834 7918 71836
rect 7672 71782 7674 71834
rect 7854 71782 7856 71834
rect 7610 71780 7616 71782
rect 7672 71780 7696 71782
rect 7752 71780 7776 71782
rect 7832 71780 7856 71782
rect 7912 71780 7918 71782
rect 7610 71771 7918 71780
rect 7610 70748 7918 70757
rect 7610 70746 7616 70748
rect 7672 70746 7696 70748
rect 7752 70746 7776 70748
rect 7832 70746 7856 70748
rect 7912 70746 7918 70748
rect 7672 70694 7674 70746
rect 7854 70694 7856 70746
rect 7610 70692 7616 70694
rect 7672 70692 7696 70694
rect 7752 70692 7776 70694
rect 7832 70692 7856 70694
rect 7912 70692 7918 70694
rect 7610 70683 7918 70692
rect 7610 69660 7918 69669
rect 7610 69658 7616 69660
rect 7672 69658 7696 69660
rect 7752 69658 7776 69660
rect 7832 69658 7856 69660
rect 7912 69658 7918 69660
rect 7672 69606 7674 69658
rect 7854 69606 7856 69658
rect 7610 69604 7616 69606
rect 7672 69604 7696 69606
rect 7752 69604 7776 69606
rect 7832 69604 7856 69606
rect 7912 69604 7918 69606
rect 7610 69595 7918 69604
rect 7472 69488 7524 69494
rect 7472 69430 7524 69436
rect 7380 54188 7432 54194
rect 7380 54130 7432 54136
rect 7380 54052 7432 54058
rect 7380 53994 7432 54000
rect 7392 48770 7420 53994
rect 7484 48890 7512 69430
rect 7610 68572 7918 68581
rect 7610 68570 7616 68572
rect 7672 68570 7696 68572
rect 7752 68570 7776 68572
rect 7832 68570 7856 68572
rect 7912 68570 7918 68572
rect 7672 68518 7674 68570
rect 7854 68518 7856 68570
rect 7610 68516 7616 68518
rect 7672 68516 7696 68518
rect 7752 68516 7776 68518
rect 7832 68516 7856 68518
rect 7912 68516 7918 68518
rect 7610 68507 7918 68516
rect 7610 67484 7918 67493
rect 7610 67482 7616 67484
rect 7672 67482 7696 67484
rect 7752 67482 7776 67484
rect 7832 67482 7856 67484
rect 7912 67482 7918 67484
rect 7672 67430 7674 67482
rect 7854 67430 7856 67482
rect 7610 67428 7616 67430
rect 7672 67428 7696 67430
rect 7752 67428 7776 67430
rect 7832 67428 7856 67430
rect 7912 67428 7918 67430
rect 7610 67419 7918 67428
rect 7610 66396 7918 66405
rect 7610 66394 7616 66396
rect 7672 66394 7696 66396
rect 7752 66394 7776 66396
rect 7832 66394 7856 66396
rect 7912 66394 7918 66396
rect 7672 66342 7674 66394
rect 7854 66342 7856 66394
rect 7610 66340 7616 66342
rect 7672 66340 7696 66342
rect 7752 66340 7776 66342
rect 7832 66340 7856 66342
rect 7912 66340 7918 66342
rect 7610 66331 7918 66340
rect 7610 65308 7918 65317
rect 7610 65306 7616 65308
rect 7672 65306 7696 65308
rect 7752 65306 7776 65308
rect 7832 65306 7856 65308
rect 7912 65306 7918 65308
rect 7672 65254 7674 65306
rect 7854 65254 7856 65306
rect 7610 65252 7616 65254
rect 7672 65252 7696 65254
rect 7752 65252 7776 65254
rect 7832 65252 7856 65254
rect 7912 65252 7918 65254
rect 7610 65243 7918 65252
rect 7932 65068 7984 65074
rect 7932 65010 7984 65016
rect 7944 64326 7972 65010
rect 7932 64320 7984 64326
rect 7932 64262 7984 64268
rect 7610 64220 7918 64229
rect 7610 64218 7616 64220
rect 7672 64218 7696 64220
rect 7752 64218 7776 64220
rect 7832 64218 7856 64220
rect 7912 64218 7918 64220
rect 7672 64166 7674 64218
rect 7854 64166 7856 64218
rect 7610 64164 7616 64166
rect 7672 64164 7696 64166
rect 7752 64164 7776 64166
rect 7832 64164 7856 64166
rect 7912 64164 7918 64166
rect 7610 64155 7918 64164
rect 7610 63132 7918 63141
rect 7610 63130 7616 63132
rect 7672 63130 7696 63132
rect 7752 63130 7776 63132
rect 7832 63130 7856 63132
rect 7912 63130 7918 63132
rect 7672 63078 7674 63130
rect 7854 63078 7856 63130
rect 7610 63076 7616 63078
rect 7672 63076 7696 63078
rect 7752 63076 7776 63078
rect 7832 63076 7856 63078
rect 7912 63076 7918 63078
rect 7610 63067 7918 63076
rect 7610 62044 7918 62053
rect 7610 62042 7616 62044
rect 7672 62042 7696 62044
rect 7752 62042 7776 62044
rect 7832 62042 7856 62044
rect 7912 62042 7918 62044
rect 7672 61990 7674 62042
rect 7854 61990 7856 62042
rect 7610 61988 7616 61990
rect 7672 61988 7696 61990
rect 7752 61988 7776 61990
rect 7832 61988 7856 61990
rect 7912 61988 7918 61990
rect 7610 61979 7918 61988
rect 7610 60956 7918 60965
rect 7610 60954 7616 60956
rect 7672 60954 7696 60956
rect 7752 60954 7776 60956
rect 7832 60954 7856 60956
rect 7912 60954 7918 60956
rect 7672 60902 7674 60954
rect 7854 60902 7856 60954
rect 7610 60900 7616 60902
rect 7672 60900 7696 60902
rect 7752 60900 7776 60902
rect 7832 60900 7856 60902
rect 7912 60900 7918 60902
rect 7610 60891 7918 60900
rect 8036 60602 8064 76214
rect 8116 75336 8168 75342
rect 8116 75278 8168 75284
rect 8128 75002 8156 75278
rect 8116 74996 8168 75002
rect 8116 74938 8168 74944
rect 8220 73710 8248 76366
rect 14660 76362 14688 76735
rect 16500 76634 16528 76774
rect 16488 76628 16540 76634
rect 16488 76570 16540 76576
rect 14924 76424 14976 76430
rect 14924 76366 14976 76372
rect 8482 76327 8484 76336
rect 8536 76327 8538 76336
rect 14648 76356 14700 76362
rect 8484 76298 8536 76304
rect 14648 76298 14700 76304
rect 8944 76288 8996 76294
rect 11244 76288 11296 76294
rect 8944 76230 8996 76236
rect 11242 76256 11244 76265
rect 11704 76288 11756 76294
rect 11296 76256 11298 76265
rect 8758 76120 8814 76129
rect 8758 76055 8814 76064
rect 8772 76022 8800 76055
rect 8760 76016 8812 76022
rect 8760 75958 8812 75964
rect 8208 73704 8260 73710
rect 8208 73646 8260 73652
rect 8116 73024 8168 73030
rect 8116 72966 8168 72972
rect 8128 64530 8156 72966
rect 8220 72758 8248 73646
rect 8208 72752 8260 72758
rect 8208 72694 8260 72700
rect 8208 71392 8260 71398
rect 8208 71334 8260 71340
rect 8116 64524 8168 64530
rect 8116 64466 8168 64472
rect 8116 64320 8168 64326
rect 8116 64262 8168 64268
rect 7944 60574 8064 60602
rect 7944 60518 7972 60574
rect 7932 60512 7984 60518
rect 7932 60454 7984 60460
rect 8024 60512 8076 60518
rect 8024 60454 8076 60460
rect 7944 60194 7972 60454
rect 8036 60314 8064 60454
rect 8024 60308 8076 60314
rect 8024 60250 8076 60256
rect 7944 60166 8064 60194
rect 8128 60178 8156 64262
rect 7610 59868 7918 59877
rect 7610 59866 7616 59868
rect 7672 59866 7696 59868
rect 7752 59866 7776 59868
rect 7832 59866 7856 59868
rect 7912 59866 7918 59868
rect 7672 59814 7674 59866
rect 7854 59814 7856 59866
rect 7610 59812 7616 59814
rect 7672 59812 7696 59814
rect 7752 59812 7776 59814
rect 7832 59812 7856 59814
rect 7912 59812 7918 59814
rect 7610 59803 7918 59812
rect 7610 58780 7918 58789
rect 7610 58778 7616 58780
rect 7672 58778 7696 58780
rect 7752 58778 7776 58780
rect 7832 58778 7856 58780
rect 7912 58778 7918 58780
rect 7672 58726 7674 58778
rect 7854 58726 7856 58778
rect 7610 58724 7616 58726
rect 7672 58724 7696 58726
rect 7752 58724 7776 58726
rect 7832 58724 7856 58726
rect 7912 58724 7918 58726
rect 7610 58715 7918 58724
rect 7610 57692 7918 57701
rect 7610 57690 7616 57692
rect 7672 57690 7696 57692
rect 7752 57690 7776 57692
rect 7832 57690 7856 57692
rect 7912 57690 7918 57692
rect 7672 57638 7674 57690
rect 7854 57638 7856 57690
rect 7610 57636 7616 57638
rect 7672 57636 7696 57638
rect 7752 57636 7776 57638
rect 7832 57636 7856 57638
rect 7912 57636 7918 57638
rect 7610 57627 7918 57636
rect 7610 56604 7918 56613
rect 7610 56602 7616 56604
rect 7672 56602 7696 56604
rect 7752 56602 7776 56604
rect 7832 56602 7856 56604
rect 7912 56602 7918 56604
rect 7672 56550 7674 56602
rect 7854 56550 7856 56602
rect 7610 56548 7616 56550
rect 7672 56548 7696 56550
rect 7752 56548 7776 56550
rect 7832 56548 7856 56550
rect 7912 56548 7918 56550
rect 7610 56539 7918 56548
rect 7610 55516 7918 55525
rect 7610 55514 7616 55516
rect 7672 55514 7696 55516
rect 7752 55514 7776 55516
rect 7832 55514 7856 55516
rect 7912 55514 7918 55516
rect 7672 55462 7674 55514
rect 7854 55462 7856 55514
rect 7610 55460 7616 55462
rect 7672 55460 7696 55462
rect 7752 55460 7776 55462
rect 7832 55460 7856 55462
rect 7912 55460 7918 55462
rect 7610 55451 7918 55460
rect 7610 54428 7918 54437
rect 7610 54426 7616 54428
rect 7672 54426 7696 54428
rect 7752 54426 7776 54428
rect 7832 54426 7856 54428
rect 7912 54426 7918 54428
rect 7672 54374 7674 54426
rect 7854 54374 7856 54426
rect 7610 54372 7616 54374
rect 7672 54372 7696 54374
rect 7752 54372 7776 54374
rect 7832 54372 7856 54374
rect 7912 54372 7918 54374
rect 7610 54363 7918 54372
rect 7610 53340 7918 53349
rect 7610 53338 7616 53340
rect 7672 53338 7696 53340
rect 7752 53338 7776 53340
rect 7832 53338 7856 53340
rect 7912 53338 7918 53340
rect 7672 53286 7674 53338
rect 7854 53286 7856 53338
rect 7610 53284 7616 53286
rect 7672 53284 7696 53286
rect 7752 53284 7776 53286
rect 7832 53284 7856 53286
rect 7912 53284 7918 53286
rect 7610 53275 7918 53284
rect 7840 53236 7892 53242
rect 7840 53178 7892 53184
rect 7852 52698 7880 53178
rect 8036 52902 8064 60166
rect 8116 60172 8168 60178
rect 8116 60114 8168 60120
rect 8116 60036 8168 60042
rect 8220 60024 8248 71334
rect 8300 69896 8352 69902
rect 8300 69838 8352 69844
rect 8312 65210 8340 69838
rect 8300 65204 8352 65210
rect 8300 65146 8352 65152
rect 8668 65068 8720 65074
rect 8668 65010 8720 65016
rect 8300 64932 8352 64938
rect 8300 64874 8352 64880
rect 8168 59996 8248 60024
rect 8116 59978 8168 59984
rect 8128 59945 8156 59978
rect 8114 59936 8170 59945
rect 8114 59871 8170 59880
rect 8312 59786 8340 64874
rect 8392 64524 8444 64530
rect 8392 64466 8444 64472
rect 8128 59758 8340 59786
rect 8128 57798 8156 59758
rect 8208 59696 8260 59702
rect 8208 59638 8260 59644
rect 8116 57792 8168 57798
rect 8116 57734 8168 57740
rect 8116 57588 8168 57594
rect 8116 57530 8168 57536
rect 8128 56370 8156 57530
rect 8116 56364 8168 56370
rect 8116 56306 8168 56312
rect 8128 54330 8156 56306
rect 8116 54324 8168 54330
rect 8116 54266 8168 54272
rect 8116 54188 8168 54194
rect 8116 54130 8168 54136
rect 8024 52896 8076 52902
rect 8024 52838 8076 52844
rect 7840 52692 7892 52698
rect 7840 52634 7892 52640
rect 7610 52252 7918 52261
rect 7610 52250 7616 52252
rect 7672 52250 7696 52252
rect 7752 52250 7776 52252
rect 7832 52250 7856 52252
rect 7912 52250 7918 52252
rect 7672 52198 7674 52250
rect 7854 52198 7856 52250
rect 7610 52196 7616 52198
rect 7672 52196 7696 52198
rect 7752 52196 7776 52198
rect 7832 52196 7856 52198
rect 7912 52196 7918 52198
rect 7610 52187 7918 52196
rect 7838 51912 7894 51921
rect 7838 51847 7894 51856
rect 7852 51610 7880 51847
rect 7840 51604 7892 51610
rect 7840 51546 7892 51552
rect 7610 51164 7918 51173
rect 7610 51162 7616 51164
rect 7672 51162 7696 51164
rect 7752 51162 7776 51164
rect 7832 51162 7856 51164
rect 7912 51162 7918 51164
rect 7672 51110 7674 51162
rect 7854 51110 7856 51162
rect 7610 51108 7616 51110
rect 7672 51108 7696 51110
rect 7752 51108 7776 51110
rect 7832 51108 7856 51110
rect 7912 51108 7918 51110
rect 7610 51099 7918 51108
rect 8024 50992 8076 50998
rect 8128 50946 8156 54130
rect 8076 50940 8156 50946
rect 8024 50934 8156 50940
rect 8036 50918 8156 50934
rect 8024 50856 8076 50862
rect 7562 50824 7618 50833
rect 8024 50798 8076 50804
rect 7562 50759 7618 50768
rect 7576 50182 7604 50759
rect 7564 50176 7616 50182
rect 7564 50118 7616 50124
rect 7610 50076 7918 50085
rect 7610 50074 7616 50076
rect 7672 50074 7696 50076
rect 7752 50074 7776 50076
rect 7832 50074 7856 50076
rect 7912 50074 7918 50076
rect 7672 50022 7674 50074
rect 7854 50022 7856 50074
rect 7610 50020 7616 50022
rect 7672 50020 7696 50022
rect 7752 50020 7776 50022
rect 7832 50020 7856 50022
rect 7912 50020 7918 50022
rect 7610 50011 7918 50020
rect 8036 49774 8064 50798
rect 8116 50788 8168 50794
rect 8116 50730 8168 50736
rect 8024 49768 8076 49774
rect 8024 49710 8076 49716
rect 8036 49230 8064 49710
rect 8024 49224 8076 49230
rect 8024 49166 8076 49172
rect 8024 49088 8076 49094
rect 8024 49030 8076 49036
rect 7610 48988 7918 48997
rect 7610 48986 7616 48988
rect 7672 48986 7696 48988
rect 7752 48986 7776 48988
rect 7832 48986 7856 48988
rect 7912 48986 7918 48988
rect 7672 48934 7674 48986
rect 7854 48934 7856 48986
rect 7610 48932 7616 48934
rect 7672 48932 7696 48934
rect 7752 48932 7776 48934
rect 7832 48932 7856 48934
rect 7912 48932 7918 48934
rect 7610 48923 7918 48932
rect 7472 48884 7524 48890
rect 7472 48826 7524 48832
rect 7392 48742 7512 48770
rect 7484 47666 7512 48742
rect 7610 47900 7918 47909
rect 7610 47898 7616 47900
rect 7672 47898 7696 47900
rect 7752 47898 7776 47900
rect 7832 47898 7856 47900
rect 7912 47898 7918 47900
rect 7672 47846 7674 47898
rect 7854 47846 7856 47898
rect 7610 47844 7616 47846
rect 7672 47844 7696 47846
rect 7752 47844 7776 47846
rect 7832 47844 7856 47846
rect 7912 47844 7918 47846
rect 7610 47835 7918 47844
rect 7656 47796 7708 47802
rect 7656 47738 7708 47744
rect 7380 47660 7432 47666
rect 7380 47602 7432 47608
rect 7472 47660 7524 47666
rect 7472 47602 7524 47608
rect 7288 46164 7340 46170
rect 7288 46106 7340 46112
rect 7288 45620 7340 45626
rect 7288 45562 7340 45568
rect 6950 45180 7258 45189
rect 6950 45178 6956 45180
rect 7012 45178 7036 45180
rect 7092 45178 7116 45180
rect 7172 45178 7196 45180
rect 7252 45178 7258 45180
rect 7012 45126 7014 45178
rect 7194 45126 7196 45178
rect 6950 45124 6956 45126
rect 7012 45124 7036 45126
rect 7092 45124 7116 45126
rect 7172 45124 7196 45126
rect 7252 45124 7258 45126
rect 6950 45115 7258 45124
rect 7300 44470 7328 45562
rect 7288 44464 7340 44470
rect 7288 44406 7340 44412
rect 6950 44092 7258 44101
rect 6950 44090 6956 44092
rect 7012 44090 7036 44092
rect 7092 44090 7116 44092
rect 7172 44090 7196 44092
rect 7252 44090 7258 44092
rect 7012 44038 7014 44090
rect 7194 44038 7196 44090
rect 6950 44036 6956 44038
rect 7012 44036 7036 44038
rect 7092 44036 7116 44038
rect 7172 44036 7196 44038
rect 7252 44036 7258 44038
rect 6950 44027 7258 44036
rect 6950 43004 7258 43013
rect 6950 43002 6956 43004
rect 7012 43002 7036 43004
rect 7092 43002 7116 43004
rect 7172 43002 7196 43004
rect 7252 43002 7258 43004
rect 7012 42950 7014 43002
rect 7194 42950 7196 43002
rect 6950 42948 6956 42950
rect 7012 42948 7036 42950
rect 7092 42948 7116 42950
rect 7172 42948 7196 42950
rect 7252 42948 7258 42950
rect 6950 42939 7258 42948
rect 7300 42226 7328 44406
rect 7288 42220 7340 42226
rect 7288 42162 7340 42168
rect 6950 41916 7258 41925
rect 6950 41914 6956 41916
rect 7012 41914 7036 41916
rect 7092 41914 7116 41916
rect 7172 41914 7196 41916
rect 7252 41914 7258 41916
rect 7012 41862 7014 41914
rect 7194 41862 7196 41914
rect 6950 41860 6956 41862
rect 7012 41860 7036 41862
rect 7092 41860 7116 41862
rect 7172 41860 7196 41862
rect 7252 41860 7258 41862
rect 6950 41851 7258 41860
rect 7196 41812 7248 41818
rect 7196 41754 7248 41760
rect 7208 40934 7236 41754
rect 7196 40928 7248 40934
rect 7196 40870 7248 40876
rect 6950 40828 7258 40837
rect 6950 40826 6956 40828
rect 7012 40826 7036 40828
rect 7092 40826 7116 40828
rect 7172 40826 7196 40828
rect 7252 40826 7258 40828
rect 7012 40774 7014 40826
rect 7194 40774 7196 40826
rect 6950 40772 6956 40774
rect 7012 40772 7036 40774
rect 7092 40772 7116 40774
rect 7172 40772 7196 40774
rect 7252 40772 7258 40774
rect 6950 40763 7258 40772
rect 6828 40044 6880 40050
rect 6828 39986 6880 39992
rect 7300 39914 7328 42162
rect 7392 41818 7420 47602
rect 7564 47524 7616 47530
rect 7564 47466 7616 47472
rect 7576 47002 7604 47466
rect 7484 46974 7604 47002
rect 7668 46986 7696 47738
rect 7748 47660 7800 47666
rect 7748 47602 7800 47608
rect 7760 47054 7788 47602
rect 7748 47048 7800 47054
rect 7748 46990 7800 46996
rect 7656 46980 7708 46986
rect 7484 42770 7512 46974
rect 7656 46922 7708 46928
rect 7610 46812 7918 46821
rect 7610 46810 7616 46812
rect 7672 46810 7696 46812
rect 7752 46810 7776 46812
rect 7832 46810 7856 46812
rect 7912 46810 7918 46812
rect 7672 46758 7674 46810
rect 7854 46758 7856 46810
rect 7610 46756 7616 46758
rect 7672 46756 7696 46758
rect 7752 46756 7776 46758
rect 7832 46756 7856 46758
rect 7912 46756 7918 46758
rect 7610 46747 7918 46756
rect 8036 46374 8064 49030
rect 8024 46368 8076 46374
rect 8024 46310 8076 46316
rect 8024 46164 8076 46170
rect 8024 46106 8076 46112
rect 7610 45724 7918 45733
rect 7610 45722 7616 45724
rect 7672 45722 7696 45724
rect 7752 45722 7776 45724
rect 7832 45722 7856 45724
rect 7912 45722 7918 45724
rect 7672 45670 7674 45722
rect 7854 45670 7856 45722
rect 7610 45668 7616 45670
rect 7672 45668 7696 45670
rect 7752 45668 7776 45670
rect 7832 45668 7856 45670
rect 7912 45668 7918 45670
rect 7610 45659 7918 45668
rect 7610 44636 7918 44645
rect 7610 44634 7616 44636
rect 7672 44634 7696 44636
rect 7752 44634 7776 44636
rect 7832 44634 7856 44636
rect 7912 44634 7918 44636
rect 7672 44582 7674 44634
rect 7854 44582 7856 44634
rect 7610 44580 7616 44582
rect 7672 44580 7696 44582
rect 7752 44580 7776 44582
rect 7832 44580 7856 44582
rect 7912 44580 7918 44582
rect 7610 44571 7918 44580
rect 7610 43548 7918 43557
rect 7610 43546 7616 43548
rect 7672 43546 7696 43548
rect 7752 43546 7776 43548
rect 7832 43546 7856 43548
rect 7912 43546 7918 43548
rect 7672 43494 7674 43546
rect 7854 43494 7856 43546
rect 7610 43492 7616 43494
rect 7672 43492 7696 43494
rect 7752 43492 7776 43494
rect 7832 43492 7856 43494
rect 7912 43492 7918 43494
rect 7610 43483 7918 43492
rect 7562 43344 7618 43353
rect 7562 43279 7618 43288
rect 7472 42764 7524 42770
rect 7472 42706 7524 42712
rect 7576 42650 7604 43279
rect 7484 42622 7604 42650
rect 7380 41812 7432 41818
rect 7380 41754 7432 41760
rect 7484 41698 7512 42622
rect 7610 42460 7918 42469
rect 7610 42458 7616 42460
rect 7672 42458 7696 42460
rect 7752 42458 7776 42460
rect 7832 42458 7856 42460
rect 7912 42458 7918 42460
rect 7672 42406 7674 42458
rect 7854 42406 7856 42458
rect 7610 42404 7616 42406
rect 7672 42404 7696 42406
rect 7752 42404 7776 42406
rect 7832 42404 7856 42406
rect 7912 42404 7918 42406
rect 7610 42395 7918 42404
rect 7392 41670 7512 41698
rect 7288 39908 7340 39914
rect 7288 39850 7340 39856
rect 6950 39740 7258 39749
rect 6950 39738 6956 39740
rect 7012 39738 7036 39740
rect 7092 39738 7116 39740
rect 7172 39738 7196 39740
rect 7252 39738 7258 39740
rect 7012 39686 7014 39738
rect 7194 39686 7196 39738
rect 6950 39684 6956 39686
rect 7012 39684 7036 39686
rect 7092 39684 7116 39686
rect 7172 39684 7196 39686
rect 7252 39684 7258 39686
rect 6950 39675 7258 39684
rect 7300 38826 7328 39850
rect 7288 38820 7340 38826
rect 7288 38762 7340 38768
rect 6828 38752 6880 38758
rect 6828 38694 6880 38700
rect 6840 35834 6868 38694
rect 6950 38652 7258 38661
rect 6950 38650 6956 38652
rect 7012 38650 7036 38652
rect 7092 38650 7116 38652
rect 7172 38650 7196 38652
rect 7252 38650 7258 38652
rect 7012 38598 7014 38650
rect 7194 38598 7196 38650
rect 6950 38596 6956 38598
rect 7012 38596 7036 38598
rect 7092 38596 7116 38598
rect 7172 38596 7196 38598
rect 7252 38596 7258 38598
rect 6950 38587 7258 38596
rect 7288 38548 7340 38554
rect 7288 38490 7340 38496
rect 6950 37564 7258 37573
rect 6950 37562 6956 37564
rect 7012 37562 7036 37564
rect 7092 37562 7116 37564
rect 7172 37562 7196 37564
rect 7252 37562 7258 37564
rect 7012 37510 7014 37562
rect 7194 37510 7196 37562
rect 6950 37508 6956 37510
rect 7012 37508 7036 37510
rect 7092 37508 7116 37510
rect 7172 37508 7196 37510
rect 7252 37508 7258 37510
rect 6950 37499 7258 37508
rect 6950 36476 7258 36485
rect 6950 36474 6956 36476
rect 7012 36474 7036 36476
rect 7092 36474 7116 36476
rect 7172 36474 7196 36476
rect 7252 36474 7258 36476
rect 7012 36422 7014 36474
rect 7194 36422 7196 36474
rect 6950 36420 6956 36422
rect 7012 36420 7036 36422
rect 7092 36420 7116 36422
rect 7172 36420 7196 36422
rect 7252 36420 7258 36422
rect 6950 36411 7258 36420
rect 6828 35828 6880 35834
rect 6828 35770 6880 35776
rect 6950 35388 7258 35397
rect 6950 35386 6956 35388
rect 7012 35386 7036 35388
rect 7092 35386 7116 35388
rect 7172 35386 7196 35388
rect 7252 35386 7258 35388
rect 7012 35334 7014 35386
rect 7194 35334 7196 35386
rect 6950 35332 6956 35334
rect 7012 35332 7036 35334
rect 7092 35332 7116 35334
rect 7172 35332 7196 35334
rect 7252 35332 7258 35334
rect 6950 35323 7258 35332
rect 7300 35170 7328 38490
rect 7208 35142 7328 35170
rect 7208 34490 7236 35142
rect 6840 34462 7236 34490
rect 7288 34536 7340 34542
rect 7288 34478 7340 34484
rect 6840 34082 6868 34462
rect 7300 34406 7328 34478
rect 7288 34400 7340 34406
rect 7288 34342 7340 34348
rect 6950 34300 7258 34309
rect 6950 34298 6956 34300
rect 7012 34298 7036 34300
rect 7092 34298 7116 34300
rect 7172 34298 7196 34300
rect 7252 34298 7258 34300
rect 7012 34246 7014 34298
rect 7194 34246 7196 34298
rect 6950 34244 6956 34246
rect 7012 34244 7036 34246
rect 7092 34244 7116 34246
rect 7172 34244 7196 34246
rect 7252 34244 7258 34246
rect 6950 34235 7258 34244
rect 6840 34054 6960 34082
rect 6932 33402 6960 34054
rect 7012 33924 7064 33930
rect 7012 33866 7064 33872
rect 6840 33374 6960 33402
rect 6736 33108 6788 33114
rect 6736 33050 6788 33056
rect 6840 32994 6868 33374
rect 7024 33318 7052 33866
rect 7012 33312 7064 33318
rect 7012 33254 7064 33260
rect 6950 33212 7258 33221
rect 6950 33210 6956 33212
rect 7012 33210 7036 33212
rect 7092 33210 7116 33212
rect 7172 33210 7196 33212
rect 7252 33210 7258 33212
rect 7012 33158 7014 33210
rect 7194 33158 7196 33210
rect 6950 33156 6956 33158
rect 7012 33156 7036 33158
rect 7092 33156 7116 33158
rect 7172 33156 7196 33158
rect 7252 33156 7258 33158
rect 6950 33147 7258 33156
rect 6840 32966 6960 32994
rect 6656 32286 6868 32314
rect 6736 32224 6788 32230
rect 6736 32166 6788 32172
rect 6644 30048 6696 30054
rect 6644 29990 6696 29996
rect 6656 29782 6684 29990
rect 6644 29776 6696 29782
rect 6644 29718 6696 29724
rect 6748 24818 6776 32166
rect 6840 31906 6868 32286
rect 6932 32230 6960 32966
rect 7300 32366 7328 34342
rect 7288 32360 7340 32366
rect 7288 32302 7340 32308
rect 6920 32224 6972 32230
rect 6920 32166 6972 32172
rect 7288 32224 7340 32230
rect 7288 32166 7340 32172
rect 6950 32124 7258 32133
rect 6950 32122 6956 32124
rect 7012 32122 7036 32124
rect 7092 32122 7116 32124
rect 7172 32122 7196 32124
rect 7252 32122 7258 32124
rect 7012 32070 7014 32122
rect 7194 32070 7196 32122
rect 6950 32068 6956 32070
rect 7012 32068 7036 32070
rect 7092 32068 7116 32070
rect 7172 32068 7196 32070
rect 7252 32068 7258 32070
rect 6950 32059 7258 32068
rect 6840 31878 6960 31906
rect 6932 31754 6960 31878
rect 6932 31726 7236 31754
rect 6920 31680 6972 31686
rect 6920 31622 6972 31628
rect 6932 31482 6960 31622
rect 6920 31476 6972 31482
rect 6920 31418 6972 31424
rect 7208 31226 7236 31726
rect 7300 31346 7328 32166
rect 7392 31346 7420 41670
rect 7472 41608 7524 41614
rect 7472 41550 7524 41556
rect 7484 32570 7512 41550
rect 7610 41372 7918 41381
rect 7610 41370 7616 41372
rect 7672 41370 7696 41372
rect 7752 41370 7776 41372
rect 7832 41370 7856 41372
rect 7912 41370 7918 41372
rect 7672 41318 7674 41370
rect 7854 41318 7856 41370
rect 7610 41316 7616 41318
rect 7672 41316 7696 41318
rect 7752 41316 7776 41318
rect 7832 41316 7856 41318
rect 7912 41316 7918 41318
rect 7610 41307 7918 41316
rect 7656 40928 7708 40934
rect 7656 40870 7708 40876
rect 7668 40390 7696 40870
rect 7656 40384 7708 40390
rect 7656 40326 7708 40332
rect 7610 40284 7918 40293
rect 7610 40282 7616 40284
rect 7672 40282 7696 40284
rect 7752 40282 7776 40284
rect 7832 40282 7856 40284
rect 7912 40282 7918 40284
rect 7672 40230 7674 40282
rect 7854 40230 7856 40282
rect 7610 40228 7616 40230
rect 7672 40228 7696 40230
rect 7752 40228 7776 40230
rect 7832 40228 7856 40230
rect 7912 40228 7918 40230
rect 7610 40219 7918 40228
rect 7610 39196 7918 39205
rect 7610 39194 7616 39196
rect 7672 39194 7696 39196
rect 7752 39194 7776 39196
rect 7832 39194 7856 39196
rect 7912 39194 7918 39196
rect 7672 39142 7674 39194
rect 7854 39142 7856 39194
rect 7610 39140 7616 39142
rect 7672 39140 7696 39142
rect 7752 39140 7776 39142
rect 7832 39140 7856 39142
rect 7912 39140 7918 39142
rect 7610 39131 7918 39140
rect 7610 38108 7918 38117
rect 7610 38106 7616 38108
rect 7672 38106 7696 38108
rect 7752 38106 7776 38108
rect 7832 38106 7856 38108
rect 7912 38106 7918 38108
rect 7672 38054 7674 38106
rect 7854 38054 7856 38106
rect 7610 38052 7616 38054
rect 7672 38052 7696 38054
rect 7752 38052 7776 38054
rect 7832 38052 7856 38054
rect 7912 38052 7918 38054
rect 7610 38043 7918 38052
rect 7610 37020 7918 37029
rect 7610 37018 7616 37020
rect 7672 37018 7696 37020
rect 7752 37018 7776 37020
rect 7832 37018 7856 37020
rect 7912 37018 7918 37020
rect 7672 36966 7674 37018
rect 7854 36966 7856 37018
rect 7610 36964 7616 36966
rect 7672 36964 7696 36966
rect 7752 36964 7776 36966
rect 7832 36964 7856 36966
rect 7912 36964 7918 36966
rect 7610 36955 7918 36964
rect 7610 35932 7918 35941
rect 7610 35930 7616 35932
rect 7672 35930 7696 35932
rect 7752 35930 7776 35932
rect 7832 35930 7856 35932
rect 7912 35930 7918 35932
rect 7672 35878 7674 35930
rect 7854 35878 7856 35930
rect 7610 35876 7616 35878
rect 7672 35876 7696 35878
rect 7752 35876 7776 35878
rect 7832 35876 7856 35878
rect 7912 35876 7918 35878
rect 7610 35867 7918 35876
rect 8036 35698 8064 46106
rect 8128 42294 8156 50730
rect 8116 42288 8168 42294
rect 8116 42230 8168 42236
rect 8116 41812 8168 41818
rect 8116 41754 8168 41760
rect 8024 35692 8076 35698
rect 8024 35634 8076 35640
rect 7610 34844 7918 34853
rect 7610 34842 7616 34844
rect 7672 34842 7696 34844
rect 7752 34842 7776 34844
rect 7832 34842 7856 34844
rect 7912 34842 7918 34844
rect 7672 34790 7674 34842
rect 7854 34790 7856 34842
rect 7610 34788 7616 34790
rect 7672 34788 7696 34790
rect 7752 34788 7776 34790
rect 7832 34788 7856 34790
rect 7912 34788 7918 34790
rect 7610 34779 7918 34788
rect 8024 34604 8076 34610
rect 8024 34546 8076 34552
rect 7610 33756 7918 33765
rect 7610 33754 7616 33756
rect 7672 33754 7696 33756
rect 7752 33754 7776 33756
rect 7832 33754 7856 33756
rect 7912 33754 7918 33756
rect 7672 33702 7674 33754
rect 7854 33702 7856 33754
rect 7610 33700 7616 33702
rect 7672 33700 7696 33702
rect 7752 33700 7776 33702
rect 7832 33700 7856 33702
rect 7912 33700 7918 33702
rect 7610 33691 7918 33700
rect 7610 32668 7918 32677
rect 7610 32666 7616 32668
rect 7672 32666 7696 32668
rect 7752 32666 7776 32668
rect 7832 32666 7856 32668
rect 7912 32666 7918 32668
rect 7672 32614 7674 32666
rect 7854 32614 7856 32666
rect 7610 32612 7616 32614
rect 7672 32612 7696 32614
rect 7752 32612 7776 32614
rect 7832 32612 7856 32614
rect 7912 32612 7918 32614
rect 7610 32603 7918 32612
rect 7472 32564 7524 32570
rect 7472 32506 7524 32512
rect 7472 32428 7524 32434
rect 7472 32370 7524 32376
rect 7288 31340 7340 31346
rect 7288 31282 7340 31288
rect 7380 31340 7432 31346
rect 7380 31282 7432 31288
rect 7208 31198 7420 31226
rect 7288 31136 7340 31142
rect 7288 31078 7340 31084
rect 6950 31036 7258 31045
rect 6950 31034 6956 31036
rect 7012 31034 7036 31036
rect 7092 31034 7116 31036
rect 7172 31034 7196 31036
rect 7252 31034 7258 31036
rect 7012 30982 7014 31034
rect 7194 30982 7196 31034
rect 6950 30980 6956 30982
rect 7012 30980 7036 30982
rect 7092 30980 7116 30982
rect 7172 30980 7196 30982
rect 7252 30980 7258 30982
rect 6950 30971 7258 30980
rect 7300 30326 7328 31078
rect 7288 30320 7340 30326
rect 7288 30262 7340 30268
rect 6950 29948 7258 29957
rect 6950 29946 6956 29948
rect 7012 29946 7036 29948
rect 7092 29946 7116 29948
rect 7172 29946 7196 29948
rect 7252 29946 7258 29948
rect 7012 29894 7014 29946
rect 7194 29894 7196 29946
rect 6950 29892 6956 29894
rect 7012 29892 7036 29894
rect 7092 29892 7116 29894
rect 7172 29892 7196 29894
rect 7252 29892 7258 29894
rect 6950 29883 7258 29892
rect 7288 29708 7340 29714
rect 7288 29650 7340 29656
rect 6950 28860 7258 28869
rect 6950 28858 6956 28860
rect 7012 28858 7036 28860
rect 7092 28858 7116 28860
rect 7172 28858 7196 28860
rect 7252 28858 7258 28860
rect 7012 28806 7014 28858
rect 7194 28806 7196 28858
rect 6950 28804 6956 28806
rect 7012 28804 7036 28806
rect 7092 28804 7116 28806
rect 7172 28804 7196 28806
rect 7252 28804 7258 28806
rect 6950 28795 7258 28804
rect 6950 27772 7258 27781
rect 6950 27770 6956 27772
rect 7012 27770 7036 27772
rect 7092 27770 7116 27772
rect 7172 27770 7196 27772
rect 7252 27770 7258 27772
rect 7012 27718 7014 27770
rect 7194 27718 7196 27770
rect 6950 27716 6956 27718
rect 7012 27716 7036 27718
rect 7092 27716 7116 27718
rect 7172 27716 7196 27718
rect 7252 27716 7258 27718
rect 6950 27707 7258 27716
rect 7300 27606 7328 29650
rect 7288 27600 7340 27606
rect 7288 27542 7340 27548
rect 6950 26684 7258 26693
rect 6950 26682 6956 26684
rect 7012 26682 7036 26684
rect 7092 26682 7116 26684
rect 7172 26682 7196 26684
rect 7252 26682 7258 26684
rect 7012 26630 7014 26682
rect 7194 26630 7196 26682
rect 6950 26628 6956 26630
rect 7012 26628 7036 26630
rect 7092 26628 7116 26630
rect 7172 26628 7196 26630
rect 7252 26628 7258 26630
rect 6950 26619 7258 26628
rect 7300 26314 7328 27542
rect 7392 26586 7420 31198
rect 7380 26580 7432 26586
rect 7380 26522 7432 26528
rect 7288 26308 7340 26314
rect 7288 26250 7340 26256
rect 6950 25596 7258 25605
rect 6950 25594 6956 25596
rect 7012 25594 7036 25596
rect 7092 25594 7116 25596
rect 7172 25594 7196 25596
rect 7252 25594 7258 25596
rect 7012 25542 7014 25594
rect 7194 25542 7196 25594
rect 6950 25540 6956 25542
rect 7012 25540 7036 25542
rect 7092 25540 7116 25542
rect 7172 25540 7196 25542
rect 7252 25540 7258 25542
rect 6950 25531 7258 25540
rect 6736 24812 6788 24818
rect 6736 24754 6788 24760
rect 6950 24508 7258 24517
rect 6950 24506 6956 24508
rect 7012 24506 7036 24508
rect 7092 24506 7116 24508
rect 7172 24506 7196 24508
rect 7252 24506 7258 24508
rect 7012 24454 7014 24506
rect 7194 24454 7196 24506
rect 6950 24452 6956 24454
rect 7012 24452 7036 24454
rect 7092 24452 7116 24454
rect 7172 24452 7196 24454
rect 7252 24452 7258 24454
rect 6950 24443 7258 24452
rect 7300 23730 7328 26250
rect 7380 26240 7432 26246
rect 7380 26182 7432 26188
rect 7392 25362 7420 26182
rect 7380 25356 7432 25362
rect 7380 25298 7432 25304
rect 7380 23792 7432 23798
rect 7380 23734 7432 23740
rect 7288 23724 7340 23730
rect 7288 23666 7340 23672
rect 6950 23420 7258 23429
rect 6950 23418 6956 23420
rect 7012 23418 7036 23420
rect 7092 23418 7116 23420
rect 7172 23418 7196 23420
rect 7252 23418 7258 23420
rect 7012 23366 7014 23418
rect 7194 23366 7196 23418
rect 6950 23364 6956 23366
rect 7012 23364 7036 23366
rect 7092 23364 7116 23366
rect 7172 23364 7196 23366
rect 7252 23364 7258 23366
rect 6950 23355 7258 23364
rect 6950 22332 7258 22341
rect 6950 22330 6956 22332
rect 7012 22330 7036 22332
rect 7092 22330 7116 22332
rect 7172 22330 7196 22332
rect 7252 22330 7258 22332
rect 7012 22278 7014 22330
rect 7194 22278 7196 22330
rect 6950 22276 6956 22278
rect 7012 22276 7036 22278
rect 7092 22276 7116 22278
rect 7172 22276 7196 22278
rect 7252 22276 7258 22278
rect 6950 22267 7258 22276
rect 7104 22092 7156 22098
rect 7104 22034 7156 22040
rect 6920 22024 6972 22030
rect 6920 21966 6972 21972
rect 6644 21888 6696 21894
rect 6644 21830 6696 21836
rect 6656 11150 6684 21830
rect 6932 21434 6960 21966
rect 7116 21894 7144 22034
rect 7300 21962 7328 23666
rect 7288 21956 7340 21962
rect 7288 21898 7340 21904
rect 7104 21888 7156 21894
rect 7104 21830 7156 21836
rect 6840 21406 6960 21434
rect 6840 21010 6868 21406
rect 6950 21244 7258 21253
rect 6950 21242 6956 21244
rect 7012 21242 7036 21244
rect 7092 21242 7116 21244
rect 7172 21242 7196 21244
rect 7252 21242 7258 21244
rect 7012 21190 7014 21242
rect 7194 21190 7196 21242
rect 6950 21188 6956 21190
rect 7012 21188 7036 21190
rect 7092 21188 7116 21190
rect 7172 21188 7196 21190
rect 7252 21188 7258 21190
rect 6950 21179 7258 21188
rect 6828 21004 6880 21010
rect 6828 20946 6880 20952
rect 6950 20156 7258 20165
rect 6950 20154 6956 20156
rect 7012 20154 7036 20156
rect 7092 20154 7116 20156
rect 7172 20154 7196 20156
rect 7252 20154 7258 20156
rect 7012 20102 7014 20154
rect 7194 20102 7196 20154
rect 6950 20100 6956 20102
rect 7012 20100 7036 20102
rect 7092 20100 7116 20102
rect 7172 20100 7196 20102
rect 7252 20100 7258 20102
rect 6950 20091 7258 20100
rect 6950 19068 7258 19077
rect 6950 19066 6956 19068
rect 7012 19066 7036 19068
rect 7092 19066 7116 19068
rect 7172 19066 7196 19068
rect 7252 19066 7258 19068
rect 7012 19014 7014 19066
rect 7194 19014 7196 19066
rect 6950 19012 6956 19014
rect 7012 19012 7036 19014
rect 7092 19012 7116 19014
rect 7172 19012 7196 19014
rect 7252 19012 7258 19014
rect 6950 19003 7258 19012
rect 6950 17980 7258 17989
rect 6950 17978 6956 17980
rect 7012 17978 7036 17980
rect 7092 17978 7116 17980
rect 7172 17978 7196 17980
rect 7252 17978 7258 17980
rect 7012 17926 7014 17978
rect 7194 17926 7196 17978
rect 6950 17924 6956 17926
rect 7012 17924 7036 17926
rect 7092 17924 7116 17926
rect 7172 17924 7196 17926
rect 7252 17924 7258 17926
rect 6950 17915 7258 17924
rect 7300 17746 7328 21898
rect 7288 17740 7340 17746
rect 7288 17682 7340 17688
rect 6950 16892 7258 16901
rect 6950 16890 6956 16892
rect 7012 16890 7036 16892
rect 7092 16890 7116 16892
rect 7172 16890 7196 16892
rect 7252 16890 7258 16892
rect 7012 16838 7014 16890
rect 7194 16838 7196 16890
rect 6950 16836 6956 16838
rect 7012 16836 7036 16838
rect 7092 16836 7116 16838
rect 7172 16836 7196 16838
rect 7252 16836 7258 16838
rect 6950 16827 7258 16836
rect 7300 16794 7328 17682
rect 7288 16788 7340 16794
rect 7288 16730 7340 16736
rect 7288 16040 7340 16046
rect 7288 15982 7340 15988
rect 6950 15804 7258 15813
rect 6950 15802 6956 15804
rect 7012 15802 7036 15804
rect 7092 15802 7116 15804
rect 7172 15802 7196 15804
rect 7252 15802 7258 15804
rect 7012 15750 7014 15802
rect 7194 15750 7196 15802
rect 6950 15748 6956 15750
rect 7012 15748 7036 15750
rect 7092 15748 7116 15750
rect 7172 15748 7196 15750
rect 7252 15748 7258 15750
rect 6950 15739 7258 15748
rect 6950 14716 7258 14725
rect 6950 14714 6956 14716
rect 7012 14714 7036 14716
rect 7092 14714 7116 14716
rect 7172 14714 7196 14716
rect 7252 14714 7258 14716
rect 7012 14662 7014 14714
rect 7194 14662 7196 14714
rect 6950 14660 6956 14662
rect 7012 14660 7036 14662
rect 7092 14660 7116 14662
rect 7172 14660 7196 14662
rect 7252 14660 7258 14662
rect 6950 14651 7258 14660
rect 6950 13628 7258 13637
rect 6950 13626 6956 13628
rect 7012 13626 7036 13628
rect 7092 13626 7116 13628
rect 7172 13626 7196 13628
rect 7252 13626 7258 13628
rect 7012 13574 7014 13626
rect 7194 13574 7196 13626
rect 6950 13572 6956 13574
rect 7012 13572 7036 13574
rect 7092 13572 7116 13574
rect 7172 13572 7196 13574
rect 7252 13572 7258 13574
rect 6950 13563 7258 13572
rect 7300 13258 7328 15982
rect 7392 14618 7420 23734
rect 7380 14612 7432 14618
rect 7380 14554 7432 14560
rect 7288 13252 7340 13258
rect 7288 13194 7340 13200
rect 6950 12540 7258 12549
rect 6950 12538 6956 12540
rect 7012 12538 7036 12540
rect 7092 12538 7116 12540
rect 7172 12538 7196 12540
rect 7252 12538 7258 12540
rect 7012 12486 7014 12538
rect 7194 12486 7196 12538
rect 6950 12484 6956 12486
rect 7012 12484 7036 12486
rect 7092 12484 7116 12486
rect 7172 12484 7196 12486
rect 7252 12484 7258 12486
rect 6950 12475 7258 12484
rect 6950 11452 7258 11461
rect 6950 11450 6956 11452
rect 7012 11450 7036 11452
rect 7092 11450 7116 11452
rect 7172 11450 7196 11452
rect 7252 11450 7258 11452
rect 7012 11398 7014 11450
rect 7194 11398 7196 11450
rect 6950 11396 6956 11398
rect 7012 11396 7036 11398
rect 7092 11396 7116 11398
rect 7172 11396 7196 11398
rect 7252 11396 7258 11398
rect 6950 11387 7258 11396
rect 6644 11144 6696 11150
rect 6644 11086 6696 11092
rect 6950 10364 7258 10373
rect 6950 10362 6956 10364
rect 7012 10362 7036 10364
rect 7092 10362 7116 10364
rect 7172 10362 7196 10364
rect 7252 10362 7258 10364
rect 7012 10310 7014 10362
rect 7194 10310 7196 10362
rect 6950 10308 6956 10310
rect 7012 10308 7036 10310
rect 7092 10308 7116 10310
rect 7172 10308 7196 10310
rect 7252 10308 7258 10310
rect 6950 10299 7258 10308
rect 6920 10260 6972 10266
rect 6920 10202 6972 10208
rect 6932 10062 6960 10202
rect 7300 10062 7328 13194
rect 7380 12436 7432 12442
rect 7484 12434 7512 32370
rect 8036 31754 8064 34546
rect 8024 31748 8076 31754
rect 8024 31690 8076 31696
rect 8128 31686 8156 41754
rect 8220 35086 8248 59638
rect 8404 57594 8432 64466
rect 8484 60784 8536 60790
rect 8484 60726 8536 60732
rect 8392 57588 8444 57594
rect 8392 57530 8444 57536
rect 8300 57248 8352 57254
rect 8300 57190 8352 57196
rect 8312 49910 8340 57190
rect 8392 54324 8444 54330
rect 8392 54266 8444 54272
rect 8300 49904 8352 49910
rect 8300 49846 8352 49852
rect 8404 47802 8432 54266
rect 8392 47796 8444 47802
rect 8392 47738 8444 47744
rect 8392 44192 8444 44198
rect 8392 44134 8444 44140
rect 8300 42288 8352 42294
rect 8300 42230 8352 42236
rect 8208 35080 8260 35086
rect 8208 35022 8260 35028
rect 8208 34944 8260 34950
rect 8208 34886 8260 34892
rect 8116 31680 8168 31686
rect 8116 31622 8168 31628
rect 7610 31580 7918 31589
rect 7610 31578 7616 31580
rect 7672 31578 7696 31580
rect 7752 31578 7776 31580
rect 7832 31578 7856 31580
rect 7912 31578 7918 31580
rect 7672 31526 7674 31578
rect 7854 31526 7856 31578
rect 7610 31524 7616 31526
rect 7672 31524 7696 31526
rect 7752 31524 7776 31526
rect 7832 31524 7856 31526
rect 7912 31524 7918 31526
rect 7610 31515 7918 31524
rect 8220 31498 8248 34886
rect 8312 32434 8340 42230
rect 8404 41818 8432 44134
rect 8392 41812 8444 41818
rect 8392 41754 8444 41760
rect 8496 40186 8524 60726
rect 8576 52896 8628 52902
rect 8576 52838 8628 52844
rect 8588 49094 8616 52838
rect 8576 49088 8628 49094
rect 8576 49030 8628 49036
rect 8576 48748 8628 48754
rect 8576 48690 8628 48696
rect 8484 40180 8536 40186
rect 8484 40122 8536 40128
rect 8392 39976 8444 39982
rect 8392 39918 8444 39924
rect 8484 39976 8536 39982
rect 8484 39918 8536 39924
rect 8404 39642 8432 39918
rect 8496 39846 8524 39918
rect 8484 39840 8536 39846
rect 8484 39782 8536 39788
rect 8392 39636 8444 39642
rect 8392 39578 8444 39584
rect 8484 39432 8536 39438
rect 8484 39374 8536 39380
rect 8392 37120 8444 37126
rect 8392 37062 8444 37068
rect 8404 36922 8432 37062
rect 8392 36916 8444 36922
rect 8392 36858 8444 36864
rect 8496 35170 8524 39374
rect 8404 35154 8524 35170
rect 8392 35148 8524 35154
rect 8444 35142 8524 35148
rect 8392 35090 8444 35096
rect 8496 33017 8524 35142
rect 8482 33008 8538 33017
rect 8482 32943 8538 32952
rect 8300 32428 8352 32434
rect 8300 32370 8352 32376
rect 8392 32360 8444 32366
rect 8392 32302 8444 32308
rect 8300 31680 8352 31686
rect 8300 31622 8352 31628
rect 8128 31470 8248 31498
rect 7610 30492 7918 30501
rect 7610 30490 7616 30492
rect 7672 30490 7696 30492
rect 7752 30490 7776 30492
rect 7832 30490 7856 30492
rect 7912 30490 7918 30492
rect 7672 30438 7674 30490
rect 7854 30438 7856 30490
rect 7610 30436 7616 30438
rect 7672 30436 7696 30438
rect 7752 30436 7776 30438
rect 7832 30436 7856 30438
rect 7912 30436 7918 30438
rect 7610 30427 7918 30436
rect 7564 30320 7616 30326
rect 7564 30262 7616 30268
rect 8024 30320 8076 30326
rect 8024 30262 8076 30268
rect 7576 29510 7604 30262
rect 7748 30252 7800 30258
rect 7748 30194 7800 30200
rect 7760 29714 7788 30194
rect 7748 29708 7800 29714
rect 7748 29650 7800 29656
rect 7564 29504 7616 29510
rect 7564 29446 7616 29452
rect 7610 29404 7918 29413
rect 7610 29402 7616 29404
rect 7672 29402 7696 29404
rect 7752 29402 7776 29404
rect 7832 29402 7856 29404
rect 7912 29402 7918 29404
rect 7672 29350 7674 29402
rect 7854 29350 7856 29402
rect 7610 29348 7616 29350
rect 7672 29348 7696 29350
rect 7752 29348 7776 29350
rect 7832 29348 7856 29350
rect 7912 29348 7918 29350
rect 7610 29339 7918 29348
rect 7932 29232 7984 29238
rect 7932 29174 7984 29180
rect 7944 28529 7972 29174
rect 7930 28520 7986 28529
rect 7930 28455 7986 28464
rect 7610 28316 7918 28325
rect 7610 28314 7616 28316
rect 7672 28314 7696 28316
rect 7752 28314 7776 28316
rect 7832 28314 7856 28316
rect 7912 28314 7918 28316
rect 7672 28262 7674 28314
rect 7854 28262 7856 28314
rect 7610 28260 7616 28262
rect 7672 28260 7696 28262
rect 7752 28260 7776 28262
rect 7832 28260 7856 28262
rect 7912 28260 7918 28262
rect 7610 28251 7918 28260
rect 7610 27228 7918 27237
rect 7610 27226 7616 27228
rect 7672 27226 7696 27228
rect 7752 27226 7776 27228
rect 7832 27226 7856 27228
rect 7912 27226 7918 27228
rect 7672 27174 7674 27226
rect 7854 27174 7856 27226
rect 7610 27172 7616 27174
rect 7672 27172 7696 27174
rect 7752 27172 7776 27174
rect 7832 27172 7856 27174
rect 7912 27172 7918 27174
rect 7610 27163 7918 27172
rect 8036 26194 8064 30262
rect 8128 26353 8156 31470
rect 8208 31340 8260 31346
rect 8208 31282 8260 31288
rect 8114 26344 8170 26353
rect 8114 26279 8170 26288
rect 8036 26166 8156 26194
rect 7610 26140 7918 26149
rect 7610 26138 7616 26140
rect 7672 26138 7696 26140
rect 7752 26138 7776 26140
rect 7832 26138 7856 26140
rect 7912 26138 7918 26140
rect 7672 26086 7674 26138
rect 7854 26086 7856 26138
rect 7610 26084 7616 26086
rect 7672 26084 7696 26086
rect 7752 26084 7776 26086
rect 7832 26084 7856 26086
rect 7912 26084 7918 26086
rect 7610 26075 7918 26084
rect 8022 26072 8078 26081
rect 8022 26007 8078 26016
rect 7610 25052 7918 25061
rect 7610 25050 7616 25052
rect 7672 25050 7696 25052
rect 7752 25050 7776 25052
rect 7832 25050 7856 25052
rect 7912 25050 7918 25052
rect 7672 24998 7674 25050
rect 7854 24998 7856 25050
rect 7610 24996 7616 24998
rect 7672 24996 7696 24998
rect 7752 24996 7776 24998
rect 7832 24996 7856 24998
rect 7912 24996 7918 24998
rect 7610 24987 7918 24996
rect 7610 23964 7918 23973
rect 7610 23962 7616 23964
rect 7672 23962 7696 23964
rect 7752 23962 7776 23964
rect 7832 23962 7856 23964
rect 7912 23962 7918 23964
rect 7672 23910 7674 23962
rect 7854 23910 7856 23962
rect 7610 23908 7616 23910
rect 7672 23908 7696 23910
rect 7752 23908 7776 23910
rect 7832 23908 7856 23910
rect 7912 23908 7918 23910
rect 7610 23899 7918 23908
rect 7610 22876 7918 22885
rect 7610 22874 7616 22876
rect 7672 22874 7696 22876
rect 7752 22874 7776 22876
rect 7832 22874 7856 22876
rect 7912 22874 7918 22876
rect 7672 22822 7674 22874
rect 7854 22822 7856 22874
rect 7610 22820 7616 22822
rect 7672 22820 7696 22822
rect 7752 22820 7776 22822
rect 7832 22820 7856 22822
rect 7912 22820 7918 22822
rect 7610 22811 7918 22820
rect 7932 22772 7984 22778
rect 7932 22714 7984 22720
rect 7944 21894 7972 22714
rect 7932 21888 7984 21894
rect 7932 21830 7984 21836
rect 7610 21788 7918 21797
rect 7610 21786 7616 21788
rect 7672 21786 7696 21788
rect 7752 21786 7776 21788
rect 7832 21786 7856 21788
rect 7912 21786 7918 21788
rect 7672 21734 7674 21786
rect 7854 21734 7856 21786
rect 7610 21732 7616 21734
rect 7672 21732 7696 21734
rect 7752 21732 7776 21734
rect 7832 21732 7856 21734
rect 7912 21732 7918 21734
rect 7610 21723 7918 21732
rect 7610 20700 7918 20709
rect 7610 20698 7616 20700
rect 7672 20698 7696 20700
rect 7752 20698 7776 20700
rect 7832 20698 7856 20700
rect 7912 20698 7918 20700
rect 7672 20646 7674 20698
rect 7854 20646 7856 20698
rect 7610 20644 7616 20646
rect 7672 20644 7696 20646
rect 7752 20644 7776 20646
rect 7832 20644 7856 20646
rect 7912 20644 7918 20646
rect 7610 20635 7918 20644
rect 7610 19612 7918 19621
rect 7610 19610 7616 19612
rect 7672 19610 7696 19612
rect 7752 19610 7776 19612
rect 7832 19610 7856 19612
rect 7912 19610 7918 19612
rect 7672 19558 7674 19610
rect 7854 19558 7856 19610
rect 7610 19556 7616 19558
rect 7672 19556 7696 19558
rect 7752 19556 7776 19558
rect 7832 19556 7856 19558
rect 7912 19556 7918 19558
rect 7610 19547 7918 19556
rect 7610 18524 7918 18533
rect 7610 18522 7616 18524
rect 7672 18522 7696 18524
rect 7752 18522 7776 18524
rect 7832 18522 7856 18524
rect 7912 18522 7918 18524
rect 7672 18470 7674 18522
rect 7854 18470 7856 18522
rect 7610 18468 7616 18470
rect 7672 18468 7696 18470
rect 7752 18468 7776 18470
rect 7832 18468 7856 18470
rect 7912 18468 7918 18470
rect 7610 18459 7918 18468
rect 7610 17436 7918 17445
rect 7610 17434 7616 17436
rect 7672 17434 7696 17436
rect 7752 17434 7776 17436
rect 7832 17434 7856 17436
rect 7912 17434 7918 17436
rect 7672 17382 7674 17434
rect 7854 17382 7856 17434
rect 7610 17380 7616 17382
rect 7672 17380 7696 17382
rect 7752 17380 7776 17382
rect 7832 17380 7856 17382
rect 7912 17380 7918 17382
rect 7610 17371 7918 17380
rect 7610 16348 7918 16357
rect 7610 16346 7616 16348
rect 7672 16346 7696 16348
rect 7752 16346 7776 16348
rect 7832 16346 7856 16348
rect 7912 16346 7918 16348
rect 7672 16294 7674 16346
rect 7854 16294 7856 16346
rect 7610 16292 7616 16294
rect 7672 16292 7696 16294
rect 7752 16292 7776 16294
rect 7832 16292 7856 16294
rect 7912 16292 7918 16294
rect 7610 16283 7918 16292
rect 7610 15260 7918 15269
rect 7610 15258 7616 15260
rect 7672 15258 7696 15260
rect 7752 15258 7776 15260
rect 7832 15258 7856 15260
rect 7912 15258 7918 15260
rect 7672 15206 7674 15258
rect 7854 15206 7856 15258
rect 7610 15204 7616 15206
rect 7672 15204 7696 15206
rect 7752 15204 7776 15206
rect 7832 15204 7856 15206
rect 7912 15204 7918 15206
rect 7610 15195 7918 15204
rect 7838 15056 7894 15065
rect 7838 14991 7894 15000
rect 7852 14414 7880 14991
rect 7840 14408 7892 14414
rect 7840 14350 7892 14356
rect 7610 14172 7918 14181
rect 7610 14170 7616 14172
rect 7672 14170 7696 14172
rect 7752 14170 7776 14172
rect 7832 14170 7856 14172
rect 7912 14170 7918 14172
rect 7672 14118 7674 14170
rect 7854 14118 7856 14170
rect 7610 14116 7616 14118
rect 7672 14116 7696 14118
rect 7752 14116 7776 14118
rect 7832 14116 7856 14118
rect 7912 14116 7918 14118
rect 7610 14107 7918 14116
rect 7610 13084 7918 13093
rect 7610 13082 7616 13084
rect 7672 13082 7696 13084
rect 7752 13082 7776 13084
rect 7832 13082 7856 13084
rect 7912 13082 7918 13084
rect 7672 13030 7674 13082
rect 7854 13030 7856 13082
rect 7610 13028 7616 13030
rect 7672 13028 7696 13030
rect 7752 13028 7776 13030
rect 7832 13028 7856 13030
rect 7912 13028 7918 13030
rect 7610 13019 7918 13028
rect 7432 12406 7512 12434
rect 7380 12378 7432 12384
rect 7392 10130 7420 12378
rect 7610 11996 7918 12005
rect 7610 11994 7616 11996
rect 7672 11994 7696 11996
rect 7752 11994 7776 11996
rect 7832 11994 7856 11996
rect 7912 11994 7918 11996
rect 7672 11942 7674 11994
rect 7854 11942 7856 11994
rect 7610 11940 7616 11942
rect 7672 11940 7696 11942
rect 7752 11940 7776 11942
rect 7832 11940 7856 11942
rect 7912 11940 7918 11942
rect 7610 11931 7918 11940
rect 7610 10908 7918 10917
rect 7610 10906 7616 10908
rect 7672 10906 7696 10908
rect 7752 10906 7776 10908
rect 7832 10906 7856 10908
rect 7912 10906 7918 10908
rect 7672 10854 7674 10906
rect 7854 10854 7856 10906
rect 7610 10852 7616 10854
rect 7672 10852 7696 10854
rect 7752 10852 7776 10854
rect 7832 10852 7856 10854
rect 7912 10852 7918 10854
rect 7610 10843 7918 10852
rect 7930 10568 7986 10577
rect 7930 10503 7986 10512
rect 7944 10130 7972 10503
rect 7380 10124 7432 10130
rect 7380 10066 7432 10072
rect 7932 10124 7984 10130
rect 7932 10066 7984 10072
rect 6920 10056 6972 10062
rect 7288 10056 7340 10062
rect 6920 9998 6972 10004
rect 7010 10024 7066 10033
rect 7288 9998 7340 10004
rect 7010 9959 7066 9968
rect 6642 9616 6698 9625
rect 6642 9551 6644 9560
rect 6696 9551 6698 9560
rect 6644 9522 6696 9528
rect 7024 9450 7052 9959
rect 7012 9444 7064 9450
rect 7012 9386 7064 9392
rect 6950 9276 7258 9285
rect 6950 9274 6956 9276
rect 7012 9274 7036 9276
rect 7092 9274 7116 9276
rect 7172 9274 7196 9276
rect 7252 9274 7258 9276
rect 7012 9222 7014 9274
rect 7194 9222 7196 9274
rect 6950 9220 6956 9222
rect 7012 9220 7036 9222
rect 7092 9220 7116 9222
rect 7172 9220 7196 9222
rect 7252 9220 7258 9222
rect 6950 9211 7258 9220
rect 6950 8188 7258 8197
rect 6950 8186 6956 8188
rect 7012 8186 7036 8188
rect 7092 8186 7116 8188
rect 7172 8186 7196 8188
rect 7252 8186 7258 8188
rect 7012 8134 7014 8186
rect 7194 8134 7196 8186
rect 6950 8132 6956 8134
rect 7012 8132 7036 8134
rect 7092 8132 7116 8134
rect 7172 8132 7196 8134
rect 7252 8132 7258 8134
rect 6950 8123 7258 8132
rect 6950 7100 7258 7109
rect 6950 7098 6956 7100
rect 7012 7098 7036 7100
rect 7092 7098 7116 7100
rect 7172 7098 7196 7100
rect 7252 7098 7258 7100
rect 7012 7046 7014 7098
rect 7194 7046 7196 7098
rect 6950 7044 6956 7046
rect 7012 7044 7036 7046
rect 7092 7044 7116 7046
rect 7172 7044 7196 7046
rect 7252 7044 7258 7046
rect 6950 7035 7258 7044
rect 6920 6928 6972 6934
rect 6920 6870 6972 6876
rect 6932 6769 6960 6870
rect 6918 6760 6974 6769
rect 6918 6695 6974 6704
rect 6950 6012 7258 6021
rect 6950 6010 6956 6012
rect 7012 6010 7036 6012
rect 7092 6010 7116 6012
rect 7172 6010 7196 6012
rect 7252 6010 7258 6012
rect 7012 5958 7014 6010
rect 7194 5958 7196 6010
rect 6950 5956 6956 5958
rect 7012 5956 7036 5958
rect 7092 5956 7116 5958
rect 7172 5956 7196 5958
rect 7252 5956 7258 5958
rect 6950 5947 7258 5956
rect 6552 5092 6604 5098
rect 6552 5034 6604 5040
rect 6950 4924 7258 4933
rect 6950 4922 6956 4924
rect 7012 4922 7036 4924
rect 7092 4922 7116 4924
rect 7172 4922 7196 4924
rect 7252 4922 7258 4924
rect 7012 4870 7014 4922
rect 7194 4870 7196 4922
rect 6950 4868 6956 4870
rect 7012 4868 7036 4870
rect 7092 4868 7116 4870
rect 7172 4868 7196 4870
rect 7252 4868 7258 4870
rect 6950 4859 7258 4868
rect 7300 4690 7328 9998
rect 7944 9926 7972 10066
rect 7932 9920 7984 9926
rect 7932 9862 7984 9868
rect 7610 9820 7918 9829
rect 7610 9818 7616 9820
rect 7672 9818 7696 9820
rect 7752 9818 7776 9820
rect 7832 9818 7856 9820
rect 7912 9818 7918 9820
rect 7672 9766 7674 9818
rect 7854 9766 7856 9818
rect 7610 9764 7616 9766
rect 7672 9764 7696 9766
rect 7752 9764 7776 9766
rect 7832 9764 7856 9766
rect 7912 9764 7918 9766
rect 7610 9755 7918 9764
rect 7932 9376 7984 9382
rect 7932 9318 7984 9324
rect 7944 9042 7972 9318
rect 7472 9036 7524 9042
rect 7472 8978 7524 8984
rect 7932 9036 7984 9042
rect 7932 8978 7984 8984
rect 7378 6896 7434 6905
rect 7484 6866 7512 8978
rect 8036 8906 8064 26007
rect 8128 9178 8156 26166
rect 8220 22778 8248 31282
rect 8312 26246 8340 31622
rect 8404 29238 8432 32302
rect 8392 29232 8444 29238
rect 8392 29174 8444 29180
rect 8392 27124 8444 27130
rect 8392 27066 8444 27072
rect 8300 26240 8352 26246
rect 8300 26182 8352 26188
rect 8298 26072 8354 26081
rect 8298 26007 8354 26016
rect 8208 22772 8260 22778
rect 8208 22714 8260 22720
rect 8208 21888 8260 21894
rect 8208 21830 8260 21836
rect 8220 10266 8248 21830
rect 8312 16046 8340 26007
rect 8404 20534 8432 27066
rect 8482 26888 8538 26897
rect 8482 26823 8538 26832
rect 8392 20528 8444 20534
rect 8392 20470 8444 20476
rect 8496 16454 8524 26823
rect 8484 16448 8536 16454
rect 8484 16390 8536 16396
rect 8300 16040 8352 16046
rect 8300 15982 8352 15988
rect 8390 15192 8446 15201
rect 8390 15127 8446 15136
rect 8404 14414 8432 15127
rect 8392 14408 8444 14414
rect 8392 14350 8444 14356
rect 8588 13530 8616 48690
rect 8680 42362 8708 65010
rect 8760 62688 8812 62694
rect 8758 62656 8760 62665
rect 8812 62656 8814 62665
rect 8758 62591 8814 62600
rect 8760 52488 8812 52494
rect 8760 52430 8812 52436
rect 8772 50794 8800 52430
rect 8760 50788 8812 50794
rect 8760 50730 8812 50736
rect 8852 47728 8904 47734
rect 8852 47670 8904 47676
rect 8760 43784 8812 43790
rect 8760 43726 8812 43732
rect 8668 42356 8720 42362
rect 8668 42298 8720 42304
rect 8680 40526 8708 42298
rect 8668 40520 8720 40526
rect 8668 40462 8720 40468
rect 8772 40202 8800 43726
rect 8864 40610 8892 47670
rect 8956 43246 8984 76230
rect 11704 76230 11756 76236
rect 11242 76191 11298 76200
rect 9220 75744 9272 75750
rect 9220 75686 9272 75692
rect 9128 70984 9180 70990
rect 9128 70926 9180 70932
rect 9036 70848 9088 70854
rect 9036 70790 9088 70796
rect 8944 43240 8996 43246
rect 8944 43182 8996 43188
rect 9048 41414 9076 70790
rect 9140 69426 9168 70926
rect 9128 69420 9180 69426
rect 9128 69362 9180 69368
rect 9140 68882 9168 69362
rect 9128 68876 9180 68882
rect 9128 68818 9180 68824
rect 9128 53100 9180 53106
rect 9128 53042 9180 53048
rect 9140 42362 9168 53042
rect 9128 42356 9180 42362
rect 9128 42298 9180 42304
rect 9048 41386 9168 41414
rect 8864 40582 9076 40610
rect 8944 40520 8996 40526
rect 8944 40462 8996 40468
rect 8772 40174 8892 40202
rect 8864 40118 8892 40174
rect 8852 40112 8904 40118
rect 8852 40054 8904 40060
rect 8760 39976 8812 39982
rect 8760 39918 8812 39924
rect 8668 39840 8720 39846
rect 8668 39782 8720 39788
rect 8680 36718 8708 39782
rect 8668 36712 8720 36718
rect 8668 36654 8720 36660
rect 8772 35086 8800 39918
rect 8760 35080 8812 35086
rect 8760 35022 8812 35028
rect 8772 34542 8800 35022
rect 8760 34536 8812 34542
rect 8760 34478 8812 34484
rect 8772 29714 8800 34478
rect 8760 29708 8812 29714
rect 8760 29650 8812 29656
rect 8760 29096 8812 29102
rect 8760 29038 8812 29044
rect 8668 26920 8720 26926
rect 8668 26862 8720 26868
rect 8680 20330 8708 26862
rect 8668 20324 8720 20330
rect 8668 20266 8720 20272
rect 8576 13524 8628 13530
rect 8576 13466 8628 13472
rect 8680 12434 8708 20266
rect 8404 12406 8708 12434
rect 8298 11112 8354 11121
rect 8298 11047 8354 11056
rect 8208 10260 8260 10266
rect 8208 10202 8260 10208
rect 8312 10146 8340 11047
rect 8220 10118 8340 10146
rect 8116 9172 8168 9178
rect 8116 9114 8168 9120
rect 8220 8974 8248 10118
rect 8116 8968 8168 8974
rect 8116 8910 8168 8916
rect 8208 8968 8260 8974
rect 8208 8910 8260 8916
rect 8024 8900 8076 8906
rect 8024 8842 8076 8848
rect 7610 8732 7918 8741
rect 7610 8730 7616 8732
rect 7672 8730 7696 8732
rect 7752 8730 7776 8732
rect 7832 8730 7856 8732
rect 7912 8730 7918 8732
rect 7672 8678 7674 8730
rect 7854 8678 7856 8730
rect 7610 8676 7616 8678
rect 7672 8676 7696 8678
rect 7752 8676 7776 8678
rect 7832 8676 7856 8678
rect 7912 8676 7918 8678
rect 7610 8667 7918 8676
rect 8128 8634 8156 8910
rect 8116 8628 8168 8634
rect 8116 8570 8168 8576
rect 7610 7644 7918 7653
rect 7610 7642 7616 7644
rect 7672 7642 7696 7644
rect 7752 7642 7776 7644
rect 7832 7642 7856 7644
rect 7912 7642 7918 7644
rect 7672 7590 7674 7642
rect 7854 7590 7856 7642
rect 7610 7588 7616 7590
rect 7672 7588 7696 7590
rect 7752 7588 7776 7590
rect 7832 7588 7856 7590
rect 7912 7588 7918 7590
rect 7610 7579 7918 7588
rect 8404 6914 8432 12406
rect 8772 7954 8800 29038
rect 8760 7948 8812 7954
rect 8760 7890 8812 7896
rect 8312 6886 8432 6914
rect 7378 6831 7380 6840
rect 7432 6831 7434 6840
rect 7472 6860 7524 6866
rect 7380 6802 7432 6808
rect 7472 6802 7524 6808
rect 7610 6556 7918 6565
rect 7610 6554 7616 6556
rect 7672 6554 7696 6556
rect 7752 6554 7776 6556
rect 7832 6554 7856 6556
rect 7912 6554 7918 6556
rect 7672 6502 7674 6554
rect 7854 6502 7856 6554
rect 7610 6500 7616 6502
rect 7672 6500 7696 6502
rect 7752 6500 7776 6502
rect 7832 6500 7856 6502
rect 7912 6500 7918 6502
rect 7610 6491 7918 6500
rect 8208 6384 8260 6390
rect 8208 6326 8260 6332
rect 7610 5468 7918 5477
rect 7610 5466 7616 5468
rect 7672 5466 7696 5468
rect 7752 5466 7776 5468
rect 7832 5466 7856 5468
rect 7912 5466 7918 5468
rect 7672 5414 7674 5466
rect 7854 5414 7856 5466
rect 7610 5412 7616 5414
rect 7672 5412 7696 5414
rect 7752 5412 7776 5414
rect 7832 5412 7856 5414
rect 7912 5412 7918 5414
rect 7610 5403 7918 5412
rect 8116 5024 8168 5030
rect 8116 4966 8168 4972
rect 7288 4684 7340 4690
rect 7288 4626 7340 4632
rect 7610 4380 7918 4389
rect 7610 4378 7616 4380
rect 7672 4378 7696 4380
rect 7752 4378 7776 4380
rect 7832 4378 7856 4380
rect 7912 4378 7918 4380
rect 7672 4326 7674 4378
rect 7854 4326 7856 4378
rect 7610 4324 7616 4326
rect 7672 4324 7696 4326
rect 7752 4324 7776 4326
rect 7832 4324 7856 4326
rect 7912 4324 7918 4326
rect 7610 4315 7918 4324
rect 6950 3836 7258 3845
rect 6950 3834 6956 3836
rect 7012 3834 7036 3836
rect 7092 3834 7116 3836
rect 7172 3834 7196 3836
rect 7252 3834 7258 3836
rect 7012 3782 7014 3834
rect 7194 3782 7196 3834
rect 6950 3780 6956 3782
rect 7012 3780 7036 3782
rect 7092 3780 7116 3782
rect 7172 3780 7196 3782
rect 7252 3780 7258 3782
rect 6950 3771 7258 3780
rect 8128 3534 8156 4966
rect 8220 4078 8248 6326
rect 8208 4072 8260 4078
rect 8208 4014 8260 4020
rect 8312 4010 8340 6886
rect 8300 4004 8352 4010
rect 8300 3946 8352 3952
rect 8116 3528 8168 3534
rect 8116 3470 8168 3476
rect 7610 3292 7918 3301
rect 7610 3290 7616 3292
rect 7672 3290 7696 3292
rect 7752 3290 7776 3292
rect 7832 3290 7856 3292
rect 7912 3290 7918 3292
rect 7672 3238 7674 3290
rect 7854 3238 7856 3290
rect 7610 3236 7616 3238
rect 7672 3236 7696 3238
rect 7752 3236 7776 3238
rect 7832 3236 7856 3238
rect 7912 3236 7918 3238
rect 7610 3227 7918 3236
rect 5632 3120 5684 3126
rect 5632 3062 5684 3068
rect 2320 2984 2372 2990
rect 2320 2926 2372 2932
rect 1950 2748 2258 2757
rect 1950 2746 1956 2748
rect 2012 2746 2036 2748
rect 2092 2746 2116 2748
rect 2172 2746 2196 2748
rect 2252 2746 2258 2748
rect 2012 2694 2014 2746
rect 2194 2694 2196 2746
rect 1950 2692 1956 2694
rect 2012 2692 2036 2694
rect 2092 2692 2116 2694
rect 2172 2692 2196 2694
rect 2252 2692 2258 2694
rect 1950 2683 2258 2692
rect 2056 870 2176 898
rect 2056 800 2084 870
rect 2042 0 2098 800
rect 2148 762 2176 870
rect 2332 762 2360 2926
rect 6950 2748 7258 2757
rect 6950 2746 6956 2748
rect 7012 2746 7036 2748
rect 7092 2746 7116 2748
rect 7172 2746 7196 2748
rect 7252 2746 7258 2748
rect 7012 2694 7014 2746
rect 7194 2694 7196 2746
rect 6950 2692 6956 2694
rect 7012 2692 7036 2694
rect 7092 2692 7116 2694
rect 7172 2692 7196 2694
rect 7252 2692 7258 2694
rect 6950 2683 7258 2692
rect 8864 2446 8892 40054
rect 8956 39574 8984 40462
rect 8944 39568 8996 39574
rect 8944 39510 8996 39516
rect 9048 37126 9076 40582
rect 9140 39370 9168 41386
rect 9128 39364 9180 39370
rect 9128 39306 9180 39312
rect 9036 37120 9088 37126
rect 9036 37062 9088 37068
rect 9128 36780 9180 36786
rect 9128 36722 9180 36728
rect 9036 33448 9088 33454
rect 9036 33390 9088 33396
rect 8942 33144 8998 33153
rect 8942 33079 8998 33088
rect 8956 27033 8984 33079
rect 8942 27024 8998 27033
rect 8942 26959 8998 26968
rect 9048 26926 9076 33390
rect 9140 30598 9168 36722
rect 9128 30592 9180 30598
rect 9128 30534 9180 30540
rect 9140 29714 9168 30534
rect 9128 29708 9180 29714
rect 9128 29650 9180 29656
rect 9140 29102 9168 29650
rect 9128 29096 9180 29102
rect 9128 29038 9180 29044
rect 9128 28620 9180 28626
rect 9128 28562 9180 28568
rect 9036 26920 9088 26926
rect 9036 26862 9088 26868
rect 8944 24608 8996 24614
rect 8944 24550 8996 24556
rect 8956 12238 8984 24550
rect 9140 21146 9168 28562
rect 9232 22166 9260 75686
rect 9404 74792 9456 74798
rect 9404 74734 9456 74740
rect 9312 69896 9364 69902
rect 9312 69838 9364 69844
rect 9324 52494 9352 69838
rect 9416 60654 9444 74734
rect 10324 74452 10376 74458
rect 10324 74394 10376 74400
rect 9864 70984 9916 70990
rect 9864 70926 9916 70932
rect 9588 68740 9640 68746
rect 9588 68682 9640 68688
rect 9496 65476 9548 65482
rect 9496 65418 9548 65424
rect 9508 60790 9536 65418
rect 9600 62830 9628 68682
rect 9680 63844 9732 63850
rect 9680 63786 9732 63792
rect 9692 63306 9720 63786
rect 9680 63300 9732 63306
rect 9680 63242 9732 63248
rect 9588 62824 9640 62830
rect 9588 62766 9640 62772
rect 9496 60784 9548 60790
rect 9496 60726 9548 60732
rect 9404 60648 9456 60654
rect 9404 60590 9456 60596
rect 9312 52488 9364 52494
rect 9312 52430 9364 52436
rect 9312 50720 9364 50726
rect 9312 50662 9364 50668
rect 9324 42566 9352 50662
rect 9312 42560 9364 42566
rect 9312 42502 9364 42508
rect 9312 42288 9364 42294
rect 9312 42230 9364 42236
rect 9324 41614 9352 42230
rect 9312 41608 9364 41614
rect 9312 41550 9364 41556
rect 9312 40180 9364 40186
rect 9312 40122 9364 40128
rect 9324 36106 9352 40122
rect 9312 36100 9364 36106
rect 9312 36042 9364 36048
rect 9324 23866 9352 36042
rect 9416 31754 9444 60590
rect 9588 59968 9640 59974
rect 9588 59910 9640 59916
rect 9496 52896 9548 52902
rect 9496 52838 9548 52844
rect 9508 52601 9536 52838
rect 9494 52592 9550 52601
rect 9494 52527 9550 52536
rect 9600 49774 9628 59910
rect 9876 53038 9904 70926
rect 9956 63776 10008 63782
rect 9956 63718 10008 63724
rect 9864 53032 9916 53038
rect 9864 52974 9916 52980
rect 9588 49768 9640 49774
rect 9588 49710 9640 49716
rect 9772 43852 9824 43858
rect 9772 43794 9824 43800
rect 9680 42560 9732 42566
rect 9680 42502 9732 42508
rect 9496 42084 9548 42090
rect 9496 42026 9548 42032
rect 9508 40497 9536 42026
rect 9494 40488 9550 40497
rect 9494 40423 9550 40432
rect 9588 37460 9640 37466
rect 9588 37402 9640 37408
rect 9496 34672 9548 34678
rect 9496 34614 9548 34620
rect 9508 31890 9536 34614
rect 9496 31884 9548 31890
rect 9496 31826 9548 31832
rect 9416 31726 9536 31754
rect 9404 29504 9456 29510
rect 9404 29446 9456 29452
rect 9312 23860 9364 23866
rect 9312 23802 9364 23808
rect 9220 22160 9272 22166
rect 9220 22102 9272 22108
rect 9128 21140 9180 21146
rect 9128 21082 9180 21088
rect 9416 21010 9444 29446
rect 9508 27130 9536 31726
rect 9496 27124 9548 27130
rect 9496 27066 9548 27072
rect 9496 22024 9548 22030
rect 9496 21966 9548 21972
rect 9404 21004 9456 21010
rect 9404 20946 9456 20952
rect 9312 20800 9364 20806
rect 9312 20742 9364 20748
rect 9034 16552 9090 16561
rect 9034 16487 9090 16496
rect 9048 16250 9076 16487
rect 9036 16244 9088 16250
rect 9036 16186 9088 16192
rect 8944 12232 8996 12238
rect 8944 12174 8996 12180
rect 9128 7744 9180 7750
rect 9128 7686 9180 7692
rect 9140 5234 9168 7686
rect 9128 5228 9180 5234
rect 9128 5170 9180 5176
rect 9324 3194 9352 20742
rect 9508 15638 9536 21966
rect 9496 15632 9548 15638
rect 9496 15574 9548 15580
rect 9600 9382 9628 37402
rect 9692 34950 9720 42502
rect 9784 42158 9812 43794
rect 9772 42152 9824 42158
rect 9772 42094 9824 42100
rect 9784 37466 9812 42094
rect 9772 37460 9824 37466
rect 9772 37402 9824 37408
rect 9772 36712 9824 36718
rect 9772 36654 9824 36660
rect 9784 36242 9812 36654
rect 9772 36236 9824 36242
rect 9772 36178 9824 36184
rect 9876 36174 9904 52974
rect 9864 36168 9916 36174
rect 9864 36110 9916 36116
rect 9772 35828 9824 35834
rect 9772 35770 9824 35776
rect 9680 34944 9732 34950
rect 9680 34886 9732 34892
rect 9784 28626 9812 35770
rect 9772 28620 9824 28626
rect 9772 28562 9824 28568
rect 9864 28484 9916 28490
rect 9864 28426 9916 28432
rect 9680 25832 9732 25838
rect 9680 25774 9732 25780
rect 9692 21078 9720 25774
rect 9770 24848 9826 24857
rect 9770 24783 9772 24792
rect 9824 24783 9826 24792
rect 9772 24754 9824 24760
rect 9876 22642 9904 28426
rect 9864 22636 9916 22642
rect 9864 22578 9916 22584
rect 9772 22160 9824 22166
rect 9772 22102 9824 22108
rect 9680 21072 9732 21078
rect 9680 21014 9732 21020
rect 9784 16250 9812 22102
rect 9772 16244 9824 16250
rect 9772 16186 9824 16192
rect 9784 15706 9812 16186
rect 9772 15700 9824 15706
rect 9772 15642 9824 15648
rect 9588 9376 9640 9382
rect 9588 9318 9640 9324
rect 9968 6914 9996 63718
rect 10048 57792 10100 57798
rect 10048 57734 10100 57740
rect 10060 48618 10088 57734
rect 10232 55616 10284 55622
rect 10232 55558 10284 55564
rect 10140 53168 10192 53174
rect 10140 53110 10192 53116
rect 10048 48612 10100 48618
rect 10048 48554 10100 48560
rect 10048 48340 10100 48346
rect 10048 48282 10100 48288
rect 10060 36417 10088 48282
rect 10046 36408 10102 36417
rect 10046 36343 10102 36352
rect 10060 36038 10088 36343
rect 10048 36032 10100 36038
rect 10048 35974 10100 35980
rect 10152 34746 10180 53110
rect 10244 48822 10272 55558
rect 10232 48816 10284 48822
rect 10232 48758 10284 48764
rect 10232 48612 10284 48618
rect 10232 48554 10284 48560
rect 10244 36378 10272 48554
rect 10232 36372 10284 36378
rect 10232 36314 10284 36320
rect 10336 35018 10364 74394
rect 10508 74180 10560 74186
rect 10508 74122 10560 74128
rect 10520 71126 10548 74122
rect 10508 71120 10560 71126
rect 10508 71062 10560 71068
rect 11060 69216 11112 69222
rect 11060 69158 11112 69164
rect 10508 68672 10560 68678
rect 10508 68614 10560 68620
rect 10416 67856 10468 67862
rect 10416 67798 10468 67804
rect 10428 55350 10456 67798
rect 10520 67697 10548 68614
rect 10506 67688 10562 67697
rect 10506 67623 10562 67632
rect 10968 60580 11020 60586
rect 10968 60522 11020 60528
rect 10508 60240 10560 60246
rect 10508 60182 10560 60188
rect 10416 55344 10468 55350
rect 10416 55286 10468 55292
rect 10416 53032 10468 53038
rect 10416 52974 10468 52980
rect 10428 51474 10456 52974
rect 10416 51468 10468 51474
rect 10416 51410 10468 51416
rect 10520 47666 10548 60182
rect 10784 60172 10836 60178
rect 10784 60114 10836 60120
rect 10600 54188 10652 54194
rect 10600 54130 10652 54136
rect 10612 52465 10640 54130
rect 10796 54126 10824 60114
rect 10980 55826 11008 60522
rect 10968 55820 11020 55826
rect 10968 55762 11020 55768
rect 10980 55214 11008 55762
rect 10888 55186 11008 55214
rect 10784 54120 10836 54126
rect 10784 54062 10836 54068
rect 10888 52902 10916 55186
rect 11072 54330 11100 69158
rect 11520 65612 11572 65618
rect 11520 65554 11572 65560
rect 11428 65476 11480 65482
rect 11428 65418 11480 65424
rect 11336 64388 11388 64394
rect 11336 64330 11388 64336
rect 11244 63980 11296 63986
rect 11244 63922 11296 63928
rect 11152 63028 11204 63034
rect 11152 62970 11204 62976
rect 11164 62422 11192 62970
rect 11152 62416 11204 62422
rect 11152 62358 11204 62364
rect 11060 54324 11112 54330
rect 11060 54266 11112 54272
rect 11060 54188 11112 54194
rect 11060 54130 11112 54136
rect 10968 54120 11020 54126
rect 10968 54062 11020 54068
rect 10876 52896 10928 52902
rect 10876 52838 10928 52844
rect 10598 52456 10654 52465
rect 10598 52391 10654 52400
rect 10600 51264 10652 51270
rect 10600 51206 10652 51212
rect 10508 47660 10560 47666
rect 10508 47602 10560 47608
rect 10612 44198 10640 51206
rect 10692 50924 10744 50930
rect 10692 50866 10744 50872
rect 10704 50726 10732 50866
rect 10692 50720 10744 50726
rect 10690 50688 10692 50697
rect 10744 50688 10746 50697
rect 10690 50623 10746 50632
rect 10784 48816 10836 48822
rect 10784 48758 10836 48764
rect 10692 48680 10744 48686
rect 10692 48622 10744 48628
rect 10704 48550 10732 48622
rect 10692 48544 10744 48550
rect 10692 48486 10744 48492
rect 10704 48346 10732 48486
rect 10692 48340 10744 48346
rect 10692 48282 10744 48288
rect 10600 44192 10652 44198
rect 10600 44134 10652 44140
rect 10414 42664 10470 42673
rect 10414 42599 10416 42608
rect 10468 42599 10470 42608
rect 10416 42570 10468 42576
rect 10508 42560 10560 42566
rect 10508 42502 10560 42508
rect 10692 42560 10744 42566
rect 10692 42502 10744 42508
rect 10520 42294 10548 42502
rect 10508 42288 10560 42294
rect 10508 42230 10560 42236
rect 10508 39364 10560 39370
rect 10508 39306 10560 39312
rect 10416 36712 10468 36718
rect 10416 36654 10468 36660
rect 10324 35012 10376 35018
rect 10324 34954 10376 34960
rect 10140 34740 10192 34746
rect 10140 34682 10192 34688
rect 10152 31754 10180 34682
rect 10152 31726 10272 31754
rect 10048 30048 10100 30054
rect 10048 29990 10100 29996
rect 10060 29102 10088 29990
rect 10048 29096 10100 29102
rect 10048 29038 10100 29044
rect 10060 7886 10088 29038
rect 10138 26072 10194 26081
rect 10138 26007 10140 26016
rect 10192 26007 10194 26016
rect 10140 25978 10192 25984
rect 10244 25294 10272 31726
rect 10322 25392 10378 25401
rect 10428 25362 10456 36654
rect 10520 28422 10548 39306
rect 10704 36922 10732 42502
rect 10692 36916 10744 36922
rect 10692 36858 10744 36864
rect 10600 36372 10652 36378
rect 10600 36314 10652 36320
rect 10612 28490 10640 36314
rect 10692 29096 10744 29102
rect 10692 29038 10744 29044
rect 10600 28484 10652 28490
rect 10600 28426 10652 28432
rect 10508 28416 10560 28422
rect 10508 28358 10560 28364
rect 10704 27962 10732 29038
rect 10796 28082 10824 48758
rect 10980 42838 11008 54062
rect 11072 48686 11100 54130
rect 11060 48680 11112 48686
rect 11060 48622 11112 48628
rect 10968 42832 11020 42838
rect 10968 42774 11020 42780
rect 11058 42800 11114 42809
rect 10980 41682 11008 42774
rect 11058 42735 11114 42744
rect 10968 41676 11020 41682
rect 10968 41618 11020 41624
rect 10968 40384 11020 40390
rect 10968 40326 11020 40332
rect 10980 40186 11008 40326
rect 10968 40180 11020 40186
rect 10968 40122 11020 40128
rect 10968 29164 11020 29170
rect 10968 29106 11020 29112
rect 10784 28076 10836 28082
rect 10784 28018 10836 28024
rect 10704 27934 10824 27962
rect 10796 25838 10824 27934
rect 10980 27878 11008 29106
rect 11072 28762 11100 42735
rect 11060 28756 11112 28762
rect 11060 28698 11112 28704
rect 10968 27872 11020 27878
rect 10968 27814 11020 27820
rect 10876 27600 10928 27606
rect 10876 27542 10928 27548
rect 10784 25832 10836 25838
rect 10784 25774 10836 25780
rect 10322 25327 10324 25336
rect 10376 25327 10378 25336
rect 10416 25356 10468 25362
rect 10324 25298 10376 25304
rect 10416 25298 10468 25304
rect 10232 25288 10284 25294
rect 10232 25230 10284 25236
rect 10244 17066 10272 25230
rect 10336 22778 10364 25298
rect 10508 25152 10560 25158
rect 10508 25094 10560 25100
rect 10324 22772 10376 22778
rect 10324 22714 10376 22720
rect 10324 18080 10376 18086
rect 10324 18022 10376 18028
rect 10232 17060 10284 17066
rect 10232 17002 10284 17008
rect 10048 7880 10100 7886
rect 10048 7822 10100 7828
rect 9876 6886 9996 6914
rect 9678 6760 9734 6769
rect 9496 6724 9548 6730
rect 9678 6695 9680 6704
rect 9496 6666 9548 6672
rect 9732 6695 9734 6704
rect 9680 6666 9732 6672
rect 9508 6458 9536 6666
rect 9496 6452 9548 6458
rect 9496 6394 9548 6400
rect 9312 3188 9364 3194
rect 9312 3130 9364 3136
rect 9876 2650 9904 6886
rect 10336 6866 10364 18022
rect 10520 10198 10548 25094
rect 10796 21690 10824 25774
rect 10784 21684 10836 21690
rect 10784 21626 10836 21632
rect 10796 20874 10824 21626
rect 10784 20868 10836 20874
rect 10784 20810 10836 20816
rect 10600 20052 10652 20058
rect 10600 19994 10652 20000
rect 10612 17746 10640 19994
rect 10600 17740 10652 17746
rect 10600 17682 10652 17688
rect 10612 13802 10640 17682
rect 10888 17678 10916 27542
rect 10876 17672 10928 17678
rect 10876 17614 10928 17620
rect 10980 16114 11008 27814
rect 11164 26217 11192 62358
rect 11256 54194 11284 63922
rect 11244 54188 11296 54194
rect 11244 54130 11296 54136
rect 11244 51264 11296 51270
rect 11244 51206 11296 51212
rect 11256 30666 11284 51206
rect 11348 40050 11376 64330
rect 11440 55865 11468 65418
rect 11426 55856 11482 55865
rect 11426 55791 11482 55800
rect 11428 54324 11480 54330
rect 11428 54266 11480 54272
rect 11440 53106 11468 54266
rect 11428 53100 11480 53106
rect 11428 53042 11480 53048
rect 11440 51377 11468 53042
rect 11426 51368 11482 51377
rect 11426 51303 11482 51312
rect 11532 47598 11560 65554
rect 11612 61736 11664 61742
rect 11612 61678 11664 61684
rect 11520 47592 11572 47598
rect 11520 47534 11572 47540
rect 11428 47184 11480 47190
rect 11428 47126 11480 47132
rect 11336 40044 11388 40050
rect 11336 39986 11388 39992
rect 11336 38208 11388 38214
rect 11336 38150 11388 38156
rect 11348 32026 11376 38150
rect 11440 35766 11468 47126
rect 11532 44810 11560 47534
rect 11520 44804 11572 44810
rect 11520 44746 11572 44752
rect 11624 42809 11652 61678
rect 11716 55894 11744 76230
rect 12610 76188 12918 76197
rect 12610 76186 12616 76188
rect 12672 76186 12696 76188
rect 12752 76186 12776 76188
rect 12832 76186 12856 76188
rect 12912 76186 12918 76188
rect 12672 76134 12674 76186
rect 12854 76134 12856 76186
rect 12610 76132 12616 76134
rect 12672 76132 12696 76134
rect 12752 76132 12776 76134
rect 12832 76132 12856 76134
rect 12912 76132 12918 76134
rect 12610 76123 12918 76132
rect 12440 76016 12492 76022
rect 12440 75958 12492 75964
rect 11950 75644 12258 75653
rect 11950 75642 11956 75644
rect 12012 75642 12036 75644
rect 12092 75642 12116 75644
rect 12172 75642 12196 75644
rect 12252 75642 12258 75644
rect 12012 75590 12014 75642
rect 12194 75590 12196 75642
rect 11950 75588 11956 75590
rect 12012 75588 12036 75590
rect 12092 75588 12116 75590
rect 12172 75588 12196 75590
rect 12252 75588 12258 75590
rect 11950 75579 12258 75588
rect 11796 75404 11848 75410
rect 11796 75346 11848 75352
rect 11808 67318 11836 75346
rect 11950 74556 12258 74565
rect 11950 74554 11956 74556
rect 12012 74554 12036 74556
rect 12092 74554 12116 74556
rect 12172 74554 12196 74556
rect 12252 74554 12258 74556
rect 12012 74502 12014 74554
rect 12194 74502 12196 74554
rect 11950 74500 11956 74502
rect 12012 74500 12036 74502
rect 12092 74500 12116 74502
rect 12172 74500 12196 74502
rect 12252 74500 12258 74502
rect 11950 74491 12258 74500
rect 12452 74118 12480 75958
rect 14096 75948 14148 75954
rect 14096 75890 14148 75896
rect 14188 75948 14240 75954
rect 14188 75890 14240 75896
rect 13728 75744 13780 75750
rect 13728 75686 13780 75692
rect 12610 75100 12918 75109
rect 12610 75098 12616 75100
rect 12672 75098 12696 75100
rect 12752 75098 12776 75100
rect 12832 75098 12856 75100
rect 12912 75098 12918 75100
rect 12672 75046 12674 75098
rect 12854 75046 12856 75098
rect 12610 75044 12616 75046
rect 12672 75044 12696 75046
rect 12752 75044 12776 75046
rect 12832 75044 12856 75046
rect 12912 75044 12918 75046
rect 12610 75035 12918 75044
rect 13740 74534 13768 75686
rect 14108 75274 14136 75890
rect 14096 75268 14148 75274
rect 14096 75210 14148 75216
rect 13556 74506 13768 74534
rect 12440 74112 12492 74118
rect 12440 74054 12492 74060
rect 13452 74112 13504 74118
rect 13452 74054 13504 74060
rect 11950 73468 12258 73477
rect 11950 73466 11956 73468
rect 12012 73466 12036 73468
rect 12092 73466 12116 73468
rect 12172 73466 12196 73468
rect 12252 73466 12258 73468
rect 12012 73414 12014 73466
rect 12194 73414 12196 73466
rect 11950 73412 11956 73414
rect 12012 73412 12036 73414
rect 12092 73412 12116 73414
rect 12172 73412 12196 73414
rect 12252 73412 12258 73414
rect 11950 73403 12258 73412
rect 12348 72684 12400 72690
rect 12348 72626 12400 72632
rect 11950 72380 12258 72389
rect 11950 72378 11956 72380
rect 12012 72378 12036 72380
rect 12092 72378 12116 72380
rect 12172 72378 12196 72380
rect 12252 72378 12258 72380
rect 12012 72326 12014 72378
rect 12194 72326 12196 72378
rect 11950 72324 11956 72326
rect 12012 72324 12036 72326
rect 12092 72324 12116 72326
rect 12172 72324 12196 72326
rect 12252 72324 12258 72326
rect 11950 72315 12258 72324
rect 11950 71292 12258 71301
rect 11950 71290 11956 71292
rect 12012 71290 12036 71292
rect 12092 71290 12116 71292
rect 12172 71290 12196 71292
rect 12252 71290 12258 71292
rect 12012 71238 12014 71290
rect 12194 71238 12196 71290
rect 11950 71236 11956 71238
rect 12012 71236 12036 71238
rect 12092 71236 12116 71238
rect 12172 71236 12196 71238
rect 12252 71236 12258 71238
rect 11950 71227 12258 71236
rect 11950 70204 12258 70213
rect 11950 70202 11956 70204
rect 12012 70202 12036 70204
rect 12092 70202 12116 70204
rect 12172 70202 12196 70204
rect 12252 70202 12258 70204
rect 12012 70150 12014 70202
rect 12194 70150 12196 70202
rect 11950 70148 11956 70150
rect 12012 70148 12036 70150
rect 12092 70148 12116 70150
rect 12172 70148 12196 70150
rect 12252 70148 12258 70150
rect 11950 70139 12258 70148
rect 11950 69116 12258 69125
rect 11950 69114 11956 69116
rect 12012 69114 12036 69116
rect 12092 69114 12116 69116
rect 12172 69114 12196 69116
rect 12252 69114 12258 69116
rect 12012 69062 12014 69114
rect 12194 69062 12196 69114
rect 11950 69060 11956 69062
rect 12012 69060 12036 69062
rect 12092 69060 12116 69062
rect 12172 69060 12196 69062
rect 12252 69060 12258 69062
rect 11950 69051 12258 69060
rect 11950 68028 12258 68037
rect 11950 68026 11956 68028
rect 12012 68026 12036 68028
rect 12092 68026 12116 68028
rect 12172 68026 12196 68028
rect 12252 68026 12258 68028
rect 12012 67974 12014 68026
rect 12194 67974 12196 68026
rect 11950 67972 11956 67974
rect 12012 67972 12036 67974
rect 12092 67972 12116 67974
rect 12172 67972 12196 67974
rect 12252 67972 12258 67974
rect 11950 67963 12258 67972
rect 12070 67688 12126 67697
rect 12070 67623 12072 67632
rect 12124 67623 12126 67632
rect 12072 67594 12124 67600
rect 11796 67312 11848 67318
rect 11796 67254 11848 67260
rect 11808 65686 11836 67254
rect 11950 66940 12258 66949
rect 11950 66938 11956 66940
rect 12012 66938 12036 66940
rect 12092 66938 12116 66940
rect 12172 66938 12196 66940
rect 12252 66938 12258 66940
rect 12012 66886 12014 66938
rect 12194 66886 12196 66938
rect 11950 66884 11956 66886
rect 12012 66884 12036 66886
rect 12092 66884 12116 66886
rect 12172 66884 12196 66886
rect 12252 66884 12258 66886
rect 11950 66875 12258 66884
rect 11950 65852 12258 65861
rect 11950 65850 11956 65852
rect 12012 65850 12036 65852
rect 12092 65850 12116 65852
rect 12172 65850 12196 65852
rect 12252 65850 12258 65852
rect 12012 65798 12014 65850
rect 12194 65798 12196 65850
rect 11950 65796 11956 65798
rect 12012 65796 12036 65798
rect 12092 65796 12116 65798
rect 12172 65796 12196 65798
rect 12252 65796 12258 65798
rect 11950 65787 12258 65796
rect 11796 65680 11848 65686
rect 11796 65622 11848 65628
rect 11796 65544 11848 65550
rect 11796 65486 11848 65492
rect 11888 65544 11940 65550
rect 11888 65486 11940 65492
rect 11808 62422 11836 65486
rect 11900 64938 11928 65486
rect 11888 64932 11940 64938
rect 11888 64874 11940 64880
rect 11950 64764 12258 64773
rect 11950 64762 11956 64764
rect 12012 64762 12036 64764
rect 12092 64762 12116 64764
rect 12172 64762 12196 64764
rect 12252 64762 12258 64764
rect 12012 64710 12014 64762
rect 12194 64710 12196 64762
rect 11950 64708 11956 64710
rect 12012 64708 12036 64710
rect 12092 64708 12116 64710
rect 12172 64708 12196 64710
rect 12252 64708 12258 64710
rect 11950 64699 12258 64708
rect 11950 63676 12258 63685
rect 11950 63674 11956 63676
rect 12012 63674 12036 63676
rect 12092 63674 12116 63676
rect 12172 63674 12196 63676
rect 12252 63674 12258 63676
rect 12012 63622 12014 63674
rect 12194 63622 12196 63674
rect 11950 63620 11956 63622
rect 12012 63620 12036 63622
rect 12092 63620 12116 63622
rect 12172 63620 12196 63622
rect 12252 63620 12258 63622
rect 11950 63611 12258 63620
rect 11950 62588 12258 62597
rect 11950 62586 11956 62588
rect 12012 62586 12036 62588
rect 12092 62586 12116 62588
rect 12172 62586 12196 62588
rect 12252 62586 12258 62588
rect 12012 62534 12014 62586
rect 12194 62534 12196 62586
rect 11950 62532 11956 62534
rect 12012 62532 12036 62534
rect 12092 62532 12116 62534
rect 12172 62532 12196 62534
rect 12252 62532 12258 62534
rect 11950 62523 12258 62532
rect 11796 62416 11848 62422
rect 11796 62358 11848 62364
rect 12360 61810 12388 72626
rect 12452 71738 12480 74054
rect 12610 74012 12918 74021
rect 12610 74010 12616 74012
rect 12672 74010 12696 74012
rect 12752 74010 12776 74012
rect 12832 74010 12856 74012
rect 12912 74010 12918 74012
rect 12672 73958 12674 74010
rect 12854 73958 12856 74010
rect 12610 73956 12616 73958
rect 12672 73956 12696 73958
rect 12752 73956 12776 73958
rect 12832 73956 12856 73958
rect 12912 73956 12918 73958
rect 12610 73947 12918 73956
rect 12610 72924 12918 72933
rect 12610 72922 12616 72924
rect 12672 72922 12696 72924
rect 12752 72922 12776 72924
rect 12832 72922 12856 72924
rect 12912 72922 12918 72924
rect 12672 72870 12674 72922
rect 12854 72870 12856 72922
rect 12610 72868 12616 72870
rect 12672 72868 12696 72870
rect 12752 72868 12776 72870
rect 12832 72868 12856 72870
rect 12912 72868 12918 72870
rect 12610 72859 12918 72868
rect 13268 72480 13320 72486
rect 13268 72422 13320 72428
rect 12610 71836 12918 71845
rect 12610 71834 12616 71836
rect 12672 71834 12696 71836
rect 12752 71834 12776 71836
rect 12832 71834 12856 71836
rect 12912 71834 12918 71836
rect 12672 71782 12674 71834
rect 12854 71782 12856 71834
rect 12610 71780 12616 71782
rect 12672 71780 12696 71782
rect 12752 71780 12776 71782
rect 12832 71780 12856 71782
rect 12912 71780 12918 71782
rect 12610 71771 12918 71780
rect 12440 71732 12492 71738
rect 12440 71674 12492 71680
rect 12610 70748 12918 70757
rect 12610 70746 12616 70748
rect 12672 70746 12696 70748
rect 12752 70746 12776 70748
rect 12832 70746 12856 70748
rect 12912 70746 12918 70748
rect 12672 70694 12674 70746
rect 12854 70694 12856 70746
rect 12610 70692 12616 70694
rect 12672 70692 12696 70694
rect 12752 70692 12776 70694
rect 12832 70692 12856 70694
rect 12912 70692 12918 70694
rect 12610 70683 12918 70692
rect 12440 69964 12492 69970
rect 12440 69906 12492 69912
rect 12452 65006 12480 69906
rect 12610 69660 12918 69669
rect 12610 69658 12616 69660
rect 12672 69658 12696 69660
rect 12752 69658 12776 69660
rect 12832 69658 12856 69660
rect 12912 69658 12918 69660
rect 12672 69606 12674 69658
rect 12854 69606 12856 69658
rect 12610 69604 12616 69606
rect 12672 69604 12696 69606
rect 12752 69604 12776 69606
rect 12832 69604 12856 69606
rect 12912 69604 12918 69606
rect 12610 69595 12918 69604
rect 13176 69556 13228 69562
rect 13176 69498 13228 69504
rect 12610 68572 12918 68581
rect 12610 68570 12616 68572
rect 12672 68570 12696 68572
rect 12752 68570 12776 68572
rect 12832 68570 12856 68572
rect 12912 68570 12918 68572
rect 12672 68518 12674 68570
rect 12854 68518 12856 68570
rect 12610 68516 12616 68518
rect 12672 68516 12696 68518
rect 12752 68516 12776 68518
rect 12832 68516 12856 68518
rect 12912 68516 12918 68518
rect 12610 68507 12918 68516
rect 12610 67484 12918 67493
rect 12610 67482 12616 67484
rect 12672 67482 12696 67484
rect 12752 67482 12776 67484
rect 12832 67482 12856 67484
rect 12912 67482 12918 67484
rect 12672 67430 12674 67482
rect 12854 67430 12856 67482
rect 12610 67428 12616 67430
rect 12672 67428 12696 67430
rect 12752 67428 12776 67430
rect 12832 67428 12856 67430
rect 12912 67428 12918 67430
rect 12610 67419 12918 67428
rect 12610 66396 12918 66405
rect 12610 66394 12616 66396
rect 12672 66394 12696 66396
rect 12752 66394 12776 66396
rect 12832 66394 12856 66396
rect 12912 66394 12918 66396
rect 12672 66342 12674 66394
rect 12854 66342 12856 66394
rect 12610 66340 12616 66342
rect 12672 66340 12696 66342
rect 12752 66340 12776 66342
rect 12832 66340 12856 66342
rect 12912 66340 12918 66342
rect 12610 66331 12918 66340
rect 12610 65308 12918 65317
rect 12610 65306 12616 65308
rect 12672 65306 12696 65308
rect 12752 65306 12776 65308
rect 12832 65306 12856 65308
rect 12912 65306 12918 65308
rect 12672 65254 12674 65306
rect 12854 65254 12856 65306
rect 12610 65252 12616 65254
rect 12672 65252 12696 65254
rect 12752 65252 12776 65254
rect 12832 65252 12856 65254
rect 12912 65252 12918 65254
rect 12610 65243 12918 65252
rect 12440 65000 12492 65006
rect 12440 64942 12492 64948
rect 12610 64220 12918 64229
rect 12610 64218 12616 64220
rect 12672 64218 12696 64220
rect 12752 64218 12776 64220
rect 12832 64218 12856 64220
rect 12912 64218 12918 64220
rect 12672 64166 12674 64218
rect 12854 64166 12856 64218
rect 12610 64164 12616 64166
rect 12672 64164 12696 64166
rect 12752 64164 12776 64166
rect 12832 64164 12856 64166
rect 12912 64164 12918 64166
rect 12610 64155 12918 64164
rect 12610 63132 12918 63141
rect 12610 63130 12616 63132
rect 12672 63130 12696 63132
rect 12752 63130 12776 63132
rect 12832 63130 12856 63132
rect 12912 63130 12918 63132
rect 12672 63078 12674 63130
rect 12854 63078 12856 63130
rect 12610 63076 12616 63078
rect 12672 63076 12696 63078
rect 12752 63076 12776 63078
rect 12832 63076 12856 63078
rect 12912 63076 12918 63078
rect 12610 63067 12918 63076
rect 12610 62044 12918 62053
rect 12610 62042 12616 62044
rect 12672 62042 12696 62044
rect 12752 62042 12776 62044
rect 12832 62042 12856 62044
rect 12912 62042 12918 62044
rect 12672 61990 12674 62042
rect 12854 61990 12856 62042
rect 12610 61988 12616 61990
rect 12672 61988 12696 61990
rect 12752 61988 12776 61990
rect 12832 61988 12856 61990
rect 12912 61988 12918 61990
rect 12610 61979 12918 61988
rect 12348 61804 12400 61810
rect 12348 61746 12400 61752
rect 11950 61500 12258 61509
rect 11950 61498 11956 61500
rect 12012 61498 12036 61500
rect 12092 61498 12116 61500
rect 12172 61498 12196 61500
rect 12252 61498 12258 61500
rect 12012 61446 12014 61498
rect 12194 61446 12196 61498
rect 11950 61444 11956 61446
rect 12012 61444 12036 61446
rect 12092 61444 12116 61446
rect 12172 61444 12196 61446
rect 12252 61444 12258 61446
rect 11950 61435 12258 61444
rect 12610 60956 12918 60965
rect 12610 60954 12616 60956
rect 12672 60954 12696 60956
rect 12752 60954 12776 60956
rect 12832 60954 12856 60956
rect 12912 60954 12918 60956
rect 12672 60902 12674 60954
rect 12854 60902 12856 60954
rect 12610 60900 12616 60902
rect 12672 60900 12696 60902
rect 12752 60900 12776 60902
rect 12832 60900 12856 60902
rect 12912 60900 12918 60902
rect 12610 60891 12918 60900
rect 11950 60412 12258 60421
rect 11950 60410 11956 60412
rect 12012 60410 12036 60412
rect 12092 60410 12116 60412
rect 12172 60410 12196 60412
rect 12252 60410 12258 60412
rect 12012 60358 12014 60410
rect 12194 60358 12196 60410
rect 11950 60356 11956 60358
rect 12012 60356 12036 60358
rect 12092 60356 12116 60358
rect 12172 60356 12196 60358
rect 12252 60356 12258 60358
rect 11950 60347 12258 60356
rect 13188 60314 13216 69498
rect 13280 64666 13308 72422
rect 13268 64660 13320 64666
rect 13268 64602 13320 64608
rect 13176 60308 13228 60314
rect 13176 60250 13228 60256
rect 13084 60036 13136 60042
rect 13084 59978 13136 59984
rect 12610 59868 12918 59877
rect 12610 59866 12616 59868
rect 12672 59866 12696 59868
rect 12752 59866 12776 59868
rect 12832 59866 12856 59868
rect 12912 59866 12918 59868
rect 12672 59814 12674 59866
rect 12854 59814 12856 59866
rect 12610 59812 12616 59814
rect 12672 59812 12696 59814
rect 12752 59812 12776 59814
rect 12832 59812 12856 59814
rect 12912 59812 12918 59814
rect 12610 59803 12918 59812
rect 11950 59324 12258 59333
rect 11950 59322 11956 59324
rect 12012 59322 12036 59324
rect 12092 59322 12116 59324
rect 12172 59322 12196 59324
rect 12252 59322 12258 59324
rect 12012 59270 12014 59322
rect 12194 59270 12196 59322
rect 11950 59268 11956 59270
rect 12012 59268 12036 59270
rect 12092 59268 12116 59270
rect 12172 59268 12196 59270
rect 12252 59268 12258 59270
rect 11950 59259 12258 59268
rect 12610 58780 12918 58789
rect 12610 58778 12616 58780
rect 12672 58778 12696 58780
rect 12752 58778 12776 58780
rect 12832 58778 12856 58780
rect 12912 58778 12918 58780
rect 12672 58726 12674 58778
rect 12854 58726 12856 58778
rect 12610 58724 12616 58726
rect 12672 58724 12696 58726
rect 12752 58724 12776 58726
rect 12832 58724 12856 58726
rect 12912 58724 12918 58726
rect 12610 58715 12918 58724
rect 11950 58236 12258 58245
rect 11950 58234 11956 58236
rect 12012 58234 12036 58236
rect 12092 58234 12116 58236
rect 12172 58234 12196 58236
rect 12252 58234 12258 58236
rect 12012 58182 12014 58234
rect 12194 58182 12196 58234
rect 11950 58180 11956 58182
rect 12012 58180 12036 58182
rect 12092 58180 12116 58182
rect 12172 58180 12196 58182
rect 12252 58180 12258 58182
rect 11950 58171 12258 58180
rect 12610 57692 12918 57701
rect 12610 57690 12616 57692
rect 12672 57690 12696 57692
rect 12752 57690 12776 57692
rect 12832 57690 12856 57692
rect 12912 57690 12918 57692
rect 12672 57638 12674 57690
rect 12854 57638 12856 57690
rect 12610 57636 12616 57638
rect 12672 57636 12696 57638
rect 12752 57636 12776 57638
rect 12832 57636 12856 57638
rect 12912 57636 12918 57638
rect 12610 57627 12918 57636
rect 11950 57148 12258 57157
rect 11950 57146 11956 57148
rect 12012 57146 12036 57148
rect 12092 57146 12116 57148
rect 12172 57146 12196 57148
rect 12252 57146 12258 57148
rect 12012 57094 12014 57146
rect 12194 57094 12196 57146
rect 11950 57092 11956 57094
rect 12012 57092 12036 57094
rect 12092 57092 12116 57094
rect 12172 57092 12196 57094
rect 12252 57092 12258 57094
rect 11950 57083 12258 57092
rect 12610 56604 12918 56613
rect 12610 56602 12616 56604
rect 12672 56602 12696 56604
rect 12752 56602 12776 56604
rect 12832 56602 12856 56604
rect 12912 56602 12918 56604
rect 12672 56550 12674 56602
rect 12854 56550 12856 56602
rect 12610 56548 12616 56550
rect 12672 56548 12696 56550
rect 12752 56548 12776 56550
rect 12832 56548 12856 56550
rect 12912 56548 12918 56550
rect 12610 56539 12918 56548
rect 12440 56296 12492 56302
rect 12440 56238 12492 56244
rect 12992 56296 13044 56302
rect 12992 56238 13044 56244
rect 11950 56060 12258 56069
rect 11950 56058 11956 56060
rect 12012 56058 12036 56060
rect 12092 56058 12116 56060
rect 12172 56058 12196 56060
rect 12252 56058 12258 56060
rect 12012 56006 12014 56058
rect 12194 56006 12196 56058
rect 11950 56004 11956 56006
rect 12012 56004 12036 56006
rect 12092 56004 12116 56006
rect 12172 56004 12196 56006
rect 12252 56004 12258 56006
rect 11950 55995 12258 56004
rect 11704 55888 11756 55894
rect 11704 55830 11756 55836
rect 11704 55752 11756 55758
rect 12452 55729 12480 56238
rect 11704 55694 11756 55700
rect 12438 55720 12494 55729
rect 11716 44878 11744 55694
rect 12438 55655 12494 55664
rect 12610 55516 12918 55525
rect 12610 55514 12616 55516
rect 12672 55514 12696 55516
rect 12752 55514 12776 55516
rect 12832 55514 12856 55516
rect 12912 55514 12918 55516
rect 12672 55462 12674 55514
rect 12854 55462 12856 55514
rect 12610 55460 12616 55462
rect 12672 55460 12696 55462
rect 12752 55460 12776 55462
rect 12832 55460 12856 55462
rect 12912 55460 12918 55462
rect 12610 55451 12918 55460
rect 11950 54972 12258 54981
rect 11950 54970 11956 54972
rect 12012 54970 12036 54972
rect 12092 54970 12116 54972
rect 12172 54970 12196 54972
rect 12252 54970 12258 54972
rect 12012 54918 12014 54970
rect 12194 54918 12196 54970
rect 11950 54916 11956 54918
rect 12012 54916 12036 54918
rect 12092 54916 12116 54918
rect 12172 54916 12196 54918
rect 12252 54916 12258 54918
rect 11950 54907 12258 54916
rect 12610 54428 12918 54437
rect 12610 54426 12616 54428
rect 12672 54426 12696 54428
rect 12752 54426 12776 54428
rect 12832 54426 12856 54428
rect 12912 54426 12918 54428
rect 12672 54374 12674 54426
rect 12854 54374 12856 54426
rect 12610 54372 12616 54374
rect 12672 54372 12696 54374
rect 12752 54372 12776 54374
rect 12832 54372 12856 54374
rect 12912 54372 12918 54374
rect 12610 54363 12918 54372
rect 12440 54188 12492 54194
rect 12440 54130 12492 54136
rect 12452 54097 12480 54130
rect 12438 54088 12494 54097
rect 12438 54023 12494 54032
rect 12532 53984 12584 53990
rect 12532 53926 12584 53932
rect 11950 53884 12258 53893
rect 11950 53882 11956 53884
rect 12012 53882 12036 53884
rect 12092 53882 12116 53884
rect 12172 53882 12196 53884
rect 12252 53882 12258 53884
rect 12012 53830 12014 53882
rect 12194 53830 12196 53882
rect 11950 53828 11956 53830
rect 12012 53828 12036 53830
rect 12092 53828 12116 53830
rect 12172 53828 12196 53830
rect 12252 53828 12258 53830
rect 11950 53819 12258 53828
rect 11950 52796 12258 52805
rect 11950 52794 11956 52796
rect 12012 52794 12036 52796
rect 12092 52794 12116 52796
rect 12172 52794 12196 52796
rect 12252 52794 12258 52796
rect 12012 52742 12014 52794
rect 12194 52742 12196 52794
rect 11950 52740 11956 52742
rect 12012 52740 12036 52742
rect 12092 52740 12116 52742
rect 12172 52740 12196 52742
rect 12252 52740 12258 52742
rect 11950 52731 12258 52740
rect 11950 51708 12258 51717
rect 11950 51706 11956 51708
rect 12012 51706 12036 51708
rect 12092 51706 12116 51708
rect 12172 51706 12196 51708
rect 12252 51706 12258 51708
rect 12012 51654 12014 51706
rect 12194 51654 12196 51706
rect 11950 51652 11956 51654
rect 12012 51652 12036 51654
rect 12092 51652 12116 51654
rect 12172 51652 12196 51654
rect 12252 51652 12258 51654
rect 11950 51643 12258 51652
rect 11950 50620 12258 50629
rect 11950 50618 11956 50620
rect 12012 50618 12036 50620
rect 12092 50618 12116 50620
rect 12172 50618 12196 50620
rect 12252 50618 12258 50620
rect 12012 50566 12014 50618
rect 12194 50566 12196 50618
rect 11950 50564 11956 50566
rect 12012 50564 12036 50566
rect 12092 50564 12116 50566
rect 12172 50564 12196 50566
rect 12252 50564 12258 50566
rect 11950 50555 12258 50564
rect 11950 49532 12258 49541
rect 11950 49530 11956 49532
rect 12012 49530 12036 49532
rect 12092 49530 12116 49532
rect 12172 49530 12196 49532
rect 12252 49530 12258 49532
rect 12012 49478 12014 49530
rect 12194 49478 12196 49530
rect 11950 49476 11956 49478
rect 12012 49476 12036 49478
rect 12092 49476 12116 49478
rect 12172 49476 12196 49478
rect 12252 49476 12258 49478
rect 11950 49467 12258 49476
rect 11950 48444 12258 48453
rect 11950 48442 11956 48444
rect 12012 48442 12036 48444
rect 12092 48442 12116 48444
rect 12172 48442 12196 48444
rect 12252 48442 12258 48444
rect 12012 48390 12014 48442
rect 12194 48390 12196 48442
rect 11950 48388 11956 48390
rect 12012 48388 12036 48390
rect 12092 48388 12116 48390
rect 12172 48388 12196 48390
rect 12252 48388 12258 48390
rect 11950 48379 12258 48388
rect 12440 47592 12492 47598
rect 12440 47534 12492 47540
rect 11950 47356 12258 47365
rect 11950 47354 11956 47356
rect 12012 47354 12036 47356
rect 12092 47354 12116 47356
rect 12172 47354 12196 47356
rect 12252 47354 12258 47356
rect 12012 47302 12014 47354
rect 12194 47302 12196 47354
rect 11950 47300 11956 47302
rect 12012 47300 12036 47302
rect 12092 47300 12116 47302
rect 12172 47300 12196 47302
rect 12252 47300 12258 47302
rect 11950 47291 12258 47300
rect 12452 46374 12480 47534
rect 12544 46646 12572 53926
rect 12610 53340 12918 53349
rect 12610 53338 12616 53340
rect 12672 53338 12696 53340
rect 12752 53338 12776 53340
rect 12832 53338 12856 53340
rect 12912 53338 12918 53340
rect 12672 53286 12674 53338
rect 12854 53286 12856 53338
rect 12610 53284 12616 53286
rect 12672 53284 12696 53286
rect 12752 53284 12776 53286
rect 12832 53284 12856 53286
rect 12912 53284 12918 53286
rect 12610 53275 12918 53284
rect 12610 52252 12918 52261
rect 12610 52250 12616 52252
rect 12672 52250 12696 52252
rect 12752 52250 12776 52252
rect 12832 52250 12856 52252
rect 12912 52250 12918 52252
rect 12672 52198 12674 52250
rect 12854 52198 12856 52250
rect 12610 52196 12616 52198
rect 12672 52196 12696 52198
rect 12752 52196 12776 52198
rect 12832 52196 12856 52198
rect 12912 52196 12918 52198
rect 12610 52187 12918 52196
rect 12610 51164 12918 51173
rect 12610 51162 12616 51164
rect 12672 51162 12696 51164
rect 12752 51162 12776 51164
rect 12832 51162 12856 51164
rect 12912 51162 12918 51164
rect 12672 51110 12674 51162
rect 12854 51110 12856 51162
rect 12610 51108 12616 51110
rect 12672 51108 12696 51110
rect 12752 51108 12776 51110
rect 12832 51108 12856 51110
rect 12912 51108 12918 51110
rect 12610 51099 12918 51108
rect 12610 50076 12918 50085
rect 12610 50074 12616 50076
rect 12672 50074 12696 50076
rect 12752 50074 12776 50076
rect 12832 50074 12856 50076
rect 12912 50074 12918 50076
rect 12672 50022 12674 50074
rect 12854 50022 12856 50074
rect 12610 50020 12616 50022
rect 12672 50020 12696 50022
rect 12752 50020 12776 50022
rect 12832 50020 12856 50022
rect 12912 50020 12918 50022
rect 12610 50011 12918 50020
rect 12610 48988 12918 48997
rect 12610 48986 12616 48988
rect 12672 48986 12696 48988
rect 12752 48986 12776 48988
rect 12832 48986 12856 48988
rect 12912 48986 12918 48988
rect 12672 48934 12674 48986
rect 12854 48934 12856 48986
rect 12610 48932 12616 48934
rect 12672 48932 12696 48934
rect 12752 48932 12776 48934
rect 12832 48932 12856 48934
rect 12912 48932 12918 48934
rect 12610 48923 12918 48932
rect 12610 47900 12918 47909
rect 12610 47898 12616 47900
rect 12672 47898 12696 47900
rect 12752 47898 12776 47900
rect 12832 47898 12856 47900
rect 12912 47898 12918 47900
rect 12672 47846 12674 47898
rect 12854 47846 12856 47898
rect 12610 47844 12616 47846
rect 12672 47844 12696 47846
rect 12752 47844 12776 47846
rect 12832 47844 12856 47846
rect 12912 47844 12918 47846
rect 12610 47835 12918 47844
rect 12610 46812 12918 46821
rect 12610 46810 12616 46812
rect 12672 46810 12696 46812
rect 12752 46810 12776 46812
rect 12832 46810 12856 46812
rect 12912 46810 12918 46812
rect 12672 46758 12674 46810
rect 12854 46758 12856 46810
rect 12610 46756 12616 46758
rect 12672 46756 12696 46758
rect 12752 46756 12776 46758
rect 12832 46756 12856 46758
rect 12912 46756 12918 46758
rect 12610 46747 12918 46756
rect 12532 46640 12584 46646
rect 12532 46582 12584 46588
rect 12440 46368 12492 46374
rect 12440 46310 12492 46316
rect 11950 46268 12258 46277
rect 11950 46266 11956 46268
rect 12012 46266 12036 46268
rect 12092 46266 12116 46268
rect 12172 46266 12196 46268
rect 12252 46266 12258 46268
rect 12012 46214 12014 46266
rect 12194 46214 12196 46266
rect 11950 46212 11956 46214
rect 12012 46212 12036 46214
rect 12092 46212 12116 46214
rect 12172 46212 12196 46214
rect 12252 46212 12258 46214
rect 11950 46203 12258 46212
rect 12452 45626 12480 46310
rect 12610 45724 12918 45733
rect 12610 45722 12616 45724
rect 12672 45722 12696 45724
rect 12752 45722 12776 45724
rect 12832 45722 12856 45724
rect 12912 45722 12918 45724
rect 12672 45670 12674 45722
rect 12854 45670 12856 45722
rect 12610 45668 12616 45670
rect 12672 45668 12696 45670
rect 12752 45668 12776 45670
rect 12832 45668 12856 45670
rect 12912 45668 12918 45670
rect 12610 45659 12918 45668
rect 12440 45620 12492 45626
rect 12440 45562 12492 45568
rect 11950 45180 12258 45189
rect 11950 45178 11956 45180
rect 12012 45178 12036 45180
rect 12092 45178 12116 45180
rect 12172 45178 12196 45180
rect 12252 45178 12258 45180
rect 12012 45126 12014 45178
rect 12194 45126 12196 45178
rect 11950 45124 11956 45126
rect 12012 45124 12036 45126
rect 12092 45124 12116 45126
rect 12172 45124 12196 45126
rect 12252 45124 12258 45126
rect 11950 45115 12258 45124
rect 12452 44946 12480 45562
rect 12440 44940 12492 44946
rect 12440 44882 12492 44888
rect 11704 44872 11756 44878
rect 11704 44814 11756 44820
rect 12610 44636 12918 44645
rect 12610 44634 12616 44636
rect 12672 44634 12696 44636
rect 12752 44634 12776 44636
rect 12832 44634 12856 44636
rect 12912 44634 12918 44636
rect 12672 44582 12674 44634
rect 12854 44582 12856 44634
rect 12610 44580 12616 44582
rect 12672 44580 12696 44582
rect 12752 44580 12776 44582
rect 12832 44580 12856 44582
rect 12912 44580 12918 44582
rect 12610 44571 12918 44580
rect 11950 44092 12258 44101
rect 11950 44090 11956 44092
rect 12012 44090 12036 44092
rect 12092 44090 12116 44092
rect 12172 44090 12196 44092
rect 12252 44090 12258 44092
rect 12012 44038 12014 44090
rect 12194 44038 12196 44090
rect 11950 44036 11956 44038
rect 12012 44036 12036 44038
rect 12092 44036 12116 44038
rect 12172 44036 12196 44038
rect 12252 44036 12258 44038
rect 11950 44027 12258 44036
rect 12610 43548 12918 43557
rect 12610 43546 12616 43548
rect 12672 43546 12696 43548
rect 12752 43546 12776 43548
rect 12832 43546 12856 43548
rect 12912 43546 12918 43548
rect 12672 43494 12674 43546
rect 12854 43494 12856 43546
rect 12610 43492 12616 43494
rect 12672 43492 12696 43494
rect 12752 43492 12776 43494
rect 12832 43492 12856 43494
rect 12912 43492 12918 43494
rect 12610 43483 12918 43492
rect 12532 43240 12584 43246
rect 12532 43182 12584 43188
rect 11950 43004 12258 43013
rect 11950 43002 11956 43004
rect 12012 43002 12036 43004
rect 12092 43002 12116 43004
rect 12172 43002 12196 43004
rect 12252 43002 12258 43004
rect 12012 42950 12014 43002
rect 12194 42950 12196 43002
rect 11950 42948 11956 42950
rect 12012 42948 12036 42950
rect 12092 42948 12116 42950
rect 12172 42948 12196 42950
rect 12252 42948 12258 42950
rect 11950 42939 12258 42948
rect 11610 42800 11666 42809
rect 11610 42735 11666 42744
rect 11624 42022 11652 42735
rect 11704 42628 11756 42634
rect 11704 42570 11756 42576
rect 11612 42016 11664 42022
rect 11612 41958 11664 41964
rect 11612 36916 11664 36922
rect 11612 36858 11664 36864
rect 11520 36032 11572 36038
rect 11520 35974 11572 35980
rect 11428 35760 11480 35766
rect 11428 35702 11480 35708
rect 11428 35624 11480 35630
rect 11428 35566 11480 35572
rect 11336 32020 11388 32026
rect 11336 31962 11388 31968
rect 11244 30660 11296 30666
rect 11244 30602 11296 30608
rect 11150 26208 11206 26217
rect 11150 26143 11206 26152
rect 11058 26072 11114 26081
rect 11058 26007 11114 26016
rect 11072 18086 11100 26007
rect 11440 24954 11468 35566
rect 11532 32298 11560 35974
rect 11520 32292 11572 32298
rect 11520 32234 11572 32240
rect 11520 32020 11572 32026
rect 11520 31962 11572 31968
rect 11532 26382 11560 31962
rect 11520 26376 11572 26382
rect 11520 26318 11572 26324
rect 11520 25220 11572 25226
rect 11520 25162 11572 25168
rect 11428 24948 11480 24954
rect 11428 24890 11480 24896
rect 11336 23520 11388 23526
rect 11336 23462 11388 23468
rect 11244 21888 11296 21894
rect 11244 21830 11296 21836
rect 11060 18080 11112 18086
rect 11060 18022 11112 18028
rect 10968 16108 11020 16114
rect 10968 16050 11020 16056
rect 11060 14068 11112 14074
rect 11060 14010 11112 14016
rect 10600 13796 10652 13802
rect 10600 13738 10652 13744
rect 10784 13796 10836 13802
rect 10784 13738 10836 13744
rect 10796 12238 10824 13738
rect 11072 12986 11100 14010
rect 11152 14000 11204 14006
rect 11152 13942 11204 13948
rect 11060 12980 11112 12986
rect 11060 12922 11112 12928
rect 11164 12434 11192 13942
rect 11256 13938 11284 21830
rect 11348 14346 11376 23462
rect 11428 21480 11480 21486
rect 11428 21422 11480 21428
rect 11440 21049 11468 21422
rect 11426 21040 11482 21049
rect 11426 20975 11482 20984
rect 11428 20392 11480 20398
rect 11428 20334 11480 20340
rect 11440 20058 11468 20334
rect 11428 20052 11480 20058
rect 11428 19994 11480 20000
rect 11428 15360 11480 15366
rect 11428 15302 11480 15308
rect 11336 14340 11388 14346
rect 11336 14282 11388 14288
rect 11244 13932 11296 13938
rect 11244 13874 11296 13880
rect 11072 12406 11192 12434
rect 11072 12238 11100 12406
rect 10692 12232 10744 12238
rect 10690 12200 10692 12209
rect 10784 12232 10836 12238
rect 10744 12200 10746 12209
rect 10784 12174 10836 12180
rect 11060 12232 11112 12238
rect 11060 12174 11112 12180
rect 10690 12135 10746 12144
rect 10508 10192 10560 10198
rect 10508 10134 10560 10140
rect 10796 8566 10824 12174
rect 10784 8560 10836 8566
rect 10784 8502 10836 8508
rect 10968 8560 11020 8566
rect 10968 8502 11020 8508
rect 10876 7880 10928 7886
rect 10876 7822 10928 7828
rect 10888 6914 10916 7822
rect 10980 7154 11008 8502
rect 10980 7126 11100 7154
rect 10888 6886 11008 6914
rect 10324 6860 10376 6866
rect 10324 6802 10376 6808
rect 10980 3738 11008 6886
rect 11072 5234 11100 7126
rect 11440 5574 11468 15302
rect 11532 8498 11560 25162
rect 11520 8492 11572 8498
rect 11520 8434 11572 8440
rect 11624 8362 11652 36858
rect 11716 12986 11744 42570
rect 11950 41916 12258 41925
rect 11950 41914 11956 41916
rect 12012 41914 12036 41916
rect 12092 41914 12116 41916
rect 12172 41914 12196 41916
rect 12252 41914 12258 41916
rect 12012 41862 12014 41914
rect 12194 41862 12196 41914
rect 11950 41860 11956 41862
rect 12012 41860 12036 41862
rect 12092 41860 12116 41862
rect 12172 41860 12196 41862
rect 12252 41860 12258 41862
rect 11950 41851 12258 41860
rect 12544 41414 12572 43182
rect 12610 42460 12918 42469
rect 12610 42458 12616 42460
rect 12672 42458 12696 42460
rect 12752 42458 12776 42460
rect 12832 42458 12856 42460
rect 12912 42458 12918 42460
rect 12672 42406 12674 42458
rect 12854 42406 12856 42458
rect 12610 42404 12616 42406
rect 12672 42404 12696 42406
rect 12752 42404 12776 42406
rect 12832 42404 12856 42406
rect 12912 42404 12918 42406
rect 12610 42395 12918 42404
rect 12452 41386 12572 41414
rect 11950 40828 12258 40837
rect 11950 40826 11956 40828
rect 12012 40826 12036 40828
rect 12092 40826 12116 40828
rect 12172 40826 12196 40828
rect 12252 40826 12258 40828
rect 12012 40774 12014 40826
rect 12194 40774 12196 40826
rect 11950 40772 11956 40774
rect 12012 40772 12036 40774
rect 12092 40772 12116 40774
rect 12172 40772 12196 40774
rect 12252 40772 12258 40774
rect 11950 40763 12258 40772
rect 11950 39740 12258 39749
rect 11950 39738 11956 39740
rect 12012 39738 12036 39740
rect 12092 39738 12116 39740
rect 12172 39738 12196 39740
rect 12252 39738 12258 39740
rect 12012 39686 12014 39738
rect 12194 39686 12196 39738
rect 11950 39684 11956 39686
rect 12012 39684 12036 39686
rect 12092 39684 12116 39686
rect 12172 39684 12196 39686
rect 12252 39684 12258 39686
rect 11950 39675 12258 39684
rect 11796 39636 11848 39642
rect 11796 39578 11848 39584
rect 11808 35630 11836 39578
rect 12348 39296 12400 39302
rect 12348 39238 12400 39244
rect 11950 38652 12258 38661
rect 11950 38650 11956 38652
rect 12012 38650 12036 38652
rect 12092 38650 12116 38652
rect 12172 38650 12196 38652
rect 12252 38650 12258 38652
rect 12012 38598 12014 38650
rect 12194 38598 12196 38650
rect 11950 38596 11956 38598
rect 12012 38596 12036 38598
rect 12092 38596 12116 38598
rect 12172 38596 12196 38598
rect 12252 38596 12258 38598
rect 11950 38587 12258 38596
rect 11950 37564 12258 37573
rect 11950 37562 11956 37564
rect 12012 37562 12036 37564
rect 12092 37562 12116 37564
rect 12172 37562 12196 37564
rect 12252 37562 12258 37564
rect 12012 37510 12014 37562
rect 12194 37510 12196 37562
rect 11950 37508 11956 37510
rect 12012 37508 12036 37510
rect 12092 37508 12116 37510
rect 12172 37508 12196 37510
rect 12252 37508 12258 37510
rect 11950 37499 12258 37508
rect 11950 36476 12258 36485
rect 11950 36474 11956 36476
rect 12012 36474 12036 36476
rect 12092 36474 12116 36476
rect 12172 36474 12196 36476
rect 12252 36474 12258 36476
rect 12012 36422 12014 36474
rect 12194 36422 12196 36474
rect 11950 36420 11956 36422
rect 12012 36420 12036 36422
rect 12092 36420 12116 36422
rect 12172 36420 12196 36422
rect 12252 36420 12258 36422
rect 11950 36411 12258 36420
rect 11888 35828 11940 35834
rect 11888 35770 11940 35776
rect 11900 35630 11928 35770
rect 11796 35624 11848 35630
rect 11796 35566 11848 35572
rect 11888 35624 11940 35630
rect 11888 35566 11940 35572
rect 11950 35388 12258 35397
rect 11950 35386 11956 35388
rect 12012 35386 12036 35388
rect 12092 35386 12116 35388
rect 12172 35386 12196 35388
rect 12252 35386 12258 35388
rect 12012 35334 12014 35386
rect 12194 35334 12196 35386
rect 11950 35332 11956 35334
rect 12012 35332 12036 35334
rect 12092 35332 12116 35334
rect 12172 35332 12196 35334
rect 12252 35332 12258 35334
rect 11950 35323 12258 35332
rect 11950 34300 12258 34309
rect 11950 34298 11956 34300
rect 12012 34298 12036 34300
rect 12092 34298 12116 34300
rect 12172 34298 12196 34300
rect 12252 34298 12258 34300
rect 12012 34246 12014 34298
rect 12194 34246 12196 34298
rect 11950 34244 11956 34246
rect 12012 34244 12036 34246
rect 12092 34244 12116 34246
rect 12172 34244 12196 34246
rect 12252 34244 12258 34246
rect 11950 34235 12258 34244
rect 11950 33212 12258 33221
rect 11950 33210 11956 33212
rect 12012 33210 12036 33212
rect 12092 33210 12116 33212
rect 12172 33210 12196 33212
rect 12252 33210 12258 33212
rect 12012 33158 12014 33210
rect 12194 33158 12196 33210
rect 11950 33156 11956 33158
rect 12012 33156 12036 33158
rect 12092 33156 12116 33158
rect 12172 33156 12196 33158
rect 12252 33156 12258 33158
rect 11950 33147 12258 33156
rect 11796 32224 11848 32230
rect 11796 32166 11848 32172
rect 11808 30190 11836 32166
rect 11950 32124 12258 32133
rect 11950 32122 11956 32124
rect 12012 32122 12036 32124
rect 12092 32122 12116 32124
rect 12172 32122 12196 32124
rect 12252 32122 12258 32124
rect 12012 32070 12014 32122
rect 12194 32070 12196 32122
rect 11950 32068 11956 32070
rect 12012 32068 12036 32070
rect 12092 32068 12116 32070
rect 12172 32068 12196 32070
rect 12252 32068 12258 32070
rect 11950 32059 12258 32068
rect 11950 31036 12258 31045
rect 11950 31034 11956 31036
rect 12012 31034 12036 31036
rect 12092 31034 12116 31036
rect 12172 31034 12196 31036
rect 12252 31034 12258 31036
rect 12012 30982 12014 31034
rect 12194 30982 12196 31034
rect 11950 30980 11956 30982
rect 12012 30980 12036 30982
rect 12092 30980 12116 30982
rect 12172 30980 12196 30982
rect 12252 30980 12258 30982
rect 11950 30971 12258 30980
rect 11796 30184 11848 30190
rect 11796 30126 11848 30132
rect 11950 29948 12258 29957
rect 11950 29946 11956 29948
rect 12012 29946 12036 29948
rect 12092 29946 12116 29948
rect 12172 29946 12196 29948
rect 12252 29946 12258 29948
rect 12012 29894 12014 29946
rect 12194 29894 12196 29946
rect 11950 29892 11956 29894
rect 12012 29892 12036 29894
rect 12092 29892 12116 29894
rect 12172 29892 12196 29894
rect 12252 29892 12258 29894
rect 11950 29883 12258 29892
rect 11950 28860 12258 28869
rect 11950 28858 11956 28860
rect 12012 28858 12036 28860
rect 12092 28858 12116 28860
rect 12172 28858 12196 28860
rect 12252 28858 12258 28860
rect 12012 28806 12014 28858
rect 12194 28806 12196 28858
rect 11950 28804 11956 28806
rect 12012 28804 12036 28806
rect 12092 28804 12116 28806
rect 12172 28804 12196 28806
rect 12252 28804 12258 28806
rect 11950 28795 12258 28804
rect 11950 27772 12258 27781
rect 11950 27770 11956 27772
rect 12012 27770 12036 27772
rect 12092 27770 12116 27772
rect 12172 27770 12196 27772
rect 12252 27770 12258 27772
rect 12012 27718 12014 27770
rect 12194 27718 12196 27770
rect 11950 27716 11956 27718
rect 12012 27716 12036 27718
rect 12092 27716 12116 27718
rect 12172 27716 12196 27718
rect 12252 27716 12258 27718
rect 11950 27707 12258 27716
rect 11796 26920 11848 26926
rect 11796 26862 11848 26868
rect 11808 15706 11836 26862
rect 11950 26684 12258 26693
rect 11950 26682 11956 26684
rect 12012 26682 12036 26684
rect 12092 26682 12116 26684
rect 12172 26682 12196 26684
rect 12252 26682 12258 26684
rect 12012 26630 12014 26682
rect 12194 26630 12196 26682
rect 11950 26628 11956 26630
rect 12012 26628 12036 26630
rect 12092 26628 12116 26630
rect 12172 26628 12196 26630
rect 12252 26628 12258 26630
rect 11950 26619 12258 26628
rect 11950 25596 12258 25605
rect 11950 25594 11956 25596
rect 12012 25594 12036 25596
rect 12092 25594 12116 25596
rect 12172 25594 12196 25596
rect 12252 25594 12258 25596
rect 12012 25542 12014 25594
rect 12194 25542 12196 25594
rect 11950 25540 11956 25542
rect 12012 25540 12036 25542
rect 12092 25540 12116 25542
rect 12172 25540 12196 25542
rect 12252 25540 12258 25542
rect 11950 25531 12258 25540
rect 11950 24508 12258 24517
rect 11950 24506 11956 24508
rect 12012 24506 12036 24508
rect 12092 24506 12116 24508
rect 12172 24506 12196 24508
rect 12252 24506 12258 24508
rect 12012 24454 12014 24506
rect 12194 24454 12196 24506
rect 11950 24452 11956 24454
rect 12012 24452 12036 24454
rect 12092 24452 12116 24454
rect 12172 24452 12196 24454
rect 12252 24452 12258 24454
rect 11950 24443 12258 24452
rect 11950 23420 12258 23429
rect 11950 23418 11956 23420
rect 12012 23418 12036 23420
rect 12092 23418 12116 23420
rect 12172 23418 12196 23420
rect 12252 23418 12258 23420
rect 12012 23366 12014 23418
rect 12194 23366 12196 23418
rect 11950 23364 11956 23366
rect 12012 23364 12036 23366
rect 12092 23364 12116 23366
rect 12172 23364 12196 23366
rect 12252 23364 12258 23366
rect 11950 23355 12258 23364
rect 11950 22332 12258 22341
rect 11950 22330 11956 22332
rect 12012 22330 12036 22332
rect 12092 22330 12116 22332
rect 12172 22330 12196 22332
rect 12252 22330 12258 22332
rect 12012 22278 12014 22330
rect 12194 22278 12196 22330
rect 11950 22276 11956 22278
rect 12012 22276 12036 22278
rect 12092 22276 12116 22278
rect 12172 22276 12196 22278
rect 12252 22276 12258 22278
rect 11950 22267 12258 22276
rect 12360 21894 12388 39238
rect 12452 37398 12480 41386
rect 12610 41372 12918 41381
rect 12610 41370 12616 41372
rect 12672 41370 12696 41372
rect 12752 41370 12776 41372
rect 12832 41370 12856 41372
rect 12912 41370 12918 41372
rect 12672 41318 12674 41370
rect 12854 41318 12856 41370
rect 12610 41316 12616 41318
rect 12672 41316 12696 41318
rect 12752 41316 12776 41318
rect 12832 41316 12856 41318
rect 12912 41316 12918 41318
rect 12610 41307 12918 41316
rect 12610 40284 12918 40293
rect 12610 40282 12616 40284
rect 12672 40282 12696 40284
rect 12752 40282 12776 40284
rect 12832 40282 12856 40284
rect 12912 40282 12918 40284
rect 12672 40230 12674 40282
rect 12854 40230 12856 40282
rect 12610 40228 12616 40230
rect 12672 40228 12696 40230
rect 12752 40228 12776 40230
rect 12832 40228 12856 40230
rect 12912 40228 12918 40230
rect 12610 40219 12918 40228
rect 12532 39500 12584 39506
rect 12532 39442 12584 39448
rect 12440 37392 12492 37398
rect 12440 37334 12492 37340
rect 12438 35592 12494 35601
rect 12438 35527 12494 35536
rect 12452 35494 12480 35527
rect 12440 35488 12492 35494
rect 12440 35430 12492 35436
rect 12544 35086 12572 39442
rect 12610 39196 12918 39205
rect 12610 39194 12616 39196
rect 12672 39194 12696 39196
rect 12752 39194 12776 39196
rect 12832 39194 12856 39196
rect 12912 39194 12918 39196
rect 12672 39142 12674 39194
rect 12854 39142 12856 39194
rect 12610 39140 12616 39142
rect 12672 39140 12696 39142
rect 12752 39140 12776 39142
rect 12832 39140 12856 39142
rect 12912 39140 12918 39142
rect 12610 39131 12918 39140
rect 12610 38108 12918 38117
rect 12610 38106 12616 38108
rect 12672 38106 12696 38108
rect 12752 38106 12776 38108
rect 12832 38106 12856 38108
rect 12912 38106 12918 38108
rect 12672 38054 12674 38106
rect 12854 38054 12856 38106
rect 12610 38052 12616 38054
rect 12672 38052 12696 38054
rect 12752 38052 12776 38054
rect 12832 38052 12856 38054
rect 12912 38052 12918 38054
rect 12610 38043 12918 38052
rect 12624 37460 12676 37466
rect 12624 37402 12676 37408
rect 12636 37194 12664 37402
rect 12624 37188 12676 37194
rect 12624 37130 12676 37136
rect 12610 37020 12918 37029
rect 12610 37018 12616 37020
rect 12672 37018 12696 37020
rect 12752 37018 12776 37020
rect 12832 37018 12856 37020
rect 12912 37018 12918 37020
rect 12672 36966 12674 37018
rect 12854 36966 12856 37018
rect 12610 36964 12616 36966
rect 12672 36964 12696 36966
rect 12752 36964 12776 36966
rect 12832 36964 12856 36966
rect 12912 36964 12918 36966
rect 12610 36955 12918 36964
rect 13004 36922 13032 56238
rect 13096 47462 13124 59978
rect 13176 57044 13228 57050
rect 13176 56986 13228 56992
rect 13188 50930 13216 56986
rect 13268 52896 13320 52902
rect 13268 52838 13320 52844
rect 13176 50924 13228 50930
rect 13176 50866 13228 50872
rect 13084 47456 13136 47462
rect 13084 47398 13136 47404
rect 13188 45554 13216 50866
rect 13096 45526 13216 45554
rect 13096 37262 13124 45526
rect 13176 42560 13228 42566
rect 13176 42502 13228 42508
rect 13188 42362 13216 42502
rect 13176 42356 13228 42362
rect 13176 42298 13228 42304
rect 13084 37256 13136 37262
rect 13084 37198 13136 37204
rect 13176 37120 13228 37126
rect 13176 37062 13228 37068
rect 12992 36916 13044 36922
rect 12992 36858 13044 36864
rect 12610 35932 12918 35941
rect 12610 35930 12616 35932
rect 12672 35930 12696 35932
rect 12752 35930 12776 35932
rect 12832 35930 12856 35932
rect 12912 35930 12918 35932
rect 12672 35878 12674 35930
rect 12854 35878 12856 35930
rect 12610 35876 12616 35878
rect 12672 35876 12696 35878
rect 12752 35876 12776 35878
rect 12832 35876 12856 35878
rect 12912 35876 12918 35878
rect 12610 35867 12918 35876
rect 12992 35556 13044 35562
rect 12992 35498 13044 35504
rect 13004 35442 13032 35498
rect 13004 35414 13124 35442
rect 12532 35080 12584 35086
rect 12532 35022 12584 35028
rect 12992 35080 13044 35086
rect 12992 35022 13044 35028
rect 12440 35012 12492 35018
rect 12440 34954 12492 34960
rect 12452 34542 12480 34954
rect 12610 34844 12918 34853
rect 12610 34842 12616 34844
rect 12672 34842 12696 34844
rect 12752 34842 12776 34844
rect 12832 34842 12856 34844
rect 12912 34842 12918 34844
rect 12672 34790 12674 34842
rect 12854 34790 12856 34842
rect 12610 34788 12616 34790
rect 12672 34788 12696 34790
rect 12752 34788 12776 34790
rect 12832 34788 12856 34790
rect 12912 34788 12918 34790
rect 12610 34779 12918 34788
rect 12440 34536 12492 34542
rect 12440 34478 12492 34484
rect 12452 25294 12480 34478
rect 13004 34474 13032 35022
rect 13096 35018 13124 35414
rect 13084 35012 13136 35018
rect 13084 34954 13136 34960
rect 12992 34468 13044 34474
rect 12992 34410 13044 34416
rect 12610 33756 12918 33765
rect 12610 33754 12616 33756
rect 12672 33754 12696 33756
rect 12752 33754 12776 33756
rect 12832 33754 12856 33756
rect 12912 33754 12918 33756
rect 12672 33702 12674 33754
rect 12854 33702 12856 33754
rect 12610 33700 12616 33702
rect 12672 33700 12696 33702
rect 12752 33700 12776 33702
rect 12832 33700 12856 33702
rect 12912 33700 12918 33702
rect 12610 33691 12918 33700
rect 12610 32668 12918 32677
rect 12610 32666 12616 32668
rect 12672 32666 12696 32668
rect 12752 32666 12776 32668
rect 12832 32666 12856 32668
rect 12912 32666 12918 32668
rect 12672 32614 12674 32666
rect 12854 32614 12856 32666
rect 12610 32612 12616 32614
rect 12672 32612 12696 32614
rect 12752 32612 12776 32614
rect 12832 32612 12856 32614
rect 12912 32612 12918 32614
rect 12610 32603 12918 32612
rect 12610 31580 12918 31589
rect 12610 31578 12616 31580
rect 12672 31578 12696 31580
rect 12752 31578 12776 31580
rect 12832 31578 12856 31580
rect 12912 31578 12918 31580
rect 12672 31526 12674 31578
rect 12854 31526 12856 31578
rect 12610 31524 12616 31526
rect 12672 31524 12696 31526
rect 12752 31524 12776 31526
rect 12832 31524 12856 31526
rect 12912 31524 12918 31526
rect 12610 31515 12918 31524
rect 12610 30492 12918 30501
rect 12610 30490 12616 30492
rect 12672 30490 12696 30492
rect 12752 30490 12776 30492
rect 12832 30490 12856 30492
rect 12912 30490 12918 30492
rect 12672 30438 12674 30490
rect 12854 30438 12856 30490
rect 12610 30436 12616 30438
rect 12672 30436 12696 30438
rect 12752 30436 12776 30438
rect 12832 30436 12856 30438
rect 12912 30436 12918 30438
rect 12610 30427 12918 30436
rect 12610 29404 12918 29413
rect 12610 29402 12616 29404
rect 12672 29402 12696 29404
rect 12752 29402 12776 29404
rect 12832 29402 12856 29404
rect 12912 29402 12918 29404
rect 12672 29350 12674 29402
rect 12854 29350 12856 29402
rect 12610 29348 12616 29350
rect 12672 29348 12696 29350
rect 12752 29348 12776 29350
rect 12832 29348 12856 29350
rect 12912 29348 12918 29350
rect 12610 29339 12918 29348
rect 12610 28316 12918 28325
rect 12610 28314 12616 28316
rect 12672 28314 12696 28316
rect 12752 28314 12776 28316
rect 12832 28314 12856 28316
rect 12912 28314 12918 28316
rect 12672 28262 12674 28314
rect 12854 28262 12856 28314
rect 12610 28260 12616 28262
rect 12672 28260 12696 28262
rect 12752 28260 12776 28262
rect 12832 28260 12856 28262
rect 12912 28260 12918 28262
rect 12610 28251 12918 28260
rect 12610 27228 12918 27237
rect 12610 27226 12616 27228
rect 12672 27226 12696 27228
rect 12752 27226 12776 27228
rect 12832 27226 12856 27228
rect 12912 27226 12918 27228
rect 12672 27174 12674 27226
rect 12854 27174 12856 27226
rect 12610 27172 12616 27174
rect 12672 27172 12696 27174
rect 12752 27172 12776 27174
rect 12832 27172 12856 27174
rect 12912 27172 12918 27174
rect 12610 27163 12918 27172
rect 12610 26140 12918 26149
rect 12610 26138 12616 26140
rect 12672 26138 12696 26140
rect 12752 26138 12776 26140
rect 12832 26138 12856 26140
rect 12912 26138 12918 26140
rect 12672 26086 12674 26138
rect 12854 26086 12856 26138
rect 12610 26084 12616 26086
rect 12672 26084 12696 26086
rect 12752 26084 12776 26086
rect 12832 26084 12856 26086
rect 12912 26084 12918 26086
rect 12610 26075 12918 26084
rect 12532 25356 12584 25362
rect 12532 25298 12584 25304
rect 12440 25288 12492 25294
rect 12440 25230 12492 25236
rect 12544 23730 12572 25298
rect 12992 25288 13044 25294
rect 12992 25230 13044 25236
rect 12610 25052 12918 25061
rect 12610 25050 12616 25052
rect 12672 25050 12696 25052
rect 12752 25050 12776 25052
rect 12832 25050 12856 25052
rect 12912 25050 12918 25052
rect 12672 24998 12674 25050
rect 12854 24998 12856 25050
rect 12610 24996 12616 24998
rect 12672 24996 12696 24998
rect 12752 24996 12776 24998
rect 12832 24996 12856 24998
rect 12912 24996 12918 24998
rect 12610 24987 12918 24996
rect 12610 23964 12918 23973
rect 12610 23962 12616 23964
rect 12672 23962 12696 23964
rect 12752 23962 12776 23964
rect 12832 23962 12856 23964
rect 12912 23962 12918 23964
rect 12672 23910 12674 23962
rect 12854 23910 12856 23962
rect 12610 23908 12616 23910
rect 12672 23908 12696 23910
rect 12752 23908 12776 23910
rect 12832 23908 12856 23910
rect 12912 23908 12918 23910
rect 12610 23899 12918 23908
rect 12532 23724 12584 23730
rect 12532 23666 12584 23672
rect 12348 21888 12400 21894
rect 12348 21830 12400 21836
rect 12348 21344 12400 21350
rect 12348 21286 12400 21292
rect 11950 21244 12258 21253
rect 11950 21242 11956 21244
rect 12012 21242 12036 21244
rect 12092 21242 12116 21244
rect 12172 21242 12196 21244
rect 12252 21242 12258 21244
rect 12012 21190 12014 21242
rect 12194 21190 12196 21242
rect 11950 21188 11956 21190
rect 12012 21188 12036 21190
rect 12092 21188 12116 21190
rect 12172 21188 12196 21190
rect 12252 21188 12258 21190
rect 11950 21179 12258 21188
rect 12360 20942 12388 21286
rect 12348 20936 12400 20942
rect 12348 20878 12400 20884
rect 11980 20596 12032 20602
rect 11980 20538 12032 20544
rect 11992 20262 12020 20538
rect 11980 20256 12032 20262
rect 11980 20198 12032 20204
rect 11950 20156 12258 20165
rect 11950 20154 11956 20156
rect 12012 20154 12036 20156
rect 12092 20154 12116 20156
rect 12172 20154 12196 20156
rect 12252 20154 12258 20156
rect 12012 20102 12014 20154
rect 12194 20102 12196 20154
rect 11950 20100 11956 20102
rect 12012 20100 12036 20102
rect 12092 20100 12116 20102
rect 12172 20100 12196 20102
rect 12252 20100 12258 20102
rect 11950 20091 12258 20100
rect 12162 19952 12218 19961
rect 12162 19887 12218 19896
rect 12176 19378 12204 19887
rect 12164 19372 12216 19378
rect 12164 19314 12216 19320
rect 11950 19068 12258 19077
rect 11950 19066 11956 19068
rect 12012 19066 12036 19068
rect 12092 19066 12116 19068
rect 12172 19066 12196 19068
rect 12252 19066 12258 19068
rect 12012 19014 12014 19066
rect 12194 19014 12196 19066
rect 11950 19012 11956 19014
rect 12012 19012 12036 19014
rect 12092 19012 12116 19014
rect 12172 19012 12196 19014
rect 12252 19012 12258 19014
rect 11950 19003 12258 19012
rect 11950 17980 12258 17989
rect 11950 17978 11956 17980
rect 12012 17978 12036 17980
rect 12092 17978 12116 17980
rect 12172 17978 12196 17980
rect 12252 17978 12258 17980
rect 12012 17926 12014 17978
rect 12194 17926 12196 17978
rect 11950 17924 11956 17926
rect 12012 17924 12036 17926
rect 12092 17924 12116 17926
rect 12172 17924 12196 17926
rect 12252 17924 12258 17926
rect 11950 17915 12258 17924
rect 12544 17610 12572 23666
rect 12610 22876 12918 22885
rect 12610 22874 12616 22876
rect 12672 22874 12696 22876
rect 12752 22874 12776 22876
rect 12832 22874 12856 22876
rect 12912 22874 12918 22876
rect 12672 22822 12674 22874
rect 12854 22822 12856 22874
rect 12610 22820 12616 22822
rect 12672 22820 12696 22822
rect 12752 22820 12776 22822
rect 12832 22820 12856 22822
rect 12912 22820 12918 22822
rect 12610 22811 12918 22820
rect 12610 21788 12918 21797
rect 12610 21786 12616 21788
rect 12672 21786 12696 21788
rect 12752 21786 12776 21788
rect 12832 21786 12856 21788
rect 12912 21786 12918 21788
rect 12672 21734 12674 21786
rect 12854 21734 12856 21786
rect 12610 21732 12616 21734
rect 12672 21732 12696 21734
rect 12752 21732 12776 21734
rect 12832 21732 12856 21734
rect 12912 21732 12918 21734
rect 12610 21723 12918 21732
rect 13004 21146 13032 25230
rect 13096 25226 13124 34954
rect 13188 34610 13216 37062
rect 13280 36718 13308 52838
rect 13360 51468 13412 51474
rect 13360 51410 13412 51416
rect 13372 42838 13400 51410
rect 13464 44962 13492 74054
rect 13556 64874 13584 74506
rect 13728 74316 13780 74322
rect 13728 74258 13780 74264
rect 13740 69970 13768 74258
rect 13728 69964 13780 69970
rect 13728 69906 13780 69912
rect 13820 68808 13872 68814
rect 13820 68750 13872 68756
rect 13636 66156 13688 66162
rect 13636 66098 13688 66104
rect 13648 66042 13676 66098
rect 13832 66042 13860 68750
rect 14004 67244 14056 67250
rect 14004 67186 14056 67192
rect 13912 66224 13964 66230
rect 13912 66166 13964 66172
rect 13648 66014 13860 66042
rect 13556 64846 13676 64874
rect 13740 64870 13768 66014
rect 13924 65498 13952 66166
rect 13832 65470 13952 65498
rect 13544 61736 13596 61742
rect 13544 61678 13596 61684
rect 13556 45082 13584 61678
rect 13648 55214 13676 64846
rect 13728 64864 13780 64870
rect 13728 64806 13780 64812
rect 13740 64462 13768 64806
rect 13728 64456 13780 64462
rect 13728 64398 13780 64404
rect 13740 62098 13768 64398
rect 13832 62490 13860 65470
rect 14016 64874 14044 67186
rect 13924 64846 14044 64874
rect 13924 64326 13952 64846
rect 13912 64320 13964 64326
rect 13912 64262 13964 64268
rect 13924 63578 13952 64262
rect 13912 63572 13964 63578
rect 13912 63514 13964 63520
rect 13820 62484 13872 62490
rect 13820 62426 13872 62432
rect 13740 62070 13860 62098
rect 13832 61198 13860 62070
rect 13820 61192 13872 61198
rect 13820 61134 13872 61140
rect 13728 58880 13780 58886
rect 13726 58848 13728 58857
rect 13780 58848 13782 58857
rect 13726 58783 13782 58792
rect 14108 55214 14136 75210
rect 13648 55186 13768 55214
rect 13636 46368 13688 46374
rect 13636 46310 13688 46316
rect 13544 45076 13596 45082
rect 13544 45018 13596 45024
rect 13464 44934 13584 44962
rect 13452 44804 13504 44810
rect 13452 44746 13504 44752
rect 13360 42832 13412 42838
rect 13360 42774 13412 42780
rect 13464 39506 13492 44746
rect 13452 39500 13504 39506
rect 13452 39442 13504 39448
rect 13556 38282 13584 44934
rect 13544 38276 13596 38282
rect 13544 38218 13596 38224
rect 13544 37800 13596 37806
rect 13544 37742 13596 37748
rect 13556 37330 13584 37742
rect 13544 37324 13596 37330
rect 13544 37266 13596 37272
rect 13452 37188 13504 37194
rect 13452 37130 13504 37136
rect 13360 36916 13412 36922
rect 13360 36858 13412 36864
rect 13268 36712 13320 36718
rect 13268 36654 13320 36660
rect 13268 34944 13320 34950
rect 13268 34886 13320 34892
rect 13280 34610 13308 34886
rect 13176 34604 13228 34610
rect 13176 34546 13228 34552
rect 13268 34604 13320 34610
rect 13268 34546 13320 34552
rect 13084 25220 13136 25226
rect 13084 25162 13136 25168
rect 13084 24132 13136 24138
rect 13084 24074 13136 24080
rect 12992 21140 13044 21146
rect 12992 21082 13044 21088
rect 12610 20700 12918 20709
rect 12610 20698 12616 20700
rect 12672 20698 12696 20700
rect 12752 20698 12776 20700
rect 12832 20698 12856 20700
rect 12912 20698 12918 20700
rect 12672 20646 12674 20698
rect 12854 20646 12856 20698
rect 12610 20644 12616 20646
rect 12672 20644 12696 20646
rect 12752 20644 12776 20646
rect 12832 20644 12856 20646
rect 12912 20644 12918 20646
rect 12610 20635 12918 20644
rect 13096 20330 13124 24074
rect 13084 20324 13136 20330
rect 13084 20266 13136 20272
rect 12610 19612 12918 19621
rect 12610 19610 12616 19612
rect 12672 19610 12696 19612
rect 12752 19610 12776 19612
rect 12832 19610 12856 19612
rect 12912 19610 12918 19612
rect 12672 19558 12674 19610
rect 12854 19558 12856 19610
rect 12610 19556 12616 19558
rect 12672 19556 12696 19558
rect 12752 19556 12776 19558
rect 12832 19556 12856 19558
rect 12912 19556 12918 19558
rect 12610 19547 12918 19556
rect 12610 18524 12918 18533
rect 12610 18522 12616 18524
rect 12672 18522 12696 18524
rect 12752 18522 12776 18524
rect 12832 18522 12856 18524
rect 12912 18522 12918 18524
rect 12672 18470 12674 18522
rect 12854 18470 12856 18522
rect 12610 18468 12616 18470
rect 12672 18468 12696 18470
rect 12752 18468 12776 18470
rect 12832 18468 12856 18470
rect 12912 18468 12918 18470
rect 12610 18459 12918 18468
rect 13096 17746 13124 20266
rect 13084 17740 13136 17746
rect 13084 17682 13136 17688
rect 12532 17604 12584 17610
rect 12532 17546 12584 17552
rect 12610 17436 12918 17445
rect 12610 17434 12616 17436
rect 12672 17434 12696 17436
rect 12752 17434 12776 17436
rect 12832 17434 12856 17436
rect 12912 17434 12918 17436
rect 12672 17382 12674 17434
rect 12854 17382 12856 17434
rect 12610 17380 12616 17382
rect 12672 17380 12696 17382
rect 12752 17380 12776 17382
rect 12832 17380 12856 17382
rect 12912 17380 12918 17382
rect 12610 17371 12918 17380
rect 11950 16892 12258 16901
rect 11950 16890 11956 16892
rect 12012 16890 12036 16892
rect 12092 16890 12116 16892
rect 12172 16890 12196 16892
rect 12252 16890 12258 16892
rect 12012 16838 12014 16890
rect 12194 16838 12196 16890
rect 11950 16836 11956 16838
rect 12012 16836 12036 16838
rect 12092 16836 12116 16838
rect 12172 16836 12196 16838
rect 12252 16836 12258 16838
rect 11950 16827 12258 16836
rect 12610 16348 12918 16357
rect 12610 16346 12616 16348
rect 12672 16346 12696 16348
rect 12752 16346 12776 16348
rect 12832 16346 12856 16348
rect 12912 16346 12918 16348
rect 12672 16294 12674 16346
rect 12854 16294 12856 16346
rect 12610 16292 12616 16294
rect 12672 16292 12696 16294
rect 12752 16292 12776 16294
rect 12832 16292 12856 16294
rect 12912 16292 12918 16294
rect 12610 16283 12918 16292
rect 11950 15804 12258 15813
rect 11950 15802 11956 15804
rect 12012 15802 12036 15804
rect 12092 15802 12116 15804
rect 12172 15802 12196 15804
rect 12252 15802 12258 15804
rect 12012 15750 12014 15802
rect 12194 15750 12196 15802
rect 11950 15748 11956 15750
rect 12012 15748 12036 15750
rect 12092 15748 12116 15750
rect 12172 15748 12196 15750
rect 12252 15748 12258 15750
rect 11950 15739 12258 15748
rect 11796 15700 11848 15706
rect 11796 15642 11848 15648
rect 12990 15600 13046 15609
rect 12990 15535 12992 15544
rect 13044 15535 13046 15544
rect 13084 15564 13136 15570
rect 12992 15506 13044 15512
rect 13084 15506 13136 15512
rect 12610 15260 12918 15269
rect 12610 15258 12616 15260
rect 12672 15258 12696 15260
rect 12752 15258 12776 15260
rect 12832 15258 12856 15260
rect 12912 15258 12918 15260
rect 12672 15206 12674 15258
rect 12854 15206 12856 15258
rect 12610 15204 12616 15206
rect 12672 15204 12696 15206
rect 12752 15204 12776 15206
rect 12832 15204 12856 15206
rect 12912 15204 12918 15206
rect 12610 15195 12918 15204
rect 11950 14716 12258 14725
rect 11950 14714 11956 14716
rect 12012 14714 12036 14716
rect 12092 14714 12116 14716
rect 12172 14714 12196 14716
rect 12252 14714 12258 14716
rect 12012 14662 12014 14714
rect 12194 14662 12196 14714
rect 11950 14660 11956 14662
rect 12012 14660 12036 14662
rect 12092 14660 12116 14662
rect 12172 14660 12196 14662
rect 12252 14660 12258 14662
rect 11950 14651 12258 14660
rect 12610 14172 12918 14181
rect 12610 14170 12616 14172
rect 12672 14170 12696 14172
rect 12752 14170 12776 14172
rect 12832 14170 12856 14172
rect 12912 14170 12918 14172
rect 12672 14118 12674 14170
rect 12854 14118 12856 14170
rect 12610 14116 12616 14118
rect 12672 14116 12696 14118
rect 12752 14116 12776 14118
rect 12832 14116 12856 14118
rect 12912 14116 12918 14118
rect 12610 14107 12918 14116
rect 11950 13628 12258 13637
rect 11950 13626 11956 13628
rect 12012 13626 12036 13628
rect 12092 13626 12116 13628
rect 12172 13626 12196 13628
rect 12252 13626 12258 13628
rect 12012 13574 12014 13626
rect 12194 13574 12196 13626
rect 11950 13572 11956 13574
rect 12012 13572 12036 13574
rect 12092 13572 12116 13574
rect 12172 13572 12196 13574
rect 12252 13572 12258 13574
rect 11950 13563 12258 13572
rect 12610 13084 12918 13093
rect 12610 13082 12616 13084
rect 12672 13082 12696 13084
rect 12752 13082 12776 13084
rect 12832 13082 12856 13084
rect 12912 13082 12918 13084
rect 12672 13030 12674 13082
rect 12854 13030 12856 13082
rect 12610 13028 12616 13030
rect 12672 13028 12696 13030
rect 12752 13028 12776 13030
rect 12832 13028 12856 13030
rect 12912 13028 12918 13030
rect 12610 13019 12918 13028
rect 11704 12980 11756 12986
rect 11704 12922 11756 12928
rect 11950 12540 12258 12549
rect 11950 12538 11956 12540
rect 12012 12538 12036 12540
rect 12092 12538 12116 12540
rect 12172 12538 12196 12540
rect 12252 12538 12258 12540
rect 12012 12486 12014 12538
rect 12194 12486 12196 12538
rect 11950 12484 11956 12486
rect 12012 12484 12036 12486
rect 12092 12484 12116 12486
rect 12172 12484 12196 12486
rect 12252 12484 12258 12486
rect 11950 12475 12258 12484
rect 12164 12368 12216 12374
rect 12162 12336 12164 12345
rect 12216 12336 12218 12345
rect 12162 12271 12218 12280
rect 12610 11996 12918 12005
rect 12610 11994 12616 11996
rect 12672 11994 12696 11996
rect 12752 11994 12776 11996
rect 12832 11994 12856 11996
rect 12912 11994 12918 11996
rect 12672 11942 12674 11994
rect 12854 11942 12856 11994
rect 12610 11940 12616 11942
rect 12672 11940 12696 11942
rect 12752 11940 12776 11942
rect 12832 11940 12856 11942
rect 12912 11940 12918 11942
rect 12610 11931 12918 11940
rect 11950 11452 12258 11461
rect 11950 11450 11956 11452
rect 12012 11450 12036 11452
rect 12092 11450 12116 11452
rect 12172 11450 12196 11452
rect 12252 11450 12258 11452
rect 12012 11398 12014 11450
rect 12194 11398 12196 11450
rect 11950 11396 11956 11398
rect 12012 11396 12036 11398
rect 12092 11396 12116 11398
rect 12172 11396 12196 11398
rect 12252 11396 12258 11398
rect 11950 11387 12258 11396
rect 12610 10908 12918 10917
rect 12610 10906 12616 10908
rect 12672 10906 12696 10908
rect 12752 10906 12776 10908
rect 12832 10906 12856 10908
rect 12912 10906 12918 10908
rect 12672 10854 12674 10906
rect 12854 10854 12856 10906
rect 12610 10852 12616 10854
rect 12672 10852 12696 10854
rect 12752 10852 12776 10854
rect 12832 10852 12856 10854
rect 12912 10852 12918 10854
rect 12610 10843 12918 10852
rect 11950 10364 12258 10373
rect 11950 10362 11956 10364
rect 12012 10362 12036 10364
rect 12092 10362 12116 10364
rect 12172 10362 12196 10364
rect 12252 10362 12258 10364
rect 12012 10310 12014 10362
rect 12194 10310 12196 10362
rect 11950 10308 11956 10310
rect 12012 10308 12036 10310
rect 12092 10308 12116 10310
rect 12172 10308 12196 10310
rect 12252 10308 12258 10310
rect 11950 10299 12258 10308
rect 12610 9820 12918 9829
rect 12610 9818 12616 9820
rect 12672 9818 12696 9820
rect 12752 9818 12776 9820
rect 12832 9818 12856 9820
rect 12912 9818 12918 9820
rect 12672 9766 12674 9818
rect 12854 9766 12856 9818
rect 12610 9764 12616 9766
rect 12672 9764 12696 9766
rect 12752 9764 12776 9766
rect 12832 9764 12856 9766
rect 12912 9764 12918 9766
rect 12610 9755 12918 9764
rect 13096 9654 13124 15506
rect 13188 14618 13216 34546
rect 13268 34468 13320 34474
rect 13268 34410 13320 34416
rect 13280 31754 13308 34410
rect 13372 32570 13400 36858
rect 13360 32564 13412 32570
rect 13360 32506 13412 32512
rect 13280 31726 13400 31754
rect 13268 30660 13320 30666
rect 13268 30602 13320 30608
rect 13280 30326 13308 30602
rect 13268 30320 13320 30326
rect 13268 30262 13320 30268
rect 13268 26988 13320 26994
rect 13268 26930 13320 26936
rect 13280 26314 13308 26930
rect 13268 26308 13320 26314
rect 13268 26250 13320 26256
rect 13372 25362 13400 31726
rect 13360 25356 13412 25362
rect 13360 25298 13412 25304
rect 13372 25242 13400 25298
rect 13280 25214 13400 25242
rect 13280 21078 13308 25214
rect 13360 22772 13412 22778
rect 13360 22714 13412 22720
rect 13268 21072 13320 21078
rect 13268 21014 13320 21020
rect 13268 20256 13320 20262
rect 13268 20198 13320 20204
rect 13176 14612 13228 14618
rect 13176 14554 13228 14560
rect 13084 9648 13136 9654
rect 13084 9590 13136 9596
rect 11950 9276 12258 9285
rect 11950 9274 11956 9276
rect 12012 9274 12036 9276
rect 12092 9274 12116 9276
rect 12172 9274 12196 9276
rect 12252 9274 12258 9276
rect 12012 9222 12014 9274
rect 12194 9222 12196 9274
rect 11950 9220 11956 9222
rect 12012 9220 12036 9222
rect 12092 9220 12116 9222
rect 12172 9220 12196 9222
rect 12252 9220 12258 9222
rect 11950 9211 12258 9220
rect 12610 8732 12918 8741
rect 12610 8730 12616 8732
rect 12672 8730 12696 8732
rect 12752 8730 12776 8732
rect 12832 8730 12856 8732
rect 12912 8730 12918 8732
rect 12672 8678 12674 8730
rect 12854 8678 12856 8730
rect 12610 8676 12616 8678
rect 12672 8676 12696 8678
rect 12752 8676 12776 8678
rect 12832 8676 12856 8678
rect 12912 8676 12918 8678
rect 12610 8667 12918 8676
rect 11612 8356 11664 8362
rect 11612 8298 11664 8304
rect 13280 8294 13308 20198
rect 13372 17678 13400 22714
rect 13360 17672 13412 17678
rect 13360 17614 13412 17620
rect 13464 16590 13492 37130
rect 13556 35154 13584 37266
rect 13544 35148 13596 35154
rect 13544 35090 13596 35096
rect 13544 34944 13596 34950
rect 13544 34886 13596 34892
rect 13556 24857 13584 34886
rect 13648 30410 13676 46310
rect 13740 44878 13768 55186
rect 14016 55186 14136 55214
rect 14016 49366 14044 55186
rect 14096 51400 14148 51406
rect 14096 51342 14148 51348
rect 14004 49360 14056 49366
rect 14004 49302 14056 49308
rect 14108 48890 14136 51342
rect 14096 48884 14148 48890
rect 14096 48826 14148 48832
rect 13820 45076 13872 45082
rect 13820 45018 13872 45024
rect 13728 44872 13780 44878
rect 13728 44814 13780 44820
rect 13728 43444 13780 43450
rect 13728 43386 13780 43392
rect 13740 42634 13768 43386
rect 13832 42770 13860 45018
rect 14004 44804 14056 44810
rect 14004 44746 14056 44752
rect 13912 42832 13964 42838
rect 13912 42774 13964 42780
rect 13820 42764 13872 42770
rect 13820 42706 13872 42712
rect 13728 42628 13780 42634
rect 13728 42570 13780 42576
rect 13740 35290 13768 42570
rect 13832 42158 13860 42706
rect 13820 42152 13872 42158
rect 13820 42094 13872 42100
rect 13820 35488 13872 35494
rect 13820 35430 13872 35436
rect 13728 35284 13780 35290
rect 13728 35226 13780 35232
rect 13728 35148 13780 35154
rect 13728 35090 13780 35096
rect 13740 30666 13768 35090
rect 13832 34678 13860 35430
rect 13820 34672 13872 34678
rect 13820 34614 13872 34620
rect 13832 32978 13860 34614
rect 13820 32972 13872 32978
rect 13820 32914 13872 32920
rect 13832 32502 13860 32914
rect 13820 32496 13872 32502
rect 13820 32438 13872 32444
rect 13728 30660 13780 30666
rect 13728 30602 13780 30608
rect 13648 30382 13768 30410
rect 13636 30320 13688 30326
rect 13636 30262 13688 30268
rect 13542 24848 13598 24857
rect 13542 24783 13598 24792
rect 13648 22094 13676 30262
rect 13740 26042 13768 30382
rect 13832 30258 13860 32438
rect 13820 30252 13872 30258
rect 13820 30194 13872 30200
rect 13832 27062 13860 30194
rect 13924 27606 13952 42774
rect 14016 38758 14044 44746
rect 14200 39642 14228 75890
rect 14464 75880 14516 75886
rect 14464 75822 14516 75828
rect 14476 74534 14504 75822
rect 14936 74866 14964 76366
rect 16868 76362 16896 77318
rect 17610 77276 17918 77285
rect 17610 77274 17616 77276
rect 17672 77274 17696 77276
rect 17752 77274 17776 77276
rect 17832 77274 17856 77276
rect 17912 77274 17918 77276
rect 17672 77222 17674 77274
rect 17854 77222 17856 77274
rect 17610 77220 17616 77222
rect 17672 77220 17696 77222
rect 17752 77220 17776 77222
rect 17832 77220 17856 77222
rect 17912 77220 17918 77222
rect 17610 77211 17918 77220
rect 18248 77081 18276 77318
rect 18234 77072 18290 77081
rect 18234 77007 18290 77016
rect 17500 76968 17552 76974
rect 17500 76910 17552 76916
rect 16950 76732 17258 76741
rect 16950 76730 16956 76732
rect 17012 76730 17036 76732
rect 17092 76730 17116 76732
rect 17172 76730 17196 76732
rect 17252 76730 17258 76732
rect 17012 76678 17014 76730
rect 17194 76678 17196 76730
rect 16950 76676 16956 76678
rect 17012 76676 17036 76678
rect 17092 76676 17116 76678
rect 17172 76676 17196 76678
rect 17252 76676 17258 76678
rect 16950 76667 17258 76676
rect 16856 76356 16908 76362
rect 16856 76298 16908 76304
rect 16304 76288 16356 76294
rect 16304 76230 16356 76236
rect 15200 75472 15252 75478
rect 15200 75414 15252 75420
rect 14924 74860 14976 74866
rect 14924 74802 14976 74808
rect 15108 74860 15160 74866
rect 15108 74802 15160 74808
rect 14384 74506 14504 74534
rect 14280 74248 14332 74254
rect 14280 74190 14332 74196
rect 14292 70990 14320 74190
rect 14280 70984 14332 70990
rect 14280 70926 14332 70932
rect 14292 68814 14320 70926
rect 14280 68808 14332 68814
rect 14280 68750 14332 68756
rect 14384 68490 14412 74506
rect 14936 74254 14964 74802
rect 14924 74248 14976 74254
rect 14924 74190 14976 74196
rect 15120 69986 15148 74802
rect 15212 71194 15240 75414
rect 16028 75200 16080 75206
rect 16028 75142 16080 75148
rect 15292 74996 15344 75002
rect 15292 74938 15344 74944
rect 15200 71188 15252 71194
rect 15200 71130 15252 71136
rect 14936 69958 15148 69986
rect 14556 68740 14608 68746
rect 14556 68682 14608 68688
rect 14292 68462 14412 68490
rect 14292 65958 14320 68462
rect 14280 65952 14332 65958
rect 14280 65894 14332 65900
rect 14292 61742 14320 65894
rect 14372 65204 14424 65210
rect 14372 65146 14424 65152
rect 14280 61736 14332 61742
rect 14280 61678 14332 61684
rect 14280 61192 14332 61198
rect 14280 61134 14332 61140
rect 14292 60110 14320 61134
rect 14280 60104 14332 60110
rect 14280 60046 14332 60052
rect 14292 53174 14320 60046
rect 14280 53168 14332 53174
rect 14280 53110 14332 53116
rect 14292 52562 14320 53110
rect 14280 52556 14332 52562
rect 14280 52498 14332 52504
rect 14280 51400 14332 51406
rect 14280 51342 14332 51348
rect 14188 39636 14240 39642
rect 14188 39578 14240 39584
rect 14004 38752 14056 38758
rect 14004 38694 14056 38700
rect 14004 36644 14056 36650
rect 14004 36586 14056 36592
rect 14016 33522 14044 36586
rect 14094 35728 14150 35737
rect 14094 35663 14150 35672
rect 14108 35562 14136 35663
rect 14096 35556 14148 35562
rect 14096 35498 14148 35504
rect 14004 33516 14056 33522
rect 14004 33458 14056 33464
rect 14186 29880 14242 29889
rect 14186 29815 14188 29824
rect 14240 29815 14242 29824
rect 14188 29786 14240 29792
rect 13912 27600 13964 27606
rect 13912 27542 13964 27548
rect 13820 27056 13872 27062
rect 13820 26998 13872 27004
rect 13728 26036 13780 26042
rect 13728 25978 13780 25984
rect 13820 24948 13872 24954
rect 13820 24890 13872 24896
rect 13728 24132 13780 24138
rect 13728 24074 13780 24080
rect 13740 23798 13768 24074
rect 13728 23792 13780 23798
rect 13728 23734 13780 23740
rect 13556 22066 13676 22094
rect 13556 20398 13584 22066
rect 13728 21004 13780 21010
rect 13728 20946 13780 20952
rect 13544 20392 13596 20398
rect 13596 20340 13676 20346
rect 13544 20334 13676 20340
rect 13556 20318 13676 20334
rect 13544 17604 13596 17610
rect 13544 17546 13596 17552
rect 13452 16584 13504 16590
rect 13452 16526 13504 16532
rect 12440 8288 12492 8294
rect 12440 8230 12492 8236
rect 13268 8288 13320 8294
rect 13268 8230 13320 8236
rect 11950 8188 12258 8197
rect 11950 8186 11956 8188
rect 12012 8186 12036 8188
rect 12092 8186 12116 8188
rect 12172 8186 12196 8188
rect 12252 8186 12258 8188
rect 12012 8134 12014 8186
rect 12194 8134 12196 8186
rect 11950 8132 11956 8134
rect 12012 8132 12036 8134
rect 12092 8132 12116 8134
rect 12172 8132 12196 8134
rect 12252 8132 12258 8134
rect 11518 8120 11574 8129
rect 11950 8123 12258 8132
rect 11518 8055 11520 8064
rect 11572 8055 11574 8064
rect 11520 8026 11572 8032
rect 12254 7984 12310 7993
rect 12452 7954 12480 8230
rect 12254 7919 12310 7928
rect 12440 7948 12492 7954
rect 12268 7886 12296 7919
rect 12440 7890 12492 7896
rect 12256 7880 12308 7886
rect 12256 7822 12308 7828
rect 12268 7546 12296 7822
rect 12610 7644 12918 7653
rect 12610 7642 12616 7644
rect 12672 7642 12696 7644
rect 12752 7642 12776 7644
rect 12832 7642 12856 7644
rect 12912 7642 12918 7644
rect 12672 7590 12674 7642
rect 12854 7590 12856 7642
rect 12610 7588 12616 7590
rect 12672 7588 12696 7590
rect 12752 7588 12776 7590
rect 12832 7588 12856 7590
rect 12912 7588 12918 7590
rect 12610 7579 12918 7588
rect 12256 7540 12308 7546
rect 12256 7482 12308 7488
rect 11950 7100 12258 7109
rect 11950 7098 11956 7100
rect 12012 7098 12036 7100
rect 12092 7098 12116 7100
rect 12172 7098 12196 7100
rect 12252 7098 12258 7100
rect 12012 7046 12014 7098
rect 12194 7046 12196 7098
rect 11950 7044 11956 7046
rect 12012 7044 12036 7046
rect 12092 7044 12116 7046
rect 12172 7044 12196 7046
rect 12252 7044 12258 7046
rect 11950 7035 12258 7044
rect 12714 6896 12770 6905
rect 12714 6831 12770 6840
rect 13358 6896 13414 6905
rect 13358 6831 13414 6840
rect 12728 6662 12756 6831
rect 12716 6656 12768 6662
rect 12716 6598 12768 6604
rect 12610 6556 12918 6565
rect 12610 6554 12616 6556
rect 12672 6554 12696 6556
rect 12752 6554 12776 6556
rect 12832 6554 12856 6556
rect 12912 6554 12918 6556
rect 12672 6502 12674 6554
rect 12854 6502 12856 6554
rect 12610 6500 12616 6502
rect 12672 6500 12696 6502
rect 12752 6500 12776 6502
rect 12832 6500 12856 6502
rect 12912 6500 12918 6502
rect 12610 6491 12918 6500
rect 11950 6012 12258 6021
rect 11950 6010 11956 6012
rect 12012 6010 12036 6012
rect 12092 6010 12116 6012
rect 12172 6010 12196 6012
rect 12252 6010 12258 6012
rect 12012 5958 12014 6010
rect 12194 5958 12196 6010
rect 11950 5956 11956 5958
rect 12012 5956 12036 5958
rect 12092 5956 12116 5958
rect 12172 5956 12196 5958
rect 12252 5956 12258 5958
rect 11950 5947 12258 5956
rect 11428 5568 11480 5574
rect 11428 5510 11480 5516
rect 12610 5468 12918 5477
rect 12610 5466 12616 5468
rect 12672 5466 12696 5468
rect 12752 5466 12776 5468
rect 12832 5466 12856 5468
rect 12912 5466 12918 5468
rect 12672 5414 12674 5466
rect 12854 5414 12856 5466
rect 12610 5412 12616 5414
rect 12672 5412 12696 5414
rect 12752 5412 12776 5414
rect 12832 5412 12856 5414
rect 12912 5412 12918 5414
rect 12610 5403 12918 5412
rect 13372 5302 13400 6831
rect 13556 6730 13584 17546
rect 13648 15570 13676 20318
rect 13740 20058 13768 20946
rect 13728 20052 13780 20058
rect 13728 19994 13780 20000
rect 13740 18290 13768 19994
rect 13728 18284 13780 18290
rect 13728 18226 13780 18232
rect 13832 17882 13860 24890
rect 14096 21888 14148 21894
rect 14096 21830 14148 21836
rect 13820 17876 13872 17882
rect 13820 17818 13872 17824
rect 13636 15564 13688 15570
rect 13636 15506 13688 15512
rect 14108 8566 14136 21830
rect 14200 20942 14228 29786
rect 14292 24682 14320 51342
rect 14384 44538 14412 65146
rect 14568 63510 14596 68682
rect 14936 68338 14964 69958
rect 15016 69896 15068 69902
rect 15016 69838 15068 69844
rect 15108 69896 15160 69902
rect 15108 69838 15160 69844
rect 15028 69057 15056 69838
rect 15014 69048 15070 69057
rect 15014 68983 15070 68992
rect 14924 68332 14976 68338
rect 14924 68274 14976 68280
rect 14832 65952 14884 65958
rect 14832 65894 14884 65900
rect 14556 63504 14608 63510
rect 14556 63446 14608 63452
rect 14462 63336 14518 63345
rect 14462 63271 14518 63280
rect 14476 63238 14504 63271
rect 14464 63232 14516 63238
rect 14464 63174 14516 63180
rect 14556 60036 14608 60042
rect 14556 59978 14608 59984
rect 14568 52154 14596 59978
rect 14556 52148 14608 52154
rect 14556 52090 14608 52096
rect 14556 50176 14608 50182
rect 14556 50118 14608 50124
rect 14568 44946 14596 50118
rect 14648 48748 14700 48754
rect 14648 48690 14700 48696
rect 14556 44940 14608 44946
rect 14556 44882 14608 44888
rect 14372 44532 14424 44538
rect 14372 44474 14424 44480
rect 14464 38752 14516 38758
rect 14464 38694 14516 38700
rect 14280 24676 14332 24682
rect 14280 24618 14332 24624
rect 14188 20936 14240 20942
rect 14188 20878 14240 20884
rect 14188 19508 14240 19514
rect 14188 19450 14240 19456
rect 14200 18358 14228 19450
rect 14188 18352 14240 18358
rect 14188 18294 14240 18300
rect 14372 10464 14424 10470
rect 14372 10406 14424 10412
rect 14096 8560 14148 8566
rect 14096 8502 14148 8508
rect 14384 8430 14412 10406
rect 14372 8424 14424 8430
rect 14372 8366 14424 8372
rect 14186 8256 14242 8265
rect 14186 8191 14242 8200
rect 14200 7478 14228 8191
rect 14188 7472 14240 7478
rect 14188 7414 14240 7420
rect 13818 7304 13874 7313
rect 13818 7239 13820 7248
rect 13872 7239 13874 7248
rect 13820 7210 13872 7216
rect 13544 6724 13596 6730
rect 13544 6666 13596 6672
rect 13360 5296 13412 5302
rect 13360 5238 13412 5244
rect 11060 5228 11112 5234
rect 11060 5170 11112 5176
rect 11704 5228 11756 5234
rect 11704 5170 11756 5176
rect 10968 3732 11020 3738
rect 10968 3674 11020 3680
rect 11716 3602 11744 5170
rect 11950 4924 12258 4933
rect 11950 4922 11956 4924
rect 12012 4922 12036 4924
rect 12092 4922 12116 4924
rect 12172 4922 12196 4924
rect 12252 4922 12258 4924
rect 12012 4870 12014 4922
rect 12194 4870 12196 4922
rect 11950 4868 11956 4870
rect 12012 4868 12036 4870
rect 12092 4868 12116 4870
rect 12172 4868 12196 4870
rect 12252 4868 12258 4870
rect 11950 4859 12258 4868
rect 14476 4622 14504 38694
rect 14660 25906 14688 48690
rect 14740 48680 14792 48686
rect 14740 48622 14792 48628
rect 14752 31482 14780 48622
rect 14844 43790 14872 65894
rect 15120 65210 15148 69838
rect 15108 65204 15160 65210
rect 15108 65146 15160 65152
rect 14924 63572 14976 63578
rect 14924 63514 14976 63520
rect 14832 43784 14884 43790
rect 14832 43726 14884 43732
rect 14832 37324 14884 37330
rect 14832 37266 14884 37272
rect 14740 31476 14792 31482
rect 14740 31418 14792 31424
rect 14648 25900 14700 25906
rect 14648 25842 14700 25848
rect 14660 25786 14688 25842
rect 14568 25758 14688 25786
rect 14568 20058 14596 25758
rect 14844 24818 14872 37266
rect 14832 24812 14884 24818
rect 14832 24754 14884 24760
rect 14740 24744 14792 24750
rect 14740 24686 14792 24692
rect 14752 24206 14780 24686
rect 14740 24200 14792 24206
rect 14740 24142 14792 24148
rect 14648 20936 14700 20942
rect 14648 20878 14700 20884
rect 14556 20052 14608 20058
rect 14556 19994 14608 20000
rect 14556 17808 14608 17814
rect 14556 17750 14608 17756
rect 14568 8566 14596 17750
rect 14660 8634 14688 20878
rect 14752 16522 14780 24142
rect 14832 20868 14884 20874
rect 14832 20810 14884 20816
rect 14740 16516 14792 16522
rect 14740 16458 14792 16464
rect 14844 11150 14872 20810
rect 14936 20534 14964 63514
rect 15200 59084 15252 59090
rect 15200 59026 15252 59032
rect 15016 48680 15068 48686
rect 15016 48622 15068 48628
rect 15028 39846 15056 48622
rect 15108 47116 15160 47122
rect 15108 47058 15160 47064
rect 15016 39840 15068 39846
rect 15016 39782 15068 39788
rect 15028 38826 15056 39782
rect 15016 38820 15068 38826
rect 15016 38762 15068 38768
rect 15016 37392 15068 37398
rect 15016 37334 15068 37340
rect 15028 34950 15056 37334
rect 15120 36582 15148 47058
rect 15212 42702 15240 59026
rect 15304 58954 15332 74938
rect 15844 74724 15896 74730
rect 15844 74666 15896 74672
rect 15568 74112 15620 74118
rect 15568 74054 15620 74060
rect 15476 69760 15528 69766
rect 15476 69702 15528 69708
rect 15384 63912 15436 63918
rect 15384 63854 15436 63860
rect 15396 60110 15424 63854
rect 15488 60178 15516 69702
rect 15580 65550 15608 74054
rect 15660 71596 15712 71602
rect 15660 71538 15712 71544
rect 15672 68678 15700 71538
rect 15752 70916 15804 70922
rect 15752 70858 15804 70864
rect 15660 68672 15712 68678
rect 15660 68614 15712 68620
rect 15568 65544 15620 65550
rect 15568 65486 15620 65492
rect 15568 63368 15620 63374
rect 15568 63310 15620 63316
rect 15476 60172 15528 60178
rect 15476 60114 15528 60120
rect 15384 60104 15436 60110
rect 15384 60046 15436 60052
rect 15396 59090 15424 60046
rect 15384 59084 15436 59090
rect 15384 59026 15436 59032
rect 15292 58948 15344 58954
rect 15292 58890 15344 58896
rect 15292 57384 15344 57390
rect 15292 57326 15344 57332
rect 15304 53242 15332 57326
rect 15292 53236 15344 53242
rect 15292 53178 15344 53184
rect 15396 48686 15424 59026
rect 15476 58948 15528 58954
rect 15476 58890 15528 58896
rect 15384 48680 15436 48686
rect 15384 48622 15436 48628
rect 15292 44736 15344 44742
rect 15292 44678 15344 44684
rect 15200 42696 15252 42702
rect 15200 42638 15252 42644
rect 15200 41540 15252 41546
rect 15200 41482 15252 41488
rect 15212 38350 15240 41482
rect 15200 38344 15252 38350
rect 15200 38286 15252 38292
rect 15200 37664 15252 37670
rect 15200 37606 15252 37612
rect 15108 36576 15160 36582
rect 15108 36518 15160 36524
rect 15016 34944 15068 34950
rect 15016 34886 15068 34892
rect 15028 34610 15056 34886
rect 15108 34740 15160 34746
rect 15108 34682 15160 34688
rect 15016 34604 15068 34610
rect 15016 34546 15068 34552
rect 15120 24750 15148 34682
rect 15108 24744 15160 24750
rect 15108 24686 15160 24692
rect 15212 22030 15240 37606
rect 15200 22024 15252 22030
rect 15200 21966 15252 21972
rect 15016 21072 15068 21078
rect 15016 21014 15068 21020
rect 14924 20528 14976 20534
rect 14924 20470 14976 20476
rect 14936 15162 14964 20470
rect 14924 15156 14976 15162
rect 14924 15098 14976 15104
rect 15028 15026 15056 21014
rect 15304 16574 15332 44678
rect 15384 37936 15436 37942
rect 15384 37878 15436 37884
rect 15396 34746 15424 37878
rect 15384 34740 15436 34746
rect 15384 34682 15436 34688
rect 15488 29510 15516 58890
rect 15580 57594 15608 63310
rect 15672 61878 15700 68614
rect 15660 61872 15712 61878
rect 15660 61814 15712 61820
rect 15568 57588 15620 57594
rect 15568 57530 15620 57536
rect 15568 52488 15620 52494
rect 15568 52430 15620 52436
rect 15580 33658 15608 52430
rect 15660 52352 15712 52358
rect 15660 52294 15712 52300
rect 15672 48550 15700 52294
rect 15660 48544 15712 48550
rect 15660 48486 15712 48492
rect 15764 37330 15792 70858
rect 15856 53106 15884 74666
rect 15936 73840 15988 73846
rect 15936 73782 15988 73788
rect 15948 53446 15976 73782
rect 16040 67182 16068 75142
rect 16316 73846 16344 76230
rect 16672 76084 16724 76090
rect 16672 76026 16724 76032
rect 16304 73840 16356 73846
rect 16304 73782 16356 73788
rect 16580 72616 16632 72622
rect 16580 72558 16632 72564
rect 16592 71942 16620 72558
rect 16684 72282 16712 76026
rect 16950 75644 17258 75653
rect 16950 75642 16956 75644
rect 17012 75642 17036 75644
rect 17092 75642 17116 75644
rect 17172 75642 17196 75644
rect 17252 75642 17258 75644
rect 17012 75590 17014 75642
rect 17194 75590 17196 75642
rect 16950 75588 16956 75590
rect 17012 75588 17036 75590
rect 17092 75588 17116 75590
rect 17172 75588 17196 75590
rect 17252 75588 17258 75590
rect 16950 75579 17258 75588
rect 16856 74860 16908 74866
rect 16856 74802 16908 74808
rect 16868 74534 16896 74802
rect 17512 74730 17540 76910
rect 17610 76188 17918 76197
rect 17610 76186 17616 76188
rect 17672 76186 17696 76188
rect 17752 76186 17776 76188
rect 17832 76186 17856 76188
rect 17912 76186 17918 76188
rect 17672 76134 17674 76186
rect 17854 76134 17856 76186
rect 17610 76132 17616 76134
rect 17672 76132 17696 76134
rect 17752 76132 17776 76134
rect 17832 76132 17856 76134
rect 17912 76132 17918 76134
rect 17610 76123 17918 76132
rect 18236 75200 18288 75206
rect 18234 75168 18236 75177
rect 18288 75168 18290 75177
rect 17610 75100 17918 75109
rect 18234 75103 18290 75112
rect 17610 75098 17616 75100
rect 17672 75098 17696 75100
rect 17752 75098 17776 75100
rect 17832 75098 17856 75100
rect 17912 75098 17918 75100
rect 17672 75046 17674 75098
rect 17854 75046 17856 75098
rect 17610 75044 17616 75046
rect 17672 75044 17696 75046
rect 17752 75044 17776 75046
rect 17832 75044 17856 75046
rect 17912 75044 17918 75046
rect 17610 75035 17918 75044
rect 17500 74724 17552 74730
rect 17500 74666 17552 74672
rect 16776 74506 16896 74534
rect 16950 74556 17258 74565
rect 16950 74554 16956 74556
rect 17012 74554 17036 74556
rect 17092 74554 17116 74556
rect 17172 74554 17196 74556
rect 17252 74554 17258 74556
rect 16672 72276 16724 72282
rect 16672 72218 16724 72224
rect 16580 71936 16632 71942
rect 16580 71878 16632 71884
rect 16672 70848 16724 70854
rect 16672 70790 16724 70796
rect 16684 70106 16712 70790
rect 16672 70100 16724 70106
rect 16672 70042 16724 70048
rect 16028 67176 16080 67182
rect 16028 67118 16080 67124
rect 16488 67176 16540 67182
rect 16488 67118 16540 67124
rect 16212 65544 16264 65550
rect 16212 65486 16264 65492
rect 16224 61402 16252 65486
rect 16500 64870 16528 67118
rect 16580 66224 16632 66230
rect 16580 66166 16632 66172
rect 16488 64864 16540 64870
rect 16488 64806 16540 64812
rect 16488 63368 16540 63374
rect 16488 63310 16540 63316
rect 16500 61946 16528 63310
rect 16488 61940 16540 61946
rect 16488 61882 16540 61888
rect 16212 61396 16264 61402
rect 16212 61338 16264 61344
rect 16212 61124 16264 61130
rect 16212 61066 16264 61072
rect 16120 59968 16172 59974
rect 16120 59910 16172 59916
rect 15936 53440 15988 53446
rect 15936 53382 15988 53388
rect 15844 53100 15896 53106
rect 15844 53042 15896 53048
rect 16028 48748 16080 48754
rect 16028 48690 16080 48696
rect 16040 48385 16068 48690
rect 16026 48376 16082 48385
rect 16026 48311 16082 48320
rect 15844 47048 15896 47054
rect 15844 46990 15896 46996
rect 15752 37324 15804 37330
rect 15752 37266 15804 37272
rect 15660 36576 15712 36582
rect 15660 36518 15712 36524
rect 15568 33652 15620 33658
rect 15568 33594 15620 33600
rect 15672 29850 15700 36518
rect 15856 35086 15884 46990
rect 16132 45554 16160 59910
rect 16040 45526 16160 45554
rect 15936 38004 15988 38010
rect 15936 37946 15988 37952
rect 15948 36786 15976 37946
rect 15936 36780 15988 36786
rect 15936 36722 15988 36728
rect 15844 35080 15896 35086
rect 15844 35022 15896 35028
rect 15752 33652 15804 33658
rect 15752 33594 15804 33600
rect 15660 29844 15712 29850
rect 15660 29786 15712 29792
rect 15476 29504 15528 29510
rect 15476 29446 15528 29452
rect 15764 22094 15792 33594
rect 16040 31754 16068 45526
rect 16120 33856 16172 33862
rect 16120 33798 16172 33804
rect 16132 32842 16160 33798
rect 16120 32836 16172 32842
rect 16120 32778 16172 32784
rect 16040 31726 16160 31754
rect 15936 30048 15988 30054
rect 15936 29990 15988 29996
rect 15948 29714 15976 29990
rect 15936 29708 15988 29714
rect 15936 29650 15988 29656
rect 16132 29510 16160 31726
rect 16028 29504 16080 29510
rect 16028 29446 16080 29452
rect 16120 29504 16172 29510
rect 16120 29446 16172 29452
rect 15844 25220 15896 25226
rect 15844 25162 15896 25168
rect 15672 22066 15792 22094
rect 15672 20806 15700 22066
rect 15660 20800 15712 20806
rect 15660 20742 15712 20748
rect 15304 16546 15424 16574
rect 15016 15020 15068 15026
rect 15016 14962 15068 14968
rect 15290 11248 15346 11257
rect 15200 11212 15252 11218
rect 15290 11183 15292 11192
rect 15200 11154 15252 11160
rect 15344 11183 15346 11192
rect 15292 11154 15344 11160
rect 14832 11144 14884 11150
rect 14832 11086 14884 11092
rect 15212 10674 15240 11154
rect 15200 10668 15252 10674
rect 15200 10610 15252 10616
rect 15396 9586 15424 16546
rect 15856 15094 15884 25162
rect 15936 20800 15988 20806
rect 15936 20742 15988 20748
rect 15844 15088 15896 15094
rect 15844 15030 15896 15036
rect 15476 14408 15528 14414
rect 15476 14350 15528 14356
rect 15488 13802 15516 14350
rect 15476 13796 15528 13802
rect 15476 13738 15528 13744
rect 15948 9994 15976 20742
rect 16040 11082 16068 29446
rect 16132 14074 16160 29446
rect 16224 22166 16252 61066
rect 16488 60240 16540 60246
rect 16488 60182 16540 60188
rect 16396 60172 16448 60178
rect 16396 60114 16448 60120
rect 16408 60081 16436 60114
rect 16394 60072 16450 60081
rect 16394 60007 16450 60016
rect 16302 49600 16358 49609
rect 16302 49535 16358 49544
rect 16316 37369 16344 49535
rect 16396 49156 16448 49162
rect 16396 49098 16448 49104
rect 16408 45082 16436 49098
rect 16500 47054 16528 60182
rect 16592 57526 16620 66166
rect 16684 58546 16712 70042
rect 16672 58540 16724 58546
rect 16672 58482 16724 58488
rect 16776 58426 16804 74506
rect 17012 74502 17014 74554
rect 17194 74502 17196 74554
rect 16950 74500 16956 74502
rect 17012 74500 17036 74502
rect 17092 74500 17116 74502
rect 17172 74500 17196 74502
rect 17252 74500 17258 74502
rect 16950 74491 17258 74500
rect 16856 74452 16908 74458
rect 16856 74394 16908 74400
rect 16868 72078 16896 74394
rect 17610 74012 17918 74021
rect 17610 74010 17616 74012
rect 17672 74010 17696 74012
rect 17752 74010 17776 74012
rect 17832 74010 17856 74012
rect 17912 74010 17918 74012
rect 17672 73958 17674 74010
rect 17854 73958 17856 74010
rect 17610 73956 17616 73958
rect 17672 73956 17696 73958
rect 17752 73956 17776 73958
rect 17832 73956 17856 73958
rect 17912 73956 17918 73958
rect 17610 73947 17918 73956
rect 17500 73704 17552 73710
rect 17500 73646 17552 73652
rect 16950 73468 17258 73477
rect 16950 73466 16956 73468
rect 17012 73466 17036 73468
rect 17092 73466 17116 73468
rect 17172 73466 17196 73468
rect 17252 73466 17258 73468
rect 17012 73414 17014 73466
rect 17194 73414 17196 73466
rect 16950 73412 16956 73414
rect 17012 73412 17036 73414
rect 17092 73412 17116 73414
rect 17172 73412 17196 73414
rect 17252 73412 17258 73414
rect 16950 73403 17258 73412
rect 16950 72380 17258 72389
rect 16950 72378 16956 72380
rect 17012 72378 17036 72380
rect 17092 72378 17116 72380
rect 17172 72378 17196 72380
rect 17252 72378 17258 72380
rect 17012 72326 17014 72378
rect 17194 72326 17196 72378
rect 16950 72324 16956 72326
rect 17012 72324 17036 72326
rect 17092 72324 17116 72326
rect 17172 72324 17196 72326
rect 17252 72324 17258 72326
rect 16950 72315 17258 72324
rect 16856 72072 16908 72078
rect 16856 72014 16908 72020
rect 16856 71936 16908 71942
rect 16856 71878 16908 71884
rect 16868 65634 16896 71878
rect 16950 71292 17258 71301
rect 16950 71290 16956 71292
rect 17012 71290 17036 71292
rect 17092 71290 17116 71292
rect 17172 71290 17196 71292
rect 17252 71290 17258 71292
rect 17012 71238 17014 71290
rect 17194 71238 17196 71290
rect 16950 71236 16956 71238
rect 17012 71236 17036 71238
rect 17092 71236 17116 71238
rect 17172 71236 17196 71238
rect 17252 71236 17258 71238
rect 16950 71227 17258 71236
rect 16950 70204 17258 70213
rect 16950 70202 16956 70204
rect 17012 70202 17036 70204
rect 17092 70202 17116 70204
rect 17172 70202 17196 70204
rect 17252 70202 17258 70204
rect 17012 70150 17014 70202
rect 17194 70150 17196 70202
rect 16950 70148 16956 70150
rect 17012 70148 17036 70150
rect 17092 70148 17116 70150
rect 17172 70148 17196 70150
rect 17252 70148 17258 70150
rect 16950 70139 17258 70148
rect 16950 69116 17258 69125
rect 16950 69114 16956 69116
rect 17012 69114 17036 69116
rect 17092 69114 17116 69116
rect 17172 69114 17196 69116
rect 17252 69114 17258 69116
rect 17012 69062 17014 69114
rect 17194 69062 17196 69114
rect 16950 69060 16956 69062
rect 17012 69060 17036 69062
rect 17092 69060 17116 69062
rect 17172 69060 17196 69062
rect 17252 69060 17258 69062
rect 16950 69051 17258 69060
rect 16950 68028 17258 68037
rect 16950 68026 16956 68028
rect 17012 68026 17036 68028
rect 17092 68026 17116 68028
rect 17172 68026 17196 68028
rect 17252 68026 17258 68028
rect 17012 67974 17014 68026
rect 17194 67974 17196 68026
rect 16950 67972 16956 67974
rect 17012 67972 17036 67974
rect 17092 67972 17116 67974
rect 17172 67972 17196 67974
rect 17252 67972 17258 67974
rect 16950 67963 17258 67972
rect 17408 67720 17460 67726
rect 17408 67662 17460 67668
rect 17316 67040 17368 67046
rect 17316 66982 17368 66988
rect 16950 66940 17258 66949
rect 16950 66938 16956 66940
rect 17012 66938 17036 66940
rect 17092 66938 17116 66940
rect 17172 66938 17196 66940
rect 17252 66938 17258 66940
rect 17012 66886 17014 66938
rect 17194 66886 17196 66938
rect 16950 66884 16956 66886
rect 17012 66884 17036 66886
rect 17092 66884 17116 66886
rect 17172 66884 17196 66886
rect 17252 66884 17258 66886
rect 16950 66875 17258 66884
rect 16950 65852 17258 65861
rect 16950 65850 16956 65852
rect 17012 65850 17036 65852
rect 17092 65850 17116 65852
rect 17172 65850 17196 65852
rect 17252 65850 17258 65852
rect 17012 65798 17014 65850
rect 17194 65798 17196 65850
rect 16950 65796 16956 65798
rect 17012 65796 17036 65798
rect 17092 65796 17116 65798
rect 17172 65796 17196 65798
rect 17252 65796 17258 65798
rect 16950 65787 17258 65796
rect 16868 65606 17080 65634
rect 17052 64938 17080 65606
rect 17328 65090 17356 66982
rect 17420 66162 17448 67662
rect 17512 66230 17540 73646
rect 18236 73568 18288 73574
rect 18236 73510 18288 73516
rect 18248 73273 18276 73510
rect 18234 73264 18290 73273
rect 18234 73199 18290 73208
rect 17610 72924 17918 72933
rect 17610 72922 17616 72924
rect 17672 72922 17696 72924
rect 17752 72922 17776 72924
rect 17832 72922 17856 72924
rect 17912 72922 17918 72924
rect 17672 72870 17674 72922
rect 17854 72870 17856 72922
rect 17610 72868 17616 72870
rect 17672 72868 17696 72870
rect 17752 72868 17776 72870
rect 17832 72868 17856 72870
rect 17912 72868 17918 72870
rect 17610 72859 17918 72868
rect 17610 71836 17918 71845
rect 17610 71834 17616 71836
rect 17672 71834 17696 71836
rect 17752 71834 17776 71836
rect 17832 71834 17856 71836
rect 17912 71834 17918 71836
rect 17672 71782 17674 71834
rect 17854 71782 17856 71834
rect 17610 71780 17616 71782
rect 17672 71780 17696 71782
rect 17752 71780 17776 71782
rect 17832 71780 17856 71782
rect 17912 71780 17918 71782
rect 17610 71771 17918 71780
rect 18236 71392 18288 71398
rect 18234 71360 18236 71369
rect 18288 71360 18290 71369
rect 18234 71295 18290 71304
rect 17610 70748 17918 70757
rect 17610 70746 17616 70748
rect 17672 70746 17696 70748
rect 17752 70746 17776 70748
rect 17832 70746 17856 70748
rect 17912 70746 17918 70748
rect 17672 70694 17674 70746
rect 17854 70694 17856 70746
rect 17610 70692 17616 70694
rect 17672 70692 17696 70694
rect 17752 70692 17776 70694
rect 17832 70692 17856 70694
rect 17912 70692 17918 70694
rect 17610 70683 17918 70692
rect 18236 69760 18288 69766
rect 18236 69702 18288 69708
rect 17610 69660 17918 69669
rect 17610 69658 17616 69660
rect 17672 69658 17696 69660
rect 17752 69658 17776 69660
rect 17832 69658 17856 69660
rect 17912 69658 17918 69660
rect 17672 69606 17674 69658
rect 17854 69606 17856 69658
rect 17610 69604 17616 69606
rect 17672 69604 17696 69606
rect 17752 69604 17776 69606
rect 17832 69604 17856 69606
rect 17912 69604 17918 69606
rect 17610 69595 17918 69604
rect 18248 69465 18276 69702
rect 18234 69456 18290 69465
rect 18234 69391 18290 69400
rect 17610 68572 17918 68581
rect 17610 68570 17616 68572
rect 17672 68570 17696 68572
rect 17752 68570 17776 68572
rect 17832 68570 17856 68572
rect 17912 68570 17918 68572
rect 17672 68518 17674 68570
rect 17854 68518 17856 68570
rect 17610 68516 17616 68518
rect 17672 68516 17696 68518
rect 17752 68516 17776 68518
rect 17832 68516 17856 68518
rect 17912 68516 17918 68518
rect 17610 68507 17918 68516
rect 18236 67856 18288 67862
rect 18236 67798 18288 67804
rect 18248 67561 18276 67798
rect 18234 67552 18290 67561
rect 17610 67484 17918 67493
rect 18234 67487 18290 67496
rect 17610 67482 17616 67484
rect 17672 67482 17696 67484
rect 17752 67482 17776 67484
rect 17832 67482 17856 67484
rect 17912 67482 17918 67484
rect 17672 67430 17674 67482
rect 17854 67430 17856 67482
rect 17610 67428 17616 67430
rect 17672 67428 17696 67430
rect 17752 67428 17776 67430
rect 17832 67428 17856 67430
rect 17912 67428 17918 67430
rect 17610 67419 17918 67428
rect 17610 66396 17918 66405
rect 17610 66394 17616 66396
rect 17672 66394 17696 66396
rect 17752 66394 17776 66396
rect 17832 66394 17856 66396
rect 17912 66394 17918 66396
rect 17672 66342 17674 66394
rect 17854 66342 17856 66394
rect 17610 66340 17616 66342
rect 17672 66340 17696 66342
rect 17752 66340 17776 66342
rect 17832 66340 17856 66342
rect 17912 66340 17918 66342
rect 17610 66331 17918 66340
rect 17500 66224 17552 66230
rect 17500 66166 17552 66172
rect 17408 66156 17460 66162
rect 17408 66098 17460 66104
rect 17420 65210 17448 66098
rect 17500 65952 17552 65958
rect 17500 65894 17552 65900
rect 17408 65204 17460 65210
rect 17408 65146 17460 65152
rect 17512 65113 17540 65894
rect 18236 65680 18288 65686
rect 18234 65648 18236 65657
rect 18288 65648 18290 65657
rect 18234 65583 18290 65592
rect 17610 65308 17918 65317
rect 17610 65306 17616 65308
rect 17672 65306 17696 65308
rect 17752 65306 17776 65308
rect 17832 65306 17856 65308
rect 17912 65306 17918 65308
rect 17672 65254 17674 65306
rect 17854 65254 17856 65306
rect 17610 65252 17616 65254
rect 17672 65252 17696 65254
rect 17752 65252 17776 65254
rect 17832 65252 17856 65254
rect 17912 65252 17918 65254
rect 17610 65243 17918 65252
rect 17592 65204 17644 65210
rect 17592 65146 17644 65152
rect 17236 65062 17356 65090
rect 17498 65104 17554 65113
rect 17040 64932 17092 64938
rect 17040 64874 17092 64880
rect 17236 64874 17264 65062
rect 17498 65039 17554 65048
rect 17408 64932 17460 64938
rect 17408 64874 17460 64880
rect 17604 64874 17632 65146
rect 16684 58398 16804 58426
rect 16868 64870 16988 64874
rect 16868 64864 17000 64870
rect 16868 64846 16948 64864
rect 16580 57520 16632 57526
rect 16580 57462 16632 57468
rect 16580 55344 16632 55350
rect 16580 55286 16632 55292
rect 16488 47048 16540 47054
rect 16488 46990 16540 46996
rect 16396 45076 16448 45082
rect 16396 45018 16448 45024
rect 16488 37868 16540 37874
rect 16488 37810 16540 37816
rect 16302 37360 16358 37369
rect 16302 37295 16358 37304
rect 16304 33992 16356 33998
rect 16304 33934 16356 33940
rect 16212 22160 16264 22166
rect 16212 22102 16264 22108
rect 16316 20330 16344 33934
rect 16500 33862 16528 37810
rect 16488 33856 16540 33862
rect 16488 33798 16540 33804
rect 16500 33658 16528 33798
rect 16488 33652 16540 33658
rect 16488 33594 16540 33600
rect 16488 33108 16540 33114
rect 16488 33050 16540 33056
rect 16500 32026 16528 33050
rect 16488 32020 16540 32026
rect 16488 31962 16540 31968
rect 16592 31906 16620 55286
rect 16684 48618 16712 58398
rect 16868 58290 16896 64846
rect 17236 64846 17356 64874
rect 16948 64806 17000 64812
rect 16950 64764 17258 64773
rect 16950 64762 16956 64764
rect 17012 64762 17036 64764
rect 17092 64762 17116 64764
rect 17172 64762 17196 64764
rect 17252 64762 17258 64764
rect 17012 64710 17014 64762
rect 17194 64710 17196 64762
rect 16950 64708 16956 64710
rect 17012 64708 17036 64710
rect 17092 64708 17116 64710
rect 17172 64708 17196 64710
rect 17252 64708 17258 64710
rect 16950 64699 17258 64708
rect 16950 63676 17258 63685
rect 16950 63674 16956 63676
rect 17012 63674 17036 63676
rect 17092 63674 17116 63676
rect 17172 63674 17196 63676
rect 17252 63674 17258 63676
rect 17012 63622 17014 63674
rect 17194 63622 17196 63674
rect 16950 63620 16956 63622
rect 17012 63620 17036 63622
rect 17092 63620 17116 63622
rect 17172 63620 17196 63622
rect 17252 63620 17258 63622
rect 16950 63611 17258 63620
rect 16950 62588 17258 62597
rect 16950 62586 16956 62588
rect 17012 62586 17036 62588
rect 17092 62586 17116 62588
rect 17172 62586 17196 62588
rect 17252 62586 17258 62588
rect 17012 62534 17014 62586
rect 17194 62534 17196 62586
rect 16950 62532 16956 62534
rect 17012 62532 17036 62534
rect 17092 62532 17116 62534
rect 17172 62532 17196 62534
rect 17252 62532 17258 62534
rect 16950 62523 17258 62532
rect 16950 61500 17258 61509
rect 16950 61498 16956 61500
rect 17012 61498 17036 61500
rect 17092 61498 17116 61500
rect 17172 61498 17196 61500
rect 17252 61498 17258 61500
rect 17012 61446 17014 61498
rect 17194 61446 17196 61498
rect 16950 61444 16956 61446
rect 17012 61444 17036 61446
rect 17092 61444 17116 61446
rect 17172 61444 17196 61446
rect 17252 61444 17258 61446
rect 16950 61435 17258 61444
rect 16950 60412 17258 60421
rect 16950 60410 16956 60412
rect 17012 60410 17036 60412
rect 17092 60410 17116 60412
rect 17172 60410 17196 60412
rect 17252 60410 17258 60412
rect 17012 60358 17014 60410
rect 17194 60358 17196 60410
rect 16950 60356 16956 60358
rect 17012 60356 17036 60358
rect 17092 60356 17116 60358
rect 17172 60356 17196 60358
rect 17252 60356 17258 60358
rect 16950 60347 17258 60356
rect 16950 59324 17258 59333
rect 16950 59322 16956 59324
rect 17012 59322 17036 59324
rect 17092 59322 17116 59324
rect 17172 59322 17196 59324
rect 17252 59322 17258 59324
rect 17012 59270 17014 59322
rect 17194 59270 17196 59322
rect 16950 59268 16956 59270
rect 17012 59268 17036 59270
rect 17092 59268 17116 59270
rect 17172 59268 17196 59270
rect 17252 59268 17258 59270
rect 16950 59259 17258 59268
rect 16776 58262 16896 58290
rect 16776 48657 16804 58262
rect 16950 58236 17258 58245
rect 16950 58234 16956 58236
rect 17012 58234 17036 58236
rect 17092 58234 17116 58236
rect 17172 58234 17196 58236
rect 17252 58234 17258 58236
rect 17012 58182 17014 58234
rect 17194 58182 17196 58234
rect 16950 58180 16956 58182
rect 17012 58180 17036 58182
rect 17092 58180 17116 58182
rect 17172 58180 17196 58182
rect 17252 58180 17258 58182
rect 16950 58171 17258 58180
rect 16856 57452 16908 57458
rect 16856 57394 16908 57400
rect 16868 55418 16896 57394
rect 16950 57148 17258 57157
rect 16950 57146 16956 57148
rect 17012 57146 17036 57148
rect 17092 57146 17116 57148
rect 17172 57146 17196 57148
rect 17252 57146 17258 57148
rect 17012 57094 17014 57146
rect 17194 57094 17196 57146
rect 16950 57092 16956 57094
rect 17012 57092 17036 57094
rect 17092 57092 17116 57094
rect 17172 57092 17196 57094
rect 17252 57092 17258 57094
rect 16950 57083 17258 57092
rect 16950 56060 17258 56069
rect 16950 56058 16956 56060
rect 17012 56058 17036 56060
rect 17092 56058 17116 56060
rect 17172 56058 17196 56060
rect 17252 56058 17258 56060
rect 17012 56006 17014 56058
rect 17194 56006 17196 56058
rect 16950 56004 16956 56006
rect 17012 56004 17036 56006
rect 17092 56004 17116 56006
rect 17172 56004 17196 56006
rect 17252 56004 17258 56006
rect 16950 55995 17258 56004
rect 17132 55684 17184 55690
rect 17132 55626 17184 55632
rect 16856 55412 16908 55418
rect 16856 55354 16908 55360
rect 16856 55276 16908 55282
rect 16856 55218 16908 55224
rect 16868 49774 16896 55218
rect 17144 55214 17172 55626
rect 17132 55208 17184 55214
rect 17132 55150 17184 55156
rect 16950 54972 17258 54981
rect 16950 54970 16956 54972
rect 17012 54970 17036 54972
rect 17092 54970 17116 54972
rect 17172 54970 17196 54972
rect 17252 54970 17258 54972
rect 17012 54918 17014 54970
rect 17194 54918 17196 54970
rect 16950 54916 16956 54918
rect 17012 54916 17036 54918
rect 17092 54916 17116 54918
rect 17172 54916 17196 54918
rect 17252 54916 17258 54918
rect 16950 54907 17258 54916
rect 16950 53884 17258 53893
rect 16950 53882 16956 53884
rect 17012 53882 17036 53884
rect 17092 53882 17116 53884
rect 17172 53882 17196 53884
rect 17252 53882 17258 53884
rect 17012 53830 17014 53882
rect 17194 53830 17196 53882
rect 16950 53828 16956 53830
rect 17012 53828 17036 53830
rect 17092 53828 17116 53830
rect 17172 53828 17196 53830
rect 17252 53828 17258 53830
rect 16950 53819 17258 53828
rect 16950 52796 17258 52805
rect 16950 52794 16956 52796
rect 17012 52794 17036 52796
rect 17092 52794 17116 52796
rect 17172 52794 17196 52796
rect 17252 52794 17258 52796
rect 17012 52742 17014 52794
rect 17194 52742 17196 52794
rect 16950 52740 16956 52742
rect 17012 52740 17036 52742
rect 17092 52740 17116 52742
rect 17172 52740 17196 52742
rect 17252 52740 17258 52742
rect 16950 52731 17258 52740
rect 16950 51708 17258 51717
rect 16950 51706 16956 51708
rect 17012 51706 17036 51708
rect 17092 51706 17116 51708
rect 17172 51706 17196 51708
rect 17252 51706 17258 51708
rect 17012 51654 17014 51706
rect 17194 51654 17196 51706
rect 16950 51652 16956 51654
rect 17012 51652 17036 51654
rect 17092 51652 17116 51654
rect 17172 51652 17196 51654
rect 17252 51652 17258 51654
rect 16950 51643 17258 51652
rect 16950 50620 17258 50629
rect 16950 50618 16956 50620
rect 17012 50618 17036 50620
rect 17092 50618 17116 50620
rect 17172 50618 17196 50620
rect 17252 50618 17258 50620
rect 17012 50566 17014 50618
rect 17194 50566 17196 50618
rect 16950 50564 16956 50566
rect 17012 50564 17036 50566
rect 17092 50564 17116 50566
rect 17172 50564 17196 50566
rect 17252 50564 17258 50566
rect 16950 50555 17258 50564
rect 16856 49768 16908 49774
rect 16856 49710 16908 49716
rect 16762 48648 16818 48657
rect 16672 48612 16724 48618
rect 16762 48583 16818 48592
rect 16672 48554 16724 48560
rect 16868 48498 16896 49710
rect 16950 49532 17258 49541
rect 16950 49530 16956 49532
rect 17012 49530 17036 49532
rect 17092 49530 17116 49532
rect 17172 49530 17196 49532
rect 17252 49530 17258 49532
rect 17012 49478 17014 49530
rect 17194 49478 17196 49530
rect 16950 49476 16956 49478
rect 17012 49476 17036 49478
rect 17092 49476 17116 49478
rect 17172 49476 17196 49478
rect 17252 49476 17258 49478
rect 16950 49467 17258 49476
rect 16408 31878 16620 31906
rect 16684 48470 16896 48498
rect 16408 30122 16436 31878
rect 16488 31816 16540 31822
rect 16488 31758 16540 31764
rect 16580 31816 16632 31822
rect 16580 31758 16632 31764
rect 16396 30116 16448 30122
rect 16396 30058 16448 30064
rect 16396 24744 16448 24750
rect 16394 24712 16396 24721
rect 16448 24712 16450 24721
rect 16394 24647 16450 24656
rect 16304 20324 16356 20330
rect 16304 20266 16356 20272
rect 16120 14068 16172 14074
rect 16120 14010 16172 14016
rect 16408 13326 16436 24647
rect 16500 20466 16528 31758
rect 16592 23662 16620 31758
rect 16684 23866 16712 48470
rect 16950 48444 17258 48453
rect 16950 48442 16956 48444
rect 17012 48442 17036 48444
rect 17092 48442 17116 48444
rect 17172 48442 17196 48444
rect 17252 48442 17258 48444
rect 17012 48390 17014 48442
rect 17194 48390 17196 48442
rect 16950 48388 16956 48390
rect 17012 48388 17036 48390
rect 17092 48388 17116 48390
rect 17172 48388 17196 48390
rect 17252 48388 17258 48390
rect 16950 48379 17258 48388
rect 16762 48240 16818 48249
rect 16762 48175 16818 48184
rect 16776 44742 16804 48175
rect 16950 47356 17258 47365
rect 16950 47354 16956 47356
rect 17012 47354 17036 47356
rect 17092 47354 17116 47356
rect 17172 47354 17196 47356
rect 17252 47354 17258 47356
rect 17012 47302 17014 47354
rect 17194 47302 17196 47354
rect 16950 47300 16956 47302
rect 17012 47300 17036 47302
rect 17092 47300 17116 47302
rect 17172 47300 17196 47302
rect 17252 47300 17258 47302
rect 16950 47291 17258 47300
rect 16856 46572 16908 46578
rect 16856 46514 16908 46520
rect 16764 44736 16816 44742
rect 16764 44678 16816 44684
rect 16764 42560 16816 42566
rect 16764 42502 16816 42508
rect 16776 39982 16804 42502
rect 16764 39976 16816 39982
rect 16764 39918 16816 39924
rect 16764 39840 16816 39846
rect 16764 39782 16816 39788
rect 16776 34241 16804 39782
rect 16762 34232 16818 34241
rect 16762 34167 16818 34176
rect 16764 34128 16816 34134
rect 16764 34070 16816 34076
rect 16776 31890 16804 34070
rect 16868 32994 16896 46514
rect 16950 46268 17258 46277
rect 16950 46266 16956 46268
rect 17012 46266 17036 46268
rect 17092 46266 17116 46268
rect 17172 46266 17196 46268
rect 17252 46266 17258 46268
rect 17012 46214 17014 46266
rect 17194 46214 17196 46266
rect 16950 46212 16956 46214
rect 17012 46212 17036 46214
rect 17092 46212 17116 46214
rect 17172 46212 17196 46214
rect 17252 46212 17258 46214
rect 16950 46203 17258 46212
rect 16950 45180 17258 45189
rect 16950 45178 16956 45180
rect 17012 45178 17036 45180
rect 17092 45178 17116 45180
rect 17172 45178 17196 45180
rect 17252 45178 17258 45180
rect 17012 45126 17014 45178
rect 17194 45126 17196 45178
rect 16950 45124 16956 45126
rect 17012 45124 17036 45126
rect 17092 45124 17116 45126
rect 17172 45124 17196 45126
rect 17252 45124 17258 45126
rect 16950 45115 17258 45124
rect 16950 44092 17258 44101
rect 16950 44090 16956 44092
rect 17012 44090 17036 44092
rect 17092 44090 17116 44092
rect 17172 44090 17196 44092
rect 17252 44090 17258 44092
rect 17012 44038 17014 44090
rect 17194 44038 17196 44090
rect 16950 44036 16956 44038
rect 17012 44036 17036 44038
rect 17092 44036 17116 44038
rect 17172 44036 17196 44038
rect 17252 44036 17258 44038
rect 16950 44027 17258 44036
rect 16950 43004 17258 43013
rect 16950 43002 16956 43004
rect 17012 43002 17036 43004
rect 17092 43002 17116 43004
rect 17172 43002 17196 43004
rect 17252 43002 17258 43004
rect 17012 42950 17014 43002
rect 17194 42950 17196 43002
rect 16950 42948 16956 42950
rect 17012 42948 17036 42950
rect 17092 42948 17116 42950
rect 17172 42948 17196 42950
rect 17252 42948 17258 42950
rect 16950 42939 17258 42948
rect 17328 42566 17356 64846
rect 17420 57322 17448 64874
rect 17512 64846 17632 64874
rect 17408 57316 17460 57322
rect 17408 57258 17460 57264
rect 17420 42650 17448 57258
rect 17512 42922 17540 64846
rect 17610 64220 17918 64229
rect 17610 64218 17616 64220
rect 17672 64218 17696 64220
rect 17752 64218 17776 64220
rect 17832 64218 17856 64220
rect 17912 64218 17918 64220
rect 17672 64166 17674 64218
rect 17854 64166 17856 64218
rect 17610 64164 17616 64166
rect 17672 64164 17696 64166
rect 17752 64164 17776 64166
rect 17832 64164 17856 64166
rect 17912 64164 17918 64166
rect 17610 64155 17918 64164
rect 18236 63776 18288 63782
rect 18234 63744 18236 63753
rect 18288 63744 18290 63753
rect 18234 63679 18290 63688
rect 17610 63132 17918 63141
rect 17610 63130 17616 63132
rect 17672 63130 17696 63132
rect 17752 63130 17776 63132
rect 17832 63130 17856 63132
rect 17912 63130 17918 63132
rect 17672 63078 17674 63130
rect 17854 63078 17856 63130
rect 17610 63076 17616 63078
rect 17672 63076 17696 63078
rect 17752 63076 17776 63078
rect 17832 63076 17856 63078
rect 17912 63076 17918 63078
rect 17610 63067 17918 63076
rect 18236 62144 18288 62150
rect 18236 62086 18288 62092
rect 17610 62044 17918 62053
rect 17610 62042 17616 62044
rect 17672 62042 17696 62044
rect 17752 62042 17776 62044
rect 17832 62042 17856 62044
rect 17912 62042 17918 62044
rect 17672 61990 17674 62042
rect 17854 61990 17856 62042
rect 17610 61988 17616 61990
rect 17672 61988 17696 61990
rect 17752 61988 17776 61990
rect 17832 61988 17856 61990
rect 17912 61988 17918 61990
rect 17610 61979 17918 61988
rect 18248 61849 18276 62086
rect 18234 61840 18290 61849
rect 18234 61775 18290 61784
rect 17960 61056 18012 61062
rect 17960 60998 18012 61004
rect 17610 60956 17918 60965
rect 17610 60954 17616 60956
rect 17672 60954 17696 60956
rect 17752 60954 17776 60956
rect 17832 60954 17856 60956
rect 17912 60954 17918 60956
rect 17672 60902 17674 60954
rect 17854 60902 17856 60954
rect 17610 60900 17616 60902
rect 17672 60900 17696 60902
rect 17752 60900 17776 60902
rect 17832 60900 17856 60902
rect 17912 60900 17918 60902
rect 17610 60891 17918 60900
rect 17610 59868 17918 59877
rect 17610 59866 17616 59868
rect 17672 59866 17696 59868
rect 17752 59866 17776 59868
rect 17832 59866 17856 59868
rect 17912 59866 17918 59868
rect 17672 59814 17674 59866
rect 17854 59814 17856 59866
rect 17610 59812 17616 59814
rect 17672 59812 17696 59814
rect 17752 59812 17776 59814
rect 17832 59812 17856 59814
rect 17912 59812 17918 59814
rect 17610 59803 17918 59812
rect 17610 58780 17918 58789
rect 17610 58778 17616 58780
rect 17672 58778 17696 58780
rect 17752 58778 17776 58780
rect 17832 58778 17856 58780
rect 17912 58778 17918 58780
rect 17672 58726 17674 58778
rect 17854 58726 17856 58778
rect 17610 58724 17616 58726
rect 17672 58724 17696 58726
rect 17752 58724 17776 58726
rect 17832 58724 17856 58726
rect 17912 58724 17918 58726
rect 17610 58715 17918 58724
rect 17610 57692 17918 57701
rect 17610 57690 17616 57692
rect 17672 57690 17696 57692
rect 17752 57690 17776 57692
rect 17832 57690 17856 57692
rect 17912 57690 17918 57692
rect 17672 57638 17674 57690
rect 17854 57638 17856 57690
rect 17610 57636 17616 57638
rect 17672 57636 17696 57638
rect 17752 57636 17776 57638
rect 17832 57636 17856 57638
rect 17912 57636 17918 57638
rect 17610 57627 17918 57636
rect 17972 56710 18000 60998
rect 18236 59968 18288 59974
rect 18234 59936 18236 59945
rect 18288 59936 18290 59945
rect 18234 59871 18290 59880
rect 18236 58336 18288 58342
rect 18236 58278 18288 58284
rect 18248 58041 18276 58278
rect 18234 58032 18290 58041
rect 18234 57967 18290 57976
rect 17960 56704 18012 56710
rect 17960 56646 18012 56652
rect 17610 56604 17918 56613
rect 17610 56602 17616 56604
rect 17672 56602 17696 56604
rect 17752 56602 17776 56604
rect 17832 56602 17856 56604
rect 17912 56602 17918 56604
rect 17672 56550 17674 56602
rect 17854 56550 17856 56602
rect 17610 56548 17616 56550
rect 17672 56548 17696 56550
rect 17752 56548 17776 56550
rect 17832 56548 17856 56550
rect 17912 56548 17918 56550
rect 17610 56539 17918 56548
rect 17610 55516 17918 55525
rect 17610 55514 17616 55516
rect 17672 55514 17696 55516
rect 17752 55514 17776 55516
rect 17832 55514 17856 55516
rect 17912 55514 17918 55516
rect 17672 55462 17674 55514
rect 17854 55462 17856 55514
rect 17610 55460 17616 55462
rect 17672 55460 17696 55462
rect 17752 55460 17776 55462
rect 17832 55460 17856 55462
rect 17912 55460 17918 55462
rect 17610 55451 17918 55460
rect 17972 55214 18000 56646
rect 18236 56160 18288 56166
rect 18234 56128 18236 56137
rect 18288 56128 18290 56137
rect 18234 56063 18290 56072
rect 17972 55186 18092 55214
rect 17610 54428 17918 54437
rect 17610 54426 17616 54428
rect 17672 54426 17696 54428
rect 17752 54426 17776 54428
rect 17832 54426 17856 54428
rect 17912 54426 17918 54428
rect 17672 54374 17674 54426
rect 17854 54374 17856 54426
rect 17610 54372 17616 54374
rect 17672 54372 17696 54374
rect 17752 54372 17776 54374
rect 17832 54372 17856 54374
rect 17912 54372 17918 54374
rect 17610 54363 17918 54372
rect 17610 53340 17918 53349
rect 17610 53338 17616 53340
rect 17672 53338 17696 53340
rect 17752 53338 17776 53340
rect 17832 53338 17856 53340
rect 17912 53338 17918 53340
rect 17672 53286 17674 53338
rect 17854 53286 17856 53338
rect 17610 53284 17616 53286
rect 17672 53284 17696 53286
rect 17752 53284 17776 53286
rect 17832 53284 17856 53286
rect 17912 53284 17918 53286
rect 17610 53275 17918 53284
rect 17960 52488 18012 52494
rect 17960 52430 18012 52436
rect 17610 52252 17918 52261
rect 17610 52250 17616 52252
rect 17672 52250 17696 52252
rect 17752 52250 17776 52252
rect 17832 52250 17856 52252
rect 17912 52250 17918 52252
rect 17672 52198 17674 52250
rect 17854 52198 17856 52250
rect 17610 52196 17616 52198
rect 17672 52196 17696 52198
rect 17752 52196 17776 52198
rect 17832 52196 17856 52198
rect 17912 52196 17918 52198
rect 17610 52187 17918 52196
rect 17610 51164 17918 51173
rect 17610 51162 17616 51164
rect 17672 51162 17696 51164
rect 17752 51162 17776 51164
rect 17832 51162 17856 51164
rect 17912 51162 17918 51164
rect 17672 51110 17674 51162
rect 17854 51110 17856 51162
rect 17610 51108 17616 51110
rect 17672 51108 17696 51110
rect 17752 51108 17776 51110
rect 17832 51108 17856 51110
rect 17912 51108 17918 51110
rect 17610 51099 17918 51108
rect 17610 50076 17918 50085
rect 17610 50074 17616 50076
rect 17672 50074 17696 50076
rect 17752 50074 17776 50076
rect 17832 50074 17856 50076
rect 17912 50074 17918 50076
rect 17672 50022 17674 50074
rect 17854 50022 17856 50074
rect 17610 50020 17616 50022
rect 17672 50020 17696 50022
rect 17752 50020 17776 50022
rect 17832 50020 17856 50022
rect 17912 50020 17918 50022
rect 17610 50011 17918 50020
rect 17610 48988 17918 48997
rect 17610 48986 17616 48988
rect 17672 48986 17696 48988
rect 17752 48986 17776 48988
rect 17832 48986 17856 48988
rect 17912 48986 17918 48988
rect 17672 48934 17674 48986
rect 17854 48934 17856 48986
rect 17610 48932 17616 48934
rect 17672 48932 17696 48934
rect 17752 48932 17776 48934
rect 17832 48932 17856 48934
rect 17912 48932 17918 48934
rect 17610 48923 17918 48932
rect 17610 47900 17918 47909
rect 17610 47898 17616 47900
rect 17672 47898 17696 47900
rect 17752 47898 17776 47900
rect 17832 47898 17856 47900
rect 17912 47898 17918 47900
rect 17672 47846 17674 47898
rect 17854 47846 17856 47898
rect 17610 47844 17616 47846
rect 17672 47844 17696 47846
rect 17752 47844 17776 47846
rect 17832 47844 17856 47846
rect 17912 47844 17918 47846
rect 17610 47835 17918 47844
rect 17610 46812 17918 46821
rect 17610 46810 17616 46812
rect 17672 46810 17696 46812
rect 17752 46810 17776 46812
rect 17832 46810 17856 46812
rect 17912 46810 17918 46812
rect 17672 46758 17674 46810
rect 17854 46758 17856 46810
rect 17610 46756 17616 46758
rect 17672 46756 17696 46758
rect 17752 46756 17776 46758
rect 17832 46756 17856 46758
rect 17912 46756 17918 46758
rect 17610 46747 17918 46756
rect 17610 45724 17918 45733
rect 17610 45722 17616 45724
rect 17672 45722 17696 45724
rect 17752 45722 17776 45724
rect 17832 45722 17856 45724
rect 17912 45722 17918 45724
rect 17672 45670 17674 45722
rect 17854 45670 17856 45722
rect 17610 45668 17616 45670
rect 17672 45668 17696 45670
rect 17752 45668 17776 45670
rect 17832 45668 17856 45670
rect 17912 45668 17918 45670
rect 17610 45659 17918 45668
rect 17610 44636 17918 44645
rect 17610 44634 17616 44636
rect 17672 44634 17696 44636
rect 17752 44634 17776 44636
rect 17832 44634 17856 44636
rect 17912 44634 17918 44636
rect 17672 44582 17674 44634
rect 17854 44582 17856 44634
rect 17610 44580 17616 44582
rect 17672 44580 17696 44582
rect 17752 44580 17776 44582
rect 17832 44580 17856 44582
rect 17912 44580 17918 44582
rect 17610 44571 17918 44580
rect 17610 43548 17918 43557
rect 17610 43546 17616 43548
rect 17672 43546 17696 43548
rect 17752 43546 17776 43548
rect 17832 43546 17856 43548
rect 17912 43546 17918 43548
rect 17672 43494 17674 43546
rect 17854 43494 17856 43546
rect 17610 43492 17616 43494
rect 17672 43492 17696 43494
rect 17752 43492 17776 43494
rect 17832 43492 17856 43494
rect 17912 43492 17918 43494
rect 17610 43483 17918 43492
rect 17512 42894 17632 42922
rect 17420 42622 17540 42650
rect 17316 42560 17368 42566
rect 17316 42502 17368 42508
rect 17408 42560 17460 42566
rect 17408 42502 17460 42508
rect 17316 42288 17368 42294
rect 17316 42230 17368 42236
rect 16950 41916 17258 41925
rect 16950 41914 16956 41916
rect 17012 41914 17036 41916
rect 17092 41914 17116 41916
rect 17172 41914 17196 41916
rect 17252 41914 17258 41916
rect 17012 41862 17014 41914
rect 17194 41862 17196 41914
rect 16950 41860 16956 41862
rect 17012 41860 17036 41862
rect 17092 41860 17116 41862
rect 17172 41860 17196 41862
rect 17252 41860 17258 41862
rect 16950 41851 17258 41860
rect 16950 40828 17258 40837
rect 16950 40826 16956 40828
rect 17012 40826 17036 40828
rect 17092 40826 17116 40828
rect 17172 40826 17196 40828
rect 17252 40826 17258 40828
rect 17012 40774 17014 40826
rect 17194 40774 17196 40826
rect 16950 40772 16956 40774
rect 17012 40772 17036 40774
rect 17092 40772 17116 40774
rect 17172 40772 17196 40774
rect 17252 40772 17258 40774
rect 16950 40763 17258 40772
rect 16946 40624 17002 40633
rect 16946 40559 17002 40568
rect 16960 39846 16988 40559
rect 16948 39840 17000 39846
rect 16948 39782 17000 39788
rect 16950 39740 17258 39749
rect 16950 39738 16956 39740
rect 17012 39738 17036 39740
rect 17092 39738 17116 39740
rect 17172 39738 17196 39740
rect 17252 39738 17258 39740
rect 17012 39686 17014 39738
rect 17194 39686 17196 39738
rect 16950 39684 16956 39686
rect 17012 39684 17036 39686
rect 17092 39684 17116 39686
rect 17172 39684 17196 39686
rect 17252 39684 17258 39686
rect 16950 39675 17258 39684
rect 17328 38962 17356 42230
rect 17316 38956 17368 38962
rect 17316 38898 17368 38904
rect 17316 38752 17368 38758
rect 17316 38694 17368 38700
rect 16950 38652 17258 38661
rect 16950 38650 16956 38652
rect 17012 38650 17036 38652
rect 17092 38650 17116 38652
rect 17172 38650 17196 38652
rect 17252 38650 17258 38652
rect 17012 38598 17014 38650
rect 17194 38598 17196 38650
rect 16950 38596 16956 38598
rect 17012 38596 17036 38598
rect 17092 38596 17116 38598
rect 17172 38596 17196 38598
rect 17252 38596 17258 38598
rect 16950 38587 17258 38596
rect 16950 37564 17258 37573
rect 16950 37562 16956 37564
rect 17012 37562 17036 37564
rect 17092 37562 17116 37564
rect 17172 37562 17196 37564
rect 17252 37562 17258 37564
rect 17012 37510 17014 37562
rect 17194 37510 17196 37562
rect 16950 37508 16956 37510
rect 17012 37508 17036 37510
rect 17092 37508 17116 37510
rect 17172 37508 17196 37510
rect 17252 37508 17258 37510
rect 16950 37499 17258 37508
rect 16950 36476 17258 36485
rect 16950 36474 16956 36476
rect 17012 36474 17036 36476
rect 17092 36474 17116 36476
rect 17172 36474 17196 36476
rect 17252 36474 17258 36476
rect 17012 36422 17014 36474
rect 17194 36422 17196 36474
rect 16950 36420 16956 36422
rect 17012 36420 17036 36422
rect 17092 36420 17116 36422
rect 17172 36420 17196 36422
rect 17252 36420 17258 36422
rect 16950 36411 17258 36420
rect 16950 35388 17258 35397
rect 16950 35386 16956 35388
rect 17012 35386 17036 35388
rect 17092 35386 17116 35388
rect 17172 35386 17196 35388
rect 17252 35386 17258 35388
rect 17012 35334 17014 35386
rect 17194 35334 17196 35386
rect 16950 35332 16956 35334
rect 17012 35332 17036 35334
rect 17092 35332 17116 35334
rect 17172 35332 17196 35334
rect 17252 35332 17258 35334
rect 16950 35323 17258 35332
rect 16950 34300 17258 34309
rect 16950 34298 16956 34300
rect 17012 34298 17036 34300
rect 17092 34298 17116 34300
rect 17172 34298 17196 34300
rect 17252 34298 17258 34300
rect 17012 34246 17014 34298
rect 17194 34246 17196 34298
rect 16950 34244 16956 34246
rect 17012 34244 17036 34246
rect 17092 34244 17116 34246
rect 17172 34244 17196 34246
rect 17252 34244 17258 34246
rect 16950 34235 17258 34244
rect 16950 33212 17258 33221
rect 16950 33210 16956 33212
rect 17012 33210 17036 33212
rect 17092 33210 17116 33212
rect 17172 33210 17196 33212
rect 17252 33210 17258 33212
rect 17012 33158 17014 33210
rect 17194 33158 17196 33210
rect 16950 33156 16956 33158
rect 17012 33156 17036 33158
rect 17092 33156 17116 33158
rect 17172 33156 17196 33158
rect 17252 33156 17258 33158
rect 16950 33147 17258 33156
rect 16868 32966 16988 32994
rect 16856 32904 16908 32910
rect 16856 32846 16908 32852
rect 16868 32434 16896 32846
rect 16856 32428 16908 32434
rect 16856 32370 16908 32376
rect 16764 31884 16816 31890
rect 16764 31826 16816 31832
rect 16762 31784 16818 31793
rect 16762 31719 16818 31728
rect 16672 23860 16724 23866
rect 16672 23802 16724 23808
rect 16776 23712 16804 31719
rect 16868 31346 16896 32370
rect 16960 32337 16988 32966
rect 16946 32328 17002 32337
rect 16946 32263 17002 32272
rect 16950 32124 17258 32133
rect 16950 32122 16956 32124
rect 17012 32122 17036 32124
rect 17092 32122 17116 32124
rect 17172 32122 17196 32124
rect 17252 32122 17258 32124
rect 17012 32070 17014 32122
rect 17194 32070 17196 32122
rect 16950 32068 16956 32070
rect 17012 32068 17036 32070
rect 17092 32068 17116 32070
rect 17172 32068 17196 32070
rect 17252 32068 17258 32070
rect 16950 32059 17258 32068
rect 16856 31340 16908 31346
rect 16856 31282 16908 31288
rect 16950 31036 17258 31045
rect 16950 31034 16956 31036
rect 17012 31034 17036 31036
rect 17092 31034 17116 31036
rect 17172 31034 17196 31036
rect 17252 31034 17258 31036
rect 17012 30982 17014 31034
rect 17194 30982 17196 31034
rect 16950 30980 16956 30982
rect 17012 30980 17036 30982
rect 17092 30980 17116 30982
rect 17172 30980 17196 30982
rect 17252 30980 17258 30982
rect 16950 30971 17258 30980
rect 16950 29948 17258 29957
rect 16950 29946 16956 29948
rect 17012 29946 17036 29948
rect 17092 29946 17116 29948
rect 17172 29946 17196 29948
rect 17252 29946 17258 29948
rect 17012 29894 17014 29946
rect 17194 29894 17196 29946
rect 16950 29892 16956 29894
rect 17012 29892 17036 29894
rect 17092 29892 17116 29894
rect 17172 29892 17196 29894
rect 17252 29892 17258 29894
rect 16950 29883 17258 29892
rect 16950 28860 17258 28869
rect 16950 28858 16956 28860
rect 17012 28858 17036 28860
rect 17092 28858 17116 28860
rect 17172 28858 17196 28860
rect 17252 28858 17258 28860
rect 17012 28806 17014 28858
rect 17194 28806 17196 28858
rect 16950 28804 16956 28806
rect 17012 28804 17036 28806
rect 17092 28804 17116 28806
rect 17172 28804 17196 28806
rect 17252 28804 17258 28806
rect 16950 28795 17258 28804
rect 16950 27772 17258 27781
rect 16950 27770 16956 27772
rect 17012 27770 17036 27772
rect 17092 27770 17116 27772
rect 17172 27770 17196 27772
rect 17252 27770 17258 27772
rect 17012 27718 17014 27770
rect 17194 27718 17196 27770
rect 16950 27716 16956 27718
rect 17012 27716 17036 27718
rect 17092 27716 17116 27718
rect 17172 27716 17196 27718
rect 17252 27716 17258 27718
rect 16950 27707 17258 27716
rect 16950 26684 17258 26693
rect 16950 26682 16956 26684
rect 17012 26682 17036 26684
rect 17092 26682 17116 26684
rect 17172 26682 17196 26684
rect 17252 26682 17258 26684
rect 17012 26630 17014 26682
rect 17194 26630 17196 26682
rect 16950 26628 16956 26630
rect 17012 26628 17036 26630
rect 17092 26628 17116 26630
rect 17172 26628 17196 26630
rect 17252 26628 17258 26630
rect 16950 26619 17258 26628
rect 16950 25596 17258 25605
rect 16950 25594 16956 25596
rect 17012 25594 17036 25596
rect 17092 25594 17116 25596
rect 17172 25594 17196 25596
rect 17252 25594 17258 25596
rect 17012 25542 17014 25594
rect 17194 25542 17196 25594
rect 16950 25540 16956 25542
rect 17012 25540 17036 25542
rect 17092 25540 17116 25542
rect 17172 25540 17196 25542
rect 17252 25540 17258 25542
rect 16950 25531 17258 25540
rect 16950 24508 17258 24517
rect 16950 24506 16956 24508
rect 17012 24506 17036 24508
rect 17092 24506 17116 24508
rect 17172 24506 17196 24508
rect 17252 24506 17258 24508
rect 17012 24454 17014 24506
rect 17194 24454 17196 24506
rect 16950 24452 16956 24454
rect 17012 24452 17036 24454
rect 17092 24452 17116 24454
rect 17172 24452 17196 24454
rect 17252 24452 17258 24454
rect 16950 24443 17258 24452
rect 16684 23684 16804 23712
rect 16580 23656 16632 23662
rect 16580 23598 16632 23604
rect 16684 23508 16712 23684
rect 16946 23624 17002 23633
rect 16946 23559 16948 23568
rect 17000 23559 17002 23568
rect 16948 23530 17000 23536
rect 16592 23480 16712 23508
rect 16764 23520 16816 23526
rect 16488 20460 16540 20466
rect 16488 20402 16540 20408
rect 16592 15434 16620 23480
rect 16764 23462 16816 23468
rect 16776 19334 16804 23462
rect 16950 23420 17258 23429
rect 16950 23418 16956 23420
rect 17012 23418 17036 23420
rect 17092 23418 17116 23420
rect 17172 23418 17196 23420
rect 17252 23418 17258 23420
rect 17012 23366 17014 23418
rect 17194 23366 17196 23418
rect 16950 23364 16956 23366
rect 17012 23364 17036 23366
rect 17092 23364 17116 23366
rect 17172 23364 17196 23366
rect 17252 23364 17258 23366
rect 16950 23355 17258 23364
rect 17222 22536 17278 22545
rect 17222 22471 17224 22480
rect 17276 22471 17278 22480
rect 17224 22442 17276 22448
rect 16950 22332 17258 22341
rect 16950 22330 16956 22332
rect 17012 22330 17036 22332
rect 17092 22330 17116 22332
rect 17172 22330 17196 22332
rect 17252 22330 17258 22332
rect 17012 22278 17014 22330
rect 17194 22278 17196 22330
rect 16950 22276 16956 22278
rect 17012 22276 17036 22278
rect 17092 22276 17116 22278
rect 17172 22276 17196 22278
rect 17252 22276 17258 22278
rect 16950 22267 17258 22276
rect 16950 21244 17258 21253
rect 16950 21242 16956 21244
rect 17012 21242 17036 21244
rect 17092 21242 17116 21244
rect 17172 21242 17196 21244
rect 17252 21242 17258 21244
rect 17012 21190 17014 21242
rect 17194 21190 17196 21242
rect 16950 21188 16956 21190
rect 17012 21188 17036 21190
rect 17092 21188 17116 21190
rect 17172 21188 17196 21190
rect 17252 21188 17258 21190
rect 16950 21179 17258 21188
rect 17222 21040 17278 21049
rect 17222 20975 17278 20984
rect 17236 20602 17264 20975
rect 17224 20596 17276 20602
rect 17224 20538 17276 20544
rect 16856 20324 16908 20330
rect 16856 20266 16908 20272
rect 16868 20058 16896 20266
rect 16950 20156 17258 20165
rect 16950 20154 16956 20156
rect 17012 20154 17036 20156
rect 17092 20154 17116 20156
rect 17172 20154 17196 20156
rect 17252 20154 17258 20156
rect 17012 20102 17014 20154
rect 17194 20102 17196 20154
rect 16950 20100 16956 20102
rect 17012 20100 17036 20102
rect 17092 20100 17116 20102
rect 17172 20100 17196 20102
rect 17252 20100 17258 20102
rect 16950 20091 17258 20100
rect 16856 20052 16908 20058
rect 16856 19994 16908 20000
rect 16684 19306 16804 19334
rect 16580 15428 16632 15434
rect 16580 15370 16632 15376
rect 16396 13320 16448 13326
rect 16396 13262 16448 13268
rect 16578 13288 16634 13297
rect 16578 13223 16634 13232
rect 16592 13190 16620 13223
rect 16580 13184 16632 13190
rect 16580 13126 16632 13132
rect 16028 11076 16080 11082
rect 16028 11018 16080 11024
rect 15936 9988 15988 9994
rect 15936 9930 15988 9936
rect 15384 9580 15436 9586
rect 15384 9522 15436 9528
rect 14648 8628 14700 8634
rect 14648 8570 14700 8576
rect 14556 8560 14608 8566
rect 14556 8502 14608 8508
rect 16210 5264 16266 5273
rect 16210 5199 16212 5208
rect 16264 5199 16266 5208
rect 16212 5170 16264 5176
rect 14464 4616 14516 4622
rect 14464 4558 14516 4564
rect 12610 4380 12918 4389
rect 12610 4378 12616 4380
rect 12672 4378 12696 4380
rect 12752 4378 12776 4380
rect 12832 4378 12856 4380
rect 12912 4378 12918 4380
rect 12672 4326 12674 4378
rect 12854 4326 12856 4378
rect 12610 4324 12616 4326
rect 12672 4324 12696 4326
rect 12752 4324 12776 4326
rect 12832 4324 12856 4326
rect 12912 4324 12918 4326
rect 12610 4315 12918 4324
rect 11950 3836 12258 3845
rect 11950 3834 11956 3836
rect 12012 3834 12036 3836
rect 12092 3834 12116 3836
rect 12172 3834 12196 3836
rect 12252 3834 12258 3836
rect 12012 3782 12014 3834
rect 12194 3782 12196 3834
rect 11950 3780 11956 3782
rect 12012 3780 12036 3782
rect 12092 3780 12116 3782
rect 12172 3780 12196 3782
rect 12252 3780 12258 3782
rect 11950 3771 12258 3780
rect 11704 3596 11756 3602
rect 11704 3538 11756 3544
rect 12610 3292 12918 3301
rect 12610 3290 12616 3292
rect 12672 3290 12696 3292
rect 12752 3290 12776 3292
rect 12832 3290 12856 3292
rect 12912 3290 12918 3292
rect 12672 3238 12674 3290
rect 12854 3238 12856 3290
rect 12610 3236 12616 3238
rect 12672 3236 12696 3238
rect 12752 3236 12776 3238
rect 12832 3236 12856 3238
rect 12912 3236 12918 3238
rect 12610 3227 12918 3236
rect 11950 2748 12258 2757
rect 11950 2746 11956 2748
rect 12012 2746 12036 2748
rect 12092 2746 12116 2748
rect 12172 2746 12196 2748
rect 12252 2746 12258 2748
rect 12012 2694 12014 2746
rect 12194 2694 12196 2746
rect 11950 2692 11956 2694
rect 12012 2692 12036 2694
rect 12092 2692 12116 2694
rect 12172 2692 12196 2694
rect 12252 2692 12258 2694
rect 11950 2683 12258 2692
rect 14476 2650 14504 4558
rect 16684 4146 16712 19306
rect 16950 19068 17258 19077
rect 16950 19066 16956 19068
rect 17012 19066 17036 19068
rect 17092 19066 17116 19068
rect 17172 19066 17196 19068
rect 17252 19066 17258 19068
rect 17012 19014 17014 19066
rect 17194 19014 17196 19066
rect 16950 19012 16956 19014
rect 17012 19012 17036 19014
rect 17092 19012 17116 19014
rect 17172 19012 17196 19014
rect 17252 19012 17258 19014
rect 16950 19003 17258 19012
rect 16950 17980 17258 17989
rect 16950 17978 16956 17980
rect 17012 17978 17036 17980
rect 17092 17978 17116 17980
rect 17172 17978 17196 17980
rect 17252 17978 17258 17980
rect 17012 17926 17014 17978
rect 17194 17926 17196 17978
rect 16950 17924 16956 17926
rect 17012 17924 17036 17926
rect 17092 17924 17116 17926
rect 17172 17924 17196 17926
rect 17252 17924 17258 17926
rect 16950 17915 17258 17924
rect 16950 16892 17258 16901
rect 16950 16890 16956 16892
rect 17012 16890 17036 16892
rect 17092 16890 17116 16892
rect 17172 16890 17196 16892
rect 17252 16890 17258 16892
rect 17012 16838 17014 16890
rect 17194 16838 17196 16890
rect 16950 16836 16956 16838
rect 17012 16836 17036 16838
rect 17092 16836 17116 16838
rect 17172 16836 17196 16838
rect 17252 16836 17258 16838
rect 16950 16827 17258 16836
rect 16950 15804 17258 15813
rect 16950 15802 16956 15804
rect 17012 15802 17036 15804
rect 17092 15802 17116 15804
rect 17172 15802 17196 15804
rect 17252 15802 17258 15804
rect 17012 15750 17014 15802
rect 17194 15750 17196 15802
rect 16950 15748 16956 15750
rect 17012 15748 17036 15750
rect 17092 15748 17116 15750
rect 17172 15748 17196 15750
rect 17252 15748 17258 15750
rect 16950 15739 17258 15748
rect 16856 15496 16908 15502
rect 16856 15438 16908 15444
rect 16868 13802 16896 15438
rect 16950 14716 17258 14725
rect 16950 14714 16956 14716
rect 17012 14714 17036 14716
rect 17092 14714 17116 14716
rect 17172 14714 17196 14716
rect 17252 14714 17258 14716
rect 17012 14662 17014 14714
rect 17194 14662 17196 14714
rect 16950 14660 16956 14662
rect 17012 14660 17036 14662
rect 17092 14660 17116 14662
rect 17172 14660 17196 14662
rect 17252 14660 17258 14662
rect 16950 14651 17258 14660
rect 16856 13796 16908 13802
rect 16856 13738 16908 13744
rect 16868 12850 16896 13738
rect 16950 13628 17258 13637
rect 16950 13626 16956 13628
rect 17012 13626 17036 13628
rect 17092 13626 17116 13628
rect 17172 13626 17196 13628
rect 17252 13626 17258 13628
rect 17012 13574 17014 13626
rect 17194 13574 17196 13626
rect 16950 13572 16956 13574
rect 17012 13572 17036 13574
rect 17092 13572 17116 13574
rect 17172 13572 17196 13574
rect 17252 13572 17258 13574
rect 16950 13563 17258 13572
rect 17328 12918 17356 38694
rect 17420 36802 17448 42502
rect 17512 36922 17540 42622
rect 17604 42566 17632 42894
rect 17592 42560 17644 42566
rect 17592 42502 17644 42508
rect 17610 42460 17918 42469
rect 17610 42458 17616 42460
rect 17672 42458 17696 42460
rect 17752 42458 17776 42460
rect 17832 42458 17856 42460
rect 17912 42458 17918 42460
rect 17672 42406 17674 42458
rect 17854 42406 17856 42458
rect 17610 42404 17616 42406
rect 17672 42404 17696 42406
rect 17752 42404 17776 42406
rect 17832 42404 17856 42406
rect 17912 42404 17918 42406
rect 17610 42395 17918 42404
rect 17610 41372 17918 41381
rect 17610 41370 17616 41372
rect 17672 41370 17696 41372
rect 17752 41370 17776 41372
rect 17832 41370 17856 41372
rect 17912 41370 17918 41372
rect 17672 41318 17674 41370
rect 17854 41318 17856 41370
rect 17610 41316 17616 41318
rect 17672 41316 17696 41318
rect 17752 41316 17776 41318
rect 17832 41316 17856 41318
rect 17912 41316 17918 41318
rect 17610 41307 17918 41316
rect 17610 40284 17918 40293
rect 17610 40282 17616 40284
rect 17672 40282 17696 40284
rect 17752 40282 17776 40284
rect 17832 40282 17856 40284
rect 17912 40282 17918 40284
rect 17672 40230 17674 40282
rect 17854 40230 17856 40282
rect 17610 40228 17616 40230
rect 17672 40228 17696 40230
rect 17752 40228 17776 40230
rect 17832 40228 17856 40230
rect 17912 40228 17918 40230
rect 17610 40219 17918 40228
rect 17610 39196 17918 39205
rect 17610 39194 17616 39196
rect 17672 39194 17696 39196
rect 17752 39194 17776 39196
rect 17832 39194 17856 39196
rect 17912 39194 17918 39196
rect 17672 39142 17674 39194
rect 17854 39142 17856 39194
rect 17610 39140 17616 39142
rect 17672 39140 17696 39142
rect 17752 39140 17776 39142
rect 17832 39140 17856 39142
rect 17912 39140 17918 39142
rect 17610 39131 17918 39140
rect 17610 38108 17918 38117
rect 17610 38106 17616 38108
rect 17672 38106 17696 38108
rect 17752 38106 17776 38108
rect 17832 38106 17856 38108
rect 17912 38106 17918 38108
rect 17672 38054 17674 38106
rect 17854 38054 17856 38106
rect 17610 38052 17616 38054
rect 17672 38052 17696 38054
rect 17752 38052 17776 38054
rect 17832 38052 17856 38054
rect 17912 38052 17918 38054
rect 17610 38043 17918 38052
rect 17610 37020 17918 37029
rect 17610 37018 17616 37020
rect 17672 37018 17696 37020
rect 17752 37018 17776 37020
rect 17832 37018 17856 37020
rect 17912 37018 17918 37020
rect 17672 36966 17674 37018
rect 17854 36966 17856 37018
rect 17610 36964 17616 36966
rect 17672 36964 17696 36966
rect 17752 36964 17776 36966
rect 17832 36964 17856 36966
rect 17912 36964 17918 36966
rect 17610 36955 17918 36964
rect 17500 36916 17552 36922
rect 17500 36858 17552 36864
rect 17420 36774 17540 36802
rect 17408 36712 17460 36718
rect 17408 36654 17460 36660
rect 17420 34474 17448 36654
rect 17408 34468 17460 34474
rect 17408 34410 17460 34416
rect 17420 34066 17448 34410
rect 17408 34060 17460 34066
rect 17408 34002 17460 34008
rect 17406 33960 17462 33969
rect 17406 33895 17462 33904
rect 17316 12912 17368 12918
rect 17316 12854 17368 12860
rect 16856 12844 16908 12850
rect 16856 12786 16908 12792
rect 16950 12540 17258 12549
rect 16950 12538 16956 12540
rect 17012 12538 17036 12540
rect 17092 12538 17116 12540
rect 17172 12538 17196 12540
rect 17252 12538 17258 12540
rect 17012 12486 17014 12538
rect 17194 12486 17196 12538
rect 16950 12484 16956 12486
rect 17012 12484 17036 12486
rect 17092 12484 17116 12486
rect 17172 12484 17196 12486
rect 17252 12484 17258 12486
rect 16950 12475 17258 12484
rect 16950 11452 17258 11461
rect 16950 11450 16956 11452
rect 17012 11450 17036 11452
rect 17092 11450 17116 11452
rect 17172 11450 17196 11452
rect 17252 11450 17258 11452
rect 17012 11398 17014 11450
rect 17194 11398 17196 11450
rect 16950 11396 16956 11398
rect 17012 11396 17036 11398
rect 17092 11396 17116 11398
rect 17172 11396 17196 11398
rect 17252 11396 17258 11398
rect 16950 11387 17258 11396
rect 16950 10364 17258 10373
rect 16950 10362 16956 10364
rect 17012 10362 17036 10364
rect 17092 10362 17116 10364
rect 17172 10362 17196 10364
rect 17252 10362 17258 10364
rect 17012 10310 17014 10362
rect 17194 10310 17196 10362
rect 16950 10308 16956 10310
rect 17012 10308 17036 10310
rect 17092 10308 17116 10310
rect 17172 10308 17196 10310
rect 17252 10308 17258 10310
rect 16950 10299 17258 10308
rect 16950 9276 17258 9285
rect 16950 9274 16956 9276
rect 17012 9274 17036 9276
rect 17092 9274 17116 9276
rect 17172 9274 17196 9276
rect 17252 9274 17258 9276
rect 17012 9222 17014 9274
rect 17194 9222 17196 9274
rect 16950 9220 16956 9222
rect 17012 9220 17036 9222
rect 17092 9220 17116 9222
rect 17172 9220 17196 9222
rect 17252 9220 17258 9222
rect 16950 9211 17258 9220
rect 17420 9178 17448 33895
rect 17512 30258 17540 36774
rect 17610 35932 17918 35941
rect 17610 35930 17616 35932
rect 17672 35930 17696 35932
rect 17752 35930 17776 35932
rect 17832 35930 17856 35932
rect 17912 35930 17918 35932
rect 17672 35878 17674 35930
rect 17854 35878 17856 35930
rect 17610 35876 17616 35878
rect 17672 35876 17696 35878
rect 17752 35876 17776 35878
rect 17832 35876 17856 35878
rect 17912 35876 17918 35878
rect 17610 35867 17918 35876
rect 17610 34844 17918 34853
rect 17610 34842 17616 34844
rect 17672 34842 17696 34844
rect 17752 34842 17776 34844
rect 17832 34842 17856 34844
rect 17912 34842 17918 34844
rect 17672 34790 17674 34842
rect 17854 34790 17856 34842
rect 17610 34788 17616 34790
rect 17672 34788 17696 34790
rect 17752 34788 17776 34790
rect 17832 34788 17856 34790
rect 17912 34788 17918 34790
rect 17610 34779 17918 34788
rect 17610 33756 17918 33765
rect 17610 33754 17616 33756
rect 17672 33754 17696 33756
rect 17752 33754 17776 33756
rect 17832 33754 17856 33756
rect 17912 33754 17918 33756
rect 17672 33702 17674 33754
rect 17854 33702 17856 33754
rect 17610 33700 17616 33702
rect 17672 33700 17696 33702
rect 17752 33700 17776 33702
rect 17832 33700 17856 33702
rect 17912 33700 17918 33702
rect 17610 33691 17918 33700
rect 17610 32668 17918 32677
rect 17610 32666 17616 32668
rect 17672 32666 17696 32668
rect 17752 32666 17776 32668
rect 17832 32666 17856 32668
rect 17912 32666 17918 32668
rect 17672 32614 17674 32666
rect 17854 32614 17856 32666
rect 17610 32612 17616 32614
rect 17672 32612 17696 32614
rect 17752 32612 17776 32614
rect 17832 32612 17856 32614
rect 17912 32612 17918 32614
rect 17610 32603 17918 32612
rect 17972 32230 18000 52430
rect 18064 37262 18092 55186
rect 18144 54664 18196 54670
rect 18144 54606 18196 54612
rect 18156 44282 18184 54606
rect 18236 54528 18288 54534
rect 18236 54470 18288 54476
rect 18248 54233 18276 54470
rect 18234 54224 18290 54233
rect 18234 54159 18290 54168
rect 18236 52624 18288 52630
rect 18236 52566 18288 52572
rect 18248 52329 18276 52566
rect 18234 52320 18290 52329
rect 18234 52255 18290 52264
rect 18236 50720 18288 50726
rect 18236 50662 18288 50668
rect 18248 50425 18276 50662
rect 18234 50416 18290 50425
rect 18234 50351 18290 50360
rect 18236 48544 18288 48550
rect 18234 48512 18236 48521
rect 18288 48512 18290 48521
rect 18234 48447 18290 48456
rect 18236 46912 18288 46918
rect 18236 46854 18288 46860
rect 18248 46617 18276 46854
rect 18234 46608 18290 46617
rect 18234 46543 18290 46552
rect 18236 44736 18288 44742
rect 18234 44704 18236 44713
rect 18288 44704 18290 44713
rect 18234 44639 18290 44648
rect 18340 44402 18368 77454
rect 18788 74656 18840 74662
rect 18788 74598 18840 74604
rect 18420 64932 18472 64938
rect 18420 64874 18472 64880
rect 18328 44396 18380 44402
rect 18328 44338 18380 44344
rect 18156 44254 18368 44282
rect 18144 44192 18196 44198
rect 18144 44134 18196 44140
rect 18052 37256 18104 37262
rect 18052 37198 18104 37204
rect 18052 36100 18104 36106
rect 18052 36042 18104 36048
rect 17960 32224 18012 32230
rect 17960 32166 18012 32172
rect 18064 31822 18092 36042
rect 18052 31816 18104 31822
rect 18052 31758 18104 31764
rect 17610 31580 17918 31589
rect 17610 31578 17616 31580
rect 17672 31578 17696 31580
rect 17752 31578 17776 31580
rect 17832 31578 17856 31580
rect 17912 31578 17918 31580
rect 17672 31526 17674 31578
rect 17854 31526 17856 31578
rect 17610 31524 17616 31526
rect 17672 31524 17696 31526
rect 17752 31524 17776 31526
rect 17832 31524 17856 31526
rect 17912 31524 17918 31526
rect 17610 31515 17918 31524
rect 17610 30492 17918 30501
rect 17610 30490 17616 30492
rect 17672 30490 17696 30492
rect 17752 30490 17776 30492
rect 17832 30490 17856 30492
rect 17912 30490 17918 30492
rect 17672 30438 17674 30490
rect 17854 30438 17856 30490
rect 17610 30436 17616 30438
rect 17672 30436 17696 30438
rect 17752 30436 17776 30438
rect 17832 30436 17856 30438
rect 17912 30436 17918 30438
rect 17610 30427 17918 30436
rect 17500 30252 17552 30258
rect 17500 30194 17552 30200
rect 17960 29708 18012 29714
rect 17960 29650 18012 29656
rect 17610 29404 17918 29413
rect 17610 29402 17616 29404
rect 17672 29402 17696 29404
rect 17752 29402 17776 29404
rect 17832 29402 17856 29404
rect 17912 29402 17918 29404
rect 17672 29350 17674 29402
rect 17854 29350 17856 29402
rect 17610 29348 17616 29350
rect 17672 29348 17696 29350
rect 17752 29348 17776 29350
rect 17832 29348 17856 29350
rect 17912 29348 17918 29350
rect 17610 29339 17918 29348
rect 17610 28316 17918 28325
rect 17610 28314 17616 28316
rect 17672 28314 17696 28316
rect 17752 28314 17776 28316
rect 17832 28314 17856 28316
rect 17912 28314 17918 28316
rect 17672 28262 17674 28314
rect 17854 28262 17856 28314
rect 17610 28260 17616 28262
rect 17672 28260 17696 28262
rect 17752 28260 17776 28262
rect 17832 28260 17856 28262
rect 17912 28260 17918 28262
rect 17610 28251 17918 28260
rect 17868 27872 17920 27878
rect 17868 27814 17920 27820
rect 17880 27577 17908 27814
rect 17866 27568 17922 27577
rect 17866 27503 17922 27512
rect 17610 27228 17918 27237
rect 17610 27226 17616 27228
rect 17672 27226 17696 27228
rect 17752 27226 17776 27228
rect 17832 27226 17856 27228
rect 17912 27226 17918 27228
rect 17672 27174 17674 27226
rect 17854 27174 17856 27226
rect 17610 27172 17616 27174
rect 17672 27172 17696 27174
rect 17752 27172 17776 27174
rect 17832 27172 17856 27174
rect 17912 27172 17918 27174
rect 17610 27163 17918 27172
rect 17610 26140 17918 26149
rect 17610 26138 17616 26140
rect 17672 26138 17696 26140
rect 17752 26138 17776 26140
rect 17832 26138 17856 26140
rect 17912 26138 17918 26140
rect 17672 26086 17674 26138
rect 17854 26086 17856 26138
rect 17610 26084 17616 26086
rect 17672 26084 17696 26086
rect 17752 26084 17776 26086
rect 17832 26084 17856 26086
rect 17912 26084 17918 26086
rect 17610 26075 17918 26084
rect 17500 26036 17552 26042
rect 17500 25978 17552 25984
rect 17408 9172 17460 9178
rect 17408 9114 17460 9120
rect 16950 8188 17258 8197
rect 16950 8186 16956 8188
rect 17012 8186 17036 8188
rect 17092 8186 17116 8188
rect 17172 8186 17196 8188
rect 17252 8186 17258 8188
rect 17012 8134 17014 8186
rect 17194 8134 17196 8186
rect 16950 8132 16956 8134
rect 17012 8132 17036 8134
rect 17092 8132 17116 8134
rect 17172 8132 17196 8134
rect 17252 8132 17258 8134
rect 16950 8123 17258 8132
rect 16950 7100 17258 7109
rect 16950 7098 16956 7100
rect 17012 7098 17036 7100
rect 17092 7098 17116 7100
rect 17172 7098 17196 7100
rect 17252 7098 17258 7100
rect 17012 7046 17014 7098
rect 17194 7046 17196 7098
rect 16950 7044 16956 7046
rect 17012 7044 17036 7046
rect 17092 7044 17116 7046
rect 17172 7044 17196 7046
rect 17252 7044 17258 7046
rect 16950 7035 17258 7044
rect 16950 6012 17258 6021
rect 16950 6010 16956 6012
rect 17012 6010 17036 6012
rect 17092 6010 17116 6012
rect 17172 6010 17196 6012
rect 17252 6010 17258 6012
rect 17012 5958 17014 6010
rect 17194 5958 17196 6010
rect 16950 5956 16956 5958
rect 17012 5956 17036 5958
rect 17092 5956 17116 5958
rect 17172 5956 17196 5958
rect 17252 5956 17258 5958
rect 16950 5947 17258 5956
rect 17512 5234 17540 25978
rect 17610 25052 17918 25061
rect 17610 25050 17616 25052
rect 17672 25050 17696 25052
rect 17752 25050 17776 25052
rect 17832 25050 17856 25052
rect 17912 25050 17918 25052
rect 17672 24998 17674 25050
rect 17854 24998 17856 25050
rect 17610 24996 17616 24998
rect 17672 24996 17696 24998
rect 17752 24996 17776 24998
rect 17832 24996 17856 24998
rect 17912 24996 17918 24998
rect 17610 24987 17918 24996
rect 17972 24818 18000 29650
rect 18156 27470 18184 44134
rect 18236 43104 18288 43110
rect 18236 43046 18288 43052
rect 18248 42809 18276 43046
rect 18234 42800 18290 42809
rect 18234 42735 18290 42744
rect 18234 42664 18290 42673
rect 18234 42599 18290 42608
rect 18248 41993 18276 42599
rect 18234 41984 18290 41993
rect 18234 41919 18290 41928
rect 18236 40928 18288 40934
rect 18234 40896 18236 40905
rect 18288 40896 18290 40905
rect 18234 40831 18290 40840
rect 18236 39296 18288 39302
rect 18236 39238 18288 39244
rect 18248 39001 18276 39238
rect 18234 38992 18290 39001
rect 18234 38927 18290 38936
rect 18340 38010 18368 44254
rect 18328 38004 18380 38010
rect 18328 37946 18380 37952
rect 18236 37120 18288 37126
rect 18234 37088 18236 37097
rect 18288 37088 18290 37097
rect 18234 37023 18290 37032
rect 18328 36576 18380 36582
rect 18328 36518 18380 36524
rect 18236 35488 18288 35494
rect 18236 35430 18288 35436
rect 18248 35193 18276 35430
rect 18234 35184 18290 35193
rect 18234 35119 18290 35128
rect 18236 33312 18288 33318
rect 18234 33280 18236 33289
rect 18288 33280 18290 33289
rect 18234 33215 18290 33224
rect 18236 31680 18288 31686
rect 18236 31622 18288 31628
rect 18248 31385 18276 31622
rect 18234 31376 18290 31385
rect 18234 31311 18290 31320
rect 18236 29504 18288 29510
rect 18234 29472 18236 29481
rect 18288 29472 18290 29481
rect 18234 29407 18290 29416
rect 18144 27464 18196 27470
rect 18144 27406 18196 27412
rect 18236 25696 18288 25702
rect 18234 25664 18236 25673
rect 18288 25664 18290 25673
rect 18234 25599 18290 25608
rect 17960 24812 18012 24818
rect 17960 24754 18012 24760
rect 18144 24744 18196 24750
rect 18144 24686 18196 24692
rect 17610 23964 17918 23973
rect 17610 23962 17616 23964
rect 17672 23962 17696 23964
rect 17752 23962 17776 23964
rect 17832 23962 17856 23964
rect 17912 23962 17918 23964
rect 17672 23910 17674 23962
rect 17854 23910 17856 23962
rect 17610 23908 17616 23910
rect 17672 23908 17696 23910
rect 17752 23908 17776 23910
rect 17832 23908 17856 23910
rect 17912 23908 17918 23910
rect 17610 23899 17918 23908
rect 18052 23316 18104 23322
rect 18052 23258 18104 23264
rect 17610 22876 17918 22885
rect 17610 22874 17616 22876
rect 17672 22874 17696 22876
rect 17752 22874 17776 22876
rect 17832 22874 17856 22876
rect 17912 22874 17918 22876
rect 17672 22822 17674 22874
rect 17854 22822 17856 22874
rect 17610 22820 17616 22822
rect 17672 22820 17696 22822
rect 17752 22820 17776 22822
rect 17832 22820 17856 22822
rect 17912 22820 17918 22822
rect 17610 22811 17918 22820
rect 18064 22574 18092 23258
rect 18052 22568 18104 22574
rect 18052 22510 18104 22516
rect 18064 22030 18092 22510
rect 18052 22024 18104 22030
rect 18052 21966 18104 21972
rect 17610 21788 17918 21797
rect 17610 21786 17616 21788
rect 17672 21786 17696 21788
rect 17752 21786 17776 21788
rect 17832 21786 17856 21788
rect 17912 21786 17918 21788
rect 17672 21734 17674 21786
rect 17854 21734 17856 21786
rect 17610 21732 17616 21734
rect 17672 21732 17696 21734
rect 17752 21732 17776 21734
rect 17832 21732 17856 21734
rect 17912 21732 17918 21734
rect 17610 21723 17918 21732
rect 17610 20700 17918 20709
rect 17610 20698 17616 20700
rect 17672 20698 17696 20700
rect 17752 20698 17776 20700
rect 17832 20698 17856 20700
rect 17912 20698 17918 20700
rect 17672 20646 17674 20698
rect 17854 20646 17856 20698
rect 17610 20644 17616 20646
rect 17672 20644 17696 20646
rect 17752 20644 17776 20646
rect 17832 20644 17856 20646
rect 17912 20644 17918 20646
rect 17610 20635 17918 20644
rect 18156 20398 18184 24686
rect 18236 24064 18288 24070
rect 18236 24006 18288 24012
rect 18248 23769 18276 24006
rect 18234 23760 18290 23769
rect 18234 23695 18290 23704
rect 18236 21888 18288 21894
rect 18234 21856 18236 21865
rect 18288 21856 18290 21865
rect 18234 21791 18290 21800
rect 18144 20392 18196 20398
rect 18144 20334 18196 20340
rect 18236 19984 18288 19990
rect 18234 19952 18236 19961
rect 18288 19952 18290 19961
rect 18234 19887 18290 19896
rect 17610 19612 17918 19621
rect 17610 19610 17616 19612
rect 17672 19610 17696 19612
rect 17752 19610 17776 19612
rect 17832 19610 17856 19612
rect 17912 19610 17918 19612
rect 17672 19558 17674 19610
rect 17854 19558 17856 19610
rect 17610 19556 17616 19558
rect 17672 19556 17696 19558
rect 17752 19556 17776 19558
rect 17832 19556 17856 19558
rect 17912 19556 17918 19558
rect 17610 19547 17918 19556
rect 17610 18524 17918 18533
rect 17610 18522 17616 18524
rect 17672 18522 17696 18524
rect 17752 18522 17776 18524
rect 17832 18522 17856 18524
rect 17912 18522 17918 18524
rect 17672 18470 17674 18522
rect 17854 18470 17856 18522
rect 17610 18468 17616 18470
rect 17672 18468 17696 18470
rect 17752 18468 17776 18470
rect 17832 18468 17856 18470
rect 17912 18468 17918 18470
rect 17610 18459 17918 18468
rect 18340 18426 18368 36518
rect 18432 32434 18460 64874
rect 18512 63980 18564 63986
rect 18512 63922 18564 63928
rect 18524 43450 18552 63922
rect 18604 62280 18656 62286
rect 18604 62222 18656 62228
rect 18512 43444 18564 43450
rect 18512 43386 18564 43392
rect 18512 43308 18564 43314
rect 18512 43250 18564 43256
rect 18420 32428 18472 32434
rect 18420 32370 18472 32376
rect 18420 32224 18472 32230
rect 18420 32166 18472 32172
rect 18432 23322 18460 32166
rect 18420 23316 18472 23322
rect 18420 23258 18472 23264
rect 18328 18420 18380 18426
rect 18328 18362 18380 18368
rect 18236 18080 18288 18086
rect 18234 18048 18236 18057
rect 18288 18048 18290 18057
rect 18234 17983 18290 17992
rect 17610 17436 17918 17445
rect 17610 17434 17616 17436
rect 17672 17434 17696 17436
rect 17752 17434 17776 17436
rect 17832 17434 17856 17436
rect 17912 17434 17918 17436
rect 17672 17382 17674 17434
rect 17854 17382 17856 17434
rect 17610 17380 17616 17382
rect 17672 17380 17696 17382
rect 17752 17380 17776 17382
rect 17832 17380 17856 17382
rect 17912 17380 17918 17382
rect 17610 17371 17918 17380
rect 17960 16788 18012 16794
rect 17960 16730 18012 16736
rect 17972 16697 18000 16730
rect 17958 16688 18014 16697
rect 17958 16623 18014 16632
rect 17610 16348 17918 16357
rect 17610 16346 17616 16348
rect 17672 16346 17696 16348
rect 17752 16346 17776 16348
rect 17832 16346 17856 16348
rect 17912 16346 17918 16348
rect 17672 16294 17674 16346
rect 17854 16294 17856 16346
rect 17610 16292 17616 16294
rect 17672 16292 17696 16294
rect 17752 16292 17776 16294
rect 17832 16292 17856 16294
rect 17912 16292 17918 16294
rect 17610 16283 17918 16292
rect 18236 16244 18288 16250
rect 18236 16186 18288 16192
rect 18248 16153 18276 16186
rect 18234 16144 18290 16153
rect 18234 16079 18290 16088
rect 18524 15366 18552 43250
rect 18616 42158 18644 62222
rect 18696 52012 18748 52018
rect 18696 51954 18748 51960
rect 18604 42152 18656 42158
rect 18604 42094 18656 42100
rect 18602 41984 18658 41993
rect 18602 41919 18658 41928
rect 18616 29646 18644 41919
rect 18708 35222 18736 51954
rect 18696 35216 18748 35222
rect 18696 35158 18748 35164
rect 18604 29640 18656 29646
rect 18604 29582 18656 29588
rect 18800 21350 18828 74598
rect 18972 71732 19024 71738
rect 18972 71674 19024 71680
rect 18880 59016 18932 59022
rect 18880 58958 18932 58964
rect 18892 30326 18920 58958
rect 18880 30320 18932 30326
rect 18880 30262 18932 30268
rect 18984 25906 19012 71674
rect 19156 65136 19208 65142
rect 19156 65078 19208 65084
rect 19064 62824 19116 62830
rect 19064 62766 19116 62772
rect 18972 25900 19024 25906
rect 18972 25842 19024 25848
rect 18788 21344 18840 21350
rect 18788 21286 18840 21292
rect 18236 15360 18288 15366
rect 18236 15302 18288 15308
rect 18512 15360 18564 15366
rect 18512 15302 18564 15308
rect 17610 15260 17918 15269
rect 17610 15258 17616 15260
rect 17672 15258 17696 15260
rect 17752 15258 17776 15260
rect 17832 15258 17856 15260
rect 17912 15258 17918 15260
rect 17672 15206 17674 15258
rect 17854 15206 17856 15258
rect 17610 15204 17616 15206
rect 17672 15204 17696 15206
rect 17752 15204 17776 15206
rect 17832 15204 17856 15206
rect 17912 15204 17918 15206
rect 17610 15195 17918 15204
rect 17682 14920 17738 14929
rect 17682 14855 17684 14864
rect 17736 14855 17738 14864
rect 17684 14826 17736 14832
rect 18248 14362 18276 15302
rect 18156 14334 18276 14362
rect 17610 14172 17918 14181
rect 17610 14170 17616 14172
rect 17672 14170 17696 14172
rect 17752 14170 17776 14172
rect 17832 14170 17856 14172
rect 17912 14170 17918 14172
rect 17672 14118 17674 14170
rect 17854 14118 17856 14170
rect 17610 14116 17616 14118
rect 17672 14116 17696 14118
rect 17752 14116 17776 14118
rect 17832 14116 17856 14118
rect 17912 14116 17918 14118
rect 17610 14107 17918 14116
rect 17610 13084 17918 13093
rect 17610 13082 17616 13084
rect 17672 13082 17696 13084
rect 17752 13082 17776 13084
rect 17832 13082 17856 13084
rect 17912 13082 17918 13084
rect 17672 13030 17674 13082
rect 17854 13030 17856 13082
rect 17610 13028 17616 13030
rect 17672 13028 17696 13030
rect 17752 13028 17776 13030
rect 17832 13028 17856 13030
rect 17912 13028 17918 13030
rect 17610 13019 17918 13028
rect 18052 12980 18104 12986
rect 18052 12922 18104 12928
rect 18064 12238 18092 12922
rect 18052 12232 18104 12238
rect 18052 12174 18104 12180
rect 17610 11996 17918 12005
rect 17610 11994 17616 11996
rect 17672 11994 17696 11996
rect 17752 11994 17776 11996
rect 17832 11994 17856 11996
rect 17912 11994 17918 11996
rect 17672 11942 17674 11994
rect 17854 11942 17856 11994
rect 17610 11940 17616 11942
rect 17672 11940 17696 11942
rect 17752 11940 17776 11942
rect 17832 11940 17856 11942
rect 17912 11940 17918 11942
rect 17610 11931 17918 11940
rect 17610 10908 17918 10917
rect 17610 10906 17616 10908
rect 17672 10906 17696 10908
rect 17752 10906 17776 10908
rect 17832 10906 17856 10908
rect 17912 10906 17918 10908
rect 17672 10854 17674 10906
rect 17854 10854 17856 10906
rect 17610 10852 17616 10854
rect 17672 10852 17696 10854
rect 17752 10852 17776 10854
rect 17832 10852 17856 10854
rect 17912 10852 17918 10854
rect 17610 10843 17918 10852
rect 17610 9820 17918 9829
rect 17610 9818 17616 9820
rect 17672 9818 17696 9820
rect 17752 9818 17776 9820
rect 17832 9818 17856 9820
rect 17912 9818 17918 9820
rect 17672 9766 17674 9818
rect 17854 9766 17856 9818
rect 17610 9764 17616 9766
rect 17672 9764 17696 9766
rect 17752 9764 17776 9766
rect 17832 9764 17856 9766
rect 17912 9764 17918 9766
rect 17610 9755 17918 9764
rect 18156 9450 18184 14334
rect 18236 14272 18288 14278
rect 18234 14240 18236 14249
rect 18288 14240 18290 14249
rect 18234 14175 18290 14184
rect 18236 12368 18288 12374
rect 18234 12336 18236 12345
rect 18288 12336 18290 12345
rect 18234 12271 18290 12280
rect 18236 10464 18288 10470
rect 18234 10432 18236 10441
rect 18288 10432 18290 10441
rect 18234 10367 18290 10376
rect 18144 9444 18196 9450
rect 18144 9386 18196 9392
rect 18236 8832 18288 8838
rect 18236 8774 18288 8780
rect 17610 8732 17918 8741
rect 17610 8730 17616 8732
rect 17672 8730 17696 8732
rect 17752 8730 17776 8732
rect 17832 8730 17856 8732
rect 17912 8730 17918 8732
rect 17672 8678 17674 8730
rect 17854 8678 17856 8730
rect 17610 8676 17616 8678
rect 17672 8676 17696 8678
rect 17752 8676 17776 8678
rect 17832 8676 17856 8678
rect 17912 8676 17918 8678
rect 17610 8667 17918 8676
rect 18052 8560 18104 8566
rect 18248 8537 18276 8774
rect 19076 8634 19104 62766
rect 19168 27606 19196 65078
rect 19340 65068 19392 65074
rect 19340 65010 19392 65016
rect 19248 60104 19300 60110
rect 19248 60046 19300 60052
rect 19260 51921 19288 60046
rect 19246 51912 19302 51921
rect 19246 51847 19302 51856
rect 19248 47456 19300 47462
rect 19248 47398 19300 47404
rect 19156 27600 19208 27606
rect 19156 27542 19208 27548
rect 19260 18290 19288 47398
rect 19352 29782 19380 65010
rect 19524 44872 19576 44878
rect 19524 44814 19576 44820
rect 19432 44124 19484 44130
rect 19432 44066 19484 44072
rect 19444 43722 19472 44066
rect 19432 43716 19484 43722
rect 19432 43658 19484 43664
rect 19444 36582 19472 43658
rect 19432 36576 19484 36582
rect 19432 36518 19484 36524
rect 19536 33114 19564 44814
rect 19800 41132 19852 41138
rect 19800 41074 19852 41080
rect 19616 38888 19668 38894
rect 19616 38830 19668 38836
rect 19524 33108 19576 33114
rect 19524 33050 19576 33056
rect 19524 30592 19576 30598
rect 19524 30534 19576 30540
rect 19340 29776 19392 29782
rect 19340 29718 19392 29724
rect 19248 18284 19300 18290
rect 19248 18226 19300 18232
rect 19536 14414 19564 30534
rect 19628 29714 19656 38830
rect 19708 35556 19760 35562
rect 19708 35498 19760 35504
rect 19616 29708 19668 29714
rect 19616 29650 19668 29656
rect 19524 14408 19576 14414
rect 19524 14350 19576 14356
rect 19064 8628 19116 8634
rect 19064 8570 19116 8576
rect 18052 8502 18104 8508
rect 18234 8528 18290 8537
rect 17610 7644 17918 7653
rect 17610 7642 17616 7644
rect 17672 7642 17696 7644
rect 17752 7642 17776 7644
rect 17832 7642 17856 7644
rect 17912 7642 17918 7644
rect 17672 7590 17674 7642
rect 17854 7590 17856 7642
rect 17610 7588 17616 7590
rect 17672 7588 17696 7590
rect 17752 7588 17776 7590
rect 17832 7588 17856 7590
rect 17912 7588 17918 7590
rect 17610 7579 17918 7588
rect 17610 6556 17918 6565
rect 17610 6554 17616 6556
rect 17672 6554 17696 6556
rect 17752 6554 17776 6556
rect 17832 6554 17856 6556
rect 17912 6554 17918 6556
rect 17672 6502 17674 6554
rect 17854 6502 17856 6554
rect 17610 6500 17616 6502
rect 17672 6500 17696 6502
rect 17752 6500 17776 6502
rect 17832 6500 17856 6502
rect 17912 6500 17918 6502
rect 17610 6491 17918 6500
rect 17610 5468 17918 5477
rect 17610 5466 17616 5468
rect 17672 5466 17696 5468
rect 17752 5466 17776 5468
rect 17832 5466 17856 5468
rect 17912 5466 17918 5468
rect 17672 5414 17674 5466
rect 17854 5414 17856 5466
rect 17610 5412 17616 5414
rect 17672 5412 17696 5414
rect 17752 5412 17776 5414
rect 17832 5412 17856 5414
rect 17912 5412 17918 5414
rect 17610 5403 17918 5412
rect 17500 5228 17552 5234
rect 17500 5170 17552 5176
rect 16950 4924 17258 4933
rect 16950 4922 16956 4924
rect 17012 4922 17036 4924
rect 17092 4922 17116 4924
rect 17172 4922 17196 4924
rect 17252 4922 17258 4924
rect 17012 4870 17014 4922
rect 17194 4870 17196 4922
rect 16950 4868 16956 4870
rect 17012 4868 17036 4870
rect 17092 4868 17116 4870
rect 17172 4868 17196 4870
rect 17252 4868 17258 4870
rect 16950 4859 17258 4868
rect 17610 4380 17918 4389
rect 17610 4378 17616 4380
rect 17672 4378 17696 4380
rect 17752 4378 17776 4380
rect 17832 4378 17856 4380
rect 17912 4378 17918 4380
rect 17672 4326 17674 4378
rect 17854 4326 17856 4378
rect 17610 4324 17616 4326
rect 17672 4324 17696 4326
rect 17752 4324 17776 4326
rect 17832 4324 17856 4326
rect 17912 4324 17918 4326
rect 17610 4315 17918 4324
rect 16672 4140 16724 4146
rect 16672 4082 16724 4088
rect 16950 3836 17258 3845
rect 16950 3834 16956 3836
rect 17012 3834 17036 3836
rect 17092 3834 17116 3836
rect 17172 3834 17196 3836
rect 17252 3834 17258 3836
rect 17012 3782 17014 3834
rect 17194 3782 17196 3834
rect 16950 3780 16956 3782
rect 17012 3780 17036 3782
rect 17092 3780 17116 3782
rect 17172 3780 17196 3782
rect 17252 3780 17258 3782
rect 16950 3771 17258 3780
rect 17610 3292 17918 3301
rect 17610 3290 17616 3292
rect 17672 3290 17696 3292
rect 17752 3290 17776 3292
rect 17832 3290 17856 3292
rect 17912 3290 17918 3292
rect 17672 3238 17674 3290
rect 17854 3238 17856 3290
rect 17610 3236 17616 3238
rect 17672 3236 17696 3238
rect 17752 3236 17776 3238
rect 17832 3236 17856 3238
rect 17912 3236 17918 3238
rect 17610 3227 17918 3236
rect 16950 2748 17258 2757
rect 16950 2746 16956 2748
rect 17012 2746 17036 2748
rect 17092 2746 17116 2748
rect 17172 2746 17196 2748
rect 17252 2746 17258 2748
rect 17012 2694 17014 2746
rect 17194 2694 17196 2746
rect 16950 2692 16956 2694
rect 17012 2692 17036 2694
rect 17092 2692 17116 2694
rect 17172 2692 17196 2694
rect 17252 2692 17258 2694
rect 16950 2683 17258 2692
rect 9864 2644 9916 2650
rect 9864 2586 9916 2592
rect 14464 2644 14516 2650
rect 14464 2586 14516 2592
rect 18064 2514 18092 8502
rect 18234 8463 18290 8472
rect 18236 6656 18288 6662
rect 18234 6624 18236 6633
rect 18288 6624 18290 6633
rect 18234 6559 18290 6568
rect 18236 5024 18288 5030
rect 18236 4966 18288 4972
rect 18248 4729 18276 4966
rect 18234 4720 18290 4729
rect 18234 4655 18290 4664
rect 19720 3058 19748 35498
rect 19812 15434 19840 41074
rect 19892 38276 19944 38282
rect 19892 38218 19944 38224
rect 19904 21690 19932 38218
rect 19892 21684 19944 21690
rect 19892 21626 19944 21632
rect 19800 15428 19852 15434
rect 19800 15370 19852 15376
rect 19708 3052 19760 3058
rect 19708 2994 19760 3000
rect 18236 2848 18288 2854
rect 18234 2816 18236 2825
rect 18288 2816 18290 2825
rect 18234 2751 18290 2760
rect 18052 2508 18104 2514
rect 18052 2450 18104 2456
rect 6000 2440 6052 2446
rect 6000 2382 6052 2388
rect 8852 2440 8904 2446
rect 8852 2382 8904 2388
rect 17868 2440 17920 2446
rect 17920 2388 18000 2394
rect 17868 2382 18000 2388
rect 2610 2204 2918 2213
rect 2610 2202 2616 2204
rect 2672 2202 2696 2204
rect 2752 2202 2776 2204
rect 2832 2202 2856 2204
rect 2912 2202 2918 2204
rect 2672 2150 2674 2202
rect 2854 2150 2856 2202
rect 2610 2148 2616 2150
rect 2672 2148 2696 2150
rect 2752 2148 2776 2150
rect 2832 2148 2856 2150
rect 2912 2148 2918 2150
rect 2610 2139 2918 2148
rect 6012 800 6040 2382
rect 13912 2372 13964 2378
rect 17880 2366 18000 2382
rect 13912 2314 13964 2320
rect 9956 2304 10008 2310
rect 9956 2246 10008 2252
rect 7610 2204 7918 2213
rect 7610 2202 7616 2204
rect 7672 2202 7696 2204
rect 7752 2202 7776 2204
rect 7832 2202 7856 2204
rect 7912 2202 7918 2204
rect 7672 2150 7674 2202
rect 7854 2150 7856 2202
rect 7610 2148 7616 2150
rect 7672 2148 7696 2150
rect 7752 2148 7776 2150
rect 7832 2148 7856 2150
rect 7912 2148 7918 2150
rect 7610 2139 7918 2148
rect 9968 800 9996 2246
rect 12610 2204 12918 2213
rect 12610 2202 12616 2204
rect 12672 2202 12696 2204
rect 12752 2202 12776 2204
rect 12832 2202 12856 2204
rect 12912 2202 12918 2204
rect 12672 2150 12674 2202
rect 12854 2150 12856 2202
rect 12610 2148 12616 2150
rect 12672 2148 12696 2150
rect 12752 2148 12776 2150
rect 12832 2148 12856 2150
rect 12912 2148 12918 2150
rect 12610 2139 12918 2148
rect 13924 800 13952 2314
rect 17610 2204 17918 2213
rect 17610 2202 17616 2204
rect 17672 2202 17696 2204
rect 17752 2202 17776 2204
rect 17832 2202 17856 2204
rect 17912 2202 17918 2204
rect 17672 2150 17674 2202
rect 17854 2150 17856 2202
rect 17610 2148 17616 2150
rect 17672 2148 17696 2150
rect 17752 2148 17776 2150
rect 17832 2148 17856 2150
rect 17912 2148 17918 2150
rect 17610 2139 17918 2148
rect 17972 1986 18000 2366
rect 17880 1958 18000 1986
rect 17880 800 17908 1958
rect 2148 734 2360 762
rect 5998 0 6054 800
rect 9954 0 10010 800
rect 13910 0 13966 800
rect 17866 0 17922 800
<< via2 >>
rect 1956 77818 2012 77820
rect 2036 77818 2092 77820
rect 2116 77818 2172 77820
rect 2196 77818 2252 77820
rect 1956 77766 2002 77818
rect 2002 77766 2012 77818
rect 2036 77766 2066 77818
rect 2066 77766 2078 77818
rect 2078 77766 2092 77818
rect 2116 77766 2130 77818
rect 2130 77766 2142 77818
rect 2142 77766 2172 77818
rect 2196 77766 2206 77818
rect 2206 77766 2252 77818
rect 1956 77764 2012 77766
rect 2036 77764 2092 77766
rect 2116 77764 2172 77766
rect 2196 77764 2252 77766
rect 6956 77818 7012 77820
rect 7036 77818 7092 77820
rect 7116 77818 7172 77820
rect 7196 77818 7252 77820
rect 6956 77766 7002 77818
rect 7002 77766 7012 77818
rect 7036 77766 7066 77818
rect 7066 77766 7078 77818
rect 7078 77766 7092 77818
rect 7116 77766 7130 77818
rect 7130 77766 7142 77818
rect 7142 77766 7172 77818
rect 7196 77766 7206 77818
rect 7206 77766 7252 77818
rect 6956 77764 7012 77766
rect 7036 77764 7092 77766
rect 7116 77764 7172 77766
rect 7196 77764 7252 77766
rect 11956 77818 12012 77820
rect 12036 77818 12092 77820
rect 12116 77818 12172 77820
rect 12196 77818 12252 77820
rect 11956 77766 12002 77818
rect 12002 77766 12012 77818
rect 12036 77766 12066 77818
rect 12066 77766 12078 77818
rect 12078 77766 12092 77818
rect 12116 77766 12130 77818
rect 12130 77766 12142 77818
rect 12142 77766 12172 77818
rect 12196 77766 12206 77818
rect 12206 77766 12252 77818
rect 11956 77764 12012 77766
rect 12036 77764 12092 77766
rect 12116 77764 12172 77766
rect 12196 77764 12252 77766
rect 16956 77818 17012 77820
rect 17036 77818 17092 77820
rect 17116 77818 17172 77820
rect 17196 77818 17252 77820
rect 16956 77766 17002 77818
rect 17002 77766 17012 77818
rect 17036 77766 17066 77818
rect 17066 77766 17078 77818
rect 17078 77766 17092 77818
rect 17116 77766 17130 77818
rect 17130 77766 17142 77818
rect 17142 77766 17172 77818
rect 17196 77766 17206 77818
rect 17206 77766 17252 77818
rect 16956 77764 17012 77766
rect 17036 77764 17092 77766
rect 17116 77764 17172 77766
rect 17196 77764 17252 77766
rect 2616 77274 2672 77276
rect 2696 77274 2752 77276
rect 2776 77274 2832 77276
rect 2856 77274 2912 77276
rect 2616 77222 2662 77274
rect 2662 77222 2672 77274
rect 2696 77222 2726 77274
rect 2726 77222 2738 77274
rect 2738 77222 2752 77274
rect 2776 77222 2790 77274
rect 2790 77222 2802 77274
rect 2802 77222 2832 77274
rect 2856 77222 2866 77274
rect 2866 77222 2912 77274
rect 2616 77220 2672 77222
rect 2696 77220 2752 77222
rect 2776 77220 2832 77222
rect 2856 77220 2912 77222
rect 7616 77274 7672 77276
rect 7696 77274 7752 77276
rect 7776 77274 7832 77276
rect 7856 77274 7912 77276
rect 7616 77222 7662 77274
rect 7662 77222 7672 77274
rect 7696 77222 7726 77274
rect 7726 77222 7738 77274
rect 7738 77222 7752 77274
rect 7776 77222 7790 77274
rect 7790 77222 7802 77274
rect 7802 77222 7832 77274
rect 7856 77222 7866 77274
rect 7866 77222 7912 77274
rect 7616 77220 7672 77222
rect 7696 77220 7752 77222
rect 7776 77220 7832 77222
rect 7856 77220 7912 77222
rect 12616 77274 12672 77276
rect 12696 77274 12752 77276
rect 12776 77274 12832 77276
rect 12856 77274 12912 77276
rect 12616 77222 12662 77274
rect 12662 77222 12672 77274
rect 12696 77222 12726 77274
rect 12726 77222 12738 77274
rect 12738 77222 12752 77274
rect 12776 77222 12790 77274
rect 12790 77222 12802 77274
rect 12802 77222 12832 77274
rect 12856 77222 12866 77274
rect 12866 77222 12912 77274
rect 12616 77220 12672 77222
rect 12696 77220 12752 77222
rect 12776 77220 12832 77222
rect 12856 77220 12912 77222
rect 14646 76780 14648 76800
rect 14648 76780 14700 76800
rect 14700 76780 14702 76800
rect 14646 76744 14702 76780
rect 1956 76730 2012 76732
rect 2036 76730 2092 76732
rect 2116 76730 2172 76732
rect 2196 76730 2252 76732
rect 1956 76678 2002 76730
rect 2002 76678 2012 76730
rect 2036 76678 2066 76730
rect 2066 76678 2078 76730
rect 2078 76678 2092 76730
rect 2116 76678 2130 76730
rect 2130 76678 2142 76730
rect 2142 76678 2172 76730
rect 2196 76678 2206 76730
rect 2206 76678 2252 76730
rect 1956 76676 2012 76678
rect 2036 76676 2092 76678
rect 2116 76676 2172 76678
rect 2196 76676 2252 76678
rect 6956 76730 7012 76732
rect 7036 76730 7092 76732
rect 7116 76730 7172 76732
rect 7196 76730 7252 76732
rect 6956 76678 7002 76730
rect 7002 76678 7012 76730
rect 7036 76678 7066 76730
rect 7066 76678 7078 76730
rect 7078 76678 7092 76730
rect 7116 76678 7130 76730
rect 7130 76678 7142 76730
rect 7142 76678 7172 76730
rect 7196 76678 7206 76730
rect 7206 76678 7252 76730
rect 6956 76676 7012 76678
rect 7036 76676 7092 76678
rect 7116 76676 7172 76678
rect 7196 76676 7252 76678
rect 15934 76780 15936 76800
rect 15936 76780 15988 76800
rect 15988 76780 15990 76800
rect 15934 76744 15990 76780
rect 11956 76730 12012 76732
rect 12036 76730 12092 76732
rect 12116 76730 12172 76732
rect 12196 76730 12252 76732
rect 11956 76678 12002 76730
rect 12002 76678 12012 76730
rect 12036 76678 12066 76730
rect 12066 76678 12078 76730
rect 12078 76678 12092 76730
rect 12116 76678 12130 76730
rect 12130 76678 12142 76730
rect 12142 76678 12172 76730
rect 12196 76678 12206 76730
rect 12206 76678 12252 76730
rect 11956 76676 12012 76678
rect 12036 76676 12092 76678
rect 12116 76676 12172 76678
rect 12196 76676 12252 76678
rect 2616 76186 2672 76188
rect 2696 76186 2752 76188
rect 2776 76186 2832 76188
rect 2856 76186 2912 76188
rect 2616 76134 2662 76186
rect 2662 76134 2672 76186
rect 2696 76134 2726 76186
rect 2726 76134 2738 76186
rect 2738 76134 2752 76186
rect 2776 76134 2790 76186
rect 2790 76134 2802 76186
rect 2802 76134 2832 76186
rect 2856 76134 2866 76186
rect 2866 76134 2912 76186
rect 2616 76132 2672 76134
rect 2696 76132 2752 76134
rect 2776 76132 2832 76134
rect 2856 76132 2912 76134
rect 1956 75642 2012 75644
rect 2036 75642 2092 75644
rect 2116 75642 2172 75644
rect 2196 75642 2252 75644
rect 1956 75590 2002 75642
rect 2002 75590 2012 75642
rect 2036 75590 2066 75642
rect 2066 75590 2078 75642
rect 2078 75590 2092 75642
rect 2116 75590 2130 75642
rect 2130 75590 2142 75642
rect 2142 75590 2172 75642
rect 2196 75590 2206 75642
rect 2206 75590 2252 75642
rect 1956 75588 2012 75590
rect 2036 75588 2092 75590
rect 2116 75588 2172 75590
rect 2196 75588 2252 75590
rect 2616 75098 2672 75100
rect 2696 75098 2752 75100
rect 2776 75098 2832 75100
rect 2856 75098 2912 75100
rect 2616 75046 2662 75098
rect 2662 75046 2672 75098
rect 2696 75046 2726 75098
rect 2726 75046 2738 75098
rect 2738 75046 2752 75098
rect 2776 75046 2790 75098
rect 2790 75046 2802 75098
rect 2802 75046 2832 75098
rect 2856 75046 2866 75098
rect 2866 75046 2912 75098
rect 2616 75044 2672 75046
rect 2696 75044 2752 75046
rect 2776 75044 2832 75046
rect 2856 75044 2912 75046
rect 1956 74554 2012 74556
rect 2036 74554 2092 74556
rect 2116 74554 2172 74556
rect 2196 74554 2252 74556
rect 1956 74502 2002 74554
rect 2002 74502 2012 74554
rect 2036 74502 2066 74554
rect 2066 74502 2078 74554
rect 2078 74502 2092 74554
rect 2116 74502 2130 74554
rect 2130 74502 2142 74554
rect 2142 74502 2172 74554
rect 2196 74502 2206 74554
rect 2206 74502 2252 74554
rect 1956 74500 2012 74502
rect 2036 74500 2092 74502
rect 2116 74500 2172 74502
rect 2196 74500 2252 74502
rect 2616 74010 2672 74012
rect 2696 74010 2752 74012
rect 2776 74010 2832 74012
rect 2856 74010 2912 74012
rect 2616 73958 2662 74010
rect 2662 73958 2672 74010
rect 2696 73958 2726 74010
rect 2726 73958 2738 74010
rect 2738 73958 2752 74010
rect 2776 73958 2790 74010
rect 2790 73958 2802 74010
rect 2802 73958 2832 74010
rect 2856 73958 2866 74010
rect 2866 73958 2912 74010
rect 2616 73956 2672 73958
rect 2696 73956 2752 73958
rect 2776 73956 2832 73958
rect 2856 73956 2912 73958
rect 1956 73466 2012 73468
rect 2036 73466 2092 73468
rect 2116 73466 2172 73468
rect 2196 73466 2252 73468
rect 1956 73414 2002 73466
rect 2002 73414 2012 73466
rect 2036 73414 2066 73466
rect 2066 73414 2078 73466
rect 2078 73414 2092 73466
rect 2116 73414 2130 73466
rect 2130 73414 2142 73466
rect 2142 73414 2172 73466
rect 2196 73414 2206 73466
rect 2206 73414 2252 73466
rect 1956 73412 2012 73414
rect 2036 73412 2092 73414
rect 2116 73412 2172 73414
rect 2196 73412 2252 73414
rect 2616 72922 2672 72924
rect 2696 72922 2752 72924
rect 2776 72922 2832 72924
rect 2856 72922 2912 72924
rect 2616 72870 2662 72922
rect 2662 72870 2672 72922
rect 2696 72870 2726 72922
rect 2726 72870 2738 72922
rect 2738 72870 2752 72922
rect 2776 72870 2790 72922
rect 2790 72870 2802 72922
rect 2802 72870 2832 72922
rect 2856 72870 2866 72922
rect 2866 72870 2912 72922
rect 2616 72868 2672 72870
rect 2696 72868 2752 72870
rect 2776 72868 2832 72870
rect 2856 72868 2912 72870
rect 1956 72378 2012 72380
rect 2036 72378 2092 72380
rect 2116 72378 2172 72380
rect 2196 72378 2252 72380
rect 1956 72326 2002 72378
rect 2002 72326 2012 72378
rect 2036 72326 2066 72378
rect 2066 72326 2078 72378
rect 2078 72326 2092 72378
rect 2116 72326 2130 72378
rect 2130 72326 2142 72378
rect 2142 72326 2172 72378
rect 2196 72326 2206 72378
rect 2206 72326 2252 72378
rect 1956 72324 2012 72326
rect 2036 72324 2092 72326
rect 2116 72324 2172 72326
rect 2196 72324 2252 72326
rect 2616 71834 2672 71836
rect 2696 71834 2752 71836
rect 2776 71834 2832 71836
rect 2856 71834 2912 71836
rect 2616 71782 2662 71834
rect 2662 71782 2672 71834
rect 2696 71782 2726 71834
rect 2726 71782 2738 71834
rect 2738 71782 2752 71834
rect 2776 71782 2790 71834
rect 2790 71782 2802 71834
rect 2802 71782 2832 71834
rect 2856 71782 2866 71834
rect 2866 71782 2912 71834
rect 2616 71780 2672 71782
rect 2696 71780 2752 71782
rect 2776 71780 2832 71782
rect 2856 71780 2912 71782
rect 1956 71290 2012 71292
rect 2036 71290 2092 71292
rect 2116 71290 2172 71292
rect 2196 71290 2252 71292
rect 1956 71238 2002 71290
rect 2002 71238 2012 71290
rect 2036 71238 2066 71290
rect 2066 71238 2078 71290
rect 2078 71238 2092 71290
rect 2116 71238 2130 71290
rect 2130 71238 2142 71290
rect 2142 71238 2172 71290
rect 2196 71238 2206 71290
rect 2206 71238 2252 71290
rect 1956 71236 2012 71238
rect 2036 71236 2092 71238
rect 2116 71236 2172 71238
rect 2196 71236 2252 71238
rect 2616 70746 2672 70748
rect 2696 70746 2752 70748
rect 2776 70746 2832 70748
rect 2856 70746 2912 70748
rect 2616 70694 2662 70746
rect 2662 70694 2672 70746
rect 2696 70694 2726 70746
rect 2726 70694 2738 70746
rect 2738 70694 2752 70746
rect 2776 70694 2790 70746
rect 2790 70694 2802 70746
rect 2802 70694 2832 70746
rect 2856 70694 2866 70746
rect 2866 70694 2912 70746
rect 2616 70692 2672 70694
rect 2696 70692 2752 70694
rect 2776 70692 2832 70694
rect 2856 70692 2912 70694
rect 1956 70202 2012 70204
rect 2036 70202 2092 70204
rect 2116 70202 2172 70204
rect 2196 70202 2252 70204
rect 1956 70150 2002 70202
rect 2002 70150 2012 70202
rect 2036 70150 2066 70202
rect 2066 70150 2078 70202
rect 2078 70150 2092 70202
rect 2116 70150 2130 70202
rect 2130 70150 2142 70202
rect 2142 70150 2172 70202
rect 2196 70150 2206 70202
rect 2206 70150 2252 70202
rect 1956 70148 2012 70150
rect 2036 70148 2092 70150
rect 2116 70148 2172 70150
rect 2196 70148 2252 70150
rect 3330 70896 3386 70952
rect 2042 69264 2098 69320
rect 1956 69114 2012 69116
rect 2036 69114 2092 69116
rect 2116 69114 2172 69116
rect 2196 69114 2252 69116
rect 1956 69062 2002 69114
rect 2002 69062 2012 69114
rect 2036 69062 2066 69114
rect 2066 69062 2078 69114
rect 2078 69062 2092 69114
rect 2116 69062 2130 69114
rect 2130 69062 2142 69114
rect 2142 69062 2172 69114
rect 2196 69062 2206 69114
rect 2206 69062 2252 69114
rect 1956 69060 2012 69062
rect 2036 69060 2092 69062
rect 2116 69060 2172 69062
rect 2196 69060 2252 69062
rect 1956 68026 2012 68028
rect 2036 68026 2092 68028
rect 2116 68026 2172 68028
rect 2196 68026 2252 68028
rect 1956 67974 2002 68026
rect 2002 67974 2012 68026
rect 2036 67974 2066 68026
rect 2066 67974 2078 68026
rect 2078 67974 2092 68026
rect 2116 67974 2130 68026
rect 2130 67974 2142 68026
rect 2142 67974 2172 68026
rect 2196 67974 2206 68026
rect 2206 67974 2252 68026
rect 1956 67972 2012 67974
rect 2036 67972 2092 67974
rect 2116 67972 2172 67974
rect 2196 67972 2252 67974
rect 1956 66938 2012 66940
rect 2036 66938 2092 66940
rect 2116 66938 2172 66940
rect 2196 66938 2252 66940
rect 1956 66886 2002 66938
rect 2002 66886 2012 66938
rect 2036 66886 2066 66938
rect 2066 66886 2078 66938
rect 2078 66886 2092 66938
rect 2116 66886 2130 66938
rect 2130 66886 2142 66938
rect 2142 66886 2172 66938
rect 2196 66886 2206 66938
rect 2206 66886 2252 66938
rect 1956 66884 2012 66886
rect 2036 66884 2092 66886
rect 2116 66884 2172 66886
rect 2196 66884 2252 66886
rect 1956 65850 2012 65852
rect 2036 65850 2092 65852
rect 2116 65850 2172 65852
rect 2196 65850 2252 65852
rect 1956 65798 2002 65850
rect 2002 65798 2012 65850
rect 2036 65798 2066 65850
rect 2066 65798 2078 65850
rect 2078 65798 2092 65850
rect 2116 65798 2130 65850
rect 2130 65798 2142 65850
rect 2142 65798 2172 65850
rect 2196 65798 2206 65850
rect 2206 65798 2252 65850
rect 1956 65796 2012 65798
rect 2036 65796 2092 65798
rect 2116 65796 2172 65798
rect 2196 65796 2252 65798
rect 1956 64762 2012 64764
rect 2036 64762 2092 64764
rect 2116 64762 2172 64764
rect 2196 64762 2252 64764
rect 1956 64710 2002 64762
rect 2002 64710 2012 64762
rect 2036 64710 2066 64762
rect 2066 64710 2078 64762
rect 2078 64710 2092 64762
rect 2116 64710 2130 64762
rect 2130 64710 2142 64762
rect 2142 64710 2172 64762
rect 2196 64710 2206 64762
rect 2206 64710 2252 64762
rect 1956 64708 2012 64710
rect 2036 64708 2092 64710
rect 2116 64708 2172 64710
rect 2196 64708 2252 64710
rect 1674 55664 1730 55720
rect 1956 63674 2012 63676
rect 2036 63674 2092 63676
rect 2116 63674 2172 63676
rect 2196 63674 2252 63676
rect 1956 63622 2002 63674
rect 2002 63622 2012 63674
rect 2036 63622 2066 63674
rect 2066 63622 2078 63674
rect 2078 63622 2092 63674
rect 2116 63622 2130 63674
rect 2130 63622 2142 63674
rect 2142 63622 2172 63674
rect 2196 63622 2206 63674
rect 2206 63622 2252 63674
rect 1956 63620 2012 63622
rect 2036 63620 2092 63622
rect 2116 63620 2172 63622
rect 2196 63620 2252 63622
rect 1956 62586 2012 62588
rect 2036 62586 2092 62588
rect 2116 62586 2172 62588
rect 2196 62586 2252 62588
rect 1956 62534 2002 62586
rect 2002 62534 2012 62586
rect 2036 62534 2066 62586
rect 2066 62534 2078 62586
rect 2078 62534 2092 62586
rect 2116 62534 2130 62586
rect 2130 62534 2142 62586
rect 2142 62534 2172 62586
rect 2196 62534 2206 62586
rect 2206 62534 2252 62586
rect 1956 62532 2012 62534
rect 2036 62532 2092 62534
rect 2116 62532 2172 62534
rect 2196 62532 2252 62534
rect 1956 61498 2012 61500
rect 2036 61498 2092 61500
rect 2116 61498 2172 61500
rect 2196 61498 2252 61500
rect 1956 61446 2002 61498
rect 2002 61446 2012 61498
rect 2036 61446 2066 61498
rect 2066 61446 2078 61498
rect 2078 61446 2092 61498
rect 2116 61446 2130 61498
rect 2130 61446 2142 61498
rect 2142 61446 2172 61498
rect 2196 61446 2206 61498
rect 2206 61446 2252 61498
rect 1956 61444 2012 61446
rect 2036 61444 2092 61446
rect 2116 61444 2172 61446
rect 2196 61444 2252 61446
rect 1956 60410 2012 60412
rect 2036 60410 2092 60412
rect 2116 60410 2172 60412
rect 2196 60410 2252 60412
rect 1956 60358 2002 60410
rect 2002 60358 2012 60410
rect 2036 60358 2066 60410
rect 2066 60358 2078 60410
rect 2078 60358 2092 60410
rect 2116 60358 2130 60410
rect 2130 60358 2142 60410
rect 2142 60358 2172 60410
rect 2196 60358 2206 60410
rect 2206 60358 2252 60410
rect 1956 60356 2012 60358
rect 2036 60356 2092 60358
rect 2116 60356 2172 60358
rect 2196 60356 2252 60358
rect 1956 59322 2012 59324
rect 2036 59322 2092 59324
rect 2116 59322 2172 59324
rect 2196 59322 2252 59324
rect 1956 59270 2002 59322
rect 2002 59270 2012 59322
rect 2036 59270 2066 59322
rect 2066 59270 2078 59322
rect 2078 59270 2092 59322
rect 2116 59270 2130 59322
rect 2130 59270 2142 59322
rect 2142 59270 2172 59322
rect 2196 59270 2206 59322
rect 2206 59270 2252 59322
rect 1956 59268 2012 59270
rect 2036 59268 2092 59270
rect 2116 59268 2172 59270
rect 2196 59268 2252 59270
rect 1956 58234 2012 58236
rect 2036 58234 2092 58236
rect 2116 58234 2172 58236
rect 2196 58234 2252 58236
rect 1956 58182 2002 58234
rect 2002 58182 2012 58234
rect 2036 58182 2066 58234
rect 2066 58182 2078 58234
rect 2078 58182 2092 58234
rect 2116 58182 2130 58234
rect 2130 58182 2142 58234
rect 2142 58182 2172 58234
rect 2196 58182 2206 58234
rect 2206 58182 2252 58234
rect 1956 58180 2012 58182
rect 2036 58180 2092 58182
rect 2116 58180 2172 58182
rect 2196 58180 2252 58182
rect 1956 57146 2012 57148
rect 2036 57146 2092 57148
rect 2116 57146 2172 57148
rect 2196 57146 2252 57148
rect 1956 57094 2002 57146
rect 2002 57094 2012 57146
rect 2036 57094 2066 57146
rect 2066 57094 2078 57146
rect 2078 57094 2092 57146
rect 2116 57094 2130 57146
rect 2130 57094 2142 57146
rect 2142 57094 2172 57146
rect 2196 57094 2206 57146
rect 2206 57094 2252 57146
rect 1956 57092 2012 57094
rect 2036 57092 2092 57094
rect 2116 57092 2172 57094
rect 2196 57092 2252 57094
rect 1956 56058 2012 56060
rect 2036 56058 2092 56060
rect 2116 56058 2172 56060
rect 2196 56058 2252 56060
rect 1956 56006 2002 56058
rect 2002 56006 2012 56058
rect 2036 56006 2066 56058
rect 2066 56006 2078 56058
rect 2078 56006 2092 56058
rect 2116 56006 2130 56058
rect 2130 56006 2142 56058
rect 2142 56006 2172 56058
rect 2196 56006 2206 56058
rect 2206 56006 2252 56058
rect 1956 56004 2012 56006
rect 2036 56004 2092 56006
rect 2116 56004 2172 56006
rect 2196 56004 2252 56006
rect 1956 54970 2012 54972
rect 2036 54970 2092 54972
rect 2116 54970 2172 54972
rect 2196 54970 2252 54972
rect 1956 54918 2002 54970
rect 2002 54918 2012 54970
rect 2036 54918 2066 54970
rect 2066 54918 2078 54970
rect 2078 54918 2092 54970
rect 2116 54918 2130 54970
rect 2130 54918 2142 54970
rect 2142 54918 2172 54970
rect 2196 54918 2206 54970
rect 2206 54918 2252 54970
rect 1956 54916 2012 54918
rect 2036 54916 2092 54918
rect 2116 54916 2172 54918
rect 2196 54916 2252 54918
rect 1956 53882 2012 53884
rect 2036 53882 2092 53884
rect 2116 53882 2172 53884
rect 2196 53882 2252 53884
rect 1956 53830 2002 53882
rect 2002 53830 2012 53882
rect 2036 53830 2066 53882
rect 2066 53830 2078 53882
rect 2078 53830 2092 53882
rect 2116 53830 2130 53882
rect 2130 53830 2142 53882
rect 2142 53830 2172 53882
rect 2196 53830 2206 53882
rect 2206 53830 2252 53882
rect 1956 53828 2012 53830
rect 2036 53828 2092 53830
rect 2116 53828 2172 53830
rect 2196 53828 2252 53830
rect 1582 40568 1638 40624
rect 1956 52794 2012 52796
rect 2036 52794 2092 52796
rect 2116 52794 2172 52796
rect 2196 52794 2252 52796
rect 1956 52742 2002 52794
rect 2002 52742 2012 52794
rect 2036 52742 2066 52794
rect 2066 52742 2078 52794
rect 2078 52742 2092 52794
rect 2116 52742 2130 52794
rect 2130 52742 2142 52794
rect 2142 52742 2172 52794
rect 2196 52742 2206 52794
rect 2206 52742 2252 52794
rect 1956 52740 2012 52742
rect 2036 52740 2092 52742
rect 2116 52740 2172 52742
rect 2196 52740 2252 52742
rect 1956 51706 2012 51708
rect 2036 51706 2092 51708
rect 2116 51706 2172 51708
rect 2196 51706 2252 51708
rect 1956 51654 2002 51706
rect 2002 51654 2012 51706
rect 2036 51654 2066 51706
rect 2066 51654 2078 51706
rect 2078 51654 2092 51706
rect 2116 51654 2130 51706
rect 2130 51654 2142 51706
rect 2142 51654 2172 51706
rect 2196 51654 2206 51706
rect 2206 51654 2252 51706
rect 1956 51652 2012 51654
rect 2036 51652 2092 51654
rect 2116 51652 2172 51654
rect 2196 51652 2252 51654
rect 1956 50618 2012 50620
rect 2036 50618 2092 50620
rect 2116 50618 2172 50620
rect 2196 50618 2252 50620
rect 1956 50566 2002 50618
rect 2002 50566 2012 50618
rect 2036 50566 2066 50618
rect 2066 50566 2078 50618
rect 2078 50566 2092 50618
rect 2116 50566 2130 50618
rect 2130 50566 2142 50618
rect 2142 50566 2172 50618
rect 2196 50566 2206 50618
rect 2206 50566 2252 50618
rect 1956 50564 2012 50566
rect 2036 50564 2092 50566
rect 2116 50564 2172 50566
rect 2196 50564 2252 50566
rect 1766 40840 1822 40896
rect 1956 49530 2012 49532
rect 2036 49530 2092 49532
rect 2116 49530 2172 49532
rect 2196 49530 2252 49532
rect 1956 49478 2002 49530
rect 2002 49478 2012 49530
rect 2036 49478 2066 49530
rect 2066 49478 2078 49530
rect 2078 49478 2092 49530
rect 2116 49478 2130 49530
rect 2130 49478 2142 49530
rect 2142 49478 2172 49530
rect 2196 49478 2206 49530
rect 2206 49478 2252 49530
rect 1956 49476 2012 49478
rect 2036 49476 2092 49478
rect 2116 49476 2172 49478
rect 2196 49476 2252 49478
rect 1956 48442 2012 48444
rect 2036 48442 2092 48444
rect 2116 48442 2172 48444
rect 2196 48442 2252 48444
rect 1956 48390 2002 48442
rect 2002 48390 2012 48442
rect 2036 48390 2066 48442
rect 2066 48390 2078 48442
rect 2078 48390 2092 48442
rect 2116 48390 2130 48442
rect 2130 48390 2142 48442
rect 2142 48390 2172 48442
rect 2196 48390 2206 48442
rect 2206 48390 2252 48442
rect 1956 48388 2012 48390
rect 2036 48388 2092 48390
rect 2116 48388 2172 48390
rect 2196 48388 2252 48390
rect 1956 47354 2012 47356
rect 2036 47354 2092 47356
rect 2116 47354 2172 47356
rect 2196 47354 2252 47356
rect 1956 47302 2002 47354
rect 2002 47302 2012 47354
rect 2036 47302 2066 47354
rect 2066 47302 2078 47354
rect 2078 47302 2092 47354
rect 2116 47302 2130 47354
rect 2130 47302 2142 47354
rect 2142 47302 2172 47354
rect 2196 47302 2206 47354
rect 2206 47302 2252 47354
rect 1956 47300 2012 47302
rect 2036 47300 2092 47302
rect 2116 47300 2172 47302
rect 2196 47300 2252 47302
rect 1956 46266 2012 46268
rect 2036 46266 2092 46268
rect 2116 46266 2172 46268
rect 2196 46266 2252 46268
rect 1956 46214 2002 46266
rect 2002 46214 2012 46266
rect 2036 46214 2066 46266
rect 2066 46214 2078 46266
rect 2078 46214 2092 46266
rect 2116 46214 2130 46266
rect 2130 46214 2142 46266
rect 2142 46214 2172 46266
rect 2196 46214 2206 46266
rect 2206 46214 2252 46266
rect 1956 46212 2012 46214
rect 2036 46212 2092 46214
rect 2116 46212 2172 46214
rect 2196 46212 2252 46214
rect 1956 45178 2012 45180
rect 2036 45178 2092 45180
rect 2116 45178 2172 45180
rect 2196 45178 2252 45180
rect 1956 45126 2002 45178
rect 2002 45126 2012 45178
rect 2036 45126 2066 45178
rect 2066 45126 2078 45178
rect 2078 45126 2092 45178
rect 2116 45126 2130 45178
rect 2130 45126 2142 45178
rect 2142 45126 2172 45178
rect 2196 45126 2206 45178
rect 2206 45126 2252 45178
rect 1956 45124 2012 45126
rect 2036 45124 2092 45126
rect 2116 45124 2172 45126
rect 2196 45124 2252 45126
rect 2616 69658 2672 69660
rect 2696 69658 2752 69660
rect 2776 69658 2832 69660
rect 2856 69658 2912 69660
rect 2616 69606 2662 69658
rect 2662 69606 2672 69658
rect 2696 69606 2726 69658
rect 2726 69606 2738 69658
rect 2738 69606 2752 69658
rect 2776 69606 2790 69658
rect 2790 69606 2802 69658
rect 2802 69606 2832 69658
rect 2856 69606 2866 69658
rect 2866 69606 2912 69658
rect 2616 69604 2672 69606
rect 2696 69604 2752 69606
rect 2776 69604 2832 69606
rect 2856 69604 2912 69606
rect 2616 68570 2672 68572
rect 2696 68570 2752 68572
rect 2776 68570 2832 68572
rect 2856 68570 2912 68572
rect 2616 68518 2662 68570
rect 2662 68518 2672 68570
rect 2696 68518 2726 68570
rect 2726 68518 2738 68570
rect 2738 68518 2752 68570
rect 2776 68518 2790 68570
rect 2790 68518 2802 68570
rect 2802 68518 2832 68570
rect 2856 68518 2866 68570
rect 2866 68518 2912 68570
rect 2616 68516 2672 68518
rect 2696 68516 2752 68518
rect 2776 68516 2832 68518
rect 2856 68516 2912 68518
rect 2616 67482 2672 67484
rect 2696 67482 2752 67484
rect 2776 67482 2832 67484
rect 2856 67482 2912 67484
rect 2616 67430 2662 67482
rect 2662 67430 2672 67482
rect 2696 67430 2726 67482
rect 2726 67430 2738 67482
rect 2738 67430 2752 67482
rect 2776 67430 2790 67482
rect 2790 67430 2802 67482
rect 2802 67430 2832 67482
rect 2856 67430 2866 67482
rect 2866 67430 2912 67482
rect 2616 67428 2672 67430
rect 2696 67428 2752 67430
rect 2776 67428 2832 67430
rect 2856 67428 2912 67430
rect 2616 66394 2672 66396
rect 2696 66394 2752 66396
rect 2776 66394 2832 66396
rect 2856 66394 2912 66396
rect 2616 66342 2662 66394
rect 2662 66342 2672 66394
rect 2696 66342 2726 66394
rect 2726 66342 2738 66394
rect 2738 66342 2752 66394
rect 2776 66342 2790 66394
rect 2790 66342 2802 66394
rect 2802 66342 2832 66394
rect 2856 66342 2866 66394
rect 2866 66342 2912 66394
rect 2616 66340 2672 66342
rect 2696 66340 2752 66342
rect 2776 66340 2832 66342
rect 2856 66340 2912 66342
rect 2616 65306 2672 65308
rect 2696 65306 2752 65308
rect 2776 65306 2832 65308
rect 2856 65306 2912 65308
rect 2616 65254 2662 65306
rect 2662 65254 2672 65306
rect 2696 65254 2726 65306
rect 2726 65254 2738 65306
rect 2738 65254 2752 65306
rect 2776 65254 2790 65306
rect 2790 65254 2802 65306
rect 2802 65254 2832 65306
rect 2856 65254 2866 65306
rect 2866 65254 2912 65306
rect 2616 65252 2672 65254
rect 2696 65252 2752 65254
rect 2776 65252 2832 65254
rect 2856 65252 2912 65254
rect 2616 64218 2672 64220
rect 2696 64218 2752 64220
rect 2776 64218 2832 64220
rect 2856 64218 2912 64220
rect 2616 64166 2662 64218
rect 2662 64166 2672 64218
rect 2696 64166 2726 64218
rect 2726 64166 2738 64218
rect 2738 64166 2752 64218
rect 2776 64166 2790 64218
rect 2790 64166 2802 64218
rect 2802 64166 2832 64218
rect 2856 64166 2866 64218
rect 2866 64166 2912 64218
rect 2616 64164 2672 64166
rect 2696 64164 2752 64166
rect 2776 64164 2832 64166
rect 2856 64164 2912 64166
rect 2616 63130 2672 63132
rect 2696 63130 2752 63132
rect 2776 63130 2832 63132
rect 2856 63130 2912 63132
rect 2616 63078 2662 63130
rect 2662 63078 2672 63130
rect 2696 63078 2726 63130
rect 2726 63078 2738 63130
rect 2738 63078 2752 63130
rect 2776 63078 2790 63130
rect 2790 63078 2802 63130
rect 2802 63078 2832 63130
rect 2856 63078 2866 63130
rect 2866 63078 2912 63130
rect 2616 63076 2672 63078
rect 2696 63076 2752 63078
rect 2776 63076 2832 63078
rect 2856 63076 2912 63078
rect 2616 62042 2672 62044
rect 2696 62042 2752 62044
rect 2776 62042 2832 62044
rect 2856 62042 2912 62044
rect 2616 61990 2662 62042
rect 2662 61990 2672 62042
rect 2696 61990 2726 62042
rect 2726 61990 2738 62042
rect 2738 61990 2752 62042
rect 2776 61990 2790 62042
rect 2790 61990 2802 62042
rect 2802 61990 2832 62042
rect 2856 61990 2866 62042
rect 2866 61990 2912 62042
rect 2616 61988 2672 61990
rect 2696 61988 2752 61990
rect 2776 61988 2832 61990
rect 2856 61988 2912 61990
rect 2616 60954 2672 60956
rect 2696 60954 2752 60956
rect 2776 60954 2832 60956
rect 2856 60954 2912 60956
rect 2616 60902 2662 60954
rect 2662 60902 2672 60954
rect 2696 60902 2726 60954
rect 2726 60902 2738 60954
rect 2738 60902 2752 60954
rect 2776 60902 2790 60954
rect 2790 60902 2802 60954
rect 2802 60902 2832 60954
rect 2856 60902 2866 60954
rect 2866 60902 2912 60954
rect 2616 60900 2672 60902
rect 2696 60900 2752 60902
rect 2776 60900 2832 60902
rect 2856 60900 2912 60902
rect 2616 59866 2672 59868
rect 2696 59866 2752 59868
rect 2776 59866 2832 59868
rect 2856 59866 2912 59868
rect 2616 59814 2662 59866
rect 2662 59814 2672 59866
rect 2696 59814 2726 59866
rect 2726 59814 2738 59866
rect 2738 59814 2752 59866
rect 2776 59814 2790 59866
rect 2790 59814 2802 59866
rect 2802 59814 2832 59866
rect 2856 59814 2866 59866
rect 2866 59814 2912 59866
rect 2616 59812 2672 59814
rect 2696 59812 2752 59814
rect 2776 59812 2832 59814
rect 2856 59812 2912 59814
rect 2616 58778 2672 58780
rect 2696 58778 2752 58780
rect 2776 58778 2832 58780
rect 2856 58778 2912 58780
rect 2616 58726 2662 58778
rect 2662 58726 2672 58778
rect 2696 58726 2726 58778
rect 2726 58726 2738 58778
rect 2738 58726 2752 58778
rect 2776 58726 2790 58778
rect 2790 58726 2802 58778
rect 2802 58726 2832 58778
rect 2856 58726 2866 58778
rect 2866 58726 2912 58778
rect 2616 58724 2672 58726
rect 2696 58724 2752 58726
rect 2776 58724 2832 58726
rect 2856 58724 2912 58726
rect 2616 57690 2672 57692
rect 2696 57690 2752 57692
rect 2776 57690 2832 57692
rect 2856 57690 2912 57692
rect 2616 57638 2662 57690
rect 2662 57638 2672 57690
rect 2696 57638 2726 57690
rect 2726 57638 2738 57690
rect 2738 57638 2752 57690
rect 2776 57638 2790 57690
rect 2790 57638 2802 57690
rect 2802 57638 2832 57690
rect 2856 57638 2866 57690
rect 2866 57638 2912 57690
rect 2616 57636 2672 57638
rect 2696 57636 2752 57638
rect 2776 57636 2832 57638
rect 2856 57636 2912 57638
rect 3054 56616 3110 56672
rect 2616 56602 2672 56604
rect 2696 56602 2752 56604
rect 2776 56602 2832 56604
rect 2856 56602 2912 56604
rect 2616 56550 2662 56602
rect 2662 56550 2672 56602
rect 2696 56550 2726 56602
rect 2726 56550 2738 56602
rect 2738 56550 2752 56602
rect 2776 56550 2790 56602
rect 2790 56550 2802 56602
rect 2802 56550 2832 56602
rect 2856 56550 2866 56602
rect 2866 56550 2912 56602
rect 2616 56548 2672 56550
rect 2696 56548 2752 56550
rect 2776 56548 2832 56550
rect 2856 56548 2912 56550
rect 2616 55514 2672 55516
rect 2696 55514 2752 55516
rect 2776 55514 2832 55516
rect 2856 55514 2912 55516
rect 2616 55462 2662 55514
rect 2662 55462 2672 55514
rect 2696 55462 2726 55514
rect 2726 55462 2738 55514
rect 2738 55462 2752 55514
rect 2776 55462 2790 55514
rect 2790 55462 2802 55514
rect 2802 55462 2832 55514
rect 2856 55462 2866 55514
rect 2866 55462 2912 55514
rect 2616 55460 2672 55462
rect 2696 55460 2752 55462
rect 2776 55460 2832 55462
rect 2856 55460 2912 55462
rect 2616 54426 2672 54428
rect 2696 54426 2752 54428
rect 2776 54426 2832 54428
rect 2856 54426 2912 54428
rect 2616 54374 2662 54426
rect 2662 54374 2672 54426
rect 2696 54374 2726 54426
rect 2726 54374 2738 54426
rect 2738 54374 2752 54426
rect 2776 54374 2790 54426
rect 2790 54374 2802 54426
rect 2802 54374 2832 54426
rect 2856 54374 2866 54426
rect 2866 54374 2912 54426
rect 2616 54372 2672 54374
rect 2696 54372 2752 54374
rect 2776 54372 2832 54374
rect 2856 54372 2912 54374
rect 2616 53338 2672 53340
rect 2696 53338 2752 53340
rect 2776 53338 2832 53340
rect 2856 53338 2912 53340
rect 2616 53286 2662 53338
rect 2662 53286 2672 53338
rect 2696 53286 2726 53338
rect 2726 53286 2738 53338
rect 2738 53286 2752 53338
rect 2776 53286 2790 53338
rect 2790 53286 2802 53338
rect 2802 53286 2832 53338
rect 2856 53286 2866 53338
rect 2866 53286 2912 53338
rect 2616 53284 2672 53286
rect 2696 53284 2752 53286
rect 2776 53284 2832 53286
rect 2856 53284 2912 53286
rect 2616 52250 2672 52252
rect 2696 52250 2752 52252
rect 2776 52250 2832 52252
rect 2856 52250 2912 52252
rect 2616 52198 2662 52250
rect 2662 52198 2672 52250
rect 2696 52198 2726 52250
rect 2726 52198 2738 52250
rect 2738 52198 2752 52250
rect 2776 52198 2790 52250
rect 2790 52198 2802 52250
rect 2802 52198 2832 52250
rect 2856 52198 2866 52250
rect 2866 52198 2912 52250
rect 2616 52196 2672 52198
rect 2696 52196 2752 52198
rect 2776 52196 2832 52198
rect 2856 52196 2912 52198
rect 2616 51162 2672 51164
rect 2696 51162 2752 51164
rect 2776 51162 2832 51164
rect 2856 51162 2912 51164
rect 2616 51110 2662 51162
rect 2662 51110 2672 51162
rect 2696 51110 2726 51162
rect 2726 51110 2738 51162
rect 2738 51110 2752 51162
rect 2776 51110 2790 51162
rect 2790 51110 2802 51162
rect 2802 51110 2832 51162
rect 2856 51110 2866 51162
rect 2866 51110 2912 51162
rect 2616 51108 2672 51110
rect 2696 51108 2752 51110
rect 2776 51108 2832 51110
rect 2856 51108 2912 51110
rect 1956 44090 2012 44092
rect 2036 44090 2092 44092
rect 2116 44090 2172 44092
rect 2196 44090 2252 44092
rect 1956 44038 2002 44090
rect 2002 44038 2012 44090
rect 2036 44038 2066 44090
rect 2066 44038 2078 44090
rect 2078 44038 2092 44090
rect 2116 44038 2130 44090
rect 2130 44038 2142 44090
rect 2142 44038 2172 44090
rect 2196 44038 2206 44090
rect 2206 44038 2252 44090
rect 1956 44036 2012 44038
rect 2036 44036 2092 44038
rect 2116 44036 2172 44038
rect 2196 44036 2252 44038
rect 1956 43002 2012 43004
rect 2036 43002 2092 43004
rect 2116 43002 2172 43004
rect 2196 43002 2252 43004
rect 1956 42950 2002 43002
rect 2002 42950 2012 43002
rect 2036 42950 2066 43002
rect 2066 42950 2078 43002
rect 2078 42950 2092 43002
rect 2116 42950 2130 43002
rect 2130 42950 2142 43002
rect 2142 42950 2172 43002
rect 2196 42950 2206 43002
rect 2206 42950 2252 43002
rect 1956 42948 2012 42950
rect 2036 42948 2092 42950
rect 2116 42948 2172 42950
rect 2196 42948 2252 42950
rect 1956 41914 2012 41916
rect 2036 41914 2092 41916
rect 2116 41914 2172 41916
rect 2196 41914 2252 41916
rect 1956 41862 2002 41914
rect 2002 41862 2012 41914
rect 2036 41862 2066 41914
rect 2066 41862 2078 41914
rect 2078 41862 2092 41914
rect 2116 41862 2130 41914
rect 2130 41862 2142 41914
rect 2142 41862 2172 41914
rect 2196 41862 2206 41914
rect 2206 41862 2252 41914
rect 1956 41860 2012 41862
rect 2036 41860 2092 41862
rect 2116 41860 2172 41862
rect 2196 41860 2252 41862
rect 1956 40826 2012 40828
rect 2036 40826 2092 40828
rect 2116 40826 2172 40828
rect 2196 40826 2252 40828
rect 1956 40774 2002 40826
rect 2002 40774 2012 40826
rect 2036 40774 2066 40826
rect 2066 40774 2078 40826
rect 2078 40774 2092 40826
rect 2116 40774 2130 40826
rect 2130 40774 2142 40826
rect 2142 40774 2172 40826
rect 2196 40774 2206 40826
rect 2206 40774 2252 40826
rect 1956 40772 2012 40774
rect 2036 40772 2092 40774
rect 2116 40772 2172 40774
rect 2196 40772 2252 40774
rect 1956 39738 2012 39740
rect 2036 39738 2092 39740
rect 2116 39738 2172 39740
rect 2196 39738 2252 39740
rect 1956 39686 2002 39738
rect 2002 39686 2012 39738
rect 2036 39686 2066 39738
rect 2066 39686 2078 39738
rect 2078 39686 2092 39738
rect 2116 39686 2130 39738
rect 2130 39686 2142 39738
rect 2142 39686 2172 39738
rect 2196 39686 2206 39738
rect 2206 39686 2252 39738
rect 1956 39684 2012 39686
rect 2036 39684 2092 39686
rect 2116 39684 2172 39686
rect 2196 39684 2252 39686
rect 1956 38650 2012 38652
rect 2036 38650 2092 38652
rect 2116 38650 2172 38652
rect 2196 38650 2252 38652
rect 1956 38598 2002 38650
rect 2002 38598 2012 38650
rect 2036 38598 2066 38650
rect 2066 38598 2078 38650
rect 2078 38598 2092 38650
rect 2116 38598 2130 38650
rect 2130 38598 2142 38650
rect 2142 38598 2172 38650
rect 2196 38598 2206 38650
rect 2206 38598 2252 38650
rect 1956 38596 2012 38598
rect 2036 38596 2092 38598
rect 2116 38596 2172 38598
rect 2196 38596 2252 38598
rect 1956 37562 2012 37564
rect 2036 37562 2092 37564
rect 2116 37562 2172 37564
rect 2196 37562 2252 37564
rect 1956 37510 2002 37562
rect 2002 37510 2012 37562
rect 2036 37510 2066 37562
rect 2066 37510 2078 37562
rect 2078 37510 2092 37562
rect 2116 37510 2130 37562
rect 2130 37510 2142 37562
rect 2142 37510 2172 37562
rect 2196 37510 2206 37562
rect 2206 37510 2252 37562
rect 1956 37508 2012 37510
rect 2036 37508 2092 37510
rect 2116 37508 2172 37510
rect 2196 37508 2252 37510
rect 1956 36474 2012 36476
rect 2036 36474 2092 36476
rect 2116 36474 2172 36476
rect 2196 36474 2252 36476
rect 1956 36422 2002 36474
rect 2002 36422 2012 36474
rect 2036 36422 2066 36474
rect 2066 36422 2078 36474
rect 2078 36422 2092 36474
rect 2116 36422 2130 36474
rect 2130 36422 2142 36474
rect 2142 36422 2172 36474
rect 2196 36422 2206 36474
rect 2206 36422 2252 36474
rect 1956 36420 2012 36422
rect 2036 36420 2092 36422
rect 2116 36420 2172 36422
rect 2196 36420 2252 36422
rect 1956 35386 2012 35388
rect 2036 35386 2092 35388
rect 2116 35386 2172 35388
rect 2196 35386 2252 35388
rect 1956 35334 2002 35386
rect 2002 35334 2012 35386
rect 2036 35334 2066 35386
rect 2066 35334 2078 35386
rect 2078 35334 2092 35386
rect 2116 35334 2130 35386
rect 2130 35334 2142 35386
rect 2142 35334 2172 35386
rect 2196 35334 2206 35386
rect 2206 35334 2252 35386
rect 1956 35332 2012 35334
rect 2036 35332 2092 35334
rect 2116 35332 2172 35334
rect 2196 35332 2252 35334
rect 1956 34298 2012 34300
rect 2036 34298 2092 34300
rect 2116 34298 2172 34300
rect 2196 34298 2252 34300
rect 1956 34246 2002 34298
rect 2002 34246 2012 34298
rect 2036 34246 2066 34298
rect 2066 34246 2078 34298
rect 2078 34246 2092 34298
rect 2116 34246 2130 34298
rect 2130 34246 2142 34298
rect 2142 34246 2172 34298
rect 2196 34246 2206 34298
rect 2206 34246 2252 34298
rect 1956 34244 2012 34246
rect 2036 34244 2092 34246
rect 2116 34244 2172 34246
rect 2196 34244 2252 34246
rect 1956 33210 2012 33212
rect 2036 33210 2092 33212
rect 2116 33210 2172 33212
rect 2196 33210 2252 33212
rect 1956 33158 2002 33210
rect 2002 33158 2012 33210
rect 2036 33158 2066 33210
rect 2066 33158 2078 33210
rect 2078 33158 2092 33210
rect 2116 33158 2130 33210
rect 2130 33158 2142 33210
rect 2142 33158 2172 33210
rect 2196 33158 2206 33210
rect 2206 33158 2252 33210
rect 1956 33156 2012 33158
rect 2036 33156 2092 33158
rect 2116 33156 2172 33158
rect 2196 33156 2252 33158
rect 1956 32122 2012 32124
rect 2036 32122 2092 32124
rect 2116 32122 2172 32124
rect 2196 32122 2252 32124
rect 1956 32070 2002 32122
rect 2002 32070 2012 32122
rect 2036 32070 2066 32122
rect 2066 32070 2078 32122
rect 2078 32070 2092 32122
rect 2116 32070 2130 32122
rect 2130 32070 2142 32122
rect 2142 32070 2172 32122
rect 2196 32070 2206 32122
rect 2206 32070 2252 32122
rect 1956 32068 2012 32070
rect 2036 32068 2092 32070
rect 2116 32068 2172 32070
rect 2196 32068 2252 32070
rect 1956 31034 2012 31036
rect 2036 31034 2092 31036
rect 2116 31034 2172 31036
rect 2196 31034 2252 31036
rect 1956 30982 2002 31034
rect 2002 30982 2012 31034
rect 2036 30982 2066 31034
rect 2066 30982 2078 31034
rect 2078 30982 2092 31034
rect 2116 30982 2130 31034
rect 2130 30982 2142 31034
rect 2142 30982 2172 31034
rect 2196 30982 2206 31034
rect 2206 30982 2252 31034
rect 1956 30980 2012 30982
rect 2036 30980 2092 30982
rect 2116 30980 2172 30982
rect 2196 30980 2252 30982
rect 1956 29946 2012 29948
rect 2036 29946 2092 29948
rect 2116 29946 2172 29948
rect 2196 29946 2252 29948
rect 1956 29894 2002 29946
rect 2002 29894 2012 29946
rect 2036 29894 2066 29946
rect 2066 29894 2078 29946
rect 2078 29894 2092 29946
rect 2116 29894 2130 29946
rect 2130 29894 2142 29946
rect 2142 29894 2172 29946
rect 2196 29894 2206 29946
rect 2206 29894 2252 29946
rect 1956 29892 2012 29894
rect 2036 29892 2092 29894
rect 2116 29892 2172 29894
rect 2196 29892 2252 29894
rect 1956 28858 2012 28860
rect 2036 28858 2092 28860
rect 2116 28858 2172 28860
rect 2196 28858 2252 28860
rect 1956 28806 2002 28858
rect 2002 28806 2012 28858
rect 2036 28806 2066 28858
rect 2066 28806 2078 28858
rect 2078 28806 2092 28858
rect 2116 28806 2130 28858
rect 2130 28806 2142 28858
rect 2142 28806 2172 28858
rect 2196 28806 2206 28858
rect 2206 28806 2252 28858
rect 1956 28804 2012 28806
rect 2036 28804 2092 28806
rect 2116 28804 2172 28806
rect 2196 28804 2252 28806
rect 1956 27770 2012 27772
rect 2036 27770 2092 27772
rect 2116 27770 2172 27772
rect 2196 27770 2252 27772
rect 1956 27718 2002 27770
rect 2002 27718 2012 27770
rect 2036 27718 2066 27770
rect 2066 27718 2078 27770
rect 2078 27718 2092 27770
rect 2116 27718 2130 27770
rect 2130 27718 2142 27770
rect 2142 27718 2172 27770
rect 2196 27718 2206 27770
rect 2206 27718 2252 27770
rect 1956 27716 2012 27718
rect 2036 27716 2092 27718
rect 2116 27716 2172 27718
rect 2196 27716 2252 27718
rect 1956 26682 2012 26684
rect 2036 26682 2092 26684
rect 2116 26682 2172 26684
rect 2196 26682 2252 26684
rect 1956 26630 2002 26682
rect 2002 26630 2012 26682
rect 2036 26630 2066 26682
rect 2066 26630 2078 26682
rect 2078 26630 2092 26682
rect 2116 26630 2130 26682
rect 2130 26630 2142 26682
rect 2142 26630 2172 26682
rect 2196 26630 2206 26682
rect 2206 26630 2252 26682
rect 1956 26628 2012 26630
rect 2036 26628 2092 26630
rect 2116 26628 2172 26630
rect 2196 26628 2252 26630
rect 1956 25594 2012 25596
rect 2036 25594 2092 25596
rect 2116 25594 2172 25596
rect 2196 25594 2252 25596
rect 1956 25542 2002 25594
rect 2002 25542 2012 25594
rect 2036 25542 2066 25594
rect 2066 25542 2078 25594
rect 2078 25542 2092 25594
rect 2116 25542 2130 25594
rect 2130 25542 2142 25594
rect 2142 25542 2172 25594
rect 2196 25542 2206 25594
rect 2206 25542 2252 25594
rect 1956 25540 2012 25542
rect 2036 25540 2092 25542
rect 2116 25540 2172 25542
rect 2196 25540 2252 25542
rect 2616 50074 2672 50076
rect 2696 50074 2752 50076
rect 2776 50074 2832 50076
rect 2856 50074 2912 50076
rect 2616 50022 2662 50074
rect 2662 50022 2672 50074
rect 2696 50022 2726 50074
rect 2726 50022 2738 50074
rect 2738 50022 2752 50074
rect 2776 50022 2790 50074
rect 2790 50022 2802 50074
rect 2802 50022 2832 50074
rect 2856 50022 2866 50074
rect 2866 50022 2912 50074
rect 2616 50020 2672 50022
rect 2696 50020 2752 50022
rect 2776 50020 2832 50022
rect 2856 50020 2912 50022
rect 2616 48986 2672 48988
rect 2696 48986 2752 48988
rect 2776 48986 2832 48988
rect 2856 48986 2912 48988
rect 2616 48934 2662 48986
rect 2662 48934 2672 48986
rect 2696 48934 2726 48986
rect 2726 48934 2738 48986
rect 2738 48934 2752 48986
rect 2776 48934 2790 48986
rect 2790 48934 2802 48986
rect 2802 48934 2832 48986
rect 2856 48934 2866 48986
rect 2866 48934 2912 48986
rect 2616 48932 2672 48934
rect 2696 48932 2752 48934
rect 2776 48932 2832 48934
rect 2856 48932 2912 48934
rect 2616 47898 2672 47900
rect 2696 47898 2752 47900
rect 2776 47898 2832 47900
rect 2856 47898 2912 47900
rect 2616 47846 2662 47898
rect 2662 47846 2672 47898
rect 2696 47846 2726 47898
rect 2726 47846 2738 47898
rect 2738 47846 2752 47898
rect 2776 47846 2790 47898
rect 2790 47846 2802 47898
rect 2802 47846 2832 47898
rect 2856 47846 2866 47898
rect 2866 47846 2912 47898
rect 2616 47844 2672 47846
rect 2696 47844 2752 47846
rect 2776 47844 2832 47846
rect 2856 47844 2912 47846
rect 3054 47232 3110 47288
rect 2616 46810 2672 46812
rect 2696 46810 2752 46812
rect 2776 46810 2832 46812
rect 2856 46810 2912 46812
rect 2616 46758 2662 46810
rect 2662 46758 2672 46810
rect 2696 46758 2726 46810
rect 2726 46758 2738 46810
rect 2738 46758 2752 46810
rect 2776 46758 2790 46810
rect 2790 46758 2802 46810
rect 2802 46758 2832 46810
rect 2856 46758 2866 46810
rect 2866 46758 2912 46810
rect 2616 46756 2672 46758
rect 2696 46756 2752 46758
rect 2776 46756 2832 46758
rect 2856 46756 2912 46758
rect 2616 45722 2672 45724
rect 2696 45722 2752 45724
rect 2776 45722 2832 45724
rect 2856 45722 2912 45724
rect 2616 45670 2662 45722
rect 2662 45670 2672 45722
rect 2696 45670 2726 45722
rect 2726 45670 2738 45722
rect 2738 45670 2752 45722
rect 2776 45670 2790 45722
rect 2790 45670 2802 45722
rect 2802 45670 2832 45722
rect 2856 45670 2866 45722
rect 2866 45670 2912 45722
rect 2616 45668 2672 45670
rect 2696 45668 2752 45670
rect 2776 45668 2832 45670
rect 2856 45668 2912 45670
rect 2616 44634 2672 44636
rect 2696 44634 2752 44636
rect 2776 44634 2832 44636
rect 2856 44634 2912 44636
rect 2616 44582 2662 44634
rect 2662 44582 2672 44634
rect 2696 44582 2726 44634
rect 2726 44582 2738 44634
rect 2738 44582 2752 44634
rect 2776 44582 2790 44634
rect 2790 44582 2802 44634
rect 2802 44582 2832 44634
rect 2856 44582 2866 44634
rect 2866 44582 2912 44634
rect 2616 44580 2672 44582
rect 2696 44580 2752 44582
rect 2776 44580 2832 44582
rect 2856 44580 2912 44582
rect 2616 43546 2672 43548
rect 2696 43546 2752 43548
rect 2776 43546 2832 43548
rect 2856 43546 2912 43548
rect 2616 43494 2662 43546
rect 2662 43494 2672 43546
rect 2696 43494 2726 43546
rect 2726 43494 2738 43546
rect 2738 43494 2752 43546
rect 2776 43494 2790 43546
rect 2790 43494 2802 43546
rect 2802 43494 2832 43546
rect 2856 43494 2866 43546
rect 2866 43494 2912 43546
rect 2616 43492 2672 43494
rect 2696 43492 2752 43494
rect 2776 43492 2832 43494
rect 2856 43492 2912 43494
rect 2616 42458 2672 42460
rect 2696 42458 2752 42460
rect 2776 42458 2832 42460
rect 2856 42458 2912 42460
rect 2616 42406 2662 42458
rect 2662 42406 2672 42458
rect 2696 42406 2726 42458
rect 2726 42406 2738 42458
rect 2738 42406 2752 42458
rect 2776 42406 2790 42458
rect 2790 42406 2802 42458
rect 2802 42406 2832 42458
rect 2856 42406 2866 42458
rect 2866 42406 2912 42458
rect 2616 42404 2672 42406
rect 2696 42404 2752 42406
rect 2776 42404 2832 42406
rect 2856 42404 2912 42406
rect 2616 41370 2672 41372
rect 2696 41370 2752 41372
rect 2776 41370 2832 41372
rect 2856 41370 2912 41372
rect 2616 41318 2662 41370
rect 2662 41318 2672 41370
rect 2696 41318 2726 41370
rect 2726 41318 2738 41370
rect 2738 41318 2752 41370
rect 2776 41318 2790 41370
rect 2790 41318 2802 41370
rect 2802 41318 2832 41370
rect 2856 41318 2866 41370
rect 2866 41318 2912 41370
rect 2616 41316 2672 41318
rect 2696 41316 2752 41318
rect 2776 41316 2832 41318
rect 2856 41316 2912 41318
rect 2616 40282 2672 40284
rect 2696 40282 2752 40284
rect 2776 40282 2832 40284
rect 2856 40282 2912 40284
rect 2616 40230 2662 40282
rect 2662 40230 2672 40282
rect 2696 40230 2726 40282
rect 2726 40230 2738 40282
rect 2738 40230 2752 40282
rect 2776 40230 2790 40282
rect 2790 40230 2802 40282
rect 2802 40230 2832 40282
rect 2856 40230 2866 40282
rect 2866 40230 2912 40282
rect 2616 40228 2672 40230
rect 2696 40228 2752 40230
rect 2776 40228 2832 40230
rect 2856 40228 2912 40230
rect 2616 39194 2672 39196
rect 2696 39194 2752 39196
rect 2776 39194 2832 39196
rect 2856 39194 2912 39196
rect 2616 39142 2662 39194
rect 2662 39142 2672 39194
rect 2696 39142 2726 39194
rect 2726 39142 2738 39194
rect 2738 39142 2752 39194
rect 2776 39142 2790 39194
rect 2790 39142 2802 39194
rect 2802 39142 2832 39194
rect 2856 39142 2866 39194
rect 2866 39142 2912 39194
rect 2616 39140 2672 39142
rect 2696 39140 2752 39142
rect 2776 39140 2832 39142
rect 2856 39140 2912 39142
rect 2616 38106 2672 38108
rect 2696 38106 2752 38108
rect 2776 38106 2832 38108
rect 2856 38106 2912 38108
rect 2616 38054 2662 38106
rect 2662 38054 2672 38106
rect 2696 38054 2726 38106
rect 2726 38054 2738 38106
rect 2738 38054 2752 38106
rect 2776 38054 2790 38106
rect 2790 38054 2802 38106
rect 2802 38054 2832 38106
rect 2856 38054 2866 38106
rect 2866 38054 2912 38106
rect 2616 38052 2672 38054
rect 2696 38052 2752 38054
rect 2776 38052 2832 38054
rect 2856 38052 2912 38054
rect 2616 37018 2672 37020
rect 2696 37018 2752 37020
rect 2776 37018 2832 37020
rect 2856 37018 2912 37020
rect 2616 36966 2662 37018
rect 2662 36966 2672 37018
rect 2696 36966 2726 37018
rect 2726 36966 2738 37018
rect 2738 36966 2752 37018
rect 2776 36966 2790 37018
rect 2790 36966 2802 37018
rect 2802 36966 2832 37018
rect 2856 36966 2866 37018
rect 2866 36966 2912 37018
rect 2616 36964 2672 36966
rect 2696 36964 2752 36966
rect 2776 36964 2832 36966
rect 2856 36964 2912 36966
rect 2616 35930 2672 35932
rect 2696 35930 2752 35932
rect 2776 35930 2832 35932
rect 2856 35930 2912 35932
rect 2616 35878 2662 35930
rect 2662 35878 2672 35930
rect 2696 35878 2726 35930
rect 2726 35878 2738 35930
rect 2738 35878 2752 35930
rect 2776 35878 2790 35930
rect 2790 35878 2802 35930
rect 2802 35878 2832 35930
rect 2856 35878 2866 35930
rect 2866 35878 2912 35930
rect 2616 35876 2672 35878
rect 2696 35876 2752 35878
rect 2776 35876 2832 35878
rect 2856 35876 2912 35878
rect 2616 34842 2672 34844
rect 2696 34842 2752 34844
rect 2776 34842 2832 34844
rect 2856 34842 2912 34844
rect 2616 34790 2662 34842
rect 2662 34790 2672 34842
rect 2696 34790 2726 34842
rect 2726 34790 2738 34842
rect 2738 34790 2752 34842
rect 2776 34790 2790 34842
rect 2790 34790 2802 34842
rect 2802 34790 2832 34842
rect 2856 34790 2866 34842
rect 2866 34790 2912 34842
rect 2616 34788 2672 34790
rect 2696 34788 2752 34790
rect 2776 34788 2832 34790
rect 2856 34788 2912 34790
rect 2616 33754 2672 33756
rect 2696 33754 2752 33756
rect 2776 33754 2832 33756
rect 2856 33754 2912 33756
rect 2616 33702 2662 33754
rect 2662 33702 2672 33754
rect 2696 33702 2726 33754
rect 2726 33702 2738 33754
rect 2738 33702 2752 33754
rect 2776 33702 2790 33754
rect 2790 33702 2802 33754
rect 2802 33702 2832 33754
rect 2856 33702 2866 33754
rect 2866 33702 2912 33754
rect 2616 33700 2672 33702
rect 2696 33700 2752 33702
rect 2776 33700 2832 33702
rect 2856 33700 2912 33702
rect 2616 32666 2672 32668
rect 2696 32666 2752 32668
rect 2776 32666 2832 32668
rect 2856 32666 2912 32668
rect 2616 32614 2662 32666
rect 2662 32614 2672 32666
rect 2696 32614 2726 32666
rect 2726 32614 2738 32666
rect 2738 32614 2752 32666
rect 2776 32614 2790 32666
rect 2790 32614 2802 32666
rect 2802 32614 2832 32666
rect 2856 32614 2866 32666
rect 2866 32614 2912 32666
rect 2616 32612 2672 32614
rect 2696 32612 2752 32614
rect 2776 32612 2832 32614
rect 2856 32612 2912 32614
rect 1956 24506 2012 24508
rect 2036 24506 2092 24508
rect 2116 24506 2172 24508
rect 2196 24506 2252 24508
rect 1956 24454 2002 24506
rect 2002 24454 2012 24506
rect 2036 24454 2066 24506
rect 2066 24454 2078 24506
rect 2078 24454 2092 24506
rect 2116 24454 2130 24506
rect 2130 24454 2142 24506
rect 2142 24454 2172 24506
rect 2196 24454 2206 24506
rect 2206 24454 2252 24506
rect 1956 24452 2012 24454
rect 2036 24452 2092 24454
rect 2116 24452 2172 24454
rect 2196 24452 2252 24454
rect 1956 23418 2012 23420
rect 2036 23418 2092 23420
rect 2116 23418 2172 23420
rect 2196 23418 2252 23420
rect 1956 23366 2002 23418
rect 2002 23366 2012 23418
rect 2036 23366 2066 23418
rect 2066 23366 2078 23418
rect 2078 23366 2092 23418
rect 2116 23366 2130 23418
rect 2130 23366 2142 23418
rect 2142 23366 2172 23418
rect 2196 23366 2206 23418
rect 2206 23366 2252 23418
rect 1956 23364 2012 23366
rect 2036 23364 2092 23366
rect 2116 23364 2172 23366
rect 2196 23364 2252 23366
rect 1956 22330 2012 22332
rect 2036 22330 2092 22332
rect 2116 22330 2172 22332
rect 2196 22330 2252 22332
rect 1956 22278 2002 22330
rect 2002 22278 2012 22330
rect 2036 22278 2066 22330
rect 2066 22278 2078 22330
rect 2078 22278 2092 22330
rect 2116 22278 2130 22330
rect 2130 22278 2142 22330
rect 2142 22278 2172 22330
rect 2196 22278 2206 22330
rect 2206 22278 2252 22330
rect 1956 22276 2012 22278
rect 2036 22276 2092 22278
rect 2116 22276 2172 22278
rect 2196 22276 2252 22278
rect 2502 31728 2558 31784
rect 1956 21242 2012 21244
rect 2036 21242 2092 21244
rect 2116 21242 2172 21244
rect 2196 21242 2252 21244
rect 1956 21190 2002 21242
rect 2002 21190 2012 21242
rect 2036 21190 2066 21242
rect 2066 21190 2078 21242
rect 2078 21190 2092 21242
rect 2116 21190 2130 21242
rect 2130 21190 2142 21242
rect 2142 21190 2172 21242
rect 2196 21190 2206 21242
rect 2206 21190 2252 21242
rect 1956 21188 2012 21190
rect 2036 21188 2092 21190
rect 2116 21188 2172 21190
rect 2196 21188 2252 21190
rect 1956 20154 2012 20156
rect 2036 20154 2092 20156
rect 2116 20154 2172 20156
rect 2196 20154 2252 20156
rect 1956 20102 2002 20154
rect 2002 20102 2012 20154
rect 2036 20102 2066 20154
rect 2066 20102 2078 20154
rect 2078 20102 2092 20154
rect 2116 20102 2130 20154
rect 2130 20102 2142 20154
rect 2142 20102 2172 20154
rect 2196 20102 2206 20154
rect 2206 20102 2252 20154
rect 1956 20100 2012 20102
rect 2036 20100 2092 20102
rect 2116 20100 2172 20102
rect 2196 20100 2252 20102
rect 1956 19066 2012 19068
rect 2036 19066 2092 19068
rect 2116 19066 2172 19068
rect 2196 19066 2252 19068
rect 1956 19014 2002 19066
rect 2002 19014 2012 19066
rect 2036 19014 2066 19066
rect 2066 19014 2078 19066
rect 2078 19014 2092 19066
rect 2116 19014 2130 19066
rect 2130 19014 2142 19066
rect 2142 19014 2172 19066
rect 2196 19014 2206 19066
rect 2206 19014 2252 19066
rect 1956 19012 2012 19014
rect 2036 19012 2092 19014
rect 2116 19012 2172 19014
rect 2196 19012 2252 19014
rect 1956 17978 2012 17980
rect 2036 17978 2092 17980
rect 2116 17978 2172 17980
rect 2196 17978 2252 17980
rect 1956 17926 2002 17978
rect 2002 17926 2012 17978
rect 2036 17926 2066 17978
rect 2066 17926 2078 17978
rect 2078 17926 2092 17978
rect 2116 17926 2130 17978
rect 2130 17926 2142 17978
rect 2142 17926 2172 17978
rect 2196 17926 2206 17978
rect 2206 17926 2252 17978
rect 1956 17924 2012 17926
rect 2036 17924 2092 17926
rect 2116 17924 2172 17926
rect 2196 17924 2252 17926
rect 1956 16890 2012 16892
rect 2036 16890 2092 16892
rect 2116 16890 2172 16892
rect 2196 16890 2252 16892
rect 1956 16838 2002 16890
rect 2002 16838 2012 16890
rect 2036 16838 2066 16890
rect 2066 16838 2078 16890
rect 2078 16838 2092 16890
rect 2116 16838 2130 16890
rect 2130 16838 2142 16890
rect 2142 16838 2172 16890
rect 2196 16838 2206 16890
rect 2206 16838 2252 16890
rect 1956 16836 2012 16838
rect 2036 16836 2092 16838
rect 2116 16836 2172 16838
rect 2196 16836 2252 16838
rect 1956 15802 2012 15804
rect 2036 15802 2092 15804
rect 2116 15802 2172 15804
rect 2196 15802 2252 15804
rect 1956 15750 2002 15802
rect 2002 15750 2012 15802
rect 2036 15750 2066 15802
rect 2066 15750 2078 15802
rect 2078 15750 2092 15802
rect 2116 15750 2130 15802
rect 2130 15750 2142 15802
rect 2142 15750 2172 15802
rect 2196 15750 2206 15802
rect 2206 15750 2252 15802
rect 1956 15748 2012 15750
rect 2036 15748 2092 15750
rect 2116 15748 2172 15750
rect 2196 15748 2252 15750
rect 1956 14714 2012 14716
rect 2036 14714 2092 14716
rect 2116 14714 2172 14716
rect 2196 14714 2252 14716
rect 1956 14662 2002 14714
rect 2002 14662 2012 14714
rect 2036 14662 2066 14714
rect 2066 14662 2078 14714
rect 2078 14662 2092 14714
rect 2116 14662 2130 14714
rect 2130 14662 2142 14714
rect 2142 14662 2172 14714
rect 2196 14662 2206 14714
rect 2206 14662 2252 14714
rect 1956 14660 2012 14662
rect 2036 14660 2092 14662
rect 2116 14660 2172 14662
rect 2196 14660 2252 14662
rect 1956 13626 2012 13628
rect 2036 13626 2092 13628
rect 2116 13626 2172 13628
rect 2196 13626 2252 13628
rect 1956 13574 2002 13626
rect 2002 13574 2012 13626
rect 2036 13574 2066 13626
rect 2066 13574 2078 13626
rect 2078 13574 2092 13626
rect 2116 13574 2130 13626
rect 2130 13574 2142 13626
rect 2142 13574 2172 13626
rect 2196 13574 2206 13626
rect 2206 13574 2252 13626
rect 1956 13572 2012 13574
rect 2036 13572 2092 13574
rect 2116 13572 2172 13574
rect 2196 13572 2252 13574
rect 1956 12538 2012 12540
rect 2036 12538 2092 12540
rect 2116 12538 2172 12540
rect 2196 12538 2252 12540
rect 1956 12486 2002 12538
rect 2002 12486 2012 12538
rect 2036 12486 2066 12538
rect 2066 12486 2078 12538
rect 2078 12486 2092 12538
rect 2116 12486 2130 12538
rect 2130 12486 2142 12538
rect 2142 12486 2172 12538
rect 2196 12486 2206 12538
rect 2206 12486 2252 12538
rect 1956 12484 2012 12486
rect 2036 12484 2092 12486
rect 2116 12484 2172 12486
rect 2196 12484 2252 12486
rect 1956 11450 2012 11452
rect 2036 11450 2092 11452
rect 2116 11450 2172 11452
rect 2196 11450 2252 11452
rect 1956 11398 2002 11450
rect 2002 11398 2012 11450
rect 2036 11398 2066 11450
rect 2066 11398 2078 11450
rect 2078 11398 2092 11450
rect 2116 11398 2130 11450
rect 2130 11398 2142 11450
rect 2142 11398 2172 11450
rect 2196 11398 2206 11450
rect 2206 11398 2252 11450
rect 1956 11396 2012 11398
rect 2036 11396 2092 11398
rect 2116 11396 2172 11398
rect 2196 11396 2252 11398
rect 1956 10362 2012 10364
rect 2036 10362 2092 10364
rect 2116 10362 2172 10364
rect 2196 10362 2252 10364
rect 1956 10310 2002 10362
rect 2002 10310 2012 10362
rect 2036 10310 2066 10362
rect 2066 10310 2078 10362
rect 2078 10310 2092 10362
rect 2116 10310 2130 10362
rect 2130 10310 2142 10362
rect 2142 10310 2172 10362
rect 2196 10310 2206 10362
rect 2206 10310 2252 10362
rect 1956 10308 2012 10310
rect 2036 10308 2092 10310
rect 2116 10308 2172 10310
rect 2196 10308 2252 10310
rect 1956 9274 2012 9276
rect 2036 9274 2092 9276
rect 2116 9274 2172 9276
rect 2196 9274 2252 9276
rect 1956 9222 2002 9274
rect 2002 9222 2012 9274
rect 2036 9222 2066 9274
rect 2066 9222 2078 9274
rect 2078 9222 2092 9274
rect 2116 9222 2130 9274
rect 2130 9222 2142 9274
rect 2142 9222 2172 9274
rect 2196 9222 2206 9274
rect 2206 9222 2252 9274
rect 1956 9220 2012 9222
rect 2036 9220 2092 9222
rect 2116 9220 2172 9222
rect 2196 9220 2252 9222
rect 2616 31578 2672 31580
rect 2696 31578 2752 31580
rect 2776 31578 2832 31580
rect 2856 31578 2912 31580
rect 2616 31526 2662 31578
rect 2662 31526 2672 31578
rect 2696 31526 2726 31578
rect 2726 31526 2738 31578
rect 2738 31526 2752 31578
rect 2776 31526 2790 31578
rect 2790 31526 2802 31578
rect 2802 31526 2832 31578
rect 2856 31526 2866 31578
rect 2866 31526 2912 31578
rect 2616 31524 2672 31526
rect 2696 31524 2752 31526
rect 2776 31524 2832 31526
rect 2856 31524 2912 31526
rect 2616 30490 2672 30492
rect 2696 30490 2752 30492
rect 2776 30490 2832 30492
rect 2856 30490 2912 30492
rect 2616 30438 2662 30490
rect 2662 30438 2672 30490
rect 2696 30438 2726 30490
rect 2726 30438 2738 30490
rect 2738 30438 2752 30490
rect 2776 30438 2790 30490
rect 2790 30438 2802 30490
rect 2802 30438 2832 30490
rect 2856 30438 2866 30490
rect 2866 30438 2912 30490
rect 2616 30436 2672 30438
rect 2696 30436 2752 30438
rect 2776 30436 2832 30438
rect 2856 30436 2912 30438
rect 2616 29402 2672 29404
rect 2696 29402 2752 29404
rect 2776 29402 2832 29404
rect 2856 29402 2912 29404
rect 2616 29350 2662 29402
rect 2662 29350 2672 29402
rect 2696 29350 2726 29402
rect 2726 29350 2738 29402
rect 2738 29350 2752 29402
rect 2776 29350 2790 29402
rect 2790 29350 2802 29402
rect 2802 29350 2832 29402
rect 2856 29350 2866 29402
rect 2866 29350 2912 29402
rect 2616 29348 2672 29350
rect 2696 29348 2752 29350
rect 2776 29348 2832 29350
rect 2856 29348 2912 29350
rect 2616 28314 2672 28316
rect 2696 28314 2752 28316
rect 2776 28314 2832 28316
rect 2856 28314 2912 28316
rect 2616 28262 2662 28314
rect 2662 28262 2672 28314
rect 2696 28262 2726 28314
rect 2726 28262 2738 28314
rect 2738 28262 2752 28314
rect 2776 28262 2790 28314
rect 2790 28262 2802 28314
rect 2802 28262 2832 28314
rect 2856 28262 2866 28314
rect 2866 28262 2912 28314
rect 2616 28260 2672 28262
rect 2696 28260 2752 28262
rect 2776 28260 2832 28262
rect 2856 28260 2912 28262
rect 2616 27226 2672 27228
rect 2696 27226 2752 27228
rect 2776 27226 2832 27228
rect 2856 27226 2912 27228
rect 2616 27174 2662 27226
rect 2662 27174 2672 27226
rect 2696 27174 2726 27226
rect 2726 27174 2738 27226
rect 2738 27174 2752 27226
rect 2776 27174 2790 27226
rect 2790 27174 2802 27226
rect 2802 27174 2832 27226
rect 2856 27174 2866 27226
rect 2866 27174 2912 27226
rect 2616 27172 2672 27174
rect 2696 27172 2752 27174
rect 2776 27172 2832 27174
rect 2856 27172 2912 27174
rect 2616 26138 2672 26140
rect 2696 26138 2752 26140
rect 2776 26138 2832 26140
rect 2856 26138 2912 26140
rect 2616 26086 2662 26138
rect 2662 26086 2672 26138
rect 2696 26086 2726 26138
rect 2726 26086 2738 26138
rect 2738 26086 2752 26138
rect 2776 26086 2790 26138
rect 2790 26086 2802 26138
rect 2802 26086 2832 26138
rect 2856 26086 2866 26138
rect 2866 26086 2912 26138
rect 2616 26084 2672 26086
rect 2696 26084 2752 26086
rect 2776 26084 2832 26086
rect 2856 26084 2912 26086
rect 2616 25050 2672 25052
rect 2696 25050 2752 25052
rect 2776 25050 2832 25052
rect 2856 25050 2912 25052
rect 2616 24998 2662 25050
rect 2662 24998 2672 25050
rect 2696 24998 2726 25050
rect 2726 24998 2738 25050
rect 2738 24998 2752 25050
rect 2776 24998 2790 25050
rect 2790 24998 2802 25050
rect 2802 24998 2832 25050
rect 2856 24998 2866 25050
rect 2866 24998 2912 25050
rect 2616 24996 2672 24998
rect 2696 24996 2752 24998
rect 2776 24996 2832 24998
rect 2856 24996 2912 24998
rect 2616 23962 2672 23964
rect 2696 23962 2752 23964
rect 2776 23962 2832 23964
rect 2856 23962 2912 23964
rect 2616 23910 2662 23962
rect 2662 23910 2672 23962
rect 2696 23910 2726 23962
rect 2726 23910 2738 23962
rect 2738 23910 2752 23962
rect 2776 23910 2790 23962
rect 2790 23910 2802 23962
rect 2802 23910 2832 23962
rect 2856 23910 2866 23962
rect 2866 23910 2912 23962
rect 2616 23908 2672 23910
rect 2696 23908 2752 23910
rect 2776 23908 2832 23910
rect 2856 23908 2912 23910
rect 2616 22874 2672 22876
rect 2696 22874 2752 22876
rect 2776 22874 2832 22876
rect 2856 22874 2912 22876
rect 2616 22822 2662 22874
rect 2662 22822 2672 22874
rect 2696 22822 2726 22874
rect 2726 22822 2738 22874
rect 2738 22822 2752 22874
rect 2776 22822 2790 22874
rect 2790 22822 2802 22874
rect 2802 22822 2832 22874
rect 2856 22822 2866 22874
rect 2866 22822 2912 22874
rect 2616 22820 2672 22822
rect 2696 22820 2752 22822
rect 2776 22820 2832 22822
rect 2856 22820 2912 22822
rect 2616 21786 2672 21788
rect 2696 21786 2752 21788
rect 2776 21786 2832 21788
rect 2856 21786 2912 21788
rect 2616 21734 2662 21786
rect 2662 21734 2672 21786
rect 2696 21734 2726 21786
rect 2726 21734 2738 21786
rect 2738 21734 2752 21786
rect 2776 21734 2790 21786
rect 2790 21734 2802 21786
rect 2802 21734 2832 21786
rect 2856 21734 2866 21786
rect 2866 21734 2912 21786
rect 2616 21732 2672 21734
rect 2696 21732 2752 21734
rect 2776 21732 2832 21734
rect 2856 21732 2912 21734
rect 2616 20698 2672 20700
rect 2696 20698 2752 20700
rect 2776 20698 2832 20700
rect 2856 20698 2912 20700
rect 2616 20646 2662 20698
rect 2662 20646 2672 20698
rect 2696 20646 2726 20698
rect 2726 20646 2738 20698
rect 2738 20646 2752 20698
rect 2776 20646 2790 20698
rect 2790 20646 2802 20698
rect 2802 20646 2832 20698
rect 2856 20646 2866 20698
rect 2866 20646 2912 20698
rect 2616 20644 2672 20646
rect 2696 20644 2752 20646
rect 2776 20644 2832 20646
rect 2856 20644 2912 20646
rect 2616 19610 2672 19612
rect 2696 19610 2752 19612
rect 2776 19610 2832 19612
rect 2856 19610 2912 19612
rect 2616 19558 2662 19610
rect 2662 19558 2672 19610
rect 2696 19558 2726 19610
rect 2726 19558 2738 19610
rect 2738 19558 2752 19610
rect 2776 19558 2790 19610
rect 2790 19558 2802 19610
rect 2802 19558 2832 19610
rect 2856 19558 2866 19610
rect 2866 19558 2912 19610
rect 2616 19556 2672 19558
rect 2696 19556 2752 19558
rect 2776 19556 2832 19558
rect 2856 19556 2912 19558
rect 2616 18522 2672 18524
rect 2696 18522 2752 18524
rect 2776 18522 2832 18524
rect 2856 18522 2912 18524
rect 2616 18470 2662 18522
rect 2662 18470 2672 18522
rect 2696 18470 2726 18522
rect 2726 18470 2738 18522
rect 2738 18470 2752 18522
rect 2776 18470 2790 18522
rect 2790 18470 2802 18522
rect 2802 18470 2832 18522
rect 2856 18470 2866 18522
rect 2866 18470 2912 18522
rect 2616 18468 2672 18470
rect 2696 18468 2752 18470
rect 2776 18468 2832 18470
rect 2856 18468 2912 18470
rect 2616 17434 2672 17436
rect 2696 17434 2752 17436
rect 2776 17434 2832 17436
rect 2856 17434 2912 17436
rect 2616 17382 2662 17434
rect 2662 17382 2672 17434
rect 2696 17382 2726 17434
rect 2726 17382 2738 17434
rect 2738 17382 2752 17434
rect 2776 17382 2790 17434
rect 2790 17382 2802 17434
rect 2802 17382 2832 17434
rect 2856 17382 2866 17434
rect 2866 17382 2912 17434
rect 2616 17380 2672 17382
rect 2696 17380 2752 17382
rect 2776 17380 2832 17382
rect 2856 17380 2912 17382
rect 2616 16346 2672 16348
rect 2696 16346 2752 16348
rect 2776 16346 2832 16348
rect 2856 16346 2912 16348
rect 2616 16294 2662 16346
rect 2662 16294 2672 16346
rect 2696 16294 2726 16346
rect 2726 16294 2738 16346
rect 2738 16294 2752 16346
rect 2776 16294 2790 16346
rect 2790 16294 2802 16346
rect 2802 16294 2832 16346
rect 2856 16294 2866 16346
rect 2866 16294 2912 16346
rect 2616 16292 2672 16294
rect 2696 16292 2752 16294
rect 2776 16292 2832 16294
rect 2856 16292 2912 16294
rect 2616 15258 2672 15260
rect 2696 15258 2752 15260
rect 2776 15258 2832 15260
rect 2856 15258 2912 15260
rect 2616 15206 2662 15258
rect 2662 15206 2672 15258
rect 2696 15206 2726 15258
rect 2726 15206 2738 15258
rect 2738 15206 2752 15258
rect 2776 15206 2790 15258
rect 2790 15206 2802 15258
rect 2802 15206 2832 15258
rect 2856 15206 2866 15258
rect 2866 15206 2912 15258
rect 2616 15204 2672 15206
rect 2696 15204 2752 15206
rect 2776 15204 2832 15206
rect 2856 15204 2912 15206
rect 2616 14170 2672 14172
rect 2696 14170 2752 14172
rect 2776 14170 2832 14172
rect 2856 14170 2912 14172
rect 2616 14118 2662 14170
rect 2662 14118 2672 14170
rect 2696 14118 2726 14170
rect 2726 14118 2738 14170
rect 2738 14118 2752 14170
rect 2776 14118 2790 14170
rect 2790 14118 2802 14170
rect 2802 14118 2832 14170
rect 2856 14118 2866 14170
rect 2866 14118 2912 14170
rect 2616 14116 2672 14118
rect 2696 14116 2752 14118
rect 2776 14116 2832 14118
rect 2856 14116 2912 14118
rect 2616 13082 2672 13084
rect 2696 13082 2752 13084
rect 2776 13082 2832 13084
rect 2856 13082 2912 13084
rect 2616 13030 2662 13082
rect 2662 13030 2672 13082
rect 2696 13030 2726 13082
rect 2726 13030 2738 13082
rect 2738 13030 2752 13082
rect 2776 13030 2790 13082
rect 2790 13030 2802 13082
rect 2802 13030 2832 13082
rect 2856 13030 2866 13082
rect 2866 13030 2912 13082
rect 2616 13028 2672 13030
rect 2696 13028 2752 13030
rect 2776 13028 2832 13030
rect 2856 13028 2912 13030
rect 2616 11994 2672 11996
rect 2696 11994 2752 11996
rect 2776 11994 2832 11996
rect 2856 11994 2912 11996
rect 2616 11942 2662 11994
rect 2662 11942 2672 11994
rect 2696 11942 2726 11994
rect 2726 11942 2738 11994
rect 2738 11942 2752 11994
rect 2776 11942 2790 11994
rect 2790 11942 2802 11994
rect 2802 11942 2832 11994
rect 2856 11942 2866 11994
rect 2866 11942 2912 11994
rect 2616 11940 2672 11942
rect 2696 11940 2752 11942
rect 2776 11940 2832 11942
rect 2856 11940 2912 11942
rect 2616 10906 2672 10908
rect 2696 10906 2752 10908
rect 2776 10906 2832 10908
rect 2856 10906 2912 10908
rect 2616 10854 2662 10906
rect 2662 10854 2672 10906
rect 2696 10854 2726 10906
rect 2726 10854 2738 10906
rect 2738 10854 2752 10906
rect 2776 10854 2790 10906
rect 2790 10854 2802 10906
rect 2802 10854 2832 10906
rect 2856 10854 2866 10906
rect 2866 10854 2912 10906
rect 2616 10852 2672 10854
rect 2696 10852 2752 10854
rect 2776 10852 2832 10854
rect 2856 10852 2912 10854
rect 2594 10684 2596 10704
rect 2596 10684 2648 10704
rect 2648 10684 2650 10704
rect 2594 10648 2650 10684
rect 2616 9818 2672 9820
rect 2696 9818 2752 9820
rect 2776 9818 2832 9820
rect 2856 9818 2912 9820
rect 2616 9766 2662 9818
rect 2662 9766 2672 9818
rect 2696 9766 2726 9818
rect 2726 9766 2738 9818
rect 2738 9766 2752 9818
rect 2776 9766 2790 9818
rect 2790 9766 2802 9818
rect 2802 9766 2832 9818
rect 2856 9766 2866 9818
rect 2866 9766 2912 9818
rect 2616 9764 2672 9766
rect 2696 9764 2752 9766
rect 2776 9764 2832 9766
rect 2856 9764 2912 9766
rect 2616 8730 2672 8732
rect 2696 8730 2752 8732
rect 2776 8730 2832 8732
rect 2856 8730 2912 8732
rect 2616 8678 2662 8730
rect 2662 8678 2672 8730
rect 2696 8678 2726 8730
rect 2726 8678 2738 8730
rect 2738 8678 2752 8730
rect 2776 8678 2790 8730
rect 2790 8678 2802 8730
rect 2802 8678 2832 8730
rect 2856 8678 2866 8730
rect 2866 8678 2912 8730
rect 2616 8676 2672 8678
rect 2696 8676 2752 8678
rect 2776 8676 2832 8678
rect 2856 8676 2912 8678
rect 1956 8186 2012 8188
rect 2036 8186 2092 8188
rect 2116 8186 2172 8188
rect 2196 8186 2252 8188
rect 1956 8134 2002 8186
rect 2002 8134 2012 8186
rect 2036 8134 2066 8186
rect 2066 8134 2078 8186
rect 2078 8134 2092 8186
rect 2116 8134 2130 8186
rect 2130 8134 2142 8186
rect 2142 8134 2172 8186
rect 2196 8134 2206 8186
rect 2206 8134 2252 8186
rect 1956 8132 2012 8134
rect 2036 8132 2092 8134
rect 2116 8132 2172 8134
rect 2196 8132 2252 8134
rect 1956 7098 2012 7100
rect 2036 7098 2092 7100
rect 2116 7098 2172 7100
rect 2196 7098 2252 7100
rect 1956 7046 2002 7098
rect 2002 7046 2012 7098
rect 2036 7046 2066 7098
rect 2066 7046 2078 7098
rect 2078 7046 2092 7098
rect 2116 7046 2130 7098
rect 2130 7046 2142 7098
rect 2142 7046 2172 7098
rect 2196 7046 2206 7098
rect 2206 7046 2252 7098
rect 1956 7044 2012 7046
rect 2036 7044 2092 7046
rect 2116 7044 2172 7046
rect 2196 7044 2252 7046
rect 1956 6010 2012 6012
rect 2036 6010 2092 6012
rect 2116 6010 2172 6012
rect 2196 6010 2252 6012
rect 1956 5958 2002 6010
rect 2002 5958 2012 6010
rect 2036 5958 2066 6010
rect 2066 5958 2078 6010
rect 2078 5958 2092 6010
rect 2116 5958 2130 6010
rect 2130 5958 2142 6010
rect 2142 5958 2172 6010
rect 2196 5958 2206 6010
rect 2206 5958 2252 6010
rect 1956 5956 2012 5958
rect 2036 5956 2092 5958
rect 2116 5956 2172 5958
rect 2196 5956 2252 5958
rect 3698 48184 3754 48240
rect 4066 65184 4122 65240
rect 2616 7642 2672 7644
rect 2696 7642 2752 7644
rect 2776 7642 2832 7644
rect 2856 7642 2912 7644
rect 2616 7590 2662 7642
rect 2662 7590 2672 7642
rect 2696 7590 2726 7642
rect 2726 7590 2738 7642
rect 2738 7590 2752 7642
rect 2776 7590 2790 7642
rect 2790 7590 2802 7642
rect 2802 7590 2832 7642
rect 2856 7590 2866 7642
rect 2866 7590 2912 7642
rect 2616 7588 2672 7590
rect 2696 7588 2752 7590
rect 2776 7588 2832 7590
rect 2856 7588 2912 7590
rect 2616 6554 2672 6556
rect 2696 6554 2752 6556
rect 2776 6554 2832 6556
rect 2856 6554 2912 6556
rect 2616 6502 2662 6554
rect 2662 6502 2672 6554
rect 2696 6502 2726 6554
rect 2726 6502 2738 6554
rect 2738 6502 2752 6554
rect 2776 6502 2790 6554
rect 2790 6502 2802 6554
rect 2802 6502 2832 6554
rect 2856 6502 2866 6554
rect 2866 6502 2912 6554
rect 2616 6500 2672 6502
rect 2696 6500 2752 6502
rect 2776 6500 2832 6502
rect 2856 6500 2912 6502
rect 4250 62212 4306 62248
rect 4250 62192 4252 62212
rect 4252 62192 4304 62212
rect 4304 62192 4306 62212
rect 4158 21936 4214 21992
rect 4434 49680 4490 49736
rect 4802 20712 4858 20768
rect 7616 76186 7672 76188
rect 7696 76186 7752 76188
rect 7776 76186 7832 76188
rect 7856 76186 7912 76188
rect 7616 76134 7662 76186
rect 7662 76134 7672 76186
rect 7696 76134 7726 76186
rect 7726 76134 7738 76186
rect 7738 76134 7752 76186
rect 7776 76134 7790 76186
rect 7790 76134 7802 76186
rect 7802 76134 7832 76186
rect 7856 76134 7866 76186
rect 7866 76134 7912 76186
rect 7616 76132 7672 76134
rect 7696 76132 7752 76134
rect 7776 76132 7832 76134
rect 7856 76132 7912 76134
rect 7562 75964 7564 75984
rect 7564 75964 7616 75984
rect 7616 75964 7618 75984
rect 7562 75928 7618 75964
rect 6550 75148 6552 75168
rect 6552 75148 6604 75168
rect 6604 75148 6606 75168
rect 6550 75112 6606 75148
rect 1956 4922 2012 4924
rect 2036 4922 2092 4924
rect 2116 4922 2172 4924
rect 2196 4922 2252 4924
rect 1956 4870 2002 4922
rect 2002 4870 2012 4922
rect 2036 4870 2066 4922
rect 2066 4870 2078 4922
rect 2078 4870 2092 4922
rect 2116 4870 2130 4922
rect 2130 4870 2142 4922
rect 2142 4870 2172 4922
rect 2196 4870 2206 4922
rect 2206 4870 2252 4922
rect 1956 4868 2012 4870
rect 2036 4868 2092 4870
rect 2116 4868 2172 4870
rect 2196 4868 2252 4870
rect 1956 3834 2012 3836
rect 2036 3834 2092 3836
rect 2116 3834 2172 3836
rect 2196 3834 2252 3836
rect 1956 3782 2002 3834
rect 2002 3782 2012 3834
rect 2036 3782 2066 3834
rect 2066 3782 2078 3834
rect 2078 3782 2092 3834
rect 2116 3782 2130 3834
rect 2130 3782 2142 3834
rect 2142 3782 2172 3834
rect 2196 3782 2206 3834
rect 2206 3782 2252 3834
rect 1956 3780 2012 3782
rect 2036 3780 2092 3782
rect 2116 3780 2172 3782
rect 2196 3780 2252 3782
rect 2616 5466 2672 5468
rect 2696 5466 2752 5468
rect 2776 5466 2832 5468
rect 2856 5466 2912 5468
rect 2616 5414 2662 5466
rect 2662 5414 2672 5466
rect 2696 5414 2726 5466
rect 2726 5414 2738 5466
rect 2738 5414 2752 5466
rect 2776 5414 2790 5466
rect 2790 5414 2802 5466
rect 2802 5414 2832 5466
rect 2856 5414 2866 5466
rect 2866 5414 2912 5466
rect 2616 5412 2672 5414
rect 2696 5412 2752 5414
rect 2776 5412 2832 5414
rect 2856 5412 2912 5414
rect 2616 4378 2672 4380
rect 2696 4378 2752 4380
rect 2776 4378 2832 4380
rect 2856 4378 2912 4380
rect 2616 4326 2662 4378
rect 2662 4326 2672 4378
rect 2696 4326 2726 4378
rect 2726 4326 2738 4378
rect 2738 4326 2752 4378
rect 2776 4326 2790 4378
rect 2790 4326 2802 4378
rect 2802 4326 2832 4378
rect 2856 4326 2866 4378
rect 2866 4326 2912 4378
rect 2616 4324 2672 4326
rect 2696 4324 2752 4326
rect 2776 4324 2832 4326
rect 2856 4324 2912 4326
rect 2616 3290 2672 3292
rect 2696 3290 2752 3292
rect 2776 3290 2832 3292
rect 2856 3290 2912 3292
rect 2616 3238 2662 3290
rect 2662 3238 2672 3290
rect 2696 3238 2726 3290
rect 2726 3238 2738 3290
rect 2738 3238 2752 3290
rect 2776 3238 2790 3290
rect 2790 3238 2802 3290
rect 2802 3238 2832 3290
rect 2856 3238 2866 3290
rect 2866 3238 2912 3290
rect 2616 3236 2672 3238
rect 2696 3236 2752 3238
rect 2776 3236 2832 3238
rect 2856 3236 2912 3238
rect 6956 75642 7012 75644
rect 7036 75642 7092 75644
rect 7116 75642 7172 75644
rect 7196 75642 7252 75644
rect 6956 75590 7002 75642
rect 7002 75590 7012 75642
rect 7036 75590 7066 75642
rect 7066 75590 7078 75642
rect 7078 75590 7092 75642
rect 7116 75590 7130 75642
rect 7130 75590 7142 75642
rect 7142 75590 7172 75642
rect 7196 75590 7206 75642
rect 7206 75590 7252 75642
rect 6956 75588 7012 75590
rect 7036 75588 7092 75590
rect 7116 75588 7172 75590
rect 7196 75588 7252 75590
rect 6956 74554 7012 74556
rect 7036 74554 7092 74556
rect 7116 74554 7172 74556
rect 7196 74554 7252 74556
rect 6956 74502 7002 74554
rect 7002 74502 7012 74554
rect 7036 74502 7066 74554
rect 7066 74502 7078 74554
rect 7078 74502 7092 74554
rect 7116 74502 7130 74554
rect 7130 74502 7142 74554
rect 7142 74502 7172 74554
rect 7196 74502 7206 74554
rect 7206 74502 7252 74554
rect 6956 74500 7012 74502
rect 7036 74500 7092 74502
rect 7116 74500 7172 74502
rect 7196 74500 7252 74502
rect 7616 75098 7672 75100
rect 7696 75098 7752 75100
rect 7776 75098 7832 75100
rect 7856 75098 7912 75100
rect 7616 75046 7662 75098
rect 7662 75046 7672 75098
rect 7696 75046 7726 75098
rect 7726 75046 7738 75098
rect 7738 75046 7752 75098
rect 7776 75046 7790 75098
rect 7790 75046 7802 75098
rect 7802 75046 7832 75098
rect 7856 75046 7866 75098
rect 7866 75046 7912 75098
rect 7616 75044 7672 75046
rect 7696 75044 7752 75046
rect 7776 75044 7832 75046
rect 7856 75044 7912 75046
rect 7616 74010 7672 74012
rect 7696 74010 7752 74012
rect 7776 74010 7832 74012
rect 7856 74010 7912 74012
rect 7616 73958 7662 74010
rect 7662 73958 7672 74010
rect 7696 73958 7726 74010
rect 7726 73958 7738 74010
rect 7738 73958 7752 74010
rect 7776 73958 7790 74010
rect 7790 73958 7802 74010
rect 7802 73958 7832 74010
rect 7856 73958 7866 74010
rect 7866 73958 7912 74010
rect 7616 73956 7672 73958
rect 7696 73956 7752 73958
rect 7776 73956 7832 73958
rect 7856 73956 7912 73958
rect 6956 73466 7012 73468
rect 7036 73466 7092 73468
rect 7116 73466 7172 73468
rect 7196 73466 7252 73468
rect 6956 73414 7002 73466
rect 7002 73414 7012 73466
rect 7036 73414 7066 73466
rect 7066 73414 7078 73466
rect 7078 73414 7092 73466
rect 7116 73414 7130 73466
rect 7130 73414 7142 73466
rect 7142 73414 7172 73466
rect 7196 73414 7206 73466
rect 7206 73414 7252 73466
rect 6956 73412 7012 73414
rect 7036 73412 7092 73414
rect 7116 73412 7172 73414
rect 7196 73412 7252 73414
rect 7616 72922 7672 72924
rect 7696 72922 7752 72924
rect 7776 72922 7832 72924
rect 7856 72922 7912 72924
rect 7616 72870 7662 72922
rect 7662 72870 7672 72922
rect 7696 72870 7726 72922
rect 7726 72870 7738 72922
rect 7738 72870 7752 72922
rect 7776 72870 7790 72922
rect 7790 72870 7802 72922
rect 7802 72870 7832 72922
rect 7856 72870 7866 72922
rect 7866 72870 7912 72922
rect 7616 72868 7672 72870
rect 7696 72868 7752 72870
rect 7776 72868 7832 72870
rect 7856 72868 7912 72870
rect 6956 72378 7012 72380
rect 7036 72378 7092 72380
rect 7116 72378 7172 72380
rect 7196 72378 7252 72380
rect 6956 72326 7002 72378
rect 7002 72326 7012 72378
rect 7036 72326 7066 72378
rect 7066 72326 7078 72378
rect 7078 72326 7092 72378
rect 7116 72326 7130 72378
rect 7130 72326 7142 72378
rect 7142 72326 7172 72378
rect 7196 72326 7206 72378
rect 7206 72326 7252 72378
rect 6956 72324 7012 72326
rect 7036 72324 7092 72326
rect 7116 72324 7172 72326
rect 7196 72324 7252 72326
rect 6956 71290 7012 71292
rect 7036 71290 7092 71292
rect 7116 71290 7172 71292
rect 7196 71290 7252 71292
rect 6956 71238 7002 71290
rect 7002 71238 7012 71290
rect 7036 71238 7066 71290
rect 7066 71238 7078 71290
rect 7078 71238 7092 71290
rect 7116 71238 7130 71290
rect 7130 71238 7142 71290
rect 7142 71238 7172 71290
rect 7196 71238 7206 71290
rect 7206 71238 7252 71290
rect 6956 71236 7012 71238
rect 7036 71236 7092 71238
rect 7116 71236 7172 71238
rect 7196 71236 7252 71238
rect 6956 70202 7012 70204
rect 7036 70202 7092 70204
rect 7116 70202 7172 70204
rect 7196 70202 7252 70204
rect 6956 70150 7002 70202
rect 7002 70150 7012 70202
rect 7036 70150 7066 70202
rect 7066 70150 7078 70202
rect 7078 70150 7092 70202
rect 7116 70150 7130 70202
rect 7130 70150 7142 70202
rect 7142 70150 7172 70202
rect 7196 70150 7206 70202
rect 7206 70150 7252 70202
rect 6956 70148 7012 70150
rect 7036 70148 7092 70150
rect 7116 70148 7172 70150
rect 7196 70148 7252 70150
rect 6956 69114 7012 69116
rect 7036 69114 7092 69116
rect 7116 69114 7172 69116
rect 7196 69114 7252 69116
rect 6956 69062 7002 69114
rect 7002 69062 7012 69114
rect 7036 69062 7066 69114
rect 7066 69062 7078 69114
rect 7078 69062 7092 69114
rect 7116 69062 7130 69114
rect 7130 69062 7142 69114
rect 7142 69062 7172 69114
rect 7196 69062 7206 69114
rect 7206 69062 7252 69114
rect 6956 69060 7012 69062
rect 7036 69060 7092 69062
rect 7116 69060 7172 69062
rect 7196 69060 7252 69062
rect 6956 68026 7012 68028
rect 7036 68026 7092 68028
rect 7116 68026 7172 68028
rect 7196 68026 7252 68028
rect 6956 67974 7002 68026
rect 7002 67974 7012 68026
rect 7036 67974 7066 68026
rect 7066 67974 7078 68026
rect 7078 67974 7092 68026
rect 7116 67974 7130 68026
rect 7130 67974 7142 68026
rect 7142 67974 7172 68026
rect 7196 67974 7206 68026
rect 7206 67974 7252 68026
rect 6956 67972 7012 67974
rect 7036 67972 7092 67974
rect 7116 67972 7172 67974
rect 7196 67972 7252 67974
rect 6956 66938 7012 66940
rect 7036 66938 7092 66940
rect 7116 66938 7172 66940
rect 7196 66938 7252 66940
rect 6956 66886 7002 66938
rect 7002 66886 7012 66938
rect 7036 66886 7066 66938
rect 7066 66886 7078 66938
rect 7078 66886 7092 66938
rect 7116 66886 7130 66938
rect 7130 66886 7142 66938
rect 7142 66886 7172 66938
rect 7196 66886 7206 66938
rect 7206 66886 7252 66938
rect 6956 66884 7012 66886
rect 7036 66884 7092 66886
rect 7116 66884 7172 66886
rect 7196 66884 7252 66886
rect 6956 65850 7012 65852
rect 7036 65850 7092 65852
rect 7116 65850 7172 65852
rect 7196 65850 7252 65852
rect 6956 65798 7002 65850
rect 7002 65798 7012 65850
rect 7036 65798 7066 65850
rect 7066 65798 7078 65850
rect 7078 65798 7092 65850
rect 7116 65798 7130 65850
rect 7130 65798 7142 65850
rect 7142 65798 7172 65850
rect 7196 65798 7206 65850
rect 7206 65798 7252 65850
rect 6956 65796 7012 65798
rect 7036 65796 7092 65798
rect 7116 65796 7172 65798
rect 7196 65796 7252 65798
rect 6956 64762 7012 64764
rect 7036 64762 7092 64764
rect 7116 64762 7172 64764
rect 7196 64762 7252 64764
rect 6956 64710 7002 64762
rect 7002 64710 7012 64762
rect 7036 64710 7066 64762
rect 7066 64710 7078 64762
rect 7078 64710 7092 64762
rect 7116 64710 7130 64762
rect 7130 64710 7142 64762
rect 7142 64710 7172 64762
rect 7196 64710 7206 64762
rect 7206 64710 7252 64762
rect 6956 64708 7012 64710
rect 7036 64708 7092 64710
rect 7116 64708 7172 64710
rect 7196 64708 7252 64710
rect 6956 63674 7012 63676
rect 7036 63674 7092 63676
rect 7116 63674 7172 63676
rect 7196 63674 7252 63676
rect 6956 63622 7002 63674
rect 7002 63622 7012 63674
rect 7036 63622 7066 63674
rect 7066 63622 7078 63674
rect 7078 63622 7092 63674
rect 7116 63622 7130 63674
rect 7130 63622 7142 63674
rect 7142 63622 7172 63674
rect 7196 63622 7206 63674
rect 7206 63622 7252 63674
rect 6956 63620 7012 63622
rect 7036 63620 7092 63622
rect 7116 63620 7172 63622
rect 7196 63620 7252 63622
rect 6956 62586 7012 62588
rect 7036 62586 7092 62588
rect 7116 62586 7172 62588
rect 7196 62586 7252 62588
rect 6956 62534 7002 62586
rect 7002 62534 7012 62586
rect 7036 62534 7066 62586
rect 7066 62534 7078 62586
rect 7078 62534 7092 62586
rect 7116 62534 7130 62586
rect 7130 62534 7142 62586
rect 7142 62534 7172 62586
rect 7196 62534 7206 62586
rect 7206 62534 7252 62586
rect 6956 62532 7012 62534
rect 7036 62532 7092 62534
rect 7116 62532 7172 62534
rect 7196 62532 7252 62534
rect 6956 61498 7012 61500
rect 7036 61498 7092 61500
rect 7116 61498 7172 61500
rect 7196 61498 7252 61500
rect 6956 61446 7002 61498
rect 7002 61446 7012 61498
rect 7036 61446 7066 61498
rect 7066 61446 7078 61498
rect 7078 61446 7092 61498
rect 7116 61446 7130 61498
rect 7130 61446 7142 61498
rect 7142 61446 7172 61498
rect 7196 61446 7206 61498
rect 7206 61446 7252 61498
rect 6956 61444 7012 61446
rect 7036 61444 7092 61446
rect 7116 61444 7172 61446
rect 7196 61444 7252 61446
rect 6956 60410 7012 60412
rect 7036 60410 7092 60412
rect 7116 60410 7172 60412
rect 7196 60410 7252 60412
rect 6956 60358 7002 60410
rect 7002 60358 7012 60410
rect 7036 60358 7066 60410
rect 7066 60358 7078 60410
rect 7078 60358 7092 60410
rect 7116 60358 7130 60410
rect 7130 60358 7142 60410
rect 7142 60358 7172 60410
rect 7196 60358 7206 60410
rect 7206 60358 7252 60410
rect 6956 60356 7012 60358
rect 7036 60356 7092 60358
rect 7116 60356 7172 60358
rect 7196 60356 7252 60358
rect 6956 59322 7012 59324
rect 7036 59322 7092 59324
rect 7116 59322 7172 59324
rect 7196 59322 7252 59324
rect 6956 59270 7002 59322
rect 7002 59270 7012 59322
rect 7036 59270 7066 59322
rect 7066 59270 7078 59322
rect 7078 59270 7092 59322
rect 7116 59270 7130 59322
rect 7130 59270 7142 59322
rect 7142 59270 7172 59322
rect 7196 59270 7206 59322
rect 7206 59270 7252 59322
rect 6956 59268 7012 59270
rect 7036 59268 7092 59270
rect 7116 59268 7172 59270
rect 7196 59268 7252 59270
rect 6956 58234 7012 58236
rect 7036 58234 7092 58236
rect 7116 58234 7172 58236
rect 7196 58234 7252 58236
rect 6956 58182 7002 58234
rect 7002 58182 7012 58234
rect 7036 58182 7066 58234
rect 7066 58182 7078 58234
rect 7078 58182 7092 58234
rect 7116 58182 7130 58234
rect 7130 58182 7142 58234
rect 7142 58182 7172 58234
rect 7196 58182 7206 58234
rect 7206 58182 7252 58234
rect 6956 58180 7012 58182
rect 7036 58180 7092 58182
rect 7116 58180 7172 58182
rect 7196 58180 7252 58182
rect 6956 57146 7012 57148
rect 7036 57146 7092 57148
rect 7116 57146 7172 57148
rect 7196 57146 7252 57148
rect 6956 57094 7002 57146
rect 7002 57094 7012 57146
rect 7036 57094 7066 57146
rect 7066 57094 7078 57146
rect 7078 57094 7092 57146
rect 7116 57094 7130 57146
rect 7130 57094 7142 57146
rect 7142 57094 7172 57146
rect 7196 57094 7206 57146
rect 7206 57094 7252 57146
rect 6956 57092 7012 57094
rect 7036 57092 7092 57094
rect 7116 57092 7172 57094
rect 7196 57092 7252 57094
rect 6956 56058 7012 56060
rect 7036 56058 7092 56060
rect 7116 56058 7172 56060
rect 7196 56058 7252 56060
rect 6956 56006 7002 56058
rect 7002 56006 7012 56058
rect 7036 56006 7066 56058
rect 7066 56006 7078 56058
rect 7078 56006 7092 56058
rect 7116 56006 7130 56058
rect 7130 56006 7142 56058
rect 7142 56006 7172 56058
rect 7196 56006 7206 56058
rect 7206 56006 7252 56058
rect 6956 56004 7012 56006
rect 7036 56004 7092 56006
rect 7116 56004 7172 56006
rect 7196 56004 7252 56006
rect 6956 54970 7012 54972
rect 7036 54970 7092 54972
rect 7116 54970 7172 54972
rect 7196 54970 7252 54972
rect 6956 54918 7002 54970
rect 7002 54918 7012 54970
rect 7036 54918 7066 54970
rect 7066 54918 7078 54970
rect 7078 54918 7092 54970
rect 7116 54918 7130 54970
rect 7130 54918 7142 54970
rect 7142 54918 7172 54970
rect 7196 54918 7206 54970
rect 7206 54918 7252 54970
rect 6956 54916 7012 54918
rect 7036 54916 7092 54918
rect 7116 54916 7172 54918
rect 7196 54916 7252 54918
rect 6956 53882 7012 53884
rect 7036 53882 7092 53884
rect 7116 53882 7172 53884
rect 7196 53882 7252 53884
rect 6956 53830 7002 53882
rect 7002 53830 7012 53882
rect 7036 53830 7066 53882
rect 7066 53830 7078 53882
rect 7078 53830 7092 53882
rect 7116 53830 7130 53882
rect 7130 53830 7142 53882
rect 7142 53830 7172 53882
rect 7196 53830 7206 53882
rect 7206 53830 7252 53882
rect 6956 53828 7012 53830
rect 7036 53828 7092 53830
rect 7116 53828 7172 53830
rect 7196 53828 7252 53830
rect 6956 52794 7012 52796
rect 7036 52794 7092 52796
rect 7116 52794 7172 52796
rect 7196 52794 7252 52796
rect 6956 52742 7002 52794
rect 7002 52742 7012 52794
rect 7036 52742 7066 52794
rect 7066 52742 7078 52794
rect 7078 52742 7092 52794
rect 7116 52742 7130 52794
rect 7130 52742 7142 52794
rect 7142 52742 7172 52794
rect 7196 52742 7206 52794
rect 7206 52742 7252 52794
rect 6956 52740 7012 52742
rect 7036 52740 7092 52742
rect 7116 52740 7172 52742
rect 7196 52740 7252 52742
rect 6956 51706 7012 51708
rect 7036 51706 7092 51708
rect 7116 51706 7172 51708
rect 7196 51706 7252 51708
rect 6956 51654 7002 51706
rect 7002 51654 7012 51706
rect 7036 51654 7066 51706
rect 7066 51654 7078 51706
rect 7078 51654 7092 51706
rect 7116 51654 7130 51706
rect 7130 51654 7142 51706
rect 7142 51654 7172 51706
rect 7196 51654 7206 51706
rect 7206 51654 7252 51706
rect 6956 51652 7012 51654
rect 7036 51652 7092 51654
rect 7116 51652 7172 51654
rect 7196 51652 7252 51654
rect 6734 42880 6790 42936
rect 6918 50768 6974 50824
rect 6956 50618 7012 50620
rect 7036 50618 7092 50620
rect 7116 50618 7172 50620
rect 7196 50618 7252 50620
rect 6956 50566 7002 50618
rect 7002 50566 7012 50618
rect 7036 50566 7066 50618
rect 7066 50566 7078 50618
rect 7078 50566 7092 50618
rect 7116 50566 7130 50618
rect 7130 50566 7142 50618
rect 7142 50566 7172 50618
rect 7196 50566 7206 50618
rect 7206 50566 7252 50618
rect 6956 50564 7012 50566
rect 7036 50564 7092 50566
rect 7116 50564 7172 50566
rect 7196 50564 7252 50566
rect 6956 49530 7012 49532
rect 7036 49530 7092 49532
rect 7116 49530 7172 49532
rect 7196 49530 7252 49532
rect 6956 49478 7002 49530
rect 7002 49478 7012 49530
rect 7036 49478 7066 49530
rect 7066 49478 7078 49530
rect 7078 49478 7092 49530
rect 7116 49478 7130 49530
rect 7130 49478 7142 49530
rect 7142 49478 7172 49530
rect 7196 49478 7206 49530
rect 7206 49478 7252 49530
rect 6956 49476 7012 49478
rect 7036 49476 7092 49478
rect 7116 49476 7172 49478
rect 7196 49476 7252 49478
rect 6956 48442 7012 48444
rect 7036 48442 7092 48444
rect 7116 48442 7172 48444
rect 7196 48442 7252 48444
rect 6956 48390 7002 48442
rect 7002 48390 7012 48442
rect 7036 48390 7066 48442
rect 7066 48390 7078 48442
rect 7078 48390 7092 48442
rect 7116 48390 7130 48442
rect 7130 48390 7142 48442
rect 7142 48390 7172 48442
rect 7196 48390 7206 48442
rect 7206 48390 7252 48442
rect 6956 48388 7012 48390
rect 7036 48388 7092 48390
rect 7116 48388 7172 48390
rect 7196 48388 7252 48390
rect 6956 47354 7012 47356
rect 7036 47354 7092 47356
rect 7116 47354 7172 47356
rect 7196 47354 7252 47356
rect 6956 47302 7002 47354
rect 7002 47302 7012 47354
rect 7036 47302 7066 47354
rect 7066 47302 7078 47354
rect 7078 47302 7092 47354
rect 7116 47302 7130 47354
rect 7130 47302 7142 47354
rect 7142 47302 7172 47354
rect 7196 47302 7206 47354
rect 7206 47302 7252 47354
rect 6956 47300 7012 47302
rect 7036 47300 7092 47302
rect 7116 47300 7172 47302
rect 7196 47300 7252 47302
rect 6956 46266 7012 46268
rect 7036 46266 7092 46268
rect 7116 46266 7172 46268
rect 7196 46266 7252 46268
rect 6956 46214 7002 46266
rect 7002 46214 7012 46266
rect 7036 46214 7066 46266
rect 7066 46214 7078 46266
rect 7078 46214 7092 46266
rect 7116 46214 7130 46266
rect 7130 46214 7142 46266
rect 7142 46214 7172 46266
rect 7196 46214 7206 46266
rect 7206 46214 7252 46266
rect 6956 46212 7012 46214
rect 7036 46212 7092 46214
rect 7116 46212 7172 46214
rect 7196 46212 7252 46214
rect 7616 71834 7672 71836
rect 7696 71834 7752 71836
rect 7776 71834 7832 71836
rect 7856 71834 7912 71836
rect 7616 71782 7662 71834
rect 7662 71782 7672 71834
rect 7696 71782 7726 71834
rect 7726 71782 7738 71834
rect 7738 71782 7752 71834
rect 7776 71782 7790 71834
rect 7790 71782 7802 71834
rect 7802 71782 7832 71834
rect 7856 71782 7866 71834
rect 7866 71782 7912 71834
rect 7616 71780 7672 71782
rect 7696 71780 7752 71782
rect 7776 71780 7832 71782
rect 7856 71780 7912 71782
rect 7616 70746 7672 70748
rect 7696 70746 7752 70748
rect 7776 70746 7832 70748
rect 7856 70746 7912 70748
rect 7616 70694 7662 70746
rect 7662 70694 7672 70746
rect 7696 70694 7726 70746
rect 7726 70694 7738 70746
rect 7738 70694 7752 70746
rect 7776 70694 7790 70746
rect 7790 70694 7802 70746
rect 7802 70694 7832 70746
rect 7856 70694 7866 70746
rect 7866 70694 7912 70746
rect 7616 70692 7672 70694
rect 7696 70692 7752 70694
rect 7776 70692 7832 70694
rect 7856 70692 7912 70694
rect 7616 69658 7672 69660
rect 7696 69658 7752 69660
rect 7776 69658 7832 69660
rect 7856 69658 7912 69660
rect 7616 69606 7662 69658
rect 7662 69606 7672 69658
rect 7696 69606 7726 69658
rect 7726 69606 7738 69658
rect 7738 69606 7752 69658
rect 7776 69606 7790 69658
rect 7790 69606 7802 69658
rect 7802 69606 7832 69658
rect 7856 69606 7866 69658
rect 7866 69606 7912 69658
rect 7616 69604 7672 69606
rect 7696 69604 7752 69606
rect 7776 69604 7832 69606
rect 7856 69604 7912 69606
rect 7616 68570 7672 68572
rect 7696 68570 7752 68572
rect 7776 68570 7832 68572
rect 7856 68570 7912 68572
rect 7616 68518 7662 68570
rect 7662 68518 7672 68570
rect 7696 68518 7726 68570
rect 7726 68518 7738 68570
rect 7738 68518 7752 68570
rect 7776 68518 7790 68570
rect 7790 68518 7802 68570
rect 7802 68518 7832 68570
rect 7856 68518 7866 68570
rect 7866 68518 7912 68570
rect 7616 68516 7672 68518
rect 7696 68516 7752 68518
rect 7776 68516 7832 68518
rect 7856 68516 7912 68518
rect 7616 67482 7672 67484
rect 7696 67482 7752 67484
rect 7776 67482 7832 67484
rect 7856 67482 7912 67484
rect 7616 67430 7662 67482
rect 7662 67430 7672 67482
rect 7696 67430 7726 67482
rect 7726 67430 7738 67482
rect 7738 67430 7752 67482
rect 7776 67430 7790 67482
rect 7790 67430 7802 67482
rect 7802 67430 7832 67482
rect 7856 67430 7866 67482
rect 7866 67430 7912 67482
rect 7616 67428 7672 67430
rect 7696 67428 7752 67430
rect 7776 67428 7832 67430
rect 7856 67428 7912 67430
rect 7616 66394 7672 66396
rect 7696 66394 7752 66396
rect 7776 66394 7832 66396
rect 7856 66394 7912 66396
rect 7616 66342 7662 66394
rect 7662 66342 7672 66394
rect 7696 66342 7726 66394
rect 7726 66342 7738 66394
rect 7738 66342 7752 66394
rect 7776 66342 7790 66394
rect 7790 66342 7802 66394
rect 7802 66342 7832 66394
rect 7856 66342 7866 66394
rect 7866 66342 7912 66394
rect 7616 66340 7672 66342
rect 7696 66340 7752 66342
rect 7776 66340 7832 66342
rect 7856 66340 7912 66342
rect 7616 65306 7672 65308
rect 7696 65306 7752 65308
rect 7776 65306 7832 65308
rect 7856 65306 7912 65308
rect 7616 65254 7662 65306
rect 7662 65254 7672 65306
rect 7696 65254 7726 65306
rect 7726 65254 7738 65306
rect 7738 65254 7752 65306
rect 7776 65254 7790 65306
rect 7790 65254 7802 65306
rect 7802 65254 7832 65306
rect 7856 65254 7866 65306
rect 7866 65254 7912 65306
rect 7616 65252 7672 65254
rect 7696 65252 7752 65254
rect 7776 65252 7832 65254
rect 7856 65252 7912 65254
rect 7616 64218 7672 64220
rect 7696 64218 7752 64220
rect 7776 64218 7832 64220
rect 7856 64218 7912 64220
rect 7616 64166 7662 64218
rect 7662 64166 7672 64218
rect 7696 64166 7726 64218
rect 7726 64166 7738 64218
rect 7738 64166 7752 64218
rect 7776 64166 7790 64218
rect 7790 64166 7802 64218
rect 7802 64166 7832 64218
rect 7856 64166 7866 64218
rect 7866 64166 7912 64218
rect 7616 64164 7672 64166
rect 7696 64164 7752 64166
rect 7776 64164 7832 64166
rect 7856 64164 7912 64166
rect 7616 63130 7672 63132
rect 7696 63130 7752 63132
rect 7776 63130 7832 63132
rect 7856 63130 7912 63132
rect 7616 63078 7662 63130
rect 7662 63078 7672 63130
rect 7696 63078 7726 63130
rect 7726 63078 7738 63130
rect 7738 63078 7752 63130
rect 7776 63078 7790 63130
rect 7790 63078 7802 63130
rect 7802 63078 7832 63130
rect 7856 63078 7866 63130
rect 7866 63078 7912 63130
rect 7616 63076 7672 63078
rect 7696 63076 7752 63078
rect 7776 63076 7832 63078
rect 7856 63076 7912 63078
rect 7616 62042 7672 62044
rect 7696 62042 7752 62044
rect 7776 62042 7832 62044
rect 7856 62042 7912 62044
rect 7616 61990 7662 62042
rect 7662 61990 7672 62042
rect 7696 61990 7726 62042
rect 7726 61990 7738 62042
rect 7738 61990 7752 62042
rect 7776 61990 7790 62042
rect 7790 61990 7802 62042
rect 7802 61990 7832 62042
rect 7856 61990 7866 62042
rect 7866 61990 7912 62042
rect 7616 61988 7672 61990
rect 7696 61988 7752 61990
rect 7776 61988 7832 61990
rect 7856 61988 7912 61990
rect 7616 60954 7672 60956
rect 7696 60954 7752 60956
rect 7776 60954 7832 60956
rect 7856 60954 7912 60956
rect 7616 60902 7662 60954
rect 7662 60902 7672 60954
rect 7696 60902 7726 60954
rect 7726 60902 7738 60954
rect 7738 60902 7752 60954
rect 7776 60902 7790 60954
rect 7790 60902 7802 60954
rect 7802 60902 7832 60954
rect 7856 60902 7866 60954
rect 7866 60902 7912 60954
rect 7616 60900 7672 60902
rect 7696 60900 7752 60902
rect 7776 60900 7832 60902
rect 7856 60900 7912 60902
rect 8482 76356 8538 76392
rect 8482 76336 8484 76356
rect 8484 76336 8536 76356
rect 8536 76336 8538 76356
rect 11242 76236 11244 76256
rect 11244 76236 11296 76256
rect 11296 76236 11298 76256
rect 8758 76064 8814 76120
rect 7616 59866 7672 59868
rect 7696 59866 7752 59868
rect 7776 59866 7832 59868
rect 7856 59866 7912 59868
rect 7616 59814 7662 59866
rect 7662 59814 7672 59866
rect 7696 59814 7726 59866
rect 7726 59814 7738 59866
rect 7738 59814 7752 59866
rect 7776 59814 7790 59866
rect 7790 59814 7802 59866
rect 7802 59814 7832 59866
rect 7856 59814 7866 59866
rect 7866 59814 7912 59866
rect 7616 59812 7672 59814
rect 7696 59812 7752 59814
rect 7776 59812 7832 59814
rect 7856 59812 7912 59814
rect 7616 58778 7672 58780
rect 7696 58778 7752 58780
rect 7776 58778 7832 58780
rect 7856 58778 7912 58780
rect 7616 58726 7662 58778
rect 7662 58726 7672 58778
rect 7696 58726 7726 58778
rect 7726 58726 7738 58778
rect 7738 58726 7752 58778
rect 7776 58726 7790 58778
rect 7790 58726 7802 58778
rect 7802 58726 7832 58778
rect 7856 58726 7866 58778
rect 7866 58726 7912 58778
rect 7616 58724 7672 58726
rect 7696 58724 7752 58726
rect 7776 58724 7832 58726
rect 7856 58724 7912 58726
rect 7616 57690 7672 57692
rect 7696 57690 7752 57692
rect 7776 57690 7832 57692
rect 7856 57690 7912 57692
rect 7616 57638 7662 57690
rect 7662 57638 7672 57690
rect 7696 57638 7726 57690
rect 7726 57638 7738 57690
rect 7738 57638 7752 57690
rect 7776 57638 7790 57690
rect 7790 57638 7802 57690
rect 7802 57638 7832 57690
rect 7856 57638 7866 57690
rect 7866 57638 7912 57690
rect 7616 57636 7672 57638
rect 7696 57636 7752 57638
rect 7776 57636 7832 57638
rect 7856 57636 7912 57638
rect 7616 56602 7672 56604
rect 7696 56602 7752 56604
rect 7776 56602 7832 56604
rect 7856 56602 7912 56604
rect 7616 56550 7662 56602
rect 7662 56550 7672 56602
rect 7696 56550 7726 56602
rect 7726 56550 7738 56602
rect 7738 56550 7752 56602
rect 7776 56550 7790 56602
rect 7790 56550 7802 56602
rect 7802 56550 7832 56602
rect 7856 56550 7866 56602
rect 7866 56550 7912 56602
rect 7616 56548 7672 56550
rect 7696 56548 7752 56550
rect 7776 56548 7832 56550
rect 7856 56548 7912 56550
rect 7616 55514 7672 55516
rect 7696 55514 7752 55516
rect 7776 55514 7832 55516
rect 7856 55514 7912 55516
rect 7616 55462 7662 55514
rect 7662 55462 7672 55514
rect 7696 55462 7726 55514
rect 7726 55462 7738 55514
rect 7738 55462 7752 55514
rect 7776 55462 7790 55514
rect 7790 55462 7802 55514
rect 7802 55462 7832 55514
rect 7856 55462 7866 55514
rect 7866 55462 7912 55514
rect 7616 55460 7672 55462
rect 7696 55460 7752 55462
rect 7776 55460 7832 55462
rect 7856 55460 7912 55462
rect 7616 54426 7672 54428
rect 7696 54426 7752 54428
rect 7776 54426 7832 54428
rect 7856 54426 7912 54428
rect 7616 54374 7662 54426
rect 7662 54374 7672 54426
rect 7696 54374 7726 54426
rect 7726 54374 7738 54426
rect 7738 54374 7752 54426
rect 7776 54374 7790 54426
rect 7790 54374 7802 54426
rect 7802 54374 7832 54426
rect 7856 54374 7866 54426
rect 7866 54374 7912 54426
rect 7616 54372 7672 54374
rect 7696 54372 7752 54374
rect 7776 54372 7832 54374
rect 7856 54372 7912 54374
rect 7616 53338 7672 53340
rect 7696 53338 7752 53340
rect 7776 53338 7832 53340
rect 7856 53338 7912 53340
rect 7616 53286 7662 53338
rect 7662 53286 7672 53338
rect 7696 53286 7726 53338
rect 7726 53286 7738 53338
rect 7738 53286 7752 53338
rect 7776 53286 7790 53338
rect 7790 53286 7802 53338
rect 7802 53286 7832 53338
rect 7856 53286 7866 53338
rect 7866 53286 7912 53338
rect 7616 53284 7672 53286
rect 7696 53284 7752 53286
rect 7776 53284 7832 53286
rect 7856 53284 7912 53286
rect 8114 59880 8170 59936
rect 7616 52250 7672 52252
rect 7696 52250 7752 52252
rect 7776 52250 7832 52252
rect 7856 52250 7912 52252
rect 7616 52198 7662 52250
rect 7662 52198 7672 52250
rect 7696 52198 7726 52250
rect 7726 52198 7738 52250
rect 7738 52198 7752 52250
rect 7776 52198 7790 52250
rect 7790 52198 7802 52250
rect 7802 52198 7832 52250
rect 7856 52198 7866 52250
rect 7866 52198 7912 52250
rect 7616 52196 7672 52198
rect 7696 52196 7752 52198
rect 7776 52196 7832 52198
rect 7856 52196 7912 52198
rect 7838 51856 7894 51912
rect 7616 51162 7672 51164
rect 7696 51162 7752 51164
rect 7776 51162 7832 51164
rect 7856 51162 7912 51164
rect 7616 51110 7662 51162
rect 7662 51110 7672 51162
rect 7696 51110 7726 51162
rect 7726 51110 7738 51162
rect 7738 51110 7752 51162
rect 7776 51110 7790 51162
rect 7790 51110 7802 51162
rect 7802 51110 7832 51162
rect 7856 51110 7866 51162
rect 7866 51110 7912 51162
rect 7616 51108 7672 51110
rect 7696 51108 7752 51110
rect 7776 51108 7832 51110
rect 7856 51108 7912 51110
rect 7562 50768 7618 50824
rect 7616 50074 7672 50076
rect 7696 50074 7752 50076
rect 7776 50074 7832 50076
rect 7856 50074 7912 50076
rect 7616 50022 7662 50074
rect 7662 50022 7672 50074
rect 7696 50022 7726 50074
rect 7726 50022 7738 50074
rect 7738 50022 7752 50074
rect 7776 50022 7790 50074
rect 7790 50022 7802 50074
rect 7802 50022 7832 50074
rect 7856 50022 7866 50074
rect 7866 50022 7912 50074
rect 7616 50020 7672 50022
rect 7696 50020 7752 50022
rect 7776 50020 7832 50022
rect 7856 50020 7912 50022
rect 7616 48986 7672 48988
rect 7696 48986 7752 48988
rect 7776 48986 7832 48988
rect 7856 48986 7912 48988
rect 7616 48934 7662 48986
rect 7662 48934 7672 48986
rect 7696 48934 7726 48986
rect 7726 48934 7738 48986
rect 7738 48934 7752 48986
rect 7776 48934 7790 48986
rect 7790 48934 7802 48986
rect 7802 48934 7832 48986
rect 7856 48934 7866 48986
rect 7866 48934 7912 48986
rect 7616 48932 7672 48934
rect 7696 48932 7752 48934
rect 7776 48932 7832 48934
rect 7856 48932 7912 48934
rect 7616 47898 7672 47900
rect 7696 47898 7752 47900
rect 7776 47898 7832 47900
rect 7856 47898 7912 47900
rect 7616 47846 7662 47898
rect 7662 47846 7672 47898
rect 7696 47846 7726 47898
rect 7726 47846 7738 47898
rect 7738 47846 7752 47898
rect 7776 47846 7790 47898
rect 7790 47846 7802 47898
rect 7802 47846 7832 47898
rect 7856 47846 7866 47898
rect 7866 47846 7912 47898
rect 7616 47844 7672 47846
rect 7696 47844 7752 47846
rect 7776 47844 7832 47846
rect 7856 47844 7912 47846
rect 6956 45178 7012 45180
rect 7036 45178 7092 45180
rect 7116 45178 7172 45180
rect 7196 45178 7252 45180
rect 6956 45126 7002 45178
rect 7002 45126 7012 45178
rect 7036 45126 7066 45178
rect 7066 45126 7078 45178
rect 7078 45126 7092 45178
rect 7116 45126 7130 45178
rect 7130 45126 7142 45178
rect 7142 45126 7172 45178
rect 7196 45126 7206 45178
rect 7206 45126 7252 45178
rect 6956 45124 7012 45126
rect 7036 45124 7092 45126
rect 7116 45124 7172 45126
rect 7196 45124 7252 45126
rect 6956 44090 7012 44092
rect 7036 44090 7092 44092
rect 7116 44090 7172 44092
rect 7196 44090 7252 44092
rect 6956 44038 7002 44090
rect 7002 44038 7012 44090
rect 7036 44038 7066 44090
rect 7066 44038 7078 44090
rect 7078 44038 7092 44090
rect 7116 44038 7130 44090
rect 7130 44038 7142 44090
rect 7142 44038 7172 44090
rect 7196 44038 7206 44090
rect 7206 44038 7252 44090
rect 6956 44036 7012 44038
rect 7036 44036 7092 44038
rect 7116 44036 7172 44038
rect 7196 44036 7252 44038
rect 6956 43002 7012 43004
rect 7036 43002 7092 43004
rect 7116 43002 7172 43004
rect 7196 43002 7252 43004
rect 6956 42950 7002 43002
rect 7002 42950 7012 43002
rect 7036 42950 7066 43002
rect 7066 42950 7078 43002
rect 7078 42950 7092 43002
rect 7116 42950 7130 43002
rect 7130 42950 7142 43002
rect 7142 42950 7172 43002
rect 7196 42950 7206 43002
rect 7206 42950 7252 43002
rect 6956 42948 7012 42950
rect 7036 42948 7092 42950
rect 7116 42948 7172 42950
rect 7196 42948 7252 42950
rect 6956 41914 7012 41916
rect 7036 41914 7092 41916
rect 7116 41914 7172 41916
rect 7196 41914 7252 41916
rect 6956 41862 7002 41914
rect 7002 41862 7012 41914
rect 7036 41862 7066 41914
rect 7066 41862 7078 41914
rect 7078 41862 7092 41914
rect 7116 41862 7130 41914
rect 7130 41862 7142 41914
rect 7142 41862 7172 41914
rect 7196 41862 7206 41914
rect 7206 41862 7252 41914
rect 6956 41860 7012 41862
rect 7036 41860 7092 41862
rect 7116 41860 7172 41862
rect 7196 41860 7252 41862
rect 6956 40826 7012 40828
rect 7036 40826 7092 40828
rect 7116 40826 7172 40828
rect 7196 40826 7252 40828
rect 6956 40774 7002 40826
rect 7002 40774 7012 40826
rect 7036 40774 7066 40826
rect 7066 40774 7078 40826
rect 7078 40774 7092 40826
rect 7116 40774 7130 40826
rect 7130 40774 7142 40826
rect 7142 40774 7172 40826
rect 7196 40774 7206 40826
rect 7206 40774 7252 40826
rect 6956 40772 7012 40774
rect 7036 40772 7092 40774
rect 7116 40772 7172 40774
rect 7196 40772 7252 40774
rect 7616 46810 7672 46812
rect 7696 46810 7752 46812
rect 7776 46810 7832 46812
rect 7856 46810 7912 46812
rect 7616 46758 7662 46810
rect 7662 46758 7672 46810
rect 7696 46758 7726 46810
rect 7726 46758 7738 46810
rect 7738 46758 7752 46810
rect 7776 46758 7790 46810
rect 7790 46758 7802 46810
rect 7802 46758 7832 46810
rect 7856 46758 7866 46810
rect 7866 46758 7912 46810
rect 7616 46756 7672 46758
rect 7696 46756 7752 46758
rect 7776 46756 7832 46758
rect 7856 46756 7912 46758
rect 7616 45722 7672 45724
rect 7696 45722 7752 45724
rect 7776 45722 7832 45724
rect 7856 45722 7912 45724
rect 7616 45670 7662 45722
rect 7662 45670 7672 45722
rect 7696 45670 7726 45722
rect 7726 45670 7738 45722
rect 7738 45670 7752 45722
rect 7776 45670 7790 45722
rect 7790 45670 7802 45722
rect 7802 45670 7832 45722
rect 7856 45670 7866 45722
rect 7866 45670 7912 45722
rect 7616 45668 7672 45670
rect 7696 45668 7752 45670
rect 7776 45668 7832 45670
rect 7856 45668 7912 45670
rect 7616 44634 7672 44636
rect 7696 44634 7752 44636
rect 7776 44634 7832 44636
rect 7856 44634 7912 44636
rect 7616 44582 7662 44634
rect 7662 44582 7672 44634
rect 7696 44582 7726 44634
rect 7726 44582 7738 44634
rect 7738 44582 7752 44634
rect 7776 44582 7790 44634
rect 7790 44582 7802 44634
rect 7802 44582 7832 44634
rect 7856 44582 7866 44634
rect 7866 44582 7912 44634
rect 7616 44580 7672 44582
rect 7696 44580 7752 44582
rect 7776 44580 7832 44582
rect 7856 44580 7912 44582
rect 7616 43546 7672 43548
rect 7696 43546 7752 43548
rect 7776 43546 7832 43548
rect 7856 43546 7912 43548
rect 7616 43494 7662 43546
rect 7662 43494 7672 43546
rect 7696 43494 7726 43546
rect 7726 43494 7738 43546
rect 7738 43494 7752 43546
rect 7776 43494 7790 43546
rect 7790 43494 7802 43546
rect 7802 43494 7832 43546
rect 7856 43494 7866 43546
rect 7866 43494 7912 43546
rect 7616 43492 7672 43494
rect 7696 43492 7752 43494
rect 7776 43492 7832 43494
rect 7856 43492 7912 43494
rect 7562 43288 7618 43344
rect 7616 42458 7672 42460
rect 7696 42458 7752 42460
rect 7776 42458 7832 42460
rect 7856 42458 7912 42460
rect 7616 42406 7662 42458
rect 7662 42406 7672 42458
rect 7696 42406 7726 42458
rect 7726 42406 7738 42458
rect 7738 42406 7752 42458
rect 7776 42406 7790 42458
rect 7790 42406 7802 42458
rect 7802 42406 7832 42458
rect 7856 42406 7866 42458
rect 7866 42406 7912 42458
rect 7616 42404 7672 42406
rect 7696 42404 7752 42406
rect 7776 42404 7832 42406
rect 7856 42404 7912 42406
rect 6956 39738 7012 39740
rect 7036 39738 7092 39740
rect 7116 39738 7172 39740
rect 7196 39738 7252 39740
rect 6956 39686 7002 39738
rect 7002 39686 7012 39738
rect 7036 39686 7066 39738
rect 7066 39686 7078 39738
rect 7078 39686 7092 39738
rect 7116 39686 7130 39738
rect 7130 39686 7142 39738
rect 7142 39686 7172 39738
rect 7196 39686 7206 39738
rect 7206 39686 7252 39738
rect 6956 39684 7012 39686
rect 7036 39684 7092 39686
rect 7116 39684 7172 39686
rect 7196 39684 7252 39686
rect 6956 38650 7012 38652
rect 7036 38650 7092 38652
rect 7116 38650 7172 38652
rect 7196 38650 7252 38652
rect 6956 38598 7002 38650
rect 7002 38598 7012 38650
rect 7036 38598 7066 38650
rect 7066 38598 7078 38650
rect 7078 38598 7092 38650
rect 7116 38598 7130 38650
rect 7130 38598 7142 38650
rect 7142 38598 7172 38650
rect 7196 38598 7206 38650
rect 7206 38598 7252 38650
rect 6956 38596 7012 38598
rect 7036 38596 7092 38598
rect 7116 38596 7172 38598
rect 7196 38596 7252 38598
rect 6956 37562 7012 37564
rect 7036 37562 7092 37564
rect 7116 37562 7172 37564
rect 7196 37562 7252 37564
rect 6956 37510 7002 37562
rect 7002 37510 7012 37562
rect 7036 37510 7066 37562
rect 7066 37510 7078 37562
rect 7078 37510 7092 37562
rect 7116 37510 7130 37562
rect 7130 37510 7142 37562
rect 7142 37510 7172 37562
rect 7196 37510 7206 37562
rect 7206 37510 7252 37562
rect 6956 37508 7012 37510
rect 7036 37508 7092 37510
rect 7116 37508 7172 37510
rect 7196 37508 7252 37510
rect 6956 36474 7012 36476
rect 7036 36474 7092 36476
rect 7116 36474 7172 36476
rect 7196 36474 7252 36476
rect 6956 36422 7002 36474
rect 7002 36422 7012 36474
rect 7036 36422 7066 36474
rect 7066 36422 7078 36474
rect 7078 36422 7092 36474
rect 7116 36422 7130 36474
rect 7130 36422 7142 36474
rect 7142 36422 7172 36474
rect 7196 36422 7206 36474
rect 7206 36422 7252 36474
rect 6956 36420 7012 36422
rect 7036 36420 7092 36422
rect 7116 36420 7172 36422
rect 7196 36420 7252 36422
rect 6956 35386 7012 35388
rect 7036 35386 7092 35388
rect 7116 35386 7172 35388
rect 7196 35386 7252 35388
rect 6956 35334 7002 35386
rect 7002 35334 7012 35386
rect 7036 35334 7066 35386
rect 7066 35334 7078 35386
rect 7078 35334 7092 35386
rect 7116 35334 7130 35386
rect 7130 35334 7142 35386
rect 7142 35334 7172 35386
rect 7196 35334 7206 35386
rect 7206 35334 7252 35386
rect 6956 35332 7012 35334
rect 7036 35332 7092 35334
rect 7116 35332 7172 35334
rect 7196 35332 7252 35334
rect 6956 34298 7012 34300
rect 7036 34298 7092 34300
rect 7116 34298 7172 34300
rect 7196 34298 7252 34300
rect 6956 34246 7002 34298
rect 7002 34246 7012 34298
rect 7036 34246 7066 34298
rect 7066 34246 7078 34298
rect 7078 34246 7092 34298
rect 7116 34246 7130 34298
rect 7130 34246 7142 34298
rect 7142 34246 7172 34298
rect 7196 34246 7206 34298
rect 7206 34246 7252 34298
rect 6956 34244 7012 34246
rect 7036 34244 7092 34246
rect 7116 34244 7172 34246
rect 7196 34244 7252 34246
rect 6956 33210 7012 33212
rect 7036 33210 7092 33212
rect 7116 33210 7172 33212
rect 7196 33210 7252 33212
rect 6956 33158 7002 33210
rect 7002 33158 7012 33210
rect 7036 33158 7066 33210
rect 7066 33158 7078 33210
rect 7078 33158 7092 33210
rect 7116 33158 7130 33210
rect 7130 33158 7142 33210
rect 7142 33158 7172 33210
rect 7196 33158 7206 33210
rect 7206 33158 7252 33210
rect 6956 33156 7012 33158
rect 7036 33156 7092 33158
rect 7116 33156 7172 33158
rect 7196 33156 7252 33158
rect 6956 32122 7012 32124
rect 7036 32122 7092 32124
rect 7116 32122 7172 32124
rect 7196 32122 7252 32124
rect 6956 32070 7002 32122
rect 7002 32070 7012 32122
rect 7036 32070 7066 32122
rect 7066 32070 7078 32122
rect 7078 32070 7092 32122
rect 7116 32070 7130 32122
rect 7130 32070 7142 32122
rect 7142 32070 7172 32122
rect 7196 32070 7206 32122
rect 7206 32070 7252 32122
rect 6956 32068 7012 32070
rect 7036 32068 7092 32070
rect 7116 32068 7172 32070
rect 7196 32068 7252 32070
rect 7616 41370 7672 41372
rect 7696 41370 7752 41372
rect 7776 41370 7832 41372
rect 7856 41370 7912 41372
rect 7616 41318 7662 41370
rect 7662 41318 7672 41370
rect 7696 41318 7726 41370
rect 7726 41318 7738 41370
rect 7738 41318 7752 41370
rect 7776 41318 7790 41370
rect 7790 41318 7802 41370
rect 7802 41318 7832 41370
rect 7856 41318 7866 41370
rect 7866 41318 7912 41370
rect 7616 41316 7672 41318
rect 7696 41316 7752 41318
rect 7776 41316 7832 41318
rect 7856 41316 7912 41318
rect 7616 40282 7672 40284
rect 7696 40282 7752 40284
rect 7776 40282 7832 40284
rect 7856 40282 7912 40284
rect 7616 40230 7662 40282
rect 7662 40230 7672 40282
rect 7696 40230 7726 40282
rect 7726 40230 7738 40282
rect 7738 40230 7752 40282
rect 7776 40230 7790 40282
rect 7790 40230 7802 40282
rect 7802 40230 7832 40282
rect 7856 40230 7866 40282
rect 7866 40230 7912 40282
rect 7616 40228 7672 40230
rect 7696 40228 7752 40230
rect 7776 40228 7832 40230
rect 7856 40228 7912 40230
rect 7616 39194 7672 39196
rect 7696 39194 7752 39196
rect 7776 39194 7832 39196
rect 7856 39194 7912 39196
rect 7616 39142 7662 39194
rect 7662 39142 7672 39194
rect 7696 39142 7726 39194
rect 7726 39142 7738 39194
rect 7738 39142 7752 39194
rect 7776 39142 7790 39194
rect 7790 39142 7802 39194
rect 7802 39142 7832 39194
rect 7856 39142 7866 39194
rect 7866 39142 7912 39194
rect 7616 39140 7672 39142
rect 7696 39140 7752 39142
rect 7776 39140 7832 39142
rect 7856 39140 7912 39142
rect 7616 38106 7672 38108
rect 7696 38106 7752 38108
rect 7776 38106 7832 38108
rect 7856 38106 7912 38108
rect 7616 38054 7662 38106
rect 7662 38054 7672 38106
rect 7696 38054 7726 38106
rect 7726 38054 7738 38106
rect 7738 38054 7752 38106
rect 7776 38054 7790 38106
rect 7790 38054 7802 38106
rect 7802 38054 7832 38106
rect 7856 38054 7866 38106
rect 7866 38054 7912 38106
rect 7616 38052 7672 38054
rect 7696 38052 7752 38054
rect 7776 38052 7832 38054
rect 7856 38052 7912 38054
rect 7616 37018 7672 37020
rect 7696 37018 7752 37020
rect 7776 37018 7832 37020
rect 7856 37018 7912 37020
rect 7616 36966 7662 37018
rect 7662 36966 7672 37018
rect 7696 36966 7726 37018
rect 7726 36966 7738 37018
rect 7738 36966 7752 37018
rect 7776 36966 7790 37018
rect 7790 36966 7802 37018
rect 7802 36966 7832 37018
rect 7856 36966 7866 37018
rect 7866 36966 7912 37018
rect 7616 36964 7672 36966
rect 7696 36964 7752 36966
rect 7776 36964 7832 36966
rect 7856 36964 7912 36966
rect 7616 35930 7672 35932
rect 7696 35930 7752 35932
rect 7776 35930 7832 35932
rect 7856 35930 7912 35932
rect 7616 35878 7662 35930
rect 7662 35878 7672 35930
rect 7696 35878 7726 35930
rect 7726 35878 7738 35930
rect 7738 35878 7752 35930
rect 7776 35878 7790 35930
rect 7790 35878 7802 35930
rect 7802 35878 7832 35930
rect 7856 35878 7866 35930
rect 7866 35878 7912 35930
rect 7616 35876 7672 35878
rect 7696 35876 7752 35878
rect 7776 35876 7832 35878
rect 7856 35876 7912 35878
rect 7616 34842 7672 34844
rect 7696 34842 7752 34844
rect 7776 34842 7832 34844
rect 7856 34842 7912 34844
rect 7616 34790 7662 34842
rect 7662 34790 7672 34842
rect 7696 34790 7726 34842
rect 7726 34790 7738 34842
rect 7738 34790 7752 34842
rect 7776 34790 7790 34842
rect 7790 34790 7802 34842
rect 7802 34790 7832 34842
rect 7856 34790 7866 34842
rect 7866 34790 7912 34842
rect 7616 34788 7672 34790
rect 7696 34788 7752 34790
rect 7776 34788 7832 34790
rect 7856 34788 7912 34790
rect 7616 33754 7672 33756
rect 7696 33754 7752 33756
rect 7776 33754 7832 33756
rect 7856 33754 7912 33756
rect 7616 33702 7662 33754
rect 7662 33702 7672 33754
rect 7696 33702 7726 33754
rect 7726 33702 7738 33754
rect 7738 33702 7752 33754
rect 7776 33702 7790 33754
rect 7790 33702 7802 33754
rect 7802 33702 7832 33754
rect 7856 33702 7866 33754
rect 7866 33702 7912 33754
rect 7616 33700 7672 33702
rect 7696 33700 7752 33702
rect 7776 33700 7832 33702
rect 7856 33700 7912 33702
rect 7616 32666 7672 32668
rect 7696 32666 7752 32668
rect 7776 32666 7832 32668
rect 7856 32666 7912 32668
rect 7616 32614 7662 32666
rect 7662 32614 7672 32666
rect 7696 32614 7726 32666
rect 7726 32614 7738 32666
rect 7738 32614 7752 32666
rect 7776 32614 7790 32666
rect 7790 32614 7802 32666
rect 7802 32614 7832 32666
rect 7856 32614 7866 32666
rect 7866 32614 7912 32666
rect 7616 32612 7672 32614
rect 7696 32612 7752 32614
rect 7776 32612 7832 32614
rect 7856 32612 7912 32614
rect 6956 31034 7012 31036
rect 7036 31034 7092 31036
rect 7116 31034 7172 31036
rect 7196 31034 7252 31036
rect 6956 30982 7002 31034
rect 7002 30982 7012 31034
rect 7036 30982 7066 31034
rect 7066 30982 7078 31034
rect 7078 30982 7092 31034
rect 7116 30982 7130 31034
rect 7130 30982 7142 31034
rect 7142 30982 7172 31034
rect 7196 30982 7206 31034
rect 7206 30982 7252 31034
rect 6956 30980 7012 30982
rect 7036 30980 7092 30982
rect 7116 30980 7172 30982
rect 7196 30980 7252 30982
rect 6956 29946 7012 29948
rect 7036 29946 7092 29948
rect 7116 29946 7172 29948
rect 7196 29946 7252 29948
rect 6956 29894 7002 29946
rect 7002 29894 7012 29946
rect 7036 29894 7066 29946
rect 7066 29894 7078 29946
rect 7078 29894 7092 29946
rect 7116 29894 7130 29946
rect 7130 29894 7142 29946
rect 7142 29894 7172 29946
rect 7196 29894 7206 29946
rect 7206 29894 7252 29946
rect 6956 29892 7012 29894
rect 7036 29892 7092 29894
rect 7116 29892 7172 29894
rect 7196 29892 7252 29894
rect 6956 28858 7012 28860
rect 7036 28858 7092 28860
rect 7116 28858 7172 28860
rect 7196 28858 7252 28860
rect 6956 28806 7002 28858
rect 7002 28806 7012 28858
rect 7036 28806 7066 28858
rect 7066 28806 7078 28858
rect 7078 28806 7092 28858
rect 7116 28806 7130 28858
rect 7130 28806 7142 28858
rect 7142 28806 7172 28858
rect 7196 28806 7206 28858
rect 7206 28806 7252 28858
rect 6956 28804 7012 28806
rect 7036 28804 7092 28806
rect 7116 28804 7172 28806
rect 7196 28804 7252 28806
rect 6956 27770 7012 27772
rect 7036 27770 7092 27772
rect 7116 27770 7172 27772
rect 7196 27770 7252 27772
rect 6956 27718 7002 27770
rect 7002 27718 7012 27770
rect 7036 27718 7066 27770
rect 7066 27718 7078 27770
rect 7078 27718 7092 27770
rect 7116 27718 7130 27770
rect 7130 27718 7142 27770
rect 7142 27718 7172 27770
rect 7196 27718 7206 27770
rect 7206 27718 7252 27770
rect 6956 27716 7012 27718
rect 7036 27716 7092 27718
rect 7116 27716 7172 27718
rect 7196 27716 7252 27718
rect 6956 26682 7012 26684
rect 7036 26682 7092 26684
rect 7116 26682 7172 26684
rect 7196 26682 7252 26684
rect 6956 26630 7002 26682
rect 7002 26630 7012 26682
rect 7036 26630 7066 26682
rect 7066 26630 7078 26682
rect 7078 26630 7092 26682
rect 7116 26630 7130 26682
rect 7130 26630 7142 26682
rect 7142 26630 7172 26682
rect 7196 26630 7206 26682
rect 7206 26630 7252 26682
rect 6956 26628 7012 26630
rect 7036 26628 7092 26630
rect 7116 26628 7172 26630
rect 7196 26628 7252 26630
rect 6956 25594 7012 25596
rect 7036 25594 7092 25596
rect 7116 25594 7172 25596
rect 7196 25594 7252 25596
rect 6956 25542 7002 25594
rect 7002 25542 7012 25594
rect 7036 25542 7066 25594
rect 7066 25542 7078 25594
rect 7078 25542 7092 25594
rect 7116 25542 7130 25594
rect 7130 25542 7142 25594
rect 7142 25542 7172 25594
rect 7196 25542 7206 25594
rect 7206 25542 7252 25594
rect 6956 25540 7012 25542
rect 7036 25540 7092 25542
rect 7116 25540 7172 25542
rect 7196 25540 7252 25542
rect 6956 24506 7012 24508
rect 7036 24506 7092 24508
rect 7116 24506 7172 24508
rect 7196 24506 7252 24508
rect 6956 24454 7002 24506
rect 7002 24454 7012 24506
rect 7036 24454 7066 24506
rect 7066 24454 7078 24506
rect 7078 24454 7092 24506
rect 7116 24454 7130 24506
rect 7130 24454 7142 24506
rect 7142 24454 7172 24506
rect 7196 24454 7206 24506
rect 7206 24454 7252 24506
rect 6956 24452 7012 24454
rect 7036 24452 7092 24454
rect 7116 24452 7172 24454
rect 7196 24452 7252 24454
rect 6956 23418 7012 23420
rect 7036 23418 7092 23420
rect 7116 23418 7172 23420
rect 7196 23418 7252 23420
rect 6956 23366 7002 23418
rect 7002 23366 7012 23418
rect 7036 23366 7066 23418
rect 7066 23366 7078 23418
rect 7078 23366 7092 23418
rect 7116 23366 7130 23418
rect 7130 23366 7142 23418
rect 7142 23366 7172 23418
rect 7196 23366 7206 23418
rect 7206 23366 7252 23418
rect 6956 23364 7012 23366
rect 7036 23364 7092 23366
rect 7116 23364 7172 23366
rect 7196 23364 7252 23366
rect 6956 22330 7012 22332
rect 7036 22330 7092 22332
rect 7116 22330 7172 22332
rect 7196 22330 7252 22332
rect 6956 22278 7002 22330
rect 7002 22278 7012 22330
rect 7036 22278 7066 22330
rect 7066 22278 7078 22330
rect 7078 22278 7092 22330
rect 7116 22278 7130 22330
rect 7130 22278 7142 22330
rect 7142 22278 7172 22330
rect 7196 22278 7206 22330
rect 7206 22278 7252 22330
rect 6956 22276 7012 22278
rect 7036 22276 7092 22278
rect 7116 22276 7172 22278
rect 7196 22276 7252 22278
rect 6956 21242 7012 21244
rect 7036 21242 7092 21244
rect 7116 21242 7172 21244
rect 7196 21242 7252 21244
rect 6956 21190 7002 21242
rect 7002 21190 7012 21242
rect 7036 21190 7066 21242
rect 7066 21190 7078 21242
rect 7078 21190 7092 21242
rect 7116 21190 7130 21242
rect 7130 21190 7142 21242
rect 7142 21190 7172 21242
rect 7196 21190 7206 21242
rect 7206 21190 7252 21242
rect 6956 21188 7012 21190
rect 7036 21188 7092 21190
rect 7116 21188 7172 21190
rect 7196 21188 7252 21190
rect 6956 20154 7012 20156
rect 7036 20154 7092 20156
rect 7116 20154 7172 20156
rect 7196 20154 7252 20156
rect 6956 20102 7002 20154
rect 7002 20102 7012 20154
rect 7036 20102 7066 20154
rect 7066 20102 7078 20154
rect 7078 20102 7092 20154
rect 7116 20102 7130 20154
rect 7130 20102 7142 20154
rect 7142 20102 7172 20154
rect 7196 20102 7206 20154
rect 7206 20102 7252 20154
rect 6956 20100 7012 20102
rect 7036 20100 7092 20102
rect 7116 20100 7172 20102
rect 7196 20100 7252 20102
rect 6956 19066 7012 19068
rect 7036 19066 7092 19068
rect 7116 19066 7172 19068
rect 7196 19066 7252 19068
rect 6956 19014 7002 19066
rect 7002 19014 7012 19066
rect 7036 19014 7066 19066
rect 7066 19014 7078 19066
rect 7078 19014 7092 19066
rect 7116 19014 7130 19066
rect 7130 19014 7142 19066
rect 7142 19014 7172 19066
rect 7196 19014 7206 19066
rect 7206 19014 7252 19066
rect 6956 19012 7012 19014
rect 7036 19012 7092 19014
rect 7116 19012 7172 19014
rect 7196 19012 7252 19014
rect 6956 17978 7012 17980
rect 7036 17978 7092 17980
rect 7116 17978 7172 17980
rect 7196 17978 7252 17980
rect 6956 17926 7002 17978
rect 7002 17926 7012 17978
rect 7036 17926 7066 17978
rect 7066 17926 7078 17978
rect 7078 17926 7092 17978
rect 7116 17926 7130 17978
rect 7130 17926 7142 17978
rect 7142 17926 7172 17978
rect 7196 17926 7206 17978
rect 7206 17926 7252 17978
rect 6956 17924 7012 17926
rect 7036 17924 7092 17926
rect 7116 17924 7172 17926
rect 7196 17924 7252 17926
rect 6956 16890 7012 16892
rect 7036 16890 7092 16892
rect 7116 16890 7172 16892
rect 7196 16890 7252 16892
rect 6956 16838 7002 16890
rect 7002 16838 7012 16890
rect 7036 16838 7066 16890
rect 7066 16838 7078 16890
rect 7078 16838 7092 16890
rect 7116 16838 7130 16890
rect 7130 16838 7142 16890
rect 7142 16838 7172 16890
rect 7196 16838 7206 16890
rect 7206 16838 7252 16890
rect 6956 16836 7012 16838
rect 7036 16836 7092 16838
rect 7116 16836 7172 16838
rect 7196 16836 7252 16838
rect 6956 15802 7012 15804
rect 7036 15802 7092 15804
rect 7116 15802 7172 15804
rect 7196 15802 7252 15804
rect 6956 15750 7002 15802
rect 7002 15750 7012 15802
rect 7036 15750 7066 15802
rect 7066 15750 7078 15802
rect 7078 15750 7092 15802
rect 7116 15750 7130 15802
rect 7130 15750 7142 15802
rect 7142 15750 7172 15802
rect 7196 15750 7206 15802
rect 7206 15750 7252 15802
rect 6956 15748 7012 15750
rect 7036 15748 7092 15750
rect 7116 15748 7172 15750
rect 7196 15748 7252 15750
rect 6956 14714 7012 14716
rect 7036 14714 7092 14716
rect 7116 14714 7172 14716
rect 7196 14714 7252 14716
rect 6956 14662 7002 14714
rect 7002 14662 7012 14714
rect 7036 14662 7066 14714
rect 7066 14662 7078 14714
rect 7078 14662 7092 14714
rect 7116 14662 7130 14714
rect 7130 14662 7142 14714
rect 7142 14662 7172 14714
rect 7196 14662 7206 14714
rect 7206 14662 7252 14714
rect 6956 14660 7012 14662
rect 7036 14660 7092 14662
rect 7116 14660 7172 14662
rect 7196 14660 7252 14662
rect 6956 13626 7012 13628
rect 7036 13626 7092 13628
rect 7116 13626 7172 13628
rect 7196 13626 7252 13628
rect 6956 13574 7002 13626
rect 7002 13574 7012 13626
rect 7036 13574 7066 13626
rect 7066 13574 7078 13626
rect 7078 13574 7092 13626
rect 7116 13574 7130 13626
rect 7130 13574 7142 13626
rect 7142 13574 7172 13626
rect 7196 13574 7206 13626
rect 7206 13574 7252 13626
rect 6956 13572 7012 13574
rect 7036 13572 7092 13574
rect 7116 13572 7172 13574
rect 7196 13572 7252 13574
rect 6956 12538 7012 12540
rect 7036 12538 7092 12540
rect 7116 12538 7172 12540
rect 7196 12538 7252 12540
rect 6956 12486 7002 12538
rect 7002 12486 7012 12538
rect 7036 12486 7066 12538
rect 7066 12486 7078 12538
rect 7078 12486 7092 12538
rect 7116 12486 7130 12538
rect 7130 12486 7142 12538
rect 7142 12486 7172 12538
rect 7196 12486 7206 12538
rect 7206 12486 7252 12538
rect 6956 12484 7012 12486
rect 7036 12484 7092 12486
rect 7116 12484 7172 12486
rect 7196 12484 7252 12486
rect 6956 11450 7012 11452
rect 7036 11450 7092 11452
rect 7116 11450 7172 11452
rect 7196 11450 7252 11452
rect 6956 11398 7002 11450
rect 7002 11398 7012 11450
rect 7036 11398 7066 11450
rect 7066 11398 7078 11450
rect 7078 11398 7092 11450
rect 7116 11398 7130 11450
rect 7130 11398 7142 11450
rect 7142 11398 7172 11450
rect 7196 11398 7206 11450
rect 7206 11398 7252 11450
rect 6956 11396 7012 11398
rect 7036 11396 7092 11398
rect 7116 11396 7172 11398
rect 7196 11396 7252 11398
rect 6956 10362 7012 10364
rect 7036 10362 7092 10364
rect 7116 10362 7172 10364
rect 7196 10362 7252 10364
rect 6956 10310 7002 10362
rect 7002 10310 7012 10362
rect 7036 10310 7066 10362
rect 7066 10310 7078 10362
rect 7078 10310 7092 10362
rect 7116 10310 7130 10362
rect 7130 10310 7142 10362
rect 7142 10310 7172 10362
rect 7196 10310 7206 10362
rect 7206 10310 7252 10362
rect 6956 10308 7012 10310
rect 7036 10308 7092 10310
rect 7116 10308 7172 10310
rect 7196 10308 7252 10310
rect 7616 31578 7672 31580
rect 7696 31578 7752 31580
rect 7776 31578 7832 31580
rect 7856 31578 7912 31580
rect 7616 31526 7662 31578
rect 7662 31526 7672 31578
rect 7696 31526 7726 31578
rect 7726 31526 7738 31578
rect 7738 31526 7752 31578
rect 7776 31526 7790 31578
rect 7790 31526 7802 31578
rect 7802 31526 7832 31578
rect 7856 31526 7866 31578
rect 7866 31526 7912 31578
rect 7616 31524 7672 31526
rect 7696 31524 7752 31526
rect 7776 31524 7832 31526
rect 7856 31524 7912 31526
rect 8482 32952 8538 33008
rect 7616 30490 7672 30492
rect 7696 30490 7752 30492
rect 7776 30490 7832 30492
rect 7856 30490 7912 30492
rect 7616 30438 7662 30490
rect 7662 30438 7672 30490
rect 7696 30438 7726 30490
rect 7726 30438 7738 30490
rect 7738 30438 7752 30490
rect 7776 30438 7790 30490
rect 7790 30438 7802 30490
rect 7802 30438 7832 30490
rect 7856 30438 7866 30490
rect 7866 30438 7912 30490
rect 7616 30436 7672 30438
rect 7696 30436 7752 30438
rect 7776 30436 7832 30438
rect 7856 30436 7912 30438
rect 7616 29402 7672 29404
rect 7696 29402 7752 29404
rect 7776 29402 7832 29404
rect 7856 29402 7912 29404
rect 7616 29350 7662 29402
rect 7662 29350 7672 29402
rect 7696 29350 7726 29402
rect 7726 29350 7738 29402
rect 7738 29350 7752 29402
rect 7776 29350 7790 29402
rect 7790 29350 7802 29402
rect 7802 29350 7832 29402
rect 7856 29350 7866 29402
rect 7866 29350 7912 29402
rect 7616 29348 7672 29350
rect 7696 29348 7752 29350
rect 7776 29348 7832 29350
rect 7856 29348 7912 29350
rect 7930 28464 7986 28520
rect 7616 28314 7672 28316
rect 7696 28314 7752 28316
rect 7776 28314 7832 28316
rect 7856 28314 7912 28316
rect 7616 28262 7662 28314
rect 7662 28262 7672 28314
rect 7696 28262 7726 28314
rect 7726 28262 7738 28314
rect 7738 28262 7752 28314
rect 7776 28262 7790 28314
rect 7790 28262 7802 28314
rect 7802 28262 7832 28314
rect 7856 28262 7866 28314
rect 7866 28262 7912 28314
rect 7616 28260 7672 28262
rect 7696 28260 7752 28262
rect 7776 28260 7832 28262
rect 7856 28260 7912 28262
rect 7616 27226 7672 27228
rect 7696 27226 7752 27228
rect 7776 27226 7832 27228
rect 7856 27226 7912 27228
rect 7616 27174 7662 27226
rect 7662 27174 7672 27226
rect 7696 27174 7726 27226
rect 7726 27174 7738 27226
rect 7738 27174 7752 27226
rect 7776 27174 7790 27226
rect 7790 27174 7802 27226
rect 7802 27174 7832 27226
rect 7856 27174 7866 27226
rect 7866 27174 7912 27226
rect 7616 27172 7672 27174
rect 7696 27172 7752 27174
rect 7776 27172 7832 27174
rect 7856 27172 7912 27174
rect 8114 26288 8170 26344
rect 7616 26138 7672 26140
rect 7696 26138 7752 26140
rect 7776 26138 7832 26140
rect 7856 26138 7912 26140
rect 7616 26086 7662 26138
rect 7662 26086 7672 26138
rect 7696 26086 7726 26138
rect 7726 26086 7738 26138
rect 7738 26086 7752 26138
rect 7776 26086 7790 26138
rect 7790 26086 7802 26138
rect 7802 26086 7832 26138
rect 7856 26086 7866 26138
rect 7866 26086 7912 26138
rect 7616 26084 7672 26086
rect 7696 26084 7752 26086
rect 7776 26084 7832 26086
rect 7856 26084 7912 26086
rect 8022 26016 8078 26072
rect 7616 25050 7672 25052
rect 7696 25050 7752 25052
rect 7776 25050 7832 25052
rect 7856 25050 7912 25052
rect 7616 24998 7662 25050
rect 7662 24998 7672 25050
rect 7696 24998 7726 25050
rect 7726 24998 7738 25050
rect 7738 24998 7752 25050
rect 7776 24998 7790 25050
rect 7790 24998 7802 25050
rect 7802 24998 7832 25050
rect 7856 24998 7866 25050
rect 7866 24998 7912 25050
rect 7616 24996 7672 24998
rect 7696 24996 7752 24998
rect 7776 24996 7832 24998
rect 7856 24996 7912 24998
rect 7616 23962 7672 23964
rect 7696 23962 7752 23964
rect 7776 23962 7832 23964
rect 7856 23962 7912 23964
rect 7616 23910 7662 23962
rect 7662 23910 7672 23962
rect 7696 23910 7726 23962
rect 7726 23910 7738 23962
rect 7738 23910 7752 23962
rect 7776 23910 7790 23962
rect 7790 23910 7802 23962
rect 7802 23910 7832 23962
rect 7856 23910 7866 23962
rect 7866 23910 7912 23962
rect 7616 23908 7672 23910
rect 7696 23908 7752 23910
rect 7776 23908 7832 23910
rect 7856 23908 7912 23910
rect 7616 22874 7672 22876
rect 7696 22874 7752 22876
rect 7776 22874 7832 22876
rect 7856 22874 7912 22876
rect 7616 22822 7662 22874
rect 7662 22822 7672 22874
rect 7696 22822 7726 22874
rect 7726 22822 7738 22874
rect 7738 22822 7752 22874
rect 7776 22822 7790 22874
rect 7790 22822 7802 22874
rect 7802 22822 7832 22874
rect 7856 22822 7866 22874
rect 7866 22822 7912 22874
rect 7616 22820 7672 22822
rect 7696 22820 7752 22822
rect 7776 22820 7832 22822
rect 7856 22820 7912 22822
rect 7616 21786 7672 21788
rect 7696 21786 7752 21788
rect 7776 21786 7832 21788
rect 7856 21786 7912 21788
rect 7616 21734 7662 21786
rect 7662 21734 7672 21786
rect 7696 21734 7726 21786
rect 7726 21734 7738 21786
rect 7738 21734 7752 21786
rect 7776 21734 7790 21786
rect 7790 21734 7802 21786
rect 7802 21734 7832 21786
rect 7856 21734 7866 21786
rect 7866 21734 7912 21786
rect 7616 21732 7672 21734
rect 7696 21732 7752 21734
rect 7776 21732 7832 21734
rect 7856 21732 7912 21734
rect 7616 20698 7672 20700
rect 7696 20698 7752 20700
rect 7776 20698 7832 20700
rect 7856 20698 7912 20700
rect 7616 20646 7662 20698
rect 7662 20646 7672 20698
rect 7696 20646 7726 20698
rect 7726 20646 7738 20698
rect 7738 20646 7752 20698
rect 7776 20646 7790 20698
rect 7790 20646 7802 20698
rect 7802 20646 7832 20698
rect 7856 20646 7866 20698
rect 7866 20646 7912 20698
rect 7616 20644 7672 20646
rect 7696 20644 7752 20646
rect 7776 20644 7832 20646
rect 7856 20644 7912 20646
rect 7616 19610 7672 19612
rect 7696 19610 7752 19612
rect 7776 19610 7832 19612
rect 7856 19610 7912 19612
rect 7616 19558 7662 19610
rect 7662 19558 7672 19610
rect 7696 19558 7726 19610
rect 7726 19558 7738 19610
rect 7738 19558 7752 19610
rect 7776 19558 7790 19610
rect 7790 19558 7802 19610
rect 7802 19558 7832 19610
rect 7856 19558 7866 19610
rect 7866 19558 7912 19610
rect 7616 19556 7672 19558
rect 7696 19556 7752 19558
rect 7776 19556 7832 19558
rect 7856 19556 7912 19558
rect 7616 18522 7672 18524
rect 7696 18522 7752 18524
rect 7776 18522 7832 18524
rect 7856 18522 7912 18524
rect 7616 18470 7662 18522
rect 7662 18470 7672 18522
rect 7696 18470 7726 18522
rect 7726 18470 7738 18522
rect 7738 18470 7752 18522
rect 7776 18470 7790 18522
rect 7790 18470 7802 18522
rect 7802 18470 7832 18522
rect 7856 18470 7866 18522
rect 7866 18470 7912 18522
rect 7616 18468 7672 18470
rect 7696 18468 7752 18470
rect 7776 18468 7832 18470
rect 7856 18468 7912 18470
rect 7616 17434 7672 17436
rect 7696 17434 7752 17436
rect 7776 17434 7832 17436
rect 7856 17434 7912 17436
rect 7616 17382 7662 17434
rect 7662 17382 7672 17434
rect 7696 17382 7726 17434
rect 7726 17382 7738 17434
rect 7738 17382 7752 17434
rect 7776 17382 7790 17434
rect 7790 17382 7802 17434
rect 7802 17382 7832 17434
rect 7856 17382 7866 17434
rect 7866 17382 7912 17434
rect 7616 17380 7672 17382
rect 7696 17380 7752 17382
rect 7776 17380 7832 17382
rect 7856 17380 7912 17382
rect 7616 16346 7672 16348
rect 7696 16346 7752 16348
rect 7776 16346 7832 16348
rect 7856 16346 7912 16348
rect 7616 16294 7662 16346
rect 7662 16294 7672 16346
rect 7696 16294 7726 16346
rect 7726 16294 7738 16346
rect 7738 16294 7752 16346
rect 7776 16294 7790 16346
rect 7790 16294 7802 16346
rect 7802 16294 7832 16346
rect 7856 16294 7866 16346
rect 7866 16294 7912 16346
rect 7616 16292 7672 16294
rect 7696 16292 7752 16294
rect 7776 16292 7832 16294
rect 7856 16292 7912 16294
rect 7616 15258 7672 15260
rect 7696 15258 7752 15260
rect 7776 15258 7832 15260
rect 7856 15258 7912 15260
rect 7616 15206 7662 15258
rect 7662 15206 7672 15258
rect 7696 15206 7726 15258
rect 7726 15206 7738 15258
rect 7738 15206 7752 15258
rect 7776 15206 7790 15258
rect 7790 15206 7802 15258
rect 7802 15206 7832 15258
rect 7856 15206 7866 15258
rect 7866 15206 7912 15258
rect 7616 15204 7672 15206
rect 7696 15204 7752 15206
rect 7776 15204 7832 15206
rect 7856 15204 7912 15206
rect 7838 15000 7894 15056
rect 7616 14170 7672 14172
rect 7696 14170 7752 14172
rect 7776 14170 7832 14172
rect 7856 14170 7912 14172
rect 7616 14118 7662 14170
rect 7662 14118 7672 14170
rect 7696 14118 7726 14170
rect 7726 14118 7738 14170
rect 7738 14118 7752 14170
rect 7776 14118 7790 14170
rect 7790 14118 7802 14170
rect 7802 14118 7832 14170
rect 7856 14118 7866 14170
rect 7866 14118 7912 14170
rect 7616 14116 7672 14118
rect 7696 14116 7752 14118
rect 7776 14116 7832 14118
rect 7856 14116 7912 14118
rect 7616 13082 7672 13084
rect 7696 13082 7752 13084
rect 7776 13082 7832 13084
rect 7856 13082 7912 13084
rect 7616 13030 7662 13082
rect 7662 13030 7672 13082
rect 7696 13030 7726 13082
rect 7726 13030 7738 13082
rect 7738 13030 7752 13082
rect 7776 13030 7790 13082
rect 7790 13030 7802 13082
rect 7802 13030 7832 13082
rect 7856 13030 7866 13082
rect 7866 13030 7912 13082
rect 7616 13028 7672 13030
rect 7696 13028 7752 13030
rect 7776 13028 7832 13030
rect 7856 13028 7912 13030
rect 7616 11994 7672 11996
rect 7696 11994 7752 11996
rect 7776 11994 7832 11996
rect 7856 11994 7912 11996
rect 7616 11942 7662 11994
rect 7662 11942 7672 11994
rect 7696 11942 7726 11994
rect 7726 11942 7738 11994
rect 7738 11942 7752 11994
rect 7776 11942 7790 11994
rect 7790 11942 7802 11994
rect 7802 11942 7832 11994
rect 7856 11942 7866 11994
rect 7866 11942 7912 11994
rect 7616 11940 7672 11942
rect 7696 11940 7752 11942
rect 7776 11940 7832 11942
rect 7856 11940 7912 11942
rect 7616 10906 7672 10908
rect 7696 10906 7752 10908
rect 7776 10906 7832 10908
rect 7856 10906 7912 10908
rect 7616 10854 7662 10906
rect 7662 10854 7672 10906
rect 7696 10854 7726 10906
rect 7726 10854 7738 10906
rect 7738 10854 7752 10906
rect 7776 10854 7790 10906
rect 7790 10854 7802 10906
rect 7802 10854 7832 10906
rect 7856 10854 7866 10906
rect 7866 10854 7912 10906
rect 7616 10852 7672 10854
rect 7696 10852 7752 10854
rect 7776 10852 7832 10854
rect 7856 10852 7912 10854
rect 7930 10512 7986 10568
rect 7010 9968 7066 10024
rect 6642 9580 6698 9616
rect 6642 9560 6644 9580
rect 6644 9560 6696 9580
rect 6696 9560 6698 9580
rect 6956 9274 7012 9276
rect 7036 9274 7092 9276
rect 7116 9274 7172 9276
rect 7196 9274 7252 9276
rect 6956 9222 7002 9274
rect 7002 9222 7012 9274
rect 7036 9222 7066 9274
rect 7066 9222 7078 9274
rect 7078 9222 7092 9274
rect 7116 9222 7130 9274
rect 7130 9222 7142 9274
rect 7142 9222 7172 9274
rect 7196 9222 7206 9274
rect 7206 9222 7252 9274
rect 6956 9220 7012 9222
rect 7036 9220 7092 9222
rect 7116 9220 7172 9222
rect 7196 9220 7252 9222
rect 6956 8186 7012 8188
rect 7036 8186 7092 8188
rect 7116 8186 7172 8188
rect 7196 8186 7252 8188
rect 6956 8134 7002 8186
rect 7002 8134 7012 8186
rect 7036 8134 7066 8186
rect 7066 8134 7078 8186
rect 7078 8134 7092 8186
rect 7116 8134 7130 8186
rect 7130 8134 7142 8186
rect 7142 8134 7172 8186
rect 7196 8134 7206 8186
rect 7206 8134 7252 8186
rect 6956 8132 7012 8134
rect 7036 8132 7092 8134
rect 7116 8132 7172 8134
rect 7196 8132 7252 8134
rect 6956 7098 7012 7100
rect 7036 7098 7092 7100
rect 7116 7098 7172 7100
rect 7196 7098 7252 7100
rect 6956 7046 7002 7098
rect 7002 7046 7012 7098
rect 7036 7046 7066 7098
rect 7066 7046 7078 7098
rect 7078 7046 7092 7098
rect 7116 7046 7130 7098
rect 7130 7046 7142 7098
rect 7142 7046 7172 7098
rect 7196 7046 7206 7098
rect 7206 7046 7252 7098
rect 6956 7044 7012 7046
rect 7036 7044 7092 7046
rect 7116 7044 7172 7046
rect 7196 7044 7252 7046
rect 6918 6704 6974 6760
rect 6956 6010 7012 6012
rect 7036 6010 7092 6012
rect 7116 6010 7172 6012
rect 7196 6010 7252 6012
rect 6956 5958 7002 6010
rect 7002 5958 7012 6010
rect 7036 5958 7066 6010
rect 7066 5958 7078 6010
rect 7078 5958 7092 6010
rect 7116 5958 7130 6010
rect 7130 5958 7142 6010
rect 7142 5958 7172 6010
rect 7196 5958 7206 6010
rect 7206 5958 7252 6010
rect 6956 5956 7012 5958
rect 7036 5956 7092 5958
rect 7116 5956 7172 5958
rect 7196 5956 7252 5958
rect 6956 4922 7012 4924
rect 7036 4922 7092 4924
rect 7116 4922 7172 4924
rect 7196 4922 7252 4924
rect 6956 4870 7002 4922
rect 7002 4870 7012 4922
rect 7036 4870 7066 4922
rect 7066 4870 7078 4922
rect 7078 4870 7092 4922
rect 7116 4870 7130 4922
rect 7130 4870 7142 4922
rect 7142 4870 7172 4922
rect 7196 4870 7206 4922
rect 7206 4870 7252 4922
rect 6956 4868 7012 4870
rect 7036 4868 7092 4870
rect 7116 4868 7172 4870
rect 7196 4868 7252 4870
rect 7616 9818 7672 9820
rect 7696 9818 7752 9820
rect 7776 9818 7832 9820
rect 7856 9818 7912 9820
rect 7616 9766 7662 9818
rect 7662 9766 7672 9818
rect 7696 9766 7726 9818
rect 7726 9766 7738 9818
rect 7738 9766 7752 9818
rect 7776 9766 7790 9818
rect 7790 9766 7802 9818
rect 7802 9766 7832 9818
rect 7856 9766 7866 9818
rect 7866 9766 7912 9818
rect 7616 9764 7672 9766
rect 7696 9764 7752 9766
rect 7776 9764 7832 9766
rect 7856 9764 7912 9766
rect 7378 6860 7434 6896
rect 8298 26016 8354 26072
rect 8482 26832 8538 26888
rect 8390 15136 8446 15192
rect 8758 62636 8760 62656
rect 8760 62636 8812 62656
rect 8812 62636 8814 62656
rect 8758 62600 8814 62636
rect 11242 76200 11298 76236
rect 8298 11056 8354 11112
rect 7616 8730 7672 8732
rect 7696 8730 7752 8732
rect 7776 8730 7832 8732
rect 7856 8730 7912 8732
rect 7616 8678 7662 8730
rect 7662 8678 7672 8730
rect 7696 8678 7726 8730
rect 7726 8678 7738 8730
rect 7738 8678 7752 8730
rect 7776 8678 7790 8730
rect 7790 8678 7802 8730
rect 7802 8678 7832 8730
rect 7856 8678 7866 8730
rect 7866 8678 7912 8730
rect 7616 8676 7672 8678
rect 7696 8676 7752 8678
rect 7776 8676 7832 8678
rect 7856 8676 7912 8678
rect 7616 7642 7672 7644
rect 7696 7642 7752 7644
rect 7776 7642 7832 7644
rect 7856 7642 7912 7644
rect 7616 7590 7662 7642
rect 7662 7590 7672 7642
rect 7696 7590 7726 7642
rect 7726 7590 7738 7642
rect 7738 7590 7752 7642
rect 7776 7590 7790 7642
rect 7790 7590 7802 7642
rect 7802 7590 7832 7642
rect 7856 7590 7866 7642
rect 7866 7590 7912 7642
rect 7616 7588 7672 7590
rect 7696 7588 7752 7590
rect 7776 7588 7832 7590
rect 7856 7588 7912 7590
rect 7378 6840 7380 6860
rect 7380 6840 7432 6860
rect 7432 6840 7434 6860
rect 7616 6554 7672 6556
rect 7696 6554 7752 6556
rect 7776 6554 7832 6556
rect 7856 6554 7912 6556
rect 7616 6502 7662 6554
rect 7662 6502 7672 6554
rect 7696 6502 7726 6554
rect 7726 6502 7738 6554
rect 7738 6502 7752 6554
rect 7776 6502 7790 6554
rect 7790 6502 7802 6554
rect 7802 6502 7832 6554
rect 7856 6502 7866 6554
rect 7866 6502 7912 6554
rect 7616 6500 7672 6502
rect 7696 6500 7752 6502
rect 7776 6500 7832 6502
rect 7856 6500 7912 6502
rect 7616 5466 7672 5468
rect 7696 5466 7752 5468
rect 7776 5466 7832 5468
rect 7856 5466 7912 5468
rect 7616 5414 7662 5466
rect 7662 5414 7672 5466
rect 7696 5414 7726 5466
rect 7726 5414 7738 5466
rect 7738 5414 7752 5466
rect 7776 5414 7790 5466
rect 7790 5414 7802 5466
rect 7802 5414 7832 5466
rect 7856 5414 7866 5466
rect 7866 5414 7912 5466
rect 7616 5412 7672 5414
rect 7696 5412 7752 5414
rect 7776 5412 7832 5414
rect 7856 5412 7912 5414
rect 7616 4378 7672 4380
rect 7696 4378 7752 4380
rect 7776 4378 7832 4380
rect 7856 4378 7912 4380
rect 7616 4326 7662 4378
rect 7662 4326 7672 4378
rect 7696 4326 7726 4378
rect 7726 4326 7738 4378
rect 7738 4326 7752 4378
rect 7776 4326 7790 4378
rect 7790 4326 7802 4378
rect 7802 4326 7832 4378
rect 7856 4326 7866 4378
rect 7866 4326 7912 4378
rect 7616 4324 7672 4326
rect 7696 4324 7752 4326
rect 7776 4324 7832 4326
rect 7856 4324 7912 4326
rect 6956 3834 7012 3836
rect 7036 3834 7092 3836
rect 7116 3834 7172 3836
rect 7196 3834 7252 3836
rect 6956 3782 7002 3834
rect 7002 3782 7012 3834
rect 7036 3782 7066 3834
rect 7066 3782 7078 3834
rect 7078 3782 7092 3834
rect 7116 3782 7130 3834
rect 7130 3782 7142 3834
rect 7142 3782 7172 3834
rect 7196 3782 7206 3834
rect 7206 3782 7252 3834
rect 6956 3780 7012 3782
rect 7036 3780 7092 3782
rect 7116 3780 7172 3782
rect 7196 3780 7252 3782
rect 7616 3290 7672 3292
rect 7696 3290 7752 3292
rect 7776 3290 7832 3292
rect 7856 3290 7912 3292
rect 7616 3238 7662 3290
rect 7662 3238 7672 3290
rect 7696 3238 7726 3290
rect 7726 3238 7738 3290
rect 7738 3238 7752 3290
rect 7776 3238 7790 3290
rect 7790 3238 7802 3290
rect 7802 3238 7832 3290
rect 7856 3238 7866 3290
rect 7866 3238 7912 3290
rect 7616 3236 7672 3238
rect 7696 3236 7752 3238
rect 7776 3236 7832 3238
rect 7856 3236 7912 3238
rect 1956 2746 2012 2748
rect 2036 2746 2092 2748
rect 2116 2746 2172 2748
rect 2196 2746 2252 2748
rect 1956 2694 2002 2746
rect 2002 2694 2012 2746
rect 2036 2694 2066 2746
rect 2066 2694 2078 2746
rect 2078 2694 2092 2746
rect 2116 2694 2130 2746
rect 2130 2694 2142 2746
rect 2142 2694 2172 2746
rect 2196 2694 2206 2746
rect 2206 2694 2252 2746
rect 1956 2692 2012 2694
rect 2036 2692 2092 2694
rect 2116 2692 2172 2694
rect 2196 2692 2252 2694
rect 6956 2746 7012 2748
rect 7036 2746 7092 2748
rect 7116 2746 7172 2748
rect 7196 2746 7252 2748
rect 6956 2694 7002 2746
rect 7002 2694 7012 2746
rect 7036 2694 7066 2746
rect 7066 2694 7078 2746
rect 7078 2694 7092 2746
rect 7116 2694 7130 2746
rect 7130 2694 7142 2746
rect 7142 2694 7172 2746
rect 7196 2694 7206 2746
rect 7206 2694 7252 2746
rect 6956 2692 7012 2694
rect 7036 2692 7092 2694
rect 7116 2692 7172 2694
rect 7196 2692 7252 2694
rect 8942 33088 8998 33144
rect 8942 26968 8998 27024
rect 9494 52536 9550 52592
rect 9494 40432 9550 40488
rect 9034 16496 9090 16552
rect 9770 24812 9826 24848
rect 9770 24792 9772 24812
rect 9772 24792 9824 24812
rect 9824 24792 9826 24812
rect 10046 36352 10102 36408
rect 10506 67632 10562 67688
rect 10598 52400 10654 52456
rect 10690 50668 10692 50688
rect 10692 50668 10744 50688
rect 10744 50668 10746 50688
rect 10690 50632 10746 50668
rect 10414 42628 10470 42664
rect 10414 42608 10416 42628
rect 10416 42608 10468 42628
rect 10468 42608 10470 42628
rect 10138 26036 10194 26072
rect 10138 26016 10140 26036
rect 10140 26016 10192 26036
rect 10192 26016 10194 26036
rect 10322 25356 10378 25392
rect 11058 42744 11114 42800
rect 10322 25336 10324 25356
rect 10324 25336 10376 25356
rect 10376 25336 10378 25356
rect 9678 6724 9734 6760
rect 9678 6704 9680 6724
rect 9680 6704 9732 6724
rect 9732 6704 9734 6724
rect 11426 55800 11482 55856
rect 11426 51312 11482 51368
rect 12616 76186 12672 76188
rect 12696 76186 12752 76188
rect 12776 76186 12832 76188
rect 12856 76186 12912 76188
rect 12616 76134 12662 76186
rect 12662 76134 12672 76186
rect 12696 76134 12726 76186
rect 12726 76134 12738 76186
rect 12738 76134 12752 76186
rect 12776 76134 12790 76186
rect 12790 76134 12802 76186
rect 12802 76134 12832 76186
rect 12856 76134 12866 76186
rect 12866 76134 12912 76186
rect 12616 76132 12672 76134
rect 12696 76132 12752 76134
rect 12776 76132 12832 76134
rect 12856 76132 12912 76134
rect 11956 75642 12012 75644
rect 12036 75642 12092 75644
rect 12116 75642 12172 75644
rect 12196 75642 12252 75644
rect 11956 75590 12002 75642
rect 12002 75590 12012 75642
rect 12036 75590 12066 75642
rect 12066 75590 12078 75642
rect 12078 75590 12092 75642
rect 12116 75590 12130 75642
rect 12130 75590 12142 75642
rect 12142 75590 12172 75642
rect 12196 75590 12206 75642
rect 12206 75590 12252 75642
rect 11956 75588 12012 75590
rect 12036 75588 12092 75590
rect 12116 75588 12172 75590
rect 12196 75588 12252 75590
rect 11956 74554 12012 74556
rect 12036 74554 12092 74556
rect 12116 74554 12172 74556
rect 12196 74554 12252 74556
rect 11956 74502 12002 74554
rect 12002 74502 12012 74554
rect 12036 74502 12066 74554
rect 12066 74502 12078 74554
rect 12078 74502 12092 74554
rect 12116 74502 12130 74554
rect 12130 74502 12142 74554
rect 12142 74502 12172 74554
rect 12196 74502 12206 74554
rect 12206 74502 12252 74554
rect 11956 74500 12012 74502
rect 12036 74500 12092 74502
rect 12116 74500 12172 74502
rect 12196 74500 12252 74502
rect 12616 75098 12672 75100
rect 12696 75098 12752 75100
rect 12776 75098 12832 75100
rect 12856 75098 12912 75100
rect 12616 75046 12662 75098
rect 12662 75046 12672 75098
rect 12696 75046 12726 75098
rect 12726 75046 12738 75098
rect 12738 75046 12752 75098
rect 12776 75046 12790 75098
rect 12790 75046 12802 75098
rect 12802 75046 12832 75098
rect 12856 75046 12866 75098
rect 12866 75046 12912 75098
rect 12616 75044 12672 75046
rect 12696 75044 12752 75046
rect 12776 75044 12832 75046
rect 12856 75044 12912 75046
rect 11956 73466 12012 73468
rect 12036 73466 12092 73468
rect 12116 73466 12172 73468
rect 12196 73466 12252 73468
rect 11956 73414 12002 73466
rect 12002 73414 12012 73466
rect 12036 73414 12066 73466
rect 12066 73414 12078 73466
rect 12078 73414 12092 73466
rect 12116 73414 12130 73466
rect 12130 73414 12142 73466
rect 12142 73414 12172 73466
rect 12196 73414 12206 73466
rect 12206 73414 12252 73466
rect 11956 73412 12012 73414
rect 12036 73412 12092 73414
rect 12116 73412 12172 73414
rect 12196 73412 12252 73414
rect 11956 72378 12012 72380
rect 12036 72378 12092 72380
rect 12116 72378 12172 72380
rect 12196 72378 12252 72380
rect 11956 72326 12002 72378
rect 12002 72326 12012 72378
rect 12036 72326 12066 72378
rect 12066 72326 12078 72378
rect 12078 72326 12092 72378
rect 12116 72326 12130 72378
rect 12130 72326 12142 72378
rect 12142 72326 12172 72378
rect 12196 72326 12206 72378
rect 12206 72326 12252 72378
rect 11956 72324 12012 72326
rect 12036 72324 12092 72326
rect 12116 72324 12172 72326
rect 12196 72324 12252 72326
rect 11956 71290 12012 71292
rect 12036 71290 12092 71292
rect 12116 71290 12172 71292
rect 12196 71290 12252 71292
rect 11956 71238 12002 71290
rect 12002 71238 12012 71290
rect 12036 71238 12066 71290
rect 12066 71238 12078 71290
rect 12078 71238 12092 71290
rect 12116 71238 12130 71290
rect 12130 71238 12142 71290
rect 12142 71238 12172 71290
rect 12196 71238 12206 71290
rect 12206 71238 12252 71290
rect 11956 71236 12012 71238
rect 12036 71236 12092 71238
rect 12116 71236 12172 71238
rect 12196 71236 12252 71238
rect 11956 70202 12012 70204
rect 12036 70202 12092 70204
rect 12116 70202 12172 70204
rect 12196 70202 12252 70204
rect 11956 70150 12002 70202
rect 12002 70150 12012 70202
rect 12036 70150 12066 70202
rect 12066 70150 12078 70202
rect 12078 70150 12092 70202
rect 12116 70150 12130 70202
rect 12130 70150 12142 70202
rect 12142 70150 12172 70202
rect 12196 70150 12206 70202
rect 12206 70150 12252 70202
rect 11956 70148 12012 70150
rect 12036 70148 12092 70150
rect 12116 70148 12172 70150
rect 12196 70148 12252 70150
rect 11956 69114 12012 69116
rect 12036 69114 12092 69116
rect 12116 69114 12172 69116
rect 12196 69114 12252 69116
rect 11956 69062 12002 69114
rect 12002 69062 12012 69114
rect 12036 69062 12066 69114
rect 12066 69062 12078 69114
rect 12078 69062 12092 69114
rect 12116 69062 12130 69114
rect 12130 69062 12142 69114
rect 12142 69062 12172 69114
rect 12196 69062 12206 69114
rect 12206 69062 12252 69114
rect 11956 69060 12012 69062
rect 12036 69060 12092 69062
rect 12116 69060 12172 69062
rect 12196 69060 12252 69062
rect 11956 68026 12012 68028
rect 12036 68026 12092 68028
rect 12116 68026 12172 68028
rect 12196 68026 12252 68028
rect 11956 67974 12002 68026
rect 12002 67974 12012 68026
rect 12036 67974 12066 68026
rect 12066 67974 12078 68026
rect 12078 67974 12092 68026
rect 12116 67974 12130 68026
rect 12130 67974 12142 68026
rect 12142 67974 12172 68026
rect 12196 67974 12206 68026
rect 12206 67974 12252 68026
rect 11956 67972 12012 67974
rect 12036 67972 12092 67974
rect 12116 67972 12172 67974
rect 12196 67972 12252 67974
rect 12070 67652 12126 67688
rect 12070 67632 12072 67652
rect 12072 67632 12124 67652
rect 12124 67632 12126 67652
rect 11956 66938 12012 66940
rect 12036 66938 12092 66940
rect 12116 66938 12172 66940
rect 12196 66938 12252 66940
rect 11956 66886 12002 66938
rect 12002 66886 12012 66938
rect 12036 66886 12066 66938
rect 12066 66886 12078 66938
rect 12078 66886 12092 66938
rect 12116 66886 12130 66938
rect 12130 66886 12142 66938
rect 12142 66886 12172 66938
rect 12196 66886 12206 66938
rect 12206 66886 12252 66938
rect 11956 66884 12012 66886
rect 12036 66884 12092 66886
rect 12116 66884 12172 66886
rect 12196 66884 12252 66886
rect 11956 65850 12012 65852
rect 12036 65850 12092 65852
rect 12116 65850 12172 65852
rect 12196 65850 12252 65852
rect 11956 65798 12002 65850
rect 12002 65798 12012 65850
rect 12036 65798 12066 65850
rect 12066 65798 12078 65850
rect 12078 65798 12092 65850
rect 12116 65798 12130 65850
rect 12130 65798 12142 65850
rect 12142 65798 12172 65850
rect 12196 65798 12206 65850
rect 12206 65798 12252 65850
rect 11956 65796 12012 65798
rect 12036 65796 12092 65798
rect 12116 65796 12172 65798
rect 12196 65796 12252 65798
rect 11956 64762 12012 64764
rect 12036 64762 12092 64764
rect 12116 64762 12172 64764
rect 12196 64762 12252 64764
rect 11956 64710 12002 64762
rect 12002 64710 12012 64762
rect 12036 64710 12066 64762
rect 12066 64710 12078 64762
rect 12078 64710 12092 64762
rect 12116 64710 12130 64762
rect 12130 64710 12142 64762
rect 12142 64710 12172 64762
rect 12196 64710 12206 64762
rect 12206 64710 12252 64762
rect 11956 64708 12012 64710
rect 12036 64708 12092 64710
rect 12116 64708 12172 64710
rect 12196 64708 12252 64710
rect 11956 63674 12012 63676
rect 12036 63674 12092 63676
rect 12116 63674 12172 63676
rect 12196 63674 12252 63676
rect 11956 63622 12002 63674
rect 12002 63622 12012 63674
rect 12036 63622 12066 63674
rect 12066 63622 12078 63674
rect 12078 63622 12092 63674
rect 12116 63622 12130 63674
rect 12130 63622 12142 63674
rect 12142 63622 12172 63674
rect 12196 63622 12206 63674
rect 12206 63622 12252 63674
rect 11956 63620 12012 63622
rect 12036 63620 12092 63622
rect 12116 63620 12172 63622
rect 12196 63620 12252 63622
rect 11956 62586 12012 62588
rect 12036 62586 12092 62588
rect 12116 62586 12172 62588
rect 12196 62586 12252 62588
rect 11956 62534 12002 62586
rect 12002 62534 12012 62586
rect 12036 62534 12066 62586
rect 12066 62534 12078 62586
rect 12078 62534 12092 62586
rect 12116 62534 12130 62586
rect 12130 62534 12142 62586
rect 12142 62534 12172 62586
rect 12196 62534 12206 62586
rect 12206 62534 12252 62586
rect 11956 62532 12012 62534
rect 12036 62532 12092 62534
rect 12116 62532 12172 62534
rect 12196 62532 12252 62534
rect 12616 74010 12672 74012
rect 12696 74010 12752 74012
rect 12776 74010 12832 74012
rect 12856 74010 12912 74012
rect 12616 73958 12662 74010
rect 12662 73958 12672 74010
rect 12696 73958 12726 74010
rect 12726 73958 12738 74010
rect 12738 73958 12752 74010
rect 12776 73958 12790 74010
rect 12790 73958 12802 74010
rect 12802 73958 12832 74010
rect 12856 73958 12866 74010
rect 12866 73958 12912 74010
rect 12616 73956 12672 73958
rect 12696 73956 12752 73958
rect 12776 73956 12832 73958
rect 12856 73956 12912 73958
rect 12616 72922 12672 72924
rect 12696 72922 12752 72924
rect 12776 72922 12832 72924
rect 12856 72922 12912 72924
rect 12616 72870 12662 72922
rect 12662 72870 12672 72922
rect 12696 72870 12726 72922
rect 12726 72870 12738 72922
rect 12738 72870 12752 72922
rect 12776 72870 12790 72922
rect 12790 72870 12802 72922
rect 12802 72870 12832 72922
rect 12856 72870 12866 72922
rect 12866 72870 12912 72922
rect 12616 72868 12672 72870
rect 12696 72868 12752 72870
rect 12776 72868 12832 72870
rect 12856 72868 12912 72870
rect 12616 71834 12672 71836
rect 12696 71834 12752 71836
rect 12776 71834 12832 71836
rect 12856 71834 12912 71836
rect 12616 71782 12662 71834
rect 12662 71782 12672 71834
rect 12696 71782 12726 71834
rect 12726 71782 12738 71834
rect 12738 71782 12752 71834
rect 12776 71782 12790 71834
rect 12790 71782 12802 71834
rect 12802 71782 12832 71834
rect 12856 71782 12866 71834
rect 12866 71782 12912 71834
rect 12616 71780 12672 71782
rect 12696 71780 12752 71782
rect 12776 71780 12832 71782
rect 12856 71780 12912 71782
rect 12616 70746 12672 70748
rect 12696 70746 12752 70748
rect 12776 70746 12832 70748
rect 12856 70746 12912 70748
rect 12616 70694 12662 70746
rect 12662 70694 12672 70746
rect 12696 70694 12726 70746
rect 12726 70694 12738 70746
rect 12738 70694 12752 70746
rect 12776 70694 12790 70746
rect 12790 70694 12802 70746
rect 12802 70694 12832 70746
rect 12856 70694 12866 70746
rect 12866 70694 12912 70746
rect 12616 70692 12672 70694
rect 12696 70692 12752 70694
rect 12776 70692 12832 70694
rect 12856 70692 12912 70694
rect 12616 69658 12672 69660
rect 12696 69658 12752 69660
rect 12776 69658 12832 69660
rect 12856 69658 12912 69660
rect 12616 69606 12662 69658
rect 12662 69606 12672 69658
rect 12696 69606 12726 69658
rect 12726 69606 12738 69658
rect 12738 69606 12752 69658
rect 12776 69606 12790 69658
rect 12790 69606 12802 69658
rect 12802 69606 12832 69658
rect 12856 69606 12866 69658
rect 12866 69606 12912 69658
rect 12616 69604 12672 69606
rect 12696 69604 12752 69606
rect 12776 69604 12832 69606
rect 12856 69604 12912 69606
rect 12616 68570 12672 68572
rect 12696 68570 12752 68572
rect 12776 68570 12832 68572
rect 12856 68570 12912 68572
rect 12616 68518 12662 68570
rect 12662 68518 12672 68570
rect 12696 68518 12726 68570
rect 12726 68518 12738 68570
rect 12738 68518 12752 68570
rect 12776 68518 12790 68570
rect 12790 68518 12802 68570
rect 12802 68518 12832 68570
rect 12856 68518 12866 68570
rect 12866 68518 12912 68570
rect 12616 68516 12672 68518
rect 12696 68516 12752 68518
rect 12776 68516 12832 68518
rect 12856 68516 12912 68518
rect 12616 67482 12672 67484
rect 12696 67482 12752 67484
rect 12776 67482 12832 67484
rect 12856 67482 12912 67484
rect 12616 67430 12662 67482
rect 12662 67430 12672 67482
rect 12696 67430 12726 67482
rect 12726 67430 12738 67482
rect 12738 67430 12752 67482
rect 12776 67430 12790 67482
rect 12790 67430 12802 67482
rect 12802 67430 12832 67482
rect 12856 67430 12866 67482
rect 12866 67430 12912 67482
rect 12616 67428 12672 67430
rect 12696 67428 12752 67430
rect 12776 67428 12832 67430
rect 12856 67428 12912 67430
rect 12616 66394 12672 66396
rect 12696 66394 12752 66396
rect 12776 66394 12832 66396
rect 12856 66394 12912 66396
rect 12616 66342 12662 66394
rect 12662 66342 12672 66394
rect 12696 66342 12726 66394
rect 12726 66342 12738 66394
rect 12738 66342 12752 66394
rect 12776 66342 12790 66394
rect 12790 66342 12802 66394
rect 12802 66342 12832 66394
rect 12856 66342 12866 66394
rect 12866 66342 12912 66394
rect 12616 66340 12672 66342
rect 12696 66340 12752 66342
rect 12776 66340 12832 66342
rect 12856 66340 12912 66342
rect 12616 65306 12672 65308
rect 12696 65306 12752 65308
rect 12776 65306 12832 65308
rect 12856 65306 12912 65308
rect 12616 65254 12662 65306
rect 12662 65254 12672 65306
rect 12696 65254 12726 65306
rect 12726 65254 12738 65306
rect 12738 65254 12752 65306
rect 12776 65254 12790 65306
rect 12790 65254 12802 65306
rect 12802 65254 12832 65306
rect 12856 65254 12866 65306
rect 12866 65254 12912 65306
rect 12616 65252 12672 65254
rect 12696 65252 12752 65254
rect 12776 65252 12832 65254
rect 12856 65252 12912 65254
rect 12616 64218 12672 64220
rect 12696 64218 12752 64220
rect 12776 64218 12832 64220
rect 12856 64218 12912 64220
rect 12616 64166 12662 64218
rect 12662 64166 12672 64218
rect 12696 64166 12726 64218
rect 12726 64166 12738 64218
rect 12738 64166 12752 64218
rect 12776 64166 12790 64218
rect 12790 64166 12802 64218
rect 12802 64166 12832 64218
rect 12856 64166 12866 64218
rect 12866 64166 12912 64218
rect 12616 64164 12672 64166
rect 12696 64164 12752 64166
rect 12776 64164 12832 64166
rect 12856 64164 12912 64166
rect 12616 63130 12672 63132
rect 12696 63130 12752 63132
rect 12776 63130 12832 63132
rect 12856 63130 12912 63132
rect 12616 63078 12662 63130
rect 12662 63078 12672 63130
rect 12696 63078 12726 63130
rect 12726 63078 12738 63130
rect 12738 63078 12752 63130
rect 12776 63078 12790 63130
rect 12790 63078 12802 63130
rect 12802 63078 12832 63130
rect 12856 63078 12866 63130
rect 12866 63078 12912 63130
rect 12616 63076 12672 63078
rect 12696 63076 12752 63078
rect 12776 63076 12832 63078
rect 12856 63076 12912 63078
rect 12616 62042 12672 62044
rect 12696 62042 12752 62044
rect 12776 62042 12832 62044
rect 12856 62042 12912 62044
rect 12616 61990 12662 62042
rect 12662 61990 12672 62042
rect 12696 61990 12726 62042
rect 12726 61990 12738 62042
rect 12738 61990 12752 62042
rect 12776 61990 12790 62042
rect 12790 61990 12802 62042
rect 12802 61990 12832 62042
rect 12856 61990 12866 62042
rect 12866 61990 12912 62042
rect 12616 61988 12672 61990
rect 12696 61988 12752 61990
rect 12776 61988 12832 61990
rect 12856 61988 12912 61990
rect 11956 61498 12012 61500
rect 12036 61498 12092 61500
rect 12116 61498 12172 61500
rect 12196 61498 12252 61500
rect 11956 61446 12002 61498
rect 12002 61446 12012 61498
rect 12036 61446 12066 61498
rect 12066 61446 12078 61498
rect 12078 61446 12092 61498
rect 12116 61446 12130 61498
rect 12130 61446 12142 61498
rect 12142 61446 12172 61498
rect 12196 61446 12206 61498
rect 12206 61446 12252 61498
rect 11956 61444 12012 61446
rect 12036 61444 12092 61446
rect 12116 61444 12172 61446
rect 12196 61444 12252 61446
rect 12616 60954 12672 60956
rect 12696 60954 12752 60956
rect 12776 60954 12832 60956
rect 12856 60954 12912 60956
rect 12616 60902 12662 60954
rect 12662 60902 12672 60954
rect 12696 60902 12726 60954
rect 12726 60902 12738 60954
rect 12738 60902 12752 60954
rect 12776 60902 12790 60954
rect 12790 60902 12802 60954
rect 12802 60902 12832 60954
rect 12856 60902 12866 60954
rect 12866 60902 12912 60954
rect 12616 60900 12672 60902
rect 12696 60900 12752 60902
rect 12776 60900 12832 60902
rect 12856 60900 12912 60902
rect 11956 60410 12012 60412
rect 12036 60410 12092 60412
rect 12116 60410 12172 60412
rect 12196 60410 12252 60412
rect 11956 60358 12002 60410
rect 12002 60358 12012 60410
rect 12036 60358 12066 60410
rect 12066 60358 12078 60410
rect 12078 60358 12092 60410
rect 12116 60358 12130 60410
rect 12130 60358 12142 60410
rect 12142 60358 12172 60410
rect 12196 60358 12206 60410
rect 12206 60358 12252 60410
rect 11956 60356 12012 60358
rect 12036 60356 12092 60358
rect 12116 60356 12172 60358
rect 12196 60356 12252 60358
rect 12616 59866 12672 59868
rect 12696 59866 12752 59868
rect 12776 59866 12832 59868
rect 12856 59866 12912 59868
rect 12616 59814 12662 59866
rect 12662 59814 12672 59866
rect 12696 59814 12726 59866
rect 12726 59814 12738 59866
rect 12738 59814 12752 59866
rect 12776 59814 12790 59866
rect 12790 59814 12802 59866
rect 12802 59814 12832 59866
rect 12856 59814 12866 59866
rect 12866 59814 12912 59866
rect 12616 59812 12672 59814
rect 12696 59812 12752 59814
rect 12776 59812 12832 59814
rect 12856 59812 12912 59814
rect 11956 59322 12012 59324
rect 12036 59322 12092 59324
rect 12116 59322 12172 59324
rect 12196 59322 12252 59324
rect 11956 59270 12002 59322
rect 12002 59270 12012 59322
rect 12036 59270 12066 59322
rect 12066 59270 12078 59322
rect 12078 59270 12092 59322
rect 12116 59270 12130 59322
rect 12130 59270 12142 59322
rect 12142 59270 12172 59322
rect 12196 59270 12206 59322
rect 12206 59270 12252 59322
rect 11956 59268 12012 59270
rect 12036 59268 12092 59270
rect 12116 59268 12172 59270
rect 12196 59268 12252 59270
rect 12616 58778 12672 58780
rect 12696 58778 12752 58780
rect 12776 58778 12832 58780
rect 12856 58778 12912 58780
rect 12616 58726 12662 58778
rect 12662 58726 12672 58778
rect 12696 58726 12726 58778
rect 12726 58726 12738 58778
rect 12738 58726 12752 58778
rect 12776 58726 12790 58778
rect 12790 58726 12802 58778
rect 12802 58726 12832 58778
rect 12856 58726 12866 58778
rect 12866 58726 12912 58778
rect 12616 58724 12672 58726
rect 12696 58724 12752 58726
rect 12776 58724 12832 58726
rect 12856 58724 12912 58726
rect 11956 58234 12012 58236
rect 12036 58234 12092 58236
rect 12116 58234 12172 58236
rect 12196 58234 12252 58236
rect 11956 58182 12002 58234
rect 12002 58182 12012 58234
rect 12036 58182 12066 58234
rect 12066 58182 12078 58234
rect 12078 58182 12092 58234
rect 12116 58182 12130 58234
rect 12130 58182 12142 58234
rect 12142 58182 12172 58234
rect 12196 58182 12206 58234
rect 12206 58182 12252 58234
rect 11956 58180 12012 58182
rect 12036 58180 12092 58182
rect 12116 58180 12172 58182
rect 12196 58180 12252 58182
rect 12616 57690 12672 57692
rect 12696 57690 12752 57692
rect 12776 57690 12832 57692
rect 12856 57690 12912 57692
rect 12616 57638 12662 57690
rect 12662 57638 12672 57690
rect 12696 57638 12726 57690
rect 12726 57638 12738 57690
rect 12738 57638 12752 57690
rect 12776 57638 12790 57690
rect 12790 57638 12802 57690
rect 12802 57638 12832 57690
rect 12856 57638 12866 57690
rect 12866 57638 12912 57690
rect 12616 57636 12672 57638
rect 12696 57636 12752 57638
rect 12776 57636 12832 57638
rect 12856 57636 12912 57638
rect 11956 57146 12012 57148
rect 12036 57146 12092 57148
rect 12116 57146 12172 57148
rect 12196 57146 12252 57148
rect 11956 57094 12002 57146
rect 12002 57094 12012 57146
rect 12036 57094 12066 57146
rect 12066 57094 12078 57146
rect 12078 57094 12092 57146
rect 12116 57094 12130 57146
rect 12130 57094 12142 57146
rect 12142 57094 12172 57146
rect 12196 57094 12206 57146
rect 12206 57094 12252 57146
rect 11956 57092 12012 57094
rect 12036 57092 12092 57094
rect 12116 57092 12172 57094
rect 12196 57092 12252 57094
rect 12616 56602 12672 56604
rect 12696 56602 12752 56604
rect 12776 56602 12832 56604
rect 12856 56602 12912 56604
rect 12616 56550 12662 56602
rect 12662 56550 12672 56602
rect 12696 56550 12726 56602
rect 12726 56550 12738 56602
rect 12738 56550 12752 56602
rect 12776 56550 12790 56602
rect 12790 56550 12802 56602
rect 12802 56550 12832 56602
rect 12856 56550 12866 56602
rect 12866 56550 12912 56602
rect 12616 56548 12672 56550
rect 12696 56548 12752 56550
rect 12776 56548 12832 56550
rect 12856 56548 12912 56550
rect 11956 56058 12012 56060
rect 12036 56058 12092 56060
rect 12116 56058 12172 56060
rect 12196 56058 12252 56060
rect 11956 56006 12002 56058
rect 12002 56006 12012 56058
rect 12036 56006 12066 56058
rect 12066 56006 12078 56058
rect 12078 56006 12092 56058
rect 12116 56006 12130 56058
rect 12130 56006 12142 56058
rect 12142 56006 12172 56058
rect 12196 56006 12206 56058
rect 12206 56006 12252 56058
rect 11956 56004 12012 56006
rect 12036 56004 12092 56006
rect 12116 56004 12172 56006
rect 12196 56004 12252 56006
rect 12438 55664 12494 55720
rect 12616 55514 12672 55516
rect 12696 55514 12752 55516
rect 12776 55514 12832 55516
rect 12856 55514 12912 55516
rect 12616 55462 12662 55514
rect 12662 55462 12672 55514
rect 12696 55462 12726 55514
rect 12726 55462 12738 55514
rect 12738 55462 12752 55514
rect 12776 55462 12790 55514
rect 12790 55462 12802 55514
rect 12802 55462 12832 55514
rect 12856 55462 12866 55514
rect 12866 55462 12912 55514
rect 12616 55460 12672 55462
rect 12696 55460 12752 55462
rect 12776 55460 12832 55462
rect 12856 55460 12912 55462
rect 11956 54970 12012 54972
rect 12036 54970 12092 54972
rect 12116 54970 12172 54972
rect 12196 54970 12252 54972
rect 11956 54918 12002 54970
rect 12002 54918 12012 54970
rect 12036 54918 12066 54970
rect 12066 54918 12078 54970
rect 12078 54918 12092 54970
rect 12116 54918 12130 54970
rect 12130 54918 12142 54970
rect 12142 54918 12172 54970
rect 12196 54918 12206 54970
rect 12206 54918 12252 54970
rect 11956 54916 12012 54918
rect 12036 54916 12092 54918
rect 12116 54916 12172 54918
rect 12196 54916 12252 54918
rect 12616 54426 12672 54428
rect 12696 54426 12752 54428
rect 12776 54426 12832 54428
rect 12856 54426 12912 54428
rect 12616 54374 12662 54426
rect 12662 54374 12672 54426
rect 12696 54374 12726 54426
rect 12726 54374 12738 54426
rect 12738 54374 12752 54426
rect 12776 54374 12790 54426
rect 12790 54374 12802 54426
rect 12802 54374 12832 54426
rect 12856 54374 12866 54426
rect 12866 54374 12912 54426
rect 12616 54372 12672 54374
rect 12696 54372 12752 54374
rect 12776 54372 12832 54374
rect 12856 54372 12912 54374
rect 12438 54032 12494 54088
rect 11956 53882 12012 53884
rect 12036 53882 12092 53884
rect 12116 53882 12172 53884
rect 12196 53882 12252 53884
rect 11956 53830 12002 53882
rect 12002 53830 12012 53882
rect 12036 53830 12066 53882
rect 12066 53830 12078 53882
rect 12078 53830 12092 53882
rect 12116 53830 12130 53882
rect 12130 53830 12142 53882
rect 12142 53830 12172 53882
rect 12196 53830 12206 53882
rect 12206 53830 12252 53882
rect 11956 53828 12012 53830
rect 12036 53828 12092 53830
rect 12116 53828 12172 53830
rect 12196 53828 12252 53830
rect 11956 52794 12012 52796
rect 12036 52794 12092 52796
rect 12116 52794 12172 52796
rect 12196 52794 12252 52796
rect 11956 52742 12002 52794
rect 12002 52742 12012 52794
rect 12036 52742 12066 52794
rect 12066 52742 12078 52794
rect 12078 52742 12092 52794
rect 12116 52742 12130 52794
rect 12130 52742 12142 52794
rect 12142 52742 12172 52794
rect 12196 52742 12206 52794
rect 12206 52742 12252 52794
rect 11956 52740 12012 52742
rect 12036 52740 12092 52742
rect 12116 52740 12172 52742
rect 12196 52740 12252 52742
rect 11956 51706 12012 51708
rect 12036 51706 12092 51708
rect 12116 51706 12172 51708
rect 12196 51706 12252 51708
rect 11956 51654 12002 51706
rect 12002 51654 12012 51706
rect 12036 51654 12066 51706
rect 12066 51654 12078 51706
rect 12078 51654 12092 51706
rect 12116 51654 12130 51706
rect 12130 51654 12142 51706
rect 12142 51654 12172 51706
rect 12196 51654 12206 51706
rect 12206 51654 12252 51706
rect 11956 51652 12012 51654
rect 12036 51652 12092 51654
rect 12116 51652 12172 51654
rect 12196 51652 12252 51654
rect 11956 50618 12012 50620
rect 12036 50618 12092 50620
rect 12116 50618 12172 50620
rect 12196 50618 12252 50620
rect 11956 50566 12002 50618
rect 12002 50566 12012 50618
rect 12036 50566 12066 50618
rect 12066 50566 12078 50618
rect 12078 50566 12092 50618
rect 12116 50566 12130 50618
rect 12130 50566 12142 50618
rect 12142 50566 12172 50618
rect 12196 50566 12206 50618
rect 12206 50566 12252 50618
rect 11956 50564 12012 50566
rect 12036 50564 12092 50566
rect 12116 50564 12172 50566
rect 12196 50564 12252 50566
rect 11956 49530 12012 49532
rect 12036 49530 12092 49532
rect 12116 49530 12172 49532
rect 12196 49530 12252 49532
rect 11956 49478 12002 49530
rect 12002 49478 12012 49530
rect 12036 49478 12066 49530
rect 12066 49478 12078 49530
rect 12078 49478 12092 49530
rect 12116 49478 12130 49530
rect 12130 49478 12142 49530
rect 12142 49478 12172 49530
rect 12196 49478 12206 49530
rect 12206 49478 12252 49530
rect 11956 49476 12012 49478
rect 12036 49476 12092 49478
rect 12116 49476 12172 49478
rect 12196 49476 12252 49478
rect 11956 48442 12012 48444
rect 12036 48442 12092 48444
rect 12116 48442 12172 48444
rect 12196 48442 12252 48444
rect 11956 48390 12002 48442
rect 12002 48390 12012 48442
rect 12036 48390 12066 48442
rect 12066 48390 12078 48442
rect 12078 48390 12092 48442
rect 12116 48390 12130 48442
rect 12130 48390 12142 48442
rect 12142 48390 12172 48442
rect 12196 48390 12206 48442
rect 12206 48390 12252 48442
rect 11956 48388 12012 48390
rect 12036 48388 12092 48390
rect 12116 48388 12172 48390
rect 12196 48388 12252 48390
rect 11956 47354 12012 47356
rect 12036 47354 12092 47356
rect 12116 47354 12172 47356
rect 12196 47354 12252 47356
rect 11956 47302 12002 47354
rect 12002 47302 12012 47354
rect 12036 47302 12066 47354
rect 12066 47302 12078 47354
rect 12078 47302 12092 47354
rect 12116 47302 12130 47354
rect 12130 47302 12142 47354
rect 12142 47302 12172 47354
rect 12196 47302 12206 47354
rect 12206 47302 12252 47354
rect 11956 47300 12012 47302
rect 12036 47300 12092 47302
rect 12116 47300 12172 47302
rect 12196 47300 12252 47302
rect 12616 53338 12672 53340
rect 12696 53338 12752 53340
rect 12776 53338 12832 53340
rect 12856 53338 12912 53340
rect 12616 53286 12662 53338
rect 12662 53286 12672 53338
rect 12696 53286 12726 53338
rect 12726 53286 12738 53338
rect 12738 53286 12752 53338
rect 12776 53286 12790 53338
rect 12790 53286 12802 53338
rect 12802 53286 12832 53338
rect 12856 53286 12866 53338
rect 12866 53286 12912 53338
rect 12616 53284 12672 53286
rect 12696 53284 12752 53286
rect 12776 53284 12832 53286
rect 12856 53284 12912 53286
rect 12616 52250 12672 52252
rect 12696 52250 12752 52252
rect 12776 52250 12832 52252
rect 12856 52250 12912 52252
rect 12616 52198 12662 52250
rect 12662 52198 12672 52250
rect 12696 52198 12726 52250
rect 12726 52198 12738 52250
rect 12738 52198 12752 52250
rect 12776 52198 12790 52250
rect 12790 52198 12802 52250
rect 12802 52198 12832 52250
rect 12856 52198 12866 52250
rect 12866 52198 12912 52250
rect 12616 52196 12672 52198
rect 12696 52196 12752 52198
rect 12776 52196 12832 52198
rect 12856 52196 12912 52198
rect 12616 51162 12672 51164
rect 12696 51162 12752 51164
rect 12776 51162 12832 51164
rect 12856 51162 12912 51164
rect 12616 51110 12662 51162
rect 12662 51110 12672 51162
rect 12696 51110 12726 51162
rect 12726 51110 12738 51162
rect 12738 51110 12752 51162
rect 12776 51110 12790 51162
rect 12790 51110 12802 51162
rect 12802 51110 12832 51162
rect 12856 51110 12866 51162
rect 12866 51110 12912 51162
rect 12616 51108 12672 51110
rect 12696 51108 12752 51110
rect 12776 51108 12832 51110
rect 12856 51108 12912 51110
rect 12616 50074 12672 50076
rect 12696 50074 12752 50076
rect 12776 50074 12832 50076
rect 12856 50074 12912 50076
rect 12616 50022 12662 50074
rect 12662 50022 12672 50074
rect 12696 50022 12726 50074
rect 12726 50022 12738 50074
rect 12738 50022 12752 50074
rect 12776 50022 12790 50074
rect 12790 50022 12802 50074
rect 12802 50022 12832 50074
rect 12856 50022 12866 50074
rect 12866 50022 12912 50074
rect 12616 50020 12672 50022
rect 12696 50020 12752 50022
rect 12776 50020 12832 50022
rect 12856 50020 12912 50022
rect 12616 48986 12672 48988
rect 12696 48986 12752 48988
rect 12776 48986 12832 48988
rect 12856 48986 12912 48988
rect 12616 48934 12662 48986
rect 12662 48934 12672 48986
rect 12696 48934 12726 48986
rect 12726 48934 12738 48986
rect 12738 48934 12752 48986
rect 12776 48934 12790 48986
rect 12790 48934 12802 48986
rect 12802 48934 12832 48986
rect 12856 48934 12866 48986
rect 12866 48934 12912 48986
rect 12616 48932 12672 48934
rect 12696 48932 12752 48934
rect 12776 48932 12832 48934
rect 12856 48932 12912 48934
rect 12616 47898 12672 47900
rect 12696 47898 12752 47900
rect 12776 47898 12832 47900
rect 12856 47898 12912 47900
rect 12616 47846 12662 47898
rect 12662 47846 12672 47898
rect 12696 47846 12726 47898
rect 12726 47846 12738 47898
rect 12738 47846 12752 47898
rect 12776 47846 12790 47898
rect 12790 47846 12802 47898
rect 12802 47846 12832 47898
rect 12856 47846 12866 47898
rect 12866 47846 12912 47898
rect 12616 47844 12672 47846
rect 12696 47844 12752 47846
rect 12776 47844 12832 47846
rect 12856 47844 12912 47846
rect 12616 46810 12672 46812
rect 12696 46810 12752 46812
rect 12776 46810 12832 46812
rect 12856 46810 12912 46812
rect 12616 46758 12662 46810
rect 12662 46758 12672 46810
rect 12696 46758 12726 46810
rect 12726 46758 12738 46810
rect 12738 46758 12752 46810
rect 12776 46758 12790 46810
rect 12790 46758 12802 46810
rect 12802 46758 12832 46810
rect 12856 46758 12866 46810
rect 12866 46758 12912 46810
rect 12616 46756 12672 46758
rect 12696 46756 12752 46758
rect 12776 46756 12832 46758
rect 12856 46756 12912 46758
rect 11956 46266 12012 46268
rect 12036 46266 12092 46268
rect 12116 46266 12172 46268
rect 12196 46266 12252 46268
rect 11956 46214 12002 46266
rect 12002 46214 12012 46266
rect 12036 46214 12066 46266
rect 12066 46214 12078 46266
rect 12078 46214 12092 46266
rect 12116 46214 12130 46266
rect 12130 46214 12142 46266
rect 12142 46214 12172 46266
rect 12196 46214 12206 46266
rect 12206 46214 12252 46266
rect 11956 46212 12012 46214
rect 12036 46212 12092 46214
rect 12116 46212 12172 46214
rect 12196 46212 12252 46214
rect 12616 45722 12672 45724
rect 12696 45722 12752 45724
rect 12776 45722 12832 45724
rect 12856 45722 12912 45724
rect 12616 45670 12662 45722
rect 12662 45670 12672 45722
rect 12696 45670 12726 45722
rect 12726 45670 12738 45722
rect 12738 45670 12752 45722
rect 12776 45670 12790 45722
rect 12790 45670 12802 45722
rect 12802 45670 12832 45722
rect 12856 45670 12866 45722
rect 12866 45670 12912 45722
rect 12616 45668 12672 45670
rect 12696 45668 12752 45670
rect 12776 45668 12832 45670
rect 12856 45668 12912 45670
rect 11956 45178 12012 45180
rect 12036 45178 12092 45180
rect 12116 45178 12172 45180
rect 12196 45178 12252 45180
rect 11956 45126 12002 45178
rect 12002 45126 12012 45178
rect 12036 45126 12066 45178
rect 12066 45126 12078 45178
rect 12078 45126 12092 45178
rect 12116 45126 12130 45178
rect 12130 45126 12142 45178
rect 12142 45126 12172 45178
rect 12196 45126 12206 45178
rect 12206 45126 12252 45178
rect 11956 45124 12012 45126
rect 12036 45124 12092 45126
rect 12116 45124 12172 45126
rect 12196 45124 12252 45126
rect 12616 44634 12672 44636
rect 12696 44634 12752 44636
rect 12776 44634 12832 44636
rect 12856 44634 12912 44636
rect 12616 44582 12662 44634
rect 12662 44582 12672 44634
rect 12696 44582 12726 44634
rect 12726 44582 12738 44634
rect 12738 44582 12752 44634
rect 12776 44582 12790 44634
rect 12790 44582 12802 44634
rect 12802 44582 12832 44634
rect 12856 44582 12866 44634
rect 12866 44582 12912 44634
rect 12616 44580 12672 44582
rect 12696 44580 12752 44582
rect 12776 44580 12832 44582
rect 12856 44580 12912 44582
rect 11956 44090 12012 44092
rect 12036 44090 12092 44092
rect 12116 44090 12172 44092
rect 12196 44090 12252 44092
rect 11956 44038 12002 44090
rect 12002 44038 12012 44090
rect 12036 44038 12066 44090
rect 12066 44038 12078 44090
rect 12078 44038 12092 44090
rect 12116 44038 12130 44090
rect 12130 44038 12142 44090
rect 12142 44038 12172 44090
rect 12196 44038 12206 44090
rect 12206 44038 12252 44090
rect 11956 44036 12012 44038
rect 12036 44036 12092 44038
rect 12116 44036 12172 44038
rect 12196 44036 12252 44038
rect 12616 43546 12672 43548
rect 12696 43546 12752 43548
rect 12776 43546 12832 43548
rect 12856 43546 12912 43548
rect 12616 43494 12662 43546
rect 12662 43494 12672 43546
rect 12696 43494 12726 43546
rect 12726 43494 12738 43546
rect 12738 43494 12752 43546
rect 12776 43494 12790 43546
rect 12790 43494 12802 43546
rect 12802 43494 12832 43546
rect 12856 43494 12866 43546
rect 12866 43494 12912 43546
rect 12616 43492 12672 43494
rect 12696 43492 12752 43494
rect 12776 43492 12832 43494
rect 12856 43492 12912 43494
rect 11956 43002 12012 43004
rect 12036 43002 12092 43004
rect 12116 43002 12172 43004
rect 12196 43002 12252 43004
rect 11956 42950 12002 43002
rect 12002 42950 12012 43002
rect 12036 42950 12066 43002
rect 12066 42950 12078 43002
rect 12078 42950 12092 43002
rect 12116 42950 12130 43002
rect 12130 42950 12142 43002
rect 12142 42950 12172 43002
rect 12196 42950 12206 43002
rect 12206 42950 12252 43002
rect 11956 42948 12012 42950
rect 12036 42948 12092 42950
rect 12116 42948 12172 42950
rect 12196 42948 12252 42950
rect 11610 42744 11666 42800
rect 11150 26152 11206 26208
rect 11058 26016 11114 26072
rect 11426 20984 11482 21040
rect 10690 12180 10692 12200
rect 10692 12180 10744 12200
rect 10744 12180 10746 12200
rect 10690 12144 10746 12180
rect 11956 41914 12012 41916
rect 12036 41914 12092 41916
rect 12116 41914 12172 41916
rect 12196 41914 12252 41916
rect 11956 41862 12002 41914
rect 12002 41862 12012 41914
rect 12036 41862 12066 41914
rect 12066 41862 12078 41914
rect 12078 41862 12092 41914
rect 12116 41862 12130 41914
rect 12130 41862 12142 41914
rect 12142 41862 12172 41914
rect 12196 41862 12206 41914
rect 12206 41862 12252 41914
rect 11956 41860 12012 41862
rect 12036 41860 12092 41862
rect 12116 41860 12172 41862
rect 12196 41860 12252 41862
rect 12616 42458 12672 42460
rect 12696 42458 12752 42460
rect 12776 42458 12832 42460
rect 12856 42458 12912 42460
rect 12616 42406 12662 42458
rect 12662 42406 12672 42458
rect 12696 42406 12726 42458
rect 12726 42406 12738 42458
rect 12738 42406 12752 42458
rect 12776 42406 12790 42458
rect 12790 42406 12802 42458
rect 12802 42406 12832 42458
rect 12856 42406 12866 42458
rect 12866 42406 12912 42458
rect 12616 42404 12672 42406
rect 12696 42404 12752 42406
rect 12776 42404 12832 42406
rect 12856 42404 12912 42406
rect 11956 40826 12012 40828
rect 12036 40826 12092 40828
rect 12116 40826 12172 40828
rect 12196 40826 12252 40828
rect 11956 40774 12002 40826
rect 12002 40774 12012 40826
rect 12036 40774 12066 40826
rect 12066 40774 12078 40826
rect 12078 40774 12092 40826
rect 12116 40774 12130 40826
rect 12130 40774 12142 40826
rect 12142 40774 12172 40826
rect 12196 40774 12206 40826
rect 12206 40774 12252 40826
rect 11956 40772 12012 40774
rect 12036 40772 12092 40774
rect 12116 40772 12172 40774
rect 12196 40772 12252 40774
rect 11956 39738 12012 39740
rect 12036 39738 12092 39740
rect 12116 39738 12172 39740
rect 12196 39738 12252 39740
rect 11956 39686 12002 39738
rect 12002 39686 12012 39738
rect 12036 39686 12066 39738
rect 12066 39686 12078 39738
rect 12078 39686 12092 39738
rect 12116 39686 12130 39738
rect 12130 39686 12142 39738
rect 12142 39686 12172 39738
rect 12196 39686 12206 39738
rect 12206 39686 12252 39738
rect 11956 39684 12012 39686
rect 12036 39684 12092 39686
rect 12116 39684 12172 39686
rect 12196 39684 12252 39686
rect 11956 38650 12012 38652
rect 12036 38650 12092 38652
rect 12116 38650 12172 38652
rect 12196 38650 12252 38652
rect 11956 38598 12002 38650
rect 12002 38598 12012 38650
rect 12036 38598 12066 38650
rect 12066 38598 12078 38650
rect 12078 38598 12092 38650
rect 12116 38598 12130 38650
rect 12130 38598 12142 38650
rect 12142 38598 12172 38650
rect 12196 38598 12206 38650
rect 12206 38598 12252 38650
rect 11956 38596 12012 38598
rect 12036 38596 12092 38598
rect 12116 38596 12172 38598
rect 12196 38596 12252 38598
rect 11956 37562 12012 37564
rect 12036 37562 12092 37564
rect 12116 37562 12172 37564
rect 12196 37562 12252 37564
rect 11956 37510 12002 37562
rect 12002 37510 12012 37562
rect 12036 37510 12066 37562
rect 12066 37510 12078 37562
rect 12078 37510 12092 37562
rect 12116 37510 12130 37562
rect 12130 37510 12142 37562
rect 12142 37510 12172 37562
rect 12196 37510 12206 37562
rect 12206 37510 12252 37562
rect 11956 37508 12012 37510
rect 12036 37508 12092 37510
rect 12116 37508 12172 37510
rect 12196 37508 12252 37510
rect 11956 36474 12012 36476
rect 12036 36474 12092 36476
rect 12116 36474 12172 36476
rect 12196 36474 12252 36476
rect 11956 36422 12002 36474
rect 12002 36422 12012 36474
rect 12036 36422 12066 36474
rect 12066 36422 12078 36474
rect 12078 36422 12092 36474
rect 12116 36422 12130 36474
rect 12130 36422 12142 36474
rect 12142 36422 12172 36474
rect 12196 36422 12206 36474
rect 12206 36422 12252 36474
rect 11956 36420 12012 36422
rect 12036 36420 12092 36422
rect 12116 36420 12172 36422
rect 12196 36420 12252 36422
rect 11956 35386 12012 35388
rect 12036 35386 12092 35388
rect 12116 35386 12172 35388
rect 12196 35386 12252 35388
rect 11956 35334 12002 35386
rect 12002 35334 12012 35386
rect 12036 35334 12066 35386
rect 12066 35334 12078 35386
rect 12078 35334 12092 35386
rect 12116 35334 12130 35386
rect 12130 35334 12142 35386
rect 12142 35334 12172 35386
rect 12196 35334 12206 35386
rect 12206 35334 12252 35386
rect 11956 35332 12012 35334
rect 12036 35332 12092 35334
rect 12116 35332 12172 35334
rect 12196 35332 12252 35334
rect 11956 34298 12012 34300
rect 12036 34298 12092 34300
rect 12116 34298 12172 34300
rect 12196 34298 12252 34300
rect 11956 34246 12002 34298
rect 12002 34246 12012 34298
rect 12036 34246 12066 34298
rect 12066 34246 12078 34298
rect 12078 34246 12092 34298
rect 12116 34246 12130 34298
rect 12130 34246 12142 34298
rect 12142 34246 12172 34298
rect 12196 34246 12206 34298
rect 12206 34246 12252 34298
rect 11956 34244 12012 34246
rect 12036 34244 12092 34246
rect 12116 34244 12172 34246
rect 12196 34244 12252 34246
rect 11956 33210 12012 33212
rect 12036 33210 12092 33212
rect 12116 33210 12172 33212
rect 12196 33210 12252 33212
rect 11956 33158 12002 33210
rect 12002 33158 12012 33210
rect 12036 33158 12066 33210
rect 12066 33158 12078 33210
rect 12078 33158 12092 33210
rect 12116 33158 12130 33210
rect 12130 33158 12142 33210
rect 12142 33158 12172 33210
rect 12196 33158 12206 33210
rect 12206 33158 12252 33210
rect 11956 33156 12012 33158
rect 12036 33156 12092 33158
rect 12116 33156 12172 33158
rect 12196 33156 12252 33158
rect 11956 32122 12012 32124
rect 12036 32122 12092 32124
rect 12116 32122 12172 32124
rect 12196 32122 12252 32124
rect 11956 32070 12002 32122
rect 12002 32070 12012 32122
rect 12036 32070 12066 32122
rect 12066 32070 12078 32122
rect 12078 32070 12092 32122
rect 12116 32070 12130 32122
rect 12130 32070 12142 32122
rect 12142 32070 12172 32122
rect 12196 32070 12206 32122
rect 12206 32070 12252 32122
rect 11956 32068 12012 32070
rect 12036 32068 12092 32070
rect 12116 32068 12172 32070
rect 12196 32068 12252 32070
rect 11956 31034 12012 31036
rect 12036 31034 12092 31036
rect 12116 31034 12172 31036
rect 12196 31034 12252 31036
rect 11956 30982 12002 31034
rect 12002 30982 12012 31034
rect 12036 30982 12066 31034
rect 12066 30982 12078 31034
rect 12078 30982 12092 31034
rect 12116 30982 12130 31034
rect 12130 30982 12142 31034
rect 12142 30982 12172 31034
rect 12196 30982 12206 31034
rect 12206 30982 12252 31034
rect 11956 30980 12012 30982
rect 12036 30980 12092 30982
rect 12116 30980 12172 30982
rect 12196 30980 12252 30982
rect 11956 29946 12012 29948
rect 12036 29946 12092 29948
rect 12116 29946 12172 29948
rect 12196 29946 12252 29948
rect 11956 29894 12002 29946
rect 12002 29894 12012 29946
rect 12036 29894 12066 29946
rect 12066 29894 12078 29946
rect 12078 29894 12092 29946
rect 12116 29894 12130 29946
rect 12130 29894 12142 29946
rect 12142 29894 12172 29946
rect 12196 29894 12206 29946
rect 12206 29894 12252 29946
rect 11956 29892 12012 29894
rect 12036 29892 12092 29894
rect 12116 29892 12172 29894
rect 12196 29892 12252 29894
rect 11956 28858 12012 28860
rect 12036 28858 12092 28860
rect 12116 28858 12172 28860
rect 12196 28858 12252 28860
rect 11956 28806 12002 28858
rect 12002 28806 12012 28858
rect 12036 28806 12066 28858
rect 12066 28806 12078 28858
rect 12078 28806 12092 28858
rect 12116 28806 12130 28858
rect 12130 28806 12142 28858
rect 12142 28806 12172 28858
rect 12196 28806 12206 28858
rect 12206 28806 12252 28858
rect 11956 28804 12012 28806
rect 12036 28804 12092 28806
rect 12116 28804 12172 28806
rect 12196 28804 12252 28806
rect 11956 27770 12012 27772
rect 12036 27770 12092 27772
rect 12116 27770 12172 27772
rect 12196 27770 12252 27772
rect 11956 27718 12002 27770
rect 12002 27718 12012 27770
rect 12036 27718 12066 27770
rect 12066 27718 12078 27770
rect 12078 27718 12092 27770
rect 12116 27718 12130 27770
rect 12130 27718 12142 27770
rect 12142 27718 12172 27770
rect 12196 27718 12206 27770
rect 12206 27718 12252 27770
rect 11956 27716 12012 27718
rect 12036 27716 12092 27718
rect 12116 27716 12172 27718
rect 12196 27716 12252 27718
rect 11956 26682 12012 26684
rect 12036 26682 12092 26684
rect 12116 26682 12172 26684
rect 12196 26682 12252 26684
rect 11956 26630 12002 26682
rect 12002 26630 12012 26682
rect 12036 26630 12066 26682
rect 12066 26630 12078 26682
rect 12078 26630 12092 26682
rect 12116 26630 12130 26682
rect 12130 26630 12142 26682
rect 12142 26630 12172 26682
rect 12196 26630 12206 26682
rect 12206 26630 12252 26682
rect 11956 26628 12012 26630
rect 12036 26628 12092 26630
rect 12116 26628 12172 26630
rect 12196 26628 12252 26630
rect 11956 25594 12012 25596
rect 12036 25594 12092 25596
rect 12116 25594 12172 25596
rect 12196 25594 12252 25596
rect 11956 25542 12002 25594
rect 12002 25542 12012 25594
rect 12036 25542 12066 25594
rect 12066 25542 12078 25594
rect 12078 25542 12092 25594
rect 12116 25542 12130 25594
rect 12130 25542 12142 25594
rect 12142 25542 12172 25594
rect 12196 25542 12206 25594
rect 12206 25542 12252 25594
rect 11956 25540 12012 25542
rect 12036 25540 12092 25542
rect 12116 25540 12172 25542
rect 12196 25540 12252 25542
rect 11956 24506 12012 24508
rect 12036 24506 12092 24508
rect 12116 24506 12172 24508
rect 12196 24506 12252 24508
rect 11956 24454 12002 24506
rect 12002 24454 12012 24506
rect 12036 24454 12066 24506
rect 12066 24454 12078 24506
rect 12078 24454 12092 24506
rect 12116 24454 12130 24506
rect 12130 24454 12142 24506
rect 12142 24454 12172 24506
rect 12196 24454 12206 24506
rect 12206 24454 12252 24506
rect 11956 24452 12012 24454
rect 12036 24452 12092 24454
rect 12116 24452 12172 24454
rect 12196 24452 12252 24454
rect 11956 23418 12012 23420
rect 12036 23418 12092 23420
rect 12116 23418 12172 23420
rect 12196 23418 12252 23420
rect 11956 23366 12002 23418
rect 12002 23366 12012 23418
rect 12036 23366 12066 23418
rect 12066 23366 12078 23418
rect 12078 23366 12092 23418
rect 12116 23366 12130 23418
rect 12130 23366 12142 23418
rect 12142 23366 12172 23418
rect 12196 23366 12206 23418
rect 12206 23366 12252 23418
rect 11956 23364 12012 23366
rect 12036 23364 12092 23366
rect 12116 23364 12172 23366
rect 12196 23364 12252 23366
rect 11956 22330 12012 22332
rect 12036 22330 12092 22332
rect 12116 22330 12172 22332
rect 12196 22330 12252 22332
rect 11956 22278 12002 22330
rect 12002 22278 12012 22330
rect 12036 22278 12066 22330
rect 12066 22278 12078 22330
rect 12078 22278 12092 22330
rect 12116 22278 12130 22330
rect 12130 22278 12142 22330
rect 12142 22278 12172 22330
rect 12196 22278 12206 22330
rect 12206 22278 12252 22330
rect 11956 22276 12012 22278
rect 12036 22276 12092 22278
rect 12116 22276 12172 22278
rect 12196 22276 12252 22278
rect 12616 41370 12672 41372
rect 12696 41370 12752 41372
rect 12776 41370 12832 41372
rect 12856 41370 12912 41372
rect 12616 41318 12662 41370
rect 12662 41318 12672 41370
rect 12696 41318 12726 41370
rect 12726 41318 12738 41370
rect 12738 41318 12752 41370
rect 12776 41318 12790 41370
rect 12790 41318 12802 41370
rect 12802 41318 12832 41370
rect 12856 41318 12866 41370
rect 12866 41318 12912 41370
rect 12616 41316 12672 41318
rect 12696 41316 12752 41318
rect 12776 41316 12832 41318
rect 12856 41316 12912 41318
rect 12616 40282 12672 40284
rect 12696 40282 12752 40284
rect 12776 40282 12832 40284
rect 12856 40282 12912 40284
rect 12616 40230 12662 40282
rect 12662 40230 12672 40282
rect 12696 40230 12726 40282
rect 12726 40230 12738 40282
rect 12738 40230 12752 40282
rect 12776 40230 12790 40282
rect 12790 40230 12802 40282
rect 12802 40230 12832 40282
rect 12856 40230 12866 40282
rect 12866 40230 12912 40282
rect 12616 40228 12672 40230
rect 12696 40228 12752 40230
rect 12776 40228 12832 40230
rect 12856 40228 12912 40230
rect 12438 35536 12494 35592
rect 12616 39194 12672 39196
rect 12696 39194 12752 39196
rect 12776 39194 12832 39196
rect 12856 39194 12912 39196
rect 12616 39142 12662 39194
rect 12662 39142 12672 39194
rect 12696 39142 12726 39194
rect 12726 39142 12738 39194
rect 12738 39142 12752 39194
rect 12776 39142 12790 39194
rect 12790 39142 12802 39194
rect 12802 39142 12832 39194
rect 12856 39142 12866 39194
rect 12866 39142 12912 39194
rect 12616 39140 12672 39142
rect 12696 39140 12752 39142
rect 12776 39140 12832 39142
rect 12856 39140 12912 39142
rect 12616 38106 12672 38108
rect 12696 38106 12752 38108
rect 12776 38106 12832 38108
rect 12856 38106 12912 38108
rect 12616 38054 12662 38106
rect 12662 38054 12672 38106
rect 12696 38054 12726 38106
rect 12726 38054 12738 38106
rect 12738 38054 12752 38106
rect 12776 38054 12790 38106
rect 12790 38054 12802 38106
rect 12802 38054 12832 38106
rect 12856 38054 12866 38106
rect 12866 38054 12912 38106
rect 12616 38052 12672 38054
rect 12696 38052 12752 38054
rect 12776 38052 12832 38054
rect 12856 38052 12912 38054
rect 12616 37018 12672 37020
rect 12696 37018 12752 37020
rect 12776 37018 12832 37020
rect 12856 37018 12912 37020
rect 12616 36966 12662 37018
rect 12662 36966 12672 37018
rect 12696 36966 12726 37018
rect 12726 36966 12738 37018
rect 12738 36966 12752 37018
rect 12776 36966 12790 37018
rect 12790 36966 12802 37018
rect 12802 36966 12832 37018
rect 12856 36966 12866 37018
rect 12866 36966 12912 37018
rect 12616 36964 12672 36966
rect 12696 36964 12752 36966
rect 12776 36964 12832 36966
rect 12856 36964 12912 36966
rect 12616 35930 12672 35932
rect 12696 35930 12752 35932
rect 12776 35930 12832 35932
rect 12856 35930 12912 35932
rect 12616 35878 12662 35930
rect 12662 35878 12672 35930
rect 12696 35878 12726 35930
rect 12726 35878 12738 35930
rect 12738 35878 12752 35930
rect 12776 35878 12790 35930
rect 12790 35878 12802 35930
rect 12802 35878 12832 35930
rect 12856 35878 12866 35930
rect 12866 35878 12912 35930
rect 12616 35876 12672 35878
rect 12696 35876 12752 35878
rect 12776 35876 12832 35878
rect 12856 35876 12912 35878
rect 12616 34842 12672 34844
rect 12696 34842 12752 34844
rect 12776 34842 12832 34844
rect 12856 34842 12912 34844
rect 12616 34790 12662 34842
rect 12662 34790 12672 34842
rect 12696 34790 12726 34842
rect 12726 34790 12738 34842
rect 12738 34790 12752 34842
rect 12776 34790 12790 34842
rect 12790 34790 12802 34842
rect 12802 34790 12832 34842
rect 12856 34790 12866 34842
rect 12866 34790 12912 34842
rect 12616 34788 12672 34790
rect 12696 34788 12752 34790
rect 12776 34788 12832 34790
rect 12856 34788 12912 34790
rect 12616 33754 12672 33756
rect 12696 33754 12752 33756
rect 12776 33754 12832 33756
rect 12856 33754 12912 33756
rect 12616 33702 12662 33754
rect 12662 33702 12672 33754
rect 12696 33702 12726 33754
rect 12726 33702 12738 33754
rect 12738 33702 12752 33754
rect 12776 33702 12790 33754
rect 12790 33702 12802 33754
rect 12802 33702 12832 33754
rect 12856 33702 12866 33754
rect 12866 33702 12912 33754
rect 12616 33700 12672 33702
rect 12696 33700 12752 33702
rect 12776 33700 12832 33702
rect 12856 33700 12912 33702
rect 12616 32666 12672 32668
rect 12696 32666 12752 32668
rect 12776 32666 12832 32668
rect 12856 32666 12912 32668
rect 12616 32614 12662 32666
rect 12662 32614 12672 32666
rect 12696 32614 12726 32666
rect 12726 32614 12738 32666
rect 12738 32614 12752 32666
rect 12776 32614 12790 32666
rect 12790 32614 12802 32666
rect 12802 32614 12832 32666
rect 12856 32614 12866 32666
rect 12866 32614 12912 32666
rect 12616 32612 12672 32614
rect 12696 32612 12752 32614
rect 12776 32612 12832 32614
rect 12856 32612 12912 32614
rect 12616 31578 12672 31580
rect 12696 31578 12752 31580
rect 12776 31578 12832 31580
rect 12856 31578 12912 31580
rect 12616 31526 12662 31578
rect 12662 31526 12672 31578
rect 12696 31526 12726 31578
rect 12726 31526 12738 31578
rect 12738 31526 12752 31578
rect 12776 31526 12790 31578
rect 12790 31526 12802 31578
rect 12802 31526 12832 31578
rect 12856 31526 12866 31578
rect 12866 31526 12912 31578
rect 12616 31524 12672 31526
rect 12696 31524 12752 31526
rect 12776 31524 12832 31526
rect 12856 31524 12912 31526
rect 12616 30490 12672 30492
rect 12696 30490 12752 30492
rect 12776 30490 12832 30492
rect 12856 30490 12912 30492
rect 12616 30438 12662 30490
rect 12662 30438 12672 30490
rect 12696 30438 12726 30490
rect 12726 30438 12738 30490
rect 12738 30438 12752 30490
rect 12776 30438 12790 30490
rect 12790 30438 12802 30490
rect 12802 30438 12832 30490
rect 12856 30438 12866 30490
rect 12866 30438 12912 30490
rect 12616 30436 12672 30438
rect 12696 30436 12752 30438
rect 12776 30436 12832 30438
rect 12856 30436 12912 30438
rect 12616 29402 12672 29404
rect 12696 29402 12752 29404
rect 12776 29402 12832 29404
rect 12856 29402 12912 29404
rect 12616 29350 12662 29402
rect 12662 29350 12672 29402
rect 12696 29350 12726 29402
rect 12726 29350 12738 29402
rect 12738 29350 12752 29402
rect 12776 29350 12790 29402
rect 12790 29350 12802 29402
rect 12802 29350 12832 29402
rect 12856 29350 12866 29402
rect 12866 29350 12912 29402
rect 12616 29348 12672 29350
rect 12696 29348 12752 29350
rect 12776 29348 12832 29350
rect 12856 29348 12912 29350
rect 12616 28314 12672 28316
rect 12696 28314 12752 28316
rect 12776 28314 12832 28316
rect 12856 28314 12912 28316
rect 12616 28262 12662 28314
rect 12662 28262 12672 28314
rect 12696 28262 12726 28314
rect 12726 28262 12738 28314
rect 12738 28262 12752 28314
rect 12776 28262 12790 28314
rect 12790 28262 12802 28314
rect 12802 28262 12832 28314
rect 12856 28262 12866 28314
rect 12866 28262 12912 28314
rect 12616 28260 12672 28262
rect 12696 28260 12752 28262
rect 12776 28260 12832 28262
rect 12856 28260 12912 28262
rect 12616 27226 12672 27228
rect 12696 27226 12752 27228
rect 12776 27226 12832 27228
rect 12856 27226 12912 27228
rect 12616 27174 12662 27226
rect 12662 27174 12672 27226
rect 12696 27174 12726 27226
rect 12726 27174 12738 27226
rect 12738 27174 12752 27226
rect 12776 27174 12790 27226
rect 12790 27174 12802 27226
rect 12802 27174 12832 27226
rect 12856 27174 12866 27226
rect 12866 27174 12912 27226
rect 12616 27172 12672 27174
rect 12696 27172 12752 27174
rect 12776 27172 12832 27174
rect 12856 27172 12912 27174
rect 12616 26138 12672 26140
rect 12696 26138 12752 26140
rect 12776 26138 12832 26140
rect 12856 26138 12912 26140
rect 12616 26086 12662 26138
rect 12662 26086 12672 26138
rect 12696 26086 12726 26138
rect 12726 26086 12738 26138
rect 12738 26086 12752 26138
rect 12776 26086 12790 26138
rect 12790 26086 12802 26138
rect 12802 26086 12832 26138
rect 12856 26086 12866 26138
rect 12866 26086 12912 26138
rect 12616 26084 12672 26086
rect 12696 26084 12752 26086
rect 12776 26084 12832 26086
rect 12856 26084 12912 26086
rect 12616 25050 12672 25052
rect 12696 25050 12752 25052
rect 12776 25050 12832 25052
rect 12856 25050 12912 25052
rect 12616 24998 12662 25050
rect 12662 24998 12672 25050
rect 12696 24998 12726 25050
rect 12726 24998 12738 25050
rect 12738 24998 12752 25050
rect 12776 24998 12790 25050
rect 12790 24998 12802 25050
rect 12802 24998 12832 25050
rect 12856 24998 12866 25050
rect 12866 24998 12912 25050
rect 12616 24996 12672 24998
rect 12696 24996 12752 24998
rect 12776 24996 12832 24998
rect 12856 24996 12912 24998
rect 12616 23962 12672 23964
rect 12696 23962 12752 23964
rect 12776 23962 12832 23964
rect 12856 23962 12912 23964
rect 12616 23910 12662 23962
rect 12662 23910 12672 23962
rect 12696 23910 12726 23962
rect 12726 23910 12738 23962
rect 12738 23910 12752 23962
rect 12776 23910 12790 23962
rect 12790 23910 12802 23962
rect 12802 23910 12832 23962
rect 12856 23910 12866 23962
rect 12866 23910 12912 23962
rect 12616 23908 12672 23910
rect 12696 23908 12752 23910
rect 12776 23908 12832 23910
rect 12856 23908 12912 23910
rect 11956 21242 12012 21244
rect 12036 21242 12092 21244
rect 12116 21242 12172 21244
rect 12196 21242 12252 21244
rect 11956 21190 12002 21242
rect 12002 21190 12012 21242
rect 12036 21190 12066 21242
rect 12066 21190 12078 21242
rect 12078 21190 12092 21242
rect 12116 21190 12130 21242
rect 12130 21190 12142 21242
rect 12142 21190 12172 21242
rect 12196 21190 12206 21242
rect 12206 21190 12252 21242
rect 11956 21188 12012 21190
rect 12036 21188 12092 21190
rect 12116 21188 12172 21190
rect 12196 21188 12252 21190
rect 11956 20154 12012 20156
rect 12036 20154 12092 20156
rect 12116 20154 12172 20156
rect 12196 20154 12252 20156
rect 11956 20102 12002 20154
rect 12002 20102 12012 20154
rect 12036 20102 12066 20154
rect 12066 20102 12078 20154
rect 12078 20102 12092 20154
rect 12116 20102 12130 20154
rect 12130 20102 12142 20154
rect 12142 20102 12172 20154
rect 12196 20102 12206 20154
rect 12206 20102 12252 20154
rect 11956 20100 12012 20102
rect 12036 20100 12092 20102
rect 12116 20100 12172 20102
rect 12196 20100 12252 20102
rect 12162 19896 12218 19952
rect 11956 19066 12012 19068
rect 12036 19066 12092 19068
rect 12116 19066 12172 19068
rect 12196 19066 12252 19068
rect 11956 19014 12002 19066
rect 12002 19014 12012 19066
rect 12036 19014 12066 19066
rect 12066 19014 12078 19066
rect 12078 19014 12092 19066
rect 12116 19014 12130 19066
rect 12130 19014 12142 19066
rect 12142 19014 12172 19066
rect 12196 19014 12206 19066
rect 12206 19014 12252 19066
rect 11956 19012 12012 19014
rect 12036 19012 12092 19014
rect 12116 19012 12172 19014
rect 12196 19012 12252 19014
rect 11956 17978 12012 17980
rect 12036 17978 12092 17980
rect 12116 17978 12172 17980
rect 12196 17978 12252 17980
rect 11956 17926 12002 17978
rect 12002 17926 12012 17978
rect 12036 17926 12066 17978
rect 12066 17926 12078 17978
rect 12078 17926 12092 17978
rect 12116 17926 12130 17978
rect 12130 17926 12142 17978
rect 12142 17926 12172 17978
rect 12196 17926 12206 17978
rect 12206 17926 12252 17978
rect 11956 17924 12012 17926
rect 12036 17924 12092 17926
rect 12116 17924 12172 17926
rect 12196 17924 12252 17926
rect 12616 22874 12672 22876
rect 12696 22874 12752 22876
rect 12776 22874 12832 22876
rect 12856 22874 12912 22876
rect 12616 22822 12662 22874
rect 12662 22822 12672 22874
rect 12696 22822 12726 22874
rect 12726 22822 12738 22874
rect 12738 22822 12752 22874
rect 12776 22822 12790 22874
rect 12790 22822 12802 22874
rect 12802 22822 12832 22874
rect 12856 22822 12866 22874
rect 12866 22822 12912 22874
rect 12616 22820 12672 22822
rect 12696 22820 12752 22822
rect 12776 22820 12832 22822
rect 12856 22820 12912 22822
rect 12616 21786 12672 21788
rect 12696 21786 12752 21788
rect 12776 21786 12832 21788
rect 12856 21786 12912 21788
rect 12616 21734 12662 21786
rect 12662 21734 12672 21786
rect 12696 21734 12726 21786
rect 12726 21734 12738 21786
rect 12738 21734 12752 21786
rect 12776 21734 12790 21786
rect 12790 21734 12802 21786
rect 12802 21734 12832 21786
rect 12856 21734 12866 21786
rect 12866 21734 12912 21786
rect 12616 21732 12672 21734
rect 12696 21732 12752 21734
rect 12776 21732 12832 21734
rect 12856 21732 12912 21734
rect 13726 58828 13728 58848
rect 13728 58828 13780 58848
rect 13780 58828 13782 58848
rect 13726 58792 13782 58828
rect 12616 20698 12672 20700
rect 12696 20698 12752 20700
rect 12776 20698 12832 20700
rect 12856 20698 12912 20700
rect 12616 20646 12662 20698
rect 12662 20646 12672 20698
rect 12696 20646 12726 20698
rect 12726 20646 12738 20698
rect 12738 20646 12752 20698
rect 12776 20646 12790 20698
rect 12790 20646 12802 20698
rect 12802 20646 12832 20698
rect 12856 20646 12866 20698
rect 12866 20646 12912 20698
rect 12616 20644 12672 20646
rect 12696 20644 12752 20646
rect 12776 20644 12832 20646
rect 12856 20644 12912 20646
rect 12616 19610 12672 19612
rect 12696 19610 12752 19612
rect 12776 19610 12832 19612
rect 12856 19610 12912 19612
rect 12616 19558 12662 19610
rect 12662 19558 12672 19610
rect 12696 19558 12726 19610
rect 12726 19558 12738 19610
rect 12738 19558 12752 19610
rect 12776 19558 12790 19610
rect 12790 19558 12802 19610
rect 12802 19558 12832 19610
rect 12856 19558 12866 19610
rect 12866 19558 12912 19610
rect 12616 19556 12672 19558
rect 12696 19556 12752 19558
rect 12776 19556 12832 19558
rect 12856 19556 12912 19558
rect 12616 18522 12672 18524
rect 12696 18522 12752 18524
rect 12776 18522 12832 18524
rect 12856 18522 12912 18524
rect 12616 18470 12662 18522
rect 12662 18470 12672 18522
rect 12696 18470 12726 18522
rect 12726 18470 12738 18522
rect 12738 18470 12752 18522
rect 12776 18470 12790 18522
rect 12790 18470 12802 18522
rect 12802 18470 12832 18522
rect 12856 18470 12866 18522
rect 12866 18470 12912 18522
rect 12616 18468 12672 18470
rect 12696 18468 12752 18470
rect 12776 18468 12832 18470
rect 12856 18468 12912 18470
rect 12616 17434 12672 17436
rect 12696 17434 12752 17436
rect 12776 17434 12832 17436
rect 12856 17434 12912 17436
rect 12616 17382 12662 17434
rect 12662 17382 12672 17434
rect 12696 17382 12726 17434
rect 12726 17382 12738 17434
rect 12738 17382 12752 17434
rect 12776 17382 12790 17434
rect 12790 17382 12802 17434
rect 12802 17382 12832 17434
rect 12856 17382 12866 17434
rect 12866 17382 12912 17434
rect 12616 17380 12672 17382
rect 12696 17380 12752 17382
rect 12776 17380 12832 17382
rect 12856 17380 12912 17382
rect 11956 16890 12012 16892
rect 12036 16890 12092 16892
rect 12116 16890 12172 16892
rect 12196 16890 12252 16892
rect 11956 16838 12002 16890
rect 12002 16838 12012 16890
rect 12036 16838 12066 16890
rect 12066 16838 12078 16890
rect 12078 16838 12092 16890
rect 12116 16838 12130 16890
rect 12130 16838 12142 16890
rect 12142 16838 12172 16890
rect 12196 16838 12206 16890
rect 12206 16838 12252 16890
rect 11956 16836 12012 16838
rect 12036 16836 12092 16838
rect 12116 16836 12172 16838
rect 12196 16836 12252 16838
rect 12616 16346 12672 16348
rect 12696 16346 12752 16348
rect 12776 16346 12832 16348
rect 12856 16346 12912 16348
rect 12616 16294 12662 16346
rect 12662 16294 12672 16346
rect 12696 16294 12726 16346
rect 12726 16294 12738 16346
rect 12738 16294 12752 16346
rect 12776 16294 12790 16346
rect 12790 16294 12802 16346
rect 12802 16294 12832 16346
rect 12856 16294 12866 16346
rect 12866 16294 12912 16346
rect 12616 16292 12672 16294
rect 12696 16292 12752 16294
rect 12776 16292 12832 16294
rect 12856 16292 12912 16294
rect 11956 15802 12012 15804
rect 12036 15802 12092 15804
rect 12116 15802 12172 15804
rect 12196 15802 12252 15804
rect 11956 15750 12002 15802
rect 12002 15750 12012 15802
rect 12036 15750 12066 15802
rect 12066 15750 12078 15802
rect 12078 15750 12092 15802
rect 12116 15750 12130 15802
rect 12130 15750 12142 15802
rect 12142 15750 12172 15802
rect 12196 15750 12206 15802
rect 12206 15750 12252 15802
rect 11956 15748 12012 15750
rect 12036 15748 12092 15750
rect 12116 15748 12172 15750
rect 12196 15748 12252 15750
rect 12990 15564 13046 15600
rect 12990 15544 12992 15564
rect 12992 15544 13044 15564
rect 13044 15544 13046 15564
rect 12616 15258 12672 15260
rect 12696 15258 12752 15260
rect 12776 15258 12832 15260
rect 12856 15258 12912 15260
rect 12616 15206 12662 15258
rect 12662 15206 12672 15258
rect 12696 15206 12726 15258
rect 12726 15206 12738 15258
rect 12738 15206 12752 15258
rect 12776 15206 12790 15258
rect 12790 15206 12802 15258
rect 12802 15206 12832 15258
rect 12856 15206 12866 15258
rect 12866 15206 12912 15258
rect 12616 15204 12672 15206
rect 12696 15204 12752 15206
rect 12776 15204 12832 15206
rect 12856 15204 12912 15206
rect 11956 14714 12012 14716
rect 12036 14714 12092 14716
rect 12116 14714 12172 14716
rect 12196 14714 12252 14716
rect 11956 14662 12002 14714
rect 12002 14662 12012 14714
rect 12036 14662 12066 14714
rect 12066 14662 12078 14714
rect 12078 14662 12092 14714
rect 12116 14662 12130 14714
rect 12130 14662 12142 14714
rect 12142 14662 12172 14714
rect 12196 14662 12206 14714
rect 12206 14662 12252 14714
rect 11956 14660 12012 14662
rect 12036 14660 12092 14662
rect 12116 14660 12172 14662
rect 12196 14660 12252 14662
rect 12616 14170 12672 14172
rect 12696 14170 12752 14172
rect 12776 14170 12832 14172
rect 12856 14170 12912 14172
rect 12616 14118 12662 14170
rect 12662 14118 12672 14170
rect 12696 14118 12726 14170
rect 12726 14118 12738 14170
rect 12738 14118 12752 14170
rect 12776 14118 12790 14170
rect 12790 14118 12802 14170
rect 12802 14118 12832 14170
rect 12856 14118 12866 14170
rect 12866 14118 12912 14170
rect 12616 14116 12672 14118
rect 12696 14116 12752 14118
rect 12776 14116 12832 14118
rect 12856 14116 12912 14118
rect 11956 13626 12012 13628
rect 12036 13626 12092 13628
rect 12116 13626 12172 13628
rect 12196 13626 12252 13628
rect 11956 13574 12002 13626
rect 12002 13574 12012 13626
rect 12036 13574 12066 13626
rect 12066 13574 12078 13626
rect 12078 13574 12092 13626
rect 12116 13574 12130 13626
rect 12130 13574 12142 13626
rect 12142 13574 12172 13626
rect 12196 13574 12206 13626
rect 12206 13574 12252 13626
rect 11956 13572 12012 13574
rect 12036 13572 12092 13574
rect 12116 13572 12172 13574
rect 12196 13572 12252 13574
rect 12616 13082 12672 13084
rect 12696 13082 12752 13084
rect 12776 13082 12832 13084
rect 12856 13082 12912 13084
rect 12616 13030 12662 13082
rect 12662 13030 12672 13082
rect 12696 13030 12726 13082
rect 12726 13030 12738 13082
rect 12738 13030 12752 13082
rect 12776 13030 12790 13082
rect 12790 13030 12802 13082
rect 12802 13030 12832 13082
rect 12856 13030 12866 13082
rect 12866 13030 12912 13082
rect 12616 13028 12672 13030
rect 12696 13028 12752 13030
rect 12776 13028 12832 13030
rect 12856 13028 12912 13030
rect 11956 12538 12012 12540
rect 12036 12538 12092 12540
rect 12116 12538 12172 12540
rect 12196 12538 12252 12540
rect 11956 12486 12002 12538
rect 12002 12486 12012 12538
rect 12036 12486 12066 12538
rect 12066 12486 12078 12538
rect 12078 12486 12092 12538
rect 12116 12486 12130 12538
rect 12130 12486 12142 12538
rect 12142 12486 12172 12538
rect 12196 12486 12206 12538
rect 12206 12486 12252 12538
rect 11956 12484 12012 12486
rect 12036 12484 12092 12486
rect 12116 12484 12172 12486
rect 12196 12484 12252 12486
rect 12162 12316 12164 12336
rect 12164 12316 12216 12336
rect 12216 12316 12218 12336
rect 12162 12280 12218 12316
rect 12616 11994 12672 11996
rect 12696 11994 12752 11996
rect 12776 11994 12832 11996
rect 12856 11994 12912 11996
rect 12616 11942 12662 11994
rect 12662 11942 12672 11994
rect 12696 11942 12726 11994
rect 12726 11942 12738 11994
rect 12738 11942 12752 11994
rect 12776 11942 12790 11994
rect 12790 11942 12802 11994
rect 12802 11942 12832 11994
rect 12856 11942 12866 11994
rect 12866 11942 12912 11994
rect 12616 11940 12672 11942
rect 12696 11940 12752 11942
rect 12776 11940 12832 11942
rect 12856 11940 12912 11942
rect 11956 11450 12012 11452
rect 12036 11450 12092 11452
rect 12116 11450 12172 11452
rect 12196 11450 12252 11452
rect 11956 11398 12002 11450
rect 12002 11398 12012 11450
rect 12036 11398 12066 11450
rect 12066 11398 12078 11450
rect 12078 11398 12092 11450
rect 12116 11398 12130 11450
rect 12130 11398 12142 11450
rect 12142 11398 12172 11450
rect 12196 11398 12206 11450
rect 12206 11398 12252 11450
rect 11956 11396 12012 11398
rect 12036 11396 12092 11398
rect 12116 11396 12172 11398
rect 12196 11396 12252 11398
rect 12616 10906 12672 10908
rect 12696 10906 12752 10908
rect 12776 10906 12832 10908
rect 12856 10906 12912 10908
rect 12616 10854 12662 10906
rect 12662 10854 12672 10906
rect 12696 10854 12726 10906
rect 12726 10854 12738 10906
rect 12738 10854 12752 10906
rect 12776 10854 12790 10906
rect 12790 10854 12802 10906
rect 12802 10854 12832 10906
rect 12856 10854 12866 10906
rect 12866 10854 12912 10906
rect 12616 10852 12672 10854
rect 12696 10852 12752 10854
rect 12776 10852 12832 10854
rect 12856 10852 12912 10854
rect 11956 10362 12012 10364
rect 12036 10362 12092 10364
rect 12116 10362 12172 10364
rect 12196 10362 12252 10364
rect 11956 10310 12002 10362
rect 12002 10310 12012 10362
rect 12036 10310 12066 10362
rect 12066 10310 12078 10362
rect 12078 10310 12092 10362
rect 12116 10310 12130 10362
rect 12130 10310 12142 10362
rect 12142 10310 12172 10362
rect 12196 10310 12206 10362
rect 12206 10310 12252 10362
rect 11956 10308 12012 10310
rect 12036 10308 12092 10310
rect 12116 10308 12172 10310
rect 12196 10308 12252 10310
rect 12616 9818 12672 9820
rect 12696 9818 12752 9820
rect 12776 9818 12832 9820
rect 12856 9818 12912 9820
rect 12616 9766 12662 9818
rect 12662 9766 12672 9818
rect 12696 9766 12726 9818
rect 12726 9766 12738 9818
rect 12738 9766 12752 9818
rect 12776 9766 12790 9818
rect 12790 9766 12802 9818
rect 12802 9766 12832 9818
rect 12856 9766 12866 9818
rect 12866 9766 12912 9818
rect 12616 9764 12672 9766
rect 12696 9764 12752 9766
rect 12776 9764 12832 9766
rect 12856 9764 12912 9766
rect 11956 9274 12012 9276
rect 12036 9274 12092 9276
rect 12116 9274 12172 9276
rect 12196 9274 12252 9276
rect 11956 9222 12002 9274
rect 12002 9222 12012 9274
rect 12036 9222 12066 9274
rect 12066 9222 12078 9274
rect 12078 9222 12092 9274
rect 12116 9222 12130 9274
rect 12130 9222 12142 9274
rect 12142 9222 12172 9274
rect 12196 9222 12206 9274
rect 12206 9222 12252 9274
rect 11956 9220 12012 9222
rect 12036 9220 12092 9222
rect 12116 9220 12172 9222
rect 12196 9220 12252 9222
rect 12616 8730 12672 8732
rect 12696 8730 12752 8732
rect 12776 8730 12832 8732
rect 12856 8730 12912 8732
rect 12616 8678 12662 8730
rect 12662 8678 12672 8730
rect 12696 8678 12726 8730
rect 12726 8678 12738 8730
rect 12738 8678 12752 8730
rect 12776 8678 12790 8730
rect 12790 8678 12802 8730
rect 12802 8678 12832 8730
rect 12856 8678 12866 8730
rect 12866 8678 12912 8730
rect 12616 8676 12672 8678
rect 12696 8676 12752 8678
rect 12776 8676 12832 8678
rect 12856 8676 12912 8678
rect 13542 24792 13598 24848
rect 17616 77274 17672 77276
rect 17696 77274 17752 77276
rect 17776 77274 17832 77276
rect 17856 77274 17912 77276
rect 17616 77222 17662 77274
rect 17662 77222 17672 77274
rect 17696 77222 17726 77274
rect 17726 77222 17738 77274
rect 17738 77222 17752 77274
rect 17776 77222 17790 77274
rect 17790 77222 17802 77274
rect 17802 77222 17832 77274
rect 17856 77222 17866 77274
rect 17866 77222 17912 77274
rect 17616 77220 17672 77222
rect 17696 77220 17752 77222
rect 17776 77220 17832 77222
rect 17856 77220 17912 77222
rect 18234 77016 18290 77072
rect 16956 76730 17012 76732
rect 17036 76730 17092 76732
rect 17116 76730 17172 76732
rect 17196 76730 17252 76732
rect 16956 76678 17002 76730
rect 17002 76678 17012 76730
rect 17036 76678 17066 76730
rect 17066 76678 17078 76730
rect 17078 76678 17092 76730
rect 17116 76678 17130 76730
rect 17130 76678 17142 76730
rect 17142 76678 17172 76730
rect 17196 76678 17206 76730
rect 17206 76678 17252 76730
rect 16956 76676 17012 76678
rect 17036 76676 17092 76678
rect 17116 76676 17172 76678
rect 17196 76676 17252 76678
rect 14094 35672 14150 35728
rect 14186 29844 14242 29880
rect 14186 29824 14188 29844
rect 14188 29824 14240 29844
rect 14240 29824 14242 29844
rect 11956 8186 12012 8188
rect 12036 8186 12092 8188
rect 12116 8186 12172 8188
rect 12196 8186 12252 8188
rect 11956 8134 12002 8186
rect 12002 8134 12012 8186
rect 12036 8134 12066 8186
rect 12066 8134 12078 8186
rect 12078 8134 12092 8186
rect 12116 8134 12130 8186
rect 12130 8134 12142 8186
rect 12142 8134 12172 8186
rect 12196 8134 12206 8186
rect 12206 8134 12252 8186
rect 11956 8132 12012 8134
rect 12036 8132 12092 8134
rect 12116 8132 12172 8134
rect 12196 8132 12252 8134
rect 11518 8084 11574 8120
rect 11518 8064 11520 8084
rect 11520 8064 11572 8084
rect 11572 8064 11574 8084
rect 12254 7928 12310 7984
rect 12616 7642 12672 7644
rect 12696 7642 12752 7644
rect 12776 7642 12832 7644
rect 12856 7642 12912 7644
rect 12616 7590 12662 7642
rect 12662 7590 12672 7642
rect 12696 7590 12726 7642
rect 12726 7590 12738 7642
rect 12738 7590 12752 7642
rect 12776 7590 12790 7642
rect 12790 7590 12802 7642
rect 12802 7590 12832 7642
rect 12856 7590 12866 7642
rect 12866 7590 12912 7642
rect 12616 7588 12672 7590
rect 12696 7588 12752 7590
rect 12776 7588 12832 7590
rect 12856 7588 12912 7590
rect 11956 7098 12012 7100
rect 12036 7098 12092 7100
rect 12116 7098 12172 7100
rect 12196 7098 12252 7100
rect 11956 7046 12002 7098
rect 12002 7046 12012 7098
rect 12036 7046 12066 7098
rect 12066 7046 12078 7098
rect 12078 7046 12092 7098
rect 12116 7046 12130 7098
rect 12130 7046 12142 7098
rect 12142 7046 12172 7098
rect 12196 7046 12206 7098
rect 12206 7046 12252 7098
rect 11956 7044 12012 7046
rect 12036 7044 12092 7046
rect 12116 7044 12172 7046
rect 12196 7044 12252 7046
rect 12714 6840 12770 6896
rect 13358 6840 13414 6896
rect 12616 6554 12672 6556
rect 12696 6554 12752 6556
rect 12776 6554 12832 6556
rect 12856 6554 12912 6556
rect 12616 6502 12662 6554
rect 12662 6502 12672 6554
rect 12696 6502 12726 6554
rect 12726 6502 12738 6554
rect 12738 6502 12752 6554
rect 12776 6502 12790 6554
rect 12790 6502 12802 6554
rect 12802 6502 12832 6554
rect 12856 6502 12866 6554
rect 12866 6502 12912 6554
rect 12616 6500 12672 6502
rect 12696 6500 12752 6502
rect 12776 6500 12832 6502
rect 12856 6500 12912 6502
rect 11956 6010 12012 6012
rect 12036 6010 12092 6012
rect 12116 6010 12172 6012
rect 12196 6010 12252 6012
rect 11956 5958 12002 6010
rect 12002 5958 12012 6010
rect 12036 5958 12066 6010
rect 12066 5958 12078 6010
rect 12078 5958 12092 6010
rect 12116 5958 12130 6010
rect 12130 5958 12142 6010
rect 12142 5958 12172 6010
rect 12196 5958 12206 6010
rect 12206 5958 12252 6010
rect 11956 5956 12012 5958
rect 12036 5956 12092 5958
rect 12116 5956 12172 5958
rect 12196 5956 12252 5958
rect 12616 5466 12672 5468
rect 12696 5466 12752 5468
rect 12776 5466 12832 5468
rect 12856 5466 12912 5468
rect 12616 5414 12662 5466
rect 12662 5414 12672 5466
rect 12696 5414 12726 5466
rect 12726 5414 12738 5466
rect 12738 5414 12752 5466
rect 12776 5414 12790 5466
rect 12790 5414 12802 5466
rect 12802 5414 12832 5466
rect 12856 5414 12866 5466
rect 12866 5414 12912 5466
rect 12616 5412 12672 5414
rect 12696 5412 12752 5414
rect 12776 5412 12832 5414
rect 12856 5412 12912 5414
rect 15014 68992 15070 69048
rect 14462 63280 14518 63336
rect 14186 8200 14242 8256
rect 13818 7268 13874 7304
rect 13818 7248 13820 7268
rect 13820 7248 13872 7268
rect 13872 7248 13874 7268
rect 11956 4922 12012 4924
rect 12036 4922 12092 4924
rect 12116 4922 12172 4924
rect 12196 4922 12252 4924
rect 11956 4870 12002 4922
rect 12002 4870 12012 4922
rect 12036 4870 12066 4922
rect 12066 4870 12078 4922
rect 12078 4870 12092 4922
rect 12116 4870 12130 4922
rect 12130 4870 12142 4922
rect 12142 4870 12172 4922
rect 12196 4870 12206 4922
rect 12206 4870 12252 4922
rect 11956 4868 12012 4870
rect 12036 4868 12092 4870
rect 12116 4868 12172 4870
rect 12196 4868 12252 4870
rect 16956 75642 17012 75644
rect 17036 75642 17092 75644
rect 17116 75642 17172 75644
rect 17196 75642 17252 75644
rect 16956 75590 17002 75642
rect 17002 75590 17012 75642
rect 17036 75590 17066 75642
rect 17066 75590 17078 75642
rect 17078 75590 17092 75642
rect 17116 75590 17130 75642
rect 17130 75590 17142 75642
rect 17142 75590 17172 75642
rect 17196 75590 17206 75642
rect 17206 75590 17252 75642
rect 16956 75588 17012 75590
rect 17036 75588 17092 75590
rect 17116 75588 17172 75590
rect 17196 75588 17252 75590
rect 17616 76186 17672 76188
rect 17696 76186 17752 76188
rect 17776 76186 17832 76188
rect 17856 76186 17912 76188
rect 17616 76134 17662 76186
rect 17662 76134 17672 76186
rect 17696 76134 17726 76186
rect 17726 76134 17738 76186
rect 17738 76134 17752 76186
rect 17776 76134 17790 76186
rect 17790 76134 17802 76186
rect 17802 76134 17832 76186
rect 17856 76134 17866 76186
rect 17866 76134 17912 76186
rect 17616 76132 17672 76134
rect 17696 76132 17752 76134
rect 17776 76132 17832 76134
rect 17856 76132 17912 76134
rect 18234 75148 18236 75168
rect 18236 75148 18288 75168
rect 18288 75148 18290 75168
rect 18234 75112 18290 75148
rect 17616 75098 17672 75100
rect 17696 75098 17752 75100
rect 17776 75098 17832 75100
rect 17856 75098 17912 75100
rect 17616 75046 17662 75098
rect 17662 75046 17672 75098
rect 17696 75046 17726 75098
rect 17726 75046 17738 75098
rect 17738 75046 17752 75098
rect 17776 75046 17790 75098
rect 17790 75046 17802 75098
rect 17802 75046 17832 75098
rect 17856 75046 17866 75098
rect 17866 75046 17912 75098
rect 17616 75044 17672 75046
rect 17696 75044 17752 75046
rect 17776 75044 17832 75046
rect 17856 75044 17912 75046
rect 16956 74554 17012 74556
rect 17036 74554 17092 74556
rect 17116 74554 17172 74556
rect 17196 74554 17252 74556
rect 16026 48320 16082 48376
rect 15290 11212 15346 11248
rect 15290 11192 15292 11212
rect 15292 11192 15344 11212
rect 15344 11192 15346 11212
rect 16394 60016 16450 60072
rect 16302 49544 16358 49600
rect 16956 74502 17002 74554
rect 17002 74502 17012 74554
rect 17036 74502 17066 74554
rect 17066 74502 17078 74554
rect 17078 74502 17092 74554
rect 17116 74502 17130 74554
rect 17130 74502 17142 74554
rect 17142 74502 17172 74554
rect 17196 74502 17206 74554
rect 17206 74502 17252 74554
rect 16956 74500 17012 74502
rect 17036 74500 17092 74502
rect 17116 74500 17172 74502
rect 17196 74500 17252 74502
rect 17616 74010 17672 74012
rect 17696 74010 17752 74012
rect 17776 74010 17832 74012
rect 17856 74010 17912 74012
rect 17616 73958 17662 74010
rect 17662 73958 17672 74010
rect 17696 73958 17726 74010
rect 17726 73958 17738 74010
rect 17738 73958 17752 74010
rect 17776 73958 17790 74010
rect 17790 73958 17802 74010
rect 17802 73958 17832 74010
rect 17856 73958 17866 74010
rect 17866 73958 17912 74010
rect 17616 73956 17672 73958
rect 17696 73956 17752 73958
rect 17776 73956 17832 73958
rect 17856 73956 17912 73958
rect 16956 73466 17012 73468
rect 17036 73466 17092 73468
rect 17116 73466 17172 73468
rect 17196 73466 17252 73468
rect 16956 73414 17002 73466
rect 17002 73414 17012 73466
rect 17036 73414 17066 73466
rect 17066 73414 17078 73466
rect 17078 73414 17092 73466
rect 17116 73414 17130 73466
rect 17130 73414 17142 73466
rect 17142 73414 17172 73466
rect 17196 73414 17206 73466
rect 17206 73414 17252 73466
rect 16956 73412 17012 73414
rect 17036 73412 17092 73414
rect 17116 73412 17172 73414
rect 17196 73412 17252 73414
rect 16956 72378 17012 72380
rect 17036 72378 17092 72380
rect 17116 72378 17172 72380
rect 17196 72378 17252 72380
rect 16956 72326 17002 72378
rect 17002 72326 17012 72378
rect 17036 72326 17066 72378
rect 17066 72326 17078 72378
rect 17078 72326 17092 72378
rect 17116 72326 17130 72378
rect 17130 72326 17142 72378
rect 17142 72326 17172 72378
rect 17196 72326 17206 72378
rect 17206 72326 17252 72378
rect 16956 72324 17012 72326
rect 17036 72324 17092 72326
rect 17116 72324 17172 72326
rect 17196 72324 17252 72326
rect 16956 71290 17012 71292
rect 17036 71290 17092 71292
rect 17116 71290 17172 71292
rect 17196 71290 17252 71292
rect 16956 71238 17002 71290
rect 17002 71238 17012 71290
rect 17036 71238 17066 71290
rect 17066 71238 17078 71290
rect 17078 71238 17092 71290
rect 17116 71238 17130 71290
rect 17130 71238 17142 71290
rect 17142 71238 17172 71290
rect 17196 71238 17206 71290
rect 17206 71238 17252 71290
rect 16956 71236 17012 71238
rect 17036 71236 17092 71238
rect 17116 71236 17172 71238
rect 17196 71236 17252 71238
rect 16956 70202 17012 70204
rect 17036 70202 17092 70204
rect 17116 70202 17172 70204
rect 17196 70202 17252 70204
rect 16956 70150 17002 70202
rect 17002 70150 17012 70202
rect 17036 70150 17066 70202
rect 17066 70150 17078 70202
rect 17078 70150 17092 70202
rect 17116 70150 17130 70202
rect 17130 70150 17142 70202
rect 17142 70150 17172 70202
rect 17196 70150 17206 70202
rect 17206 70150 17252 70202
rect 16956 70148 17012 70150
rect 17036 70148 17092 70150
rect 17116 70148 17172 70150
rect 17196 70148 17252 70150
rect 16956 69114 17012 69116
rect 17036 69114 17092 69116
rect 17116 69114 17172 69116
rect 17196 69114 17252 69116
rect 16956 69062 17002 69114
rect 17002 69062 17012 69114
rect 17036 69062 17066 69114
rect 17066 69062 17078 69114
rect 17078 69062 17092 69114
rect 17116 69062 17130 69114
rect 17130 69062 17142 69114
rect 17142 69062 17172 69114
rect 17196 69062 17206 69114
rect 17206 69062 17252 69114
rect 16956 69060 17012 69062
rect 17036 69060 17092 69062
rect 17116 69060 17172 69062
rect 17196 69060 17252 69062
rect 16956 68026 17012 68028
rect 17036 68026 17092 68028
rect 17116 68026 17172 68028
rect 17196 68026 17252 68028
rect 16956 67974 17002 68026
rect 17002 67974 17012 68026
rect 17036 67974 17066 68026
rect 17066 67974 17078 68026
rect 17078 67974 17092 68026
rect 17116 67974 17130 68026
rect 17130 67974 17142 68026
rect 17142 67974 17172 68026
rect 17196 67974 17206 68026
rect 17206 67974 17252 68026
rect 16956 67972 17012 67974
rect 17036 67972 17092 67974
rect 17116 67972 17172 67974
rect 17196 67972 17252 67974
rect 16956 66938 17012 66940
rect 17036 66938 17092 66940
rect 17116 66938 17172 66940
rect 17196 66938 17252 66940
rect 16956 66886 17002 66938
rect 17002 66886 17012 66938
rect 17036 66886 17066 66938
rect 17066 66886 17078 66938
rect 17078 66886 17092 66938
rect 17116 66886 17130 66938
rect 17130 66886 17142 66938
rect 17142 66886 17172 66938
rect 17196 66886 17206 66938
rect 17206 66886 17252 66938
rect 16956 66884 17012 66886
rect 17036 66884 17092 66886
rect 17116 66884 17172 66886
rect 17196 66884 17252 66886
rect 16956 65850 17012 65852
rect 17036 65850 17092 65852
rect 17116 65850 17172 65852
rect 17196 65850 17252 65852
rect 16956 65798 17002 65850
rect 17002 65798 17012 65850
rect 17036 65798 17066 65850
rect 17066 65798 17078 65850
rect 17078 65798 17092 65850
rect 17116 65798 17130 65850
rect 17130 65798 17142 65850
rect 17142 65798 17172 65850
rect 17196 65798 17206 65850
rect 17206 65798 17252 65850
rect 16956 65796 17012 65798
rect 17036 65796 17092 65798
rect 17116 65796 17172 65798
rect 17196 65796 17252 65798
rect 18234 73208 18290 73264
rect 17616 72922 17672 72924
rect 17696 72922 17752 72924
rect 17776 72922 17832 72924
rect 17856 72922 17912 72924
rect 17616 72870 17662 72922
rect 17662 72870 17672 72922
rect 17696 72870 17726 72922
rect 17726 72870 17738 72922
rect 17738 72870 17752 72922
rect 17776 72870 17790 72922
rect 17790 72870 17802 72922
rect 17802 72870 17832 72922
rect 17856 72870 17866 72922
rect 17866 72870 17912 72922
rect 17616 72868 17672 72870
rect 17696 72868 17752 72870
rect 17776 72868 17832 72870
rect 17856 72868 17912 72870
rect 17616 71834 17672 71836
rect 17696 71834 17752 71836
rect 17776 71834 17832 71836
rect 17856 71834 17912 71836
rect 17616 71782 17662 71834
rect 17662 71782 17672 71834
rect 17696 71782 17726 71834
rect 17726 71782 17738 71834
rect 17738 71782 17752 71834
rect 17776 71782 17790 71834
rect 17790 71782 17802 71834
rect 17802 71782 17832 71834
rect 17856 71782 17866 71834
rect 17866 71782 17912 71834
rect 17616 71780 17672 71782
rect 17696 71780 17752 71782
rect 17776 71780 17832 71782
rect 17856 71780 17912 71782
rect 18234 71340 18236 71360
rect 18236 71340 18288 71360
rect 18288 71340 18290 71360
rect 18234 71304 18290 71340
rect 17616 70746 17672 70748
rect 17696 70746 17752 70748
rect 17776 70746 17832 70748
rect 17856 70746 17912 70748
rect 17616 70694 17662 70746
rect 17662 70694 17672 70746
rect 17696 70694 17726 70746
rect 17726 70694 17738 70746
rect 17738 70694 17752 70746
rect 17776 70694 17790 70746
rect 17790 70694 17802 70746
rect 17802 70694 17832 70746
rect 17856 70694 17866 70746
rect 17866 70694 17912 70746
rect 17616 70692 17672 70694
rect 17696 70692 17752 70694
rect 17776 70692 17832 70694
rect 17856 70692 17912 70694
rect 17616 69658 17672 69660
rect 17696 69658 17752 69660
rect 17776 69658 17832 69660
rect 17856 69658 17912 69660
rect 17616 69606 17662 69658
rect 17662 69606 17672 69658
rect 17696 69606 17726 69658
rect 17726 69606 17738 69658
rect 17738 69606 17752 69658
rect 17776 69606 17790 69658
rect 17790 69606 17802 69658
rect 17802 69606 17832 69658
rect 17856 69606 17866 69658
rect 17866 69606 17912 69658
rect 17616 69604 17672 69606
rect 17696 69604 17752 69606
rect 17776 69604 17832 69606
rect 17856 69604 17912 69606
rect 18234 69400 18290 69456
rect 17616 68570 17672 68572
rect 17696 68570 17752 68572
rect 17776 68570 17832 68572
rect 17856 68570 17912 68572
rect 17616 68518 17662 68570
rect 17662 68518 17672 68570
rect 17696 68518 17726 68570
rect 17726 68518 17738 68570
rect 17738 68518 17752 68570
rect 17776 68518 17790 68570
rect 17790 68518 17802 68570
rect 17802 68518 17832 68570
rect 17856 68518 17866 68570
rect 17866 68518 17912 68570
rect 17616 68516 17672 68518
rect 17696 68516 17752 68518
rect 17776 68516 17832 68518
rect 17856 68516 17912 68518
rect 18234 67496 18290 67552
rect 17616 67482 17672 67484
rect 17696 67482 17752 67484
rect 17776 67482 17832 67484
rect 17856 67482 17912 67484
rect 17616 67430 17662 67482
rect 17662 67430 17672 67482
rect 17696 67430 17726 67482
rect 17726 67430 17738 67482
rect 17738 67430 17752 67482
rect 17776 67430 17790 67482
rect 17790 67430 17802 67482
rect 17802 67430 17832 67482
rect 17856 67430 17866 67482
rect 17866 67430 17912 67482
rect 17616 67428 17672 67430
rect 17696 67428 17752 67430
rect 17776 67428 17832 67430
rect 17856 67428 17912 67430
rect 17616 66394 17672 66396
rect 17696 66394 17752 66396
rect 17776 66394 17832 66396
rect 17856 66394 17912 66396
rect 17616 66342 17662 66394
rect 17662 66342 17672 66394
rect 17696 66342 17726 66394
rect 17726 66342 17738 66394
rect 17738 66342 17752 66394
rect 17776 66342 17790 66394
rect 17790 66342 17802 66394
rect 17802 66342 17832 66394
rect 17856 66342 17866 66394
rect 17866 66342 17912 66394
rect 17616 66340 17672 66342
rect 17696 66340 17752 66342
rect 17776 66340 17832 66342
rect 17856 66340 17912 66342
rect 18234 65628 18236 65648
rect 18236 65628 18288 65648
rect 18288 65628 18290 65648
rect 18234 65592 18290 65628
rect 17616 65306 17672 65308
rect 17696 65306 17752 65308
rect 17776 65306 17832 65308
rect 17856 65306 17912 65308
rect 17616 65254 17662 65306
rect 17662 65254 17672 65306
rect 17696 65254 17726 65306
rect 17726 65254 17738 65306
rect 17738 65254 17752 65306
rect 17776 65254 17790 65306
rect 17790 65254 17802 65306
rect 17802 65254 17832 65306
rect 17856 65254 17866 65306
rect 17866 65254 17912 65306
rect 17616 65252 17672 65254
rect 17696 65252 17752 65254
rect 17776 65252 17832 65254
rect 17856 65252 17912 65254
rect 17498 65048 17554 65104
rect 16302 37304 16358 37360
rect 16956 64762 17012 64764
rect 17036 64762 17092 64764
rect 17116 64762 17172 64764
rect 17196 64762 17252 64764
rect 16956 64710 17002 64762
rect 17002 64710 17012 64762
rect 17036 64710 17066 64762
rect 17066 64710 17078 64762
rect 17078 64710 17092 64762
rect 17116 64710 17130 64762
rect 17130 64710 17142 64762
rect 17142 64710 17172 64762
rect 17196 64710 17206 64762
rect 17206 64710 17252 64762
rect 16956 64708 17012 64710
rect 17036 64708 17092 64710
rect 17116 64708 17172 64710
rect 17196 64708 17252 64710
rect 16956 63674 17012 63676
rect 17036 63674 17092 63676
rect 17116 63674 17172 63676
rect 17196 63674 17252 63676
rect 16956 63622 17002 63674
rect 17002 63622 17012 63674
rect 17036 63622 17066 63674
rect 17066 63622 17078 63674
rect 17078 63622 17092 63674
rect 17116 63622 17130 63674
rect 17130 63622 17142 63674
rect 17142 63622 17172 63674
rect 17196 63622 17206 63674
rect 17206 63622 17252 63674
rect 16956 63620 17012 63622
rect 17036 63620 17092 63622
rect 17116 63620 17172 63622
rect 17196 63620 17252 63622
rect 16956 62586 17012 62588
rect 17036 62586 17092 62588
rect 17116 62586 17172 62588
rect 17196 62586 17252 62588
rect 16956 62534 17002 62586
rect 17002 62534 17012 62586
rect 17036 62534 17066 62586
rect 17066 62534 17078 62586
rect 17078 62534 17092 62586
rect 17116 62534 17130 62586
rect 17130 62534 17142 62586
rect 17142 62534 17172 62586
rect 17196 62534 17206 62586
rect 17206 62534 17252 62586
rect 16956 62532 17012 62534
rect 17036 62532 17092 62534
rect 17116 62532 17172 62534
rect 17196 62532 17252 62534
rect 16956 61498 17012 61500
rect 17036 61498 17092 61500
rect 17116 61498 17172 61500
rect 17196 61498 17252 61500
rect 16956 61446 17002 61498
rect 17002 61446 17012 61498
rect 17036 61446 17066 61498
rect 17066 61446 17078 61498
rect 17078 61446 17092 61498
rect 17116 61446 17130 61498
rect 17130 61446 17142 61498
rect 17142 61446 17172 61498
rect 17196 61446 17206 61498
rect 17206 61446 17252 61498
rect 16956 61444 17012 61446
rect 17036 61444 17092 61446
rect 17116 61444 17172 61446
rect 17196 61444 17252 61446
rect 16956 60410 17012 60412
rect 17036 60410 17092 60412
rect 17116 60410 17172 60412
rect 17196 60410 17252 60412
rect 16956 60358 17002 60410
rect 17002 60358 17012 60410
rect 17036 60358 17066 60410
rect 17066 60358 17078 60410
rect 17078 60358 17092 60410
rect 17116 60358 17130 60410
rect 17130 60358 17142 60410
rect 17142 60358 17172 60410
rect 17196 60358 17206 60410
rect 17206 60358 17252 60410
rect 16956 60356 17012 60358
rect 17036 60356 17092 60358
rect 17116 60356 17172 60358
rect 17196 60356 17252 60358
rect 16956 59322 17012 59324
rect 17036 59322 17092 59324
rect 17116 59322 17172 59324
rect 17196 59322 17252 59324
rect 16956 59270 17002 59322
rect 17002 59270 17012 59322
rect 17036 59270 17066 59322
rect 17066 59270 17078 59322
rect 17078 59270 17092 59322
rect 17116 59270 17130 59322
rect 17130 59270 17142 59322
rect 17142 59270 17172 59322
rect 17196 59270 17206 59322
rect 17206 59270 17252 59322
rect 16956 59268 17012 59270
rect 17036 59268 17092 59270
rect 17116 59268 17172 59270
rect 17196 59268 17252 59270
rect 16956 58234 17012 58236
rect 17036 58234 17092 58236
rect 17116 58234 17172 58236
rect 17196 58234 17252 58236
rect 16956 58182 17002 58234
rect 17002 58182 17012 58234
rect 17036 58182 17066 58234
rect 17066 58182 17078 58234
rect 17078 58182 17092 58234
rect 17116 58182 17130 58234
rect 17130 58182 17142 58234
rect 17142 58182 17172 58234
rect 17196 58182 17206 58234
rect 17206 58182 17252 58234
rect 16956 58180 17012 58182
rect 17036 58180 17092 58182
rect 17116 58180 17172 58182
rect 17196 58180 17252 58182
rect 16956 57146 17012 57148
rect 17036 57146 17092 57148
rect 17116 57146 17172 57148
rect 17196 57146 17252 57148
rect 16956 57094 17002 57146
rect 17002 57094 17012 57146
rect 17036 57094 17066 57146
rect 17066 57094 17078 57146
rect 17078 57094 17092 57146
rect 17116 57094 17130 57146
rect 17130 57094 17142 57146
rect 17142 57094 17172 57146
rect 17196 57094 17206 57146
rect 17206 57094 17252 57146
rect 16956 57092 17012 57094
rect 17036 57092 17092 57094
rect 17116 57092 17172 57094
rect 17196 57092 17252 57094
rect 16956 56058 17012 56060
rect 17036 56058 17092 56060
rect 17116 56058 17172 56060
rect 17196 56058 17252 56060
rect 16956 56006 17002 56058
rect 17002 56006 17012 56058
rect 17036 56006 17066 56058
rect 17066 56006 17078 56058
rect 17078 56006 17092 56058
rect 17116 56006 17130 56058
rect 17130 56006 17142 56058
rect 17142 56006 17172 56058
rect 17196 56006 17206 56058
rect 17206 56006 17252 56058
rect 16956 56004 17012 56006
rect 17036 56004 17092 56006
rect 17116 56004 17172 56006
rect 17196 56004 17252 56006
rect 16956 54970 17012 54972
rect 17036 54970 17092 54972
rect 17116 54970 17172 54972
rect 17196 54970 17252 54972
rect 16956 54918 17002 54970
rect 17002 54918 17012 54970
rect 17036 54918 17066 54970
rect 17066 54918 17078 54970
rect 17078 54918 17092 54970
rect 17116 54918 17130 54970
rect 17130 54918 17142 54970
rect 17142 54918 17172 54970
rect 17196 54918 17206 54970
rect 17206 54918 17252 54970
rect 16956 54916 17012 54918
rect 17036 54916 17092 54918
rect 17116 54916 17172 54918
rect 17196 54916 17252 54918
rect 16956 53882 17012 53884
rect 17036 53882 17092 53884
rect 17116 53882 17172 53884
rect 17196 53882 17252 53884
rect 16956 53830 17002 53882
rect 17002 53830 17012 53882
rect 17036 53830 17066 53882
rect 17066 53830 17078 53882
rect 17078 53830 17092 53882
rect 17116 53830 17130 53882
rect 17130 53830 17142 53882
rect 17142 53830 17172 53882
rect 17196 53830 17206 53882
rect 17206 53830 17252 53882
rect 16956 53828 17012 53830
rect 17036 53828 17092 53830
rect 17116 53828 17172 53830
rect 17196 53828 17252 53830
rect 16956 52794 17012 52796
rect 17036 52794 17092 52796
rect 17116 52794 17172 52796
rect 17196 52794 17252 52796
rect 16956 52742 17002 52794
rect 17002 52742 17012 52794
rect 17036 52742 17066 52794
rect 17066 52742 17078 52794
rect 17078 52742 17092 52794
rect 17116 52742 17130 52794
rect 17130 52742 17142 52794
rect 17142 52742 17172 52794
rect 17196 52742 17206 52794
rect 17206 52742 17252 52794
rect 16956 52740 17012 52742
rect 17036 52740 17092 52742
rect 17116 52740 17172 52742
rect 17196 52740 17252 52742
rect 16956 51706 17012 51708
rect 17036 51706 17092 51708
rect 17116 51706 17172 51708
rect 17196 51706 17252 51708
rect 16956 51654 17002 51706
rect 17002 51654 17012 51706
rect 17036 51654 17066 51706
rect 17066 51654 17078 51706
rect 17078 51654 17092 51706
rect 17116 51654 17130 51706
rect 17130 51654 17142 51706
rect 17142 51654 17172 51706
rect 17196 51654 17206 51706
rect 17206 51654 17252 51706
rect 16956 51652 17012 51654
rect 17036 51652 17092 51654
rect 17116 51652 17172 51654
rect 17196 51652 17252 51654
rect 16956 50618 17012 50620
rect 17036 50618 17092 50620
rect 17116 50618 17172 50620
rect 17196 50618 17252 50620
rect 16956 50566 17002 50618
rect 17002 50566 17012 50618
rect 17036 50566 17066 50618
rect 17066 50566 17078 50618
rect 17078 50566 17092 50618
rect 17116 50566 17130 50618
rect 17130 50566 17142 50618
rect 17142 50566 17172 50618
rect 17196 50566 17206 50618
rect 17206 50566 17252 50618
rect 16956 50564 17012 50566
rect 17036 50564 17092 50566
rect 17116 50564 17172 50566
rect 17196 50564 17252 50566
rect 16762 48592 16818 48648
rect 16956 49530 17012 49532
rect 17036 49530 17092 49532
rect 17116 49530 17172 49532
rect 17196 49530 17252 49532
rect 16956 49478 17002 49530
rect 17002 49478 17012 49530
rect 17036 49478 17066 49530
rect 17066 49478 17078 49530
rect 17078 49478 17092 49530
rect 17116 49478 17130 49530
rect 17130 49478 17142 49530
rect 17142 49478 17172 49530
rect 17196 49478 17206 49530
rect 17206 49478 17252 49530
rect 16956 49476 17012 49478
rect 17036 49476 17092 49478
rect 17116 49476 17172 49478
rect 17196 49476 17252 49478
rect 16394 24692 16396 24712
rect 16396 24692 16448 24712
rect 16448 24692 16450 24712
rect 16394 24656 16450 24692
rect 16956 48442 17012 48444
rect 17036 48442 17092 48444
rect 17116 48442 17172 48444
rect 17196 48442 17252 48444
rect 16956 48390 17002 48442
rect 17002 48390 17012 48442
rect 17036 48390 17066 48442
rect 17066 48390 17078 48442
rect 17078 48390 17092 48442
rect 17116 48390 17130 48442
rect 17130 48390 17142 48442
rect 17142 48390 17172 48442
rect 17196 48390 17206 48442
rect 17206 48390 17252 48442
rect 16956 48388 17012 48390
rect 17036 48388 17092 48390
rect 17116 48388 17172 48390
rect 17196 48388 17252 48390
rect 16762 48184 16818 48240
rect 16956 47354 17012 47356
rect 17036 47354 17092 47356
rect 17116 47354 17172 47356
rect 17196 47354 17252 47356
rect 16956 47302 17002 47354
rect 17002 47302 17012 47354
rect 17036 47302 17066 47354
rect 17066 47302 17078 47354
rect 17078 47302 17092 47354
rect 17116 47302 17130 47354
rect 17130 47302 17142 47354
rect 17142 47302 17172 47354
rect 17196 47302 17206 47354
rect 17206 47302 17252 47354
rect 16956 47300 17012 47302
rect 17036 47300 17092 47302
rect 17116 47300 17172 47302
rect 17196 47300 17252 47302
rect 16762 34176 16818 34232
rect 16956 46266 17012 46268
rect 17036 46266 17092 46268
rect 17116 46266 17172 46268
rect 17196 46266 17252 46268
rect 16956 46214 17002 46266
rect 17002 46214 17012 46266
rect 17036 46214 17066 46266
rect 17066 46214 17078 46266
rect 17078 46214 17092 46266
rect 17116 46214 17130 46266
rect 17130 46214 17142 46266
rect 17142 46214 17172 46266
rect 17196 46214 17206 46266
rect 17206 46214 17252 46266
rect 16956 46212 17012 46214
rect 17036 46212 17092 46214
rect 17116 46212 17172 46214
rect 17196 46212 17252 46214
rect 16956 45178 17012 45180
rect 17036 45178 17092 45180
rect 17116 45178 17172 45180
rect 17196 45178 17252 45180
rect 16956 45126 17002 45178
rect 17002 45126 17012 45178
rect 17036 45126 17066 45178
rect 17066 45126 17078 45178
rect 17078 45126 17092 45178
rect 17116 45126 17130 45178
rect 17130 45126 17142 45178
rect 17142 45126 17172 45178
rect 17196 45126 17206 45178
rect 17206 45126 17252 45178
rect 16956 45124 17012 45126
rect 17036 45124 17092 45126
rect 17116 45124 17172 45126
rect 17196 45124 17252 45126
rect 16956 44090 17012 44092
rect 17036 44090 17092 44092
rect 17116 44090 17172 44092
rect 17196 44090 17252 44092
rect 16956 44038 17002 44090
rect 17002 44038 17012 44090
rect 17036 44038 17066 44090
rect 17066 44038 17078 44090
rect 17078 44038 17092 44090
rect 17116 44038 17130 44090
rect 17130 44038 17142 44090
rect 17142 44038 17172 44090
rect 17196 44038 17206 44090
rect 17206 44038 17252 44090
rect 16956 44036 17012 44038
rect 17036 44036 17092 44038
rect 17116 44036 17172 44038
rect 17196 44036 17252 44038
rect 16956 43002 17012 43004
rect 17036 43002 17092 43004
rect 17116 43002 17172 43004
rect 17196 43002 17252 43004
rect 16956 42950 17002 43002
rect 17002 42950 17012 43002
rect 17036 42950 17066 43002
rect 17066 42950 17078 43002
rect 17078 42950 17092 43002
rect 17116 42950 17130 43002
rect 17130 42950 17142 43002
rect 17142 42950 17172 43002
rect 17196 42950 17206 43002
rect 17206 42950 17252 43002
rect 16956 42948 17012 42950
rect 17036 42948 17092 42950
rect 17116 42948 17172 42950
rect 17196 42948 17252 42950
rect 17616 64218 17672 64220
rect 17696 64218 17752 64220
rect 17776 64218 17832 64220
rect 17856 64218 17912 64220
rect 17616 64166 17662 64218
rect 17662 64166 17672 64218
rect 17696 64166 17726 64218
rect 17726 64166 17738 64218
rect 17738 64166 17752 64218
rect 17776 64166 17790 64218
rect 17790 64166 17802 64218
rect 17802 64166 17832 64218
rect 17856 64166 17866 64218
rect 17866 64166 17912 64218
rect 17616 64164 17672 64166
rect 17696 64164 17752 64166
rect 17776 64164 17832 64166
rect 17856 64164 17912 64166
rect 18234 63724 18236 63744
rect 18236 63724 18288 63744
rect 18288 63724 18290 63744
rect 18234 63688 18290 63724
rect 17616 63130 17672 63132
rect 17696 63130 17752 63132
rect 17776 63130 17832 63132
rect 17856 63130 17912 63132
rect 17616 63078 17662 63130
rect 17662 63078 17672 63130
rect 17696 63078 17726 63130
rect 17726 63078 17738 63130
rect 17738 63078 17752 63130
rect 17776 63078 17790 63130
rect 17790 63078 17802 63130
rect 17802 63078 17832 63130
rect 17856 63078 17866 63130
rect 17866 63078 17912 63130
rect 17616 63076 17672 63078
rect 17696 63076 17752 63078
rect 17776 63076 17832 63078
rect 17856 63076 17912 63078
rect 17616 62042 17672 62044
rect 17696 62042 17752 62044
rect 17776 62042 17832 62044
rect 17856 62042 17912 62044
rect 17616 61990 17662 62042
rect 17662 61990 17672 62042
rect 17696 61990 17726 62042
rect 17726 61990 17738 62042
rect 17738 61990 17752 62042
rect 17776 61990 17790 62042
rect 17790 61990 17802 62042
rect 17802 61990 17832 62042
rect 17856 61990 17866 62042
rect 17866 61990 17912 62042
rect 17616 61988 17672 61990
rect 17696 61988 17752 61990
rect 17776 61988 17832 61990
rect 17856 61988 17912 61990
rect 18234 61784 18290 61840
rect 17616 60954 17672 60956
rect 17696 60954 17752 60956
rect 17776 60954 17832 60956
rect 17856 60954 17912 60956
rect 17616 60902 17662 60954
rect 17662 60902 17672 60954
rect 17696 60902 17726 60954
rect 17726 60902 17738 60954
rect 17738 60902 17752 60954
rect 17776 60902 17790 60954
rect 17790 60902 17802 60954
rect 17802 60902 17832 60954
rect 17856 60902 17866 60954
rect 17866 60902 17912 60954
rect 17616 60900 17672 60902
rect 17696 60900 17752 60902
rect 17776 60900 17832 60902
rect 17856 60900 17912 60902
rect 17616 59866 17672 59868
rect 17696 59866 17752 59868
rect 17776 59866 17832 59868
rect 17856 59866 17912 59868
rect 17616 59814 17662 59866
rect 17662 59814 17672 59866
rect 17696 59814 17726 59866
rect 17726 59814 17738 59866
rect 17738 59814 17752 59866
rect 17776 59814 17790 59866
rect 17790 59814 17802 59866
rect 17802 59814 17832 59866
rect 17856 59814 17866 59866
rect 17866 59814 17912 59866
rect 17616 59812 17672 59814
rect 17696 59812 17752 59814
rect 17776 59812 17832 59814
rect 17856 59812 17912 59814
rect 17616 58778 17672 58780
rect 17696 58778 17752 58780
rect 17776 58778 17832 58780
rect 17856 58778 17912 58780
rect 17616 58726 17662 58778
rect 17662 58726 17672 58778
rect 17696 58726 17726 58778
rect 17726 58726 17738 58778
rect 17738 58726 17752 58778
rect 17776 58726 17790 58778
rect 17790 58726 17802 58778
rect 17802 58726 17832 58778
rect 17856 58726 17866 58778
rect 17866 58726 17912 58778
rect 17616 58724 17672 58726
rect 17696 58724 17752 58726
rect 17776 58724 17832 58726
rect 17856 58724 17912 58726
rect 17616 57690 17672 57692
rect 17696 57690 17752 57692
rect 17776 57690 17832 57692
rect 17856 57690 17912 57692
rect 17616 57638 17662 57690
rect 17662 57638 17672 57690
rect 17696 57638 17726 57690
rect 17726 57638 17738 57690
rect 17738 57638 17752 57690
rect 17776 57638 17790 57690
rect 17790 57638 17802 57690
rect 17802 57638 17832 57690
rect 17856 57638 17866 57690
rect 17866 57638 17912 57690
rect 17616 57636 17672 57638
rect 17696 57636 17752 57638
rect 17776 57636 17832 57638
rect 17856 57636 17912 57638
rect 18234 59916 18236 59936
rect 18236 59916 18288 59936
rect 18288 59916 18290 59936
rect 18234 59880 18290 59916
rect 18234 57976 18290 58032
rect 17616 56602 17672 56604
rect 17696 56602 17752 56604
rect 17776 56602 17832 56604
rect 17856 56602 17912 56604
rect 17616 56550 17662 56602
rect 17662 56550 17672 56602
rect 17696 56550 17726 56602
rect 17726 56550 17738 56602
rect 17738 56550 17752 56602
rect 17776 56550 17790 56602
rect 17790 56550 17802 56602
rect 17802 56550 17832 56602
rect 17856 56550 17866 56602
rect 17866 56550 17912 56602
rect 17616 56548 17672 56550
rect 17696 56548 17752 56550
rect 17776 56548 17832 56550
rect 17856 56548 17912 56550
rect 17616 55514 17672 55516
rect 17696 55514 17752 55516
rect 17776 55514 17832 55516
rect 17856 55514 17912 55516
rect 17616 55462 17662 55514
rect 17662 55462 17672 55514
rect 17696 55462 17726 55514
rect 17726 55462 17738 55514
rect 17738 55462 17752 55514
rect 17776 55462 17790 55514
rect 17790 55462 17802 55514
rect 17802 55462 17832 55514
rect 17856 55462 17866 55514
rect 17866 55462 17912 55514
rect 17616 55460 17672 55462
rect 17696 55460 17752 55462
rect 17776 55460 17832 55462
rect 17856 55460 17912 55462
rect 18234 56108 18236 56128
rect 18236 56108 18288 56128
rect 18288 56108 18290 56128
rect 18234 56072 18290 56108
rect 17616 54426 17672 54428
rect 17696 54426 17752 54428
rect 17776 54426 17832 54428
rect 17856 54426 17912 54428
rect 17616 54374 17662 54426
rect 17662 54374 17672 54426
rect 17696 54374 17726 54426
rect 17726 54374 17738 54426
rect 17738 54374 17752 54426
rect 17776 54374 17790 54426
rect 17790 54374 17802 54426
rect 17802 54374 17832 54426
rect 17856 54374 17866 54426
rect 17866 54374 17912 54426
rect 17616 54372 17672 54374
rect 17696 54372 17752 54374
rect 17776 54372 17832 54374
rect 17856 54372 17912 54374
rect 17616 53338 17672 53340
rect 17696 53338 17752 53340
rect 17776 53338 17832 53340
rect 17856 53338 17912 53340
rect 17616 53286 17662 53338
rect 17662 53286 17672 53338
rect 17696 53286 17726 53338
rect 17726 53286 17738 53338
rect 17738 53286 17752 53338
rect 17776 53286 17790 53338
rect 17790 53286 17802 53338
rect 17802 53286 17832 53338
rect 17856 53286 17866 53338
rect 17866 53286 17912 53338
rect 17616 53284 17672 53286
rect 17696 53284 17752 53286
rect 17776 53284 17832 53286
rect 17856 53284 17912 53286
rect 17616 52250 17672 52252
rect 17696 52250 17752 52252
rect 17776 52250 17832 52252
rect 17856 52250 17912 52252
rect 17616 52198 17662 52250
rect 17662 52198 17672 52250
rect 17696 52198 17726 52250
rect 17726 52198 17738 52250
rect 17738 52198 17752 52250
rect 17776 52198 17790 52250
rect 17790 52198 17802 52250
rect 17802 52198 17832 52250
rect 17856 52198 17866 52250
rect 17866 52198 17912 52250
rect 17616 52196 17672 52198
rect 17696 52196 17752 52198
rect 17776 52196 17832 52198
rect 17856 52196 17912 52198
rect 17616 51162 17672 51164
rect 17696 51162 17752 51164
rect 17776 51162 17832 51164
rect 17856 51162 17912 51164
rect 17616 51110 17662 51162
rect 17662 51110 17672 51162
rect 17696 51110 17726 51162
rect 17726 51110 17738 51162
rect 17738 51110 17752 51162
rect 17776 51110 17790 51162
rect 17790 51110 17802 51162
rect 17802 51110 17832 51162
rect 17856 51110 17866 51162
rect 17866 51110 17912 51162
rect 17616 51108 17672 51110
rect 17696 51108 17752 51110
rect 17776 51108 17832 51110
rect 17856 51108 17912 51110
rect 17616 50074 17672 50076
rect 17696 50074 17752 50076
rect 17776 50074 17832 50076
rect 17856 50074 17912 50076
rect 17616 50022 17662 50074
rect 17662 50022 17672 50074
rect 17696 50022 17726 50074
rect 17726 50022 17738 50074
rect 17738 50022 17752 50074
rect 17776 50022 17790 50074
rect 17790 50022 17802 50074
rect 17802 50022 17832 50074
rect 17856 50022 17866 50074
rect 17866 50022 17912 50074
rect 17616 50020 17672 50022
rect 17696 50020 17752 50022
rect 17776 50020 17832 50022
rect 17856 50020 17912 50022
rect 17616 48986 17672 48988
rect 17696 48986 17752 48988
rect 17776 48986 17832 48988
rect 17856 48986 17912 48988
rect 17616 48934 17662 48986
rect 17662 48934 17672 48986
rect 17696 48934 17726 48986
rect 17726 48934 17738 48986
rect 17738 48934 17752 48986
rect 17776 48934 17790 48986
rect 17790 48934 17802 48986
rect 17802 48934 17832 48986
rect 17856 48934 17866 48986
rect 17866 48934 17912 48986
rect 17616 48932 17672 48934
rect 17696 48932 17752 48934
rect 17776 48932 17832 48934
rect 17856 48932 17912 48934
rect 17616 47898 17672 47900
rect 17696 47898 17752 47900
rect 17776 47898 17832 47900
rect 17856 47898 17912 47900
rect 17616 47846 17662 47898
rect 17662 47846 17672 47898
rect 17696 47846 17726 47898
rect 17726 47846 17738 47898
rect 17738 47846 17752 47898
rect 17776 47846 17790 47898
rect 17790 47846 17802 47898
rect 17802 47846 17832 47898
rect 17856 47846 17866 47898
rect 17866 47846 17912 47898
rect 17616 47844 17672 47846
rect 17696 47844 17752 47846
rect 17776 47844 17832 47846
rect 17856 47844 17912 47846
rect 17616 46810 17672 46812
rect 17696 46810 17752 46812
rect 17776 46810 17832 46812
rect 17856 46810 17912 46812
rect 17616 46758 17662 46810
rect 17662 46758 17672 46810
rect 17696 46758 17726 46810
rect 17726 46758 17738 46810
rect 17738 46758 17752 46810
rect 17776 46758 17790 46810
rect 17790 46758 17802 46810
rect 17802 46758 17832 46810
rect 17856 46758 17866 46810
rect 17866 46758 17912 46810
rect 17616 46756 17672 46758
rect 17696 46756 17752 46758
rect 17776 46756 17832 46758
rect 17856 46756 17912 46758
rect 17616 45722 17672 45724
rect 17696 45722 17752 45724
rect 17776 45722 17832 45724
rect 17856 45722 17912 45724
rect 17616 45670 17662 45722
rect 17662 45670 17672 45722
rect 17696 45670 17726 45722
rect 17726 45670 17738 45722
rect 17738 45670 17752 45722
rect 17776 45670 17790 45722
rect 17790 45670 17802 45722
rect 17802 45670 17832 45722
rect 17856 45670 17866 45722
rect 17866 45670 17912 45722
rect 17616 45668 17672 45670
rect 17696 45668 17752 45670
rect 17776 45668 17832 45670
rect 17856 45668 17912 45670
rect 17616 44634 17672 44636
rect 17696 44634 17752 44636
rect 17776 44634 17832 44636
rect 17856 44634 17912 44636
rect 17616 44582 17662 44634
rect 17662 44582 17672 44634
rect 17696 44582 17726 44634
rect 17726 44582 17738 44634
rect 17738 44582 17752 44634
rect 17776 44582 17790 44634
rect 17790 44582 17802 44634
rect 17802 44582 17832 44634
rect 17856 44582 17866 44634
rect 17866 44582 17912 44634
rect 17616 44580 17672 44582
rect 17696 44580 17752 44582
rect 17776 44580 17832 44582
rect 17856 44580 17912 44582
rect 17616 43546 17672 43548
rect 17696 43546 17752 43548
rect 17776 43546 17832 43548
rect 17856 43546 17912 43548
rect 17616 43494 17662 43546
rect 17662 43494 17672 43546
rect 17696 43494 17726 43546
rect 17726 43494 17738 43546
rect 17738 43494 17752 43546
rect 17776 43494 17790 43546
rect 17790 43494 17802 43546
rect 17802 43494 17832 43546
rect 17856 43494 17866 43546
rect 17866 43494 17912 43546
rect 17616 43492 17672 43494
rect 17696 43492 17752 43494
rect 17776 43492 17832 43494
rect 17856 43492 17912 43494
rect 16956 41914 17012 41916
rect 17036 41914 17092 41916
rect 17116 41914 17172 41916
rect 17196 41914 17252 41916
rect 16956 41862 17002 41914
rect 17002 41862 17012 41914
rect 17036 41862 17066 41914
rect 17066 41862 17078 41914
rect 17078 41862 17092 41914
rect 17116 41862 17130 41914
rect 17130 41862 17142 41914
rect 17142 41862 17172 41914
rect 17196 41862 17206 41914
rect 17206 41862 17252 41914
rect 16956 41860 17012 41862
rect 17036 41860 17092 41862
rect 17116 41860 17172 41862
rect 17196 41860 17252 41862
rect 16956 40826 17012 40828
rect 17036 40826 17092 40828
rect 17116 40826 17172 40828
rect 17196 40826 17252 40828
rect 16956 40774 17002 40826
rect 17002 40774 17012 40826
rect 17036 40774 17066 40826
rect 17066 40774 17078 40826
rect 17078 40774 17092 40826
rect 17116 40774 17130 40826
rect 17130 40774 17142 40826
rect 17142 40774 17172 40826
rect 17196 40774 17206 40826
rect 17206 40774 17252 40826
rect 16956 40772 17012 40774
rect 17036 40772 17092 40774
rect 17116 40772 17172 40774
rect 17196 40772 17252 40774
rect 16946 40568 17002 40624
rect 16956 39738 17012 39740
rect 17036 39738 17092 39740
rect 17116 39738 17172 39740
rect 17196 39738 17252 39740
rect 16956 39686 17002 39738
rect 17002 39686 17012 39738
rect 17036 39686 17066 39738
rect 17066 39686 17078 39738
rect 17078 39686 17092 39738
rect 17116 39686 17130 39738
rect 17130 39686 17142 39738
rect 17142 39686 17172 39738
rect 17196 39686 17206 39738
rect 17206 39686 17252 39738
rect 16956 39684 17012 39686
rect 17036 39684 17092 39686
rect 17116 39684 17172 39686
rect 17196 39684 17252 39686
rect 16956 38650 17012 38652
rect 17036 38650 17092 38652
rect 17116 38650 17172 38652
rect 17196 38650 17252 38652
rect 16956 38598 17002 38650
rect 17002 38598 17012 38650
rect 17036 38598 17066 38650
rect 17066 38598 17078 38650
rect 17078 38598 17092 38650
rect 17116 38598 17130 38650
rect 17130 38598 17142 38650
rect 17142 38598 17172 38650
rect 17196 38598 17206 38650
rect 17206 38598 17252 38650
rect 16956 38596 17012 38598
rect 17036 38596 17092 38598
rect 17116 38596 17172 38598
rect 17196 38596 17252 38598
rect 16956 37562 17012 37564
rect 17036 37562 17092 37564
rect 17116 37562 17172 37564
rect 17196 37562 17252 37564
rect 16956 37510 17002 37562
rect 17002 37510 17012 37562
rect 17036 37510 17066 37562
rect 17066 37510 17078 37562
rect 17078 37510 17092 37562
rect 17116 37510 17130 37562
rect 17130 37510 17142 37562
rect 17142 37510 17172 37562
rect 17196 37510 17206 37562
rect 17206 37510 17252 37562
rect 16956 37508 17012 37510
rect 17036 37508 17092 37510
rect 17116 37508 17172 37510
rect 17196 37508 17252 37510
rect 16956 36474 17012 36476
rect 17036 36474 17092 36476
rect 17116 36474 17172 36476
rect 17196 36474 17252 36476
rect 16956 36422 17002 36474
rect 17002 36422 17012 36474
rect 17036 36422 17066 36474
rect 17066 36422 17078 36474
rect 17078 36422 17092 36474
rect 17116 36422 17130 36474
rect 17130 36422 17142 36474
rect 17142 36422 17172 36474
rect 17196 36422 17206 36474
rect 17206 36422 17252 36474
rect 16956 36420 17012 36422
rect 17036 36420 17092 36422
rect 17116 36420 17172 36422
rect 17196 36420 17252 36422
rect 16956 35386 17012 35388
rect 17036 35386 17092 35388
rect 17116 35386 17172 35388
rect 17196 35386 17252 35388
rect 16956 35334 17002 35386
rect 17002 35334 17012 35386
rect 17036 35334 17066 35386
rect 17066 35334 17078 35386
rect 17078 35334 17092 35386
rect 17116 35334 17130 35386
rect 17130 35334 17142 35386
rect 17142 35334 17172 35386
rect 17196 35334 17206 35386
rect 17206 35334 17252 35386
rect 16956 35332 17012 35334
rect 17036 35332 17092 35334
rect 17116 35332 17172 35334
rect 17196 35332 17252 35334
rect 16956 34298 17012 34300
rect 17036 34298 17092 34300
rect 17116 34298 17172 34300
rect 17196 34298 17252 34300
rect 16956 34246 17002 34298
rect 17002 34246 17012 34298
rect 17036 34246 17066 34298
rect 17066 34246 17078 34298
rect 17078 34246 17092 34298
rect 17116 34246 17130 34298
rect 17130 34246 17142 34298
rect 17142 34246 17172 34298
rect 17196 34246 17206 34298
rect 17206 34246 17252 34298
rect 16956 34244 17012 34246
rect 17036 34244 17092 34246
rect 17116 34244 17172 34246
rect 17196 34244 17252 34246
rect 16956 33210 17012 33212
rect 17036 33210 17092 33212
rect 17116 33210 17172 33212
rect 17196 33210 17252 33212
rect 16956 33158 17002 33210
rect 17002 33158 17012 33210
rect 17036 33158 17066 33210
rect 17066 33158 17078 33210
rect 17078 33158 17092 33210
rect 17116 33158 17130 33210
rect 17130 33158 17142 33210
rect 17142 33158 17172 33210
rect 17196 33158 17206 33210
rect 17206 33158 17252 33210
rect 16956 33156 17012 33158
rect 17036 33156 17092 33158
rect 17116 33156 17172 33158
rect 17196 33156 17252 33158
rect 16762 31728 16818 31784
rect 16946 32272 17002 32328
rect 16956 32122 17012 32124
rect 17036 32122 17092 32124
rect 17116 32122 17172 32124
rect 17196 32122 17252 32124
rect 16956 32070 17002 32122
rect 17002 32070 17012 32122
rect 17036 32070 17066 32122
rect 17066 32070 17078 32122
rect 17078 32070 17092 32122
rect 17116 32070 17130 32122
rect 17130 32070 17142 32122
rect 17142 32070 17172 32122
rect 17196 32070 17206 32122
rect 17206 32070 17252 32122
rect 16956 32068 17012 32070
rect 17036 32068 17092 32070
rect 17116 32068 17172 32070
rect 17196 32068 17252 32070
rect 16956 31034 17012 31036
rect 17036 31034 17092 31036
rect 17116 31034 17172 31036
rect 17196 31034 17252 31036
rect 16956 30982 17002 31034
rect 17002 30982 17012 31034
rect 17036 30982 17066 31034
rect 17066 30982 17078 31034
rect 17078 30982 17092 31034
rect 17116 30982 17130 31034
rect 17130 30982 17142 31034
rect 17142 30982 17172 31034
rect 17196 30982 17206 31034
rect 17206 30982 17252 31034
rect 16956 30980 17012 30982
rect 17036 30980 17092 30982
rect 17116 30980 17172 30982
rect 17196 30980 17252 30982
rect 16956 29946 17012 29948
rect 17036 29946 17092 29948
rect 17116 29946 17172 29948
rect 17196 29946 17252 29948
rect 16956 29894 17002 29946
rect 17002 29894 17012 29946
rect 17036 29894 17066 29946
rect 17066 29894 17078 29946
rect 17078 29894 17092 29946
rect 17116 29894 17130 29946
rect 17130 29894 17142 29946
rect 17142 29894 17172 29946
rect 17196 29894 17206 29946
rect 17206 29894 17252 29946
rect 16956 29892 17012 29894
rect 17036 29892 17092 29894
rect 17116 29892 17172 29894
rect 17196 29892 17252 29894
rect 16956 28858 17012 28860
rect 17036 28858 17092 28860
rect 17116 28858 17172 28860
rect 17196 28858 17252 28860
rect 16956 28806 17002 28858
rect 17002 28806 17012 28858
rect 17036 28806 17066 28858
rect 17066 28806 17078 28858
rect 17078 28806 17092 28858
rect 17116 28806 17130 28858
rect 17130 28806 17142 28858
rect 17142 28806 17172 28858
rect 17196 28806 17206 28858
rect 17206 28806 17252 28858
rect 16956 28804 17012 28806
rect 17036 28804 17092 28806
rect 17116 28804 17172 28806
rect 17196 28804 17252 28806
rect 16956 27770 17012 27772
rect 17036 27770 17092 27772
rect 17116 27770 17172 27772
rect 17196 27770 17252 27772
rect 16956 27718 17002 27770
rect 17002 27718 17012 27770
rect 17036 27718 17066 27770
rect 17066 27718 17078 27770
rect 17078 27718 17092 27770
rect 17116 27718 17130 27770
rect 17130 27718 17142 27770
rect 17142 27718 17172 27770
rect 17196 27718 17206 27770
rect 17206 27718 17252 27770
rect 16956 27716 17012 27718
rect 17036 27716 17092 27718
rect 17116 27716 17172 27718
rect 17196 27716 17252 27718
rect 16956 26682 17012 26684
rect 17036 26682 17092 26684
rect 17116 26682 17172 26684
rect 17196 26682 17252 26684
rect 16956 26630 17002 26682
rect 17002 26630 17012 26682
rect 17036 26630 17066 26682
rect 17066 26630 17078 26682
rect 17078 26630 17092 26682
rect 17116 26630 17130 26682
rect 17130 26630 17142 26682
rect 17142 26630 17172 26682
rect 17196 26630 17206 26682
rect 17206 26630 17252 26682
rect 16956 26628 17012 26630
rect 17036 26628 17092 26630
rect 17116 26628 17172 26630
rect 17196 26628 17252 26630
rect 16956 25594 17012 25596
rect 17036 25594 17092 25596
rect 17116 25594 17172 25596
rect 17196 25594 17252 25596
rect 16956 25542 17002 25594
rect 17002 25542 17012 25594
rect 17036 25542 17066 25594
rect 17066 25542 17078 25594
rect 17078 25542 17092 25594
rect 17116 25542 17130 25594
rect 17130 25542 17142 25594
rect 17142 25542 17172 25594
rect 17196 25542 17206 25594
rect 17206 25542 17252 25594
rect 16956 25540 17012 25542
rect 17036 25540 17092 25542
rect 17116 25540 17172 25542
rect 17196 25540 17252 25542
rect 16956 24506 17012 24508
rect 17036 24506 17092 24508
rect 17116 24506 17172 24508
rect 17196 24506 17252 24508
rect 16956 24454 17002 24506
rect 17002 24454 17012 24506
rect 17036 24454 17066 24506
rect 17066 24454 17078 24506
rect 17078 24454 17092 24506
rect 17116 24454 17130 24506
rect 17130 24454 17142 24506
rect 17142 24454 17172 24506
rect 17196 24454 17206 24506
rect 17206 24454 17252 24506
rect 16956 24452 17012 24454
rect 17036 24452 17092 24454
rect 17116 24452 17172 24454
rect 17196 24452 17252 24454
rect 16946 23588 17002 23624
rect 16946 23568 16948 23588
rect 16948 23568 17000 23588
rect 17000 23568 17002 23588
rect 16956 23418 17012 23420
rect 17036 23418 17092 23420
rect 17116 23418 17172 23420
rect 17196 23418 17252 23420
rect 16956 23366 17002 23418
rect 17002 23366 17012 23418
rect 17036 23366 17066 23418
rect 17066 23366 17078 23418
rect 17078 23366 17092 23418
rect 17116 23366 17130 23418
rect 17130 23366 17142 23418
rect 17142 23366 17172 23418
rect 17196 23366 17206 23418
rect 17206 23366 17252 23418
rect 16956 23364 17012 23366
rect 17036 23364 17092 23366
rect 17116 23364 17172 23366
rect 17196 23364 17252 23366
rect 17222 22500 17278 22536
rect 17222 22480 17224 22500
rect 17224 22480 17276 22500
rect 17276 22480 17278 22500
rect 16956 22330 17012 22332
rect 17036 22330 17092 22332
rect 17116 22330 17172 22332
rect 17196 22330 17252 22332
rect 16956 22278 17002 22330
rect 17002 22278 17012 22330
rect 17036 22278 17066 22330
rect 17066 22278 17078 22330
rect 17078 22278 17092 22330
rect 17116 22278 17130 22330
rect 17130 22278 17142 22330
rect 17142 22278 17172 22330
rect 17196 22278 17206 22330
rect 17206 22278 17252 22330
rect 16956 22276 17012 22278
rect 17036 22276 17092 22278
rect 17116 22276 17172 22278
rect 17196 22276 17252 22278
rect 16956 21242 17012 21244
rect 17036 21242 17092 21244
rect 17116 21242 17172 21244
rect 17196 21242 17252 21244
rect 16956 21190 17002 21242
rect 17002 21190 17012 21242
rect 17036 21190 17066 21242
rect 17066 21190 17078 21242
rect 17078 21190 17092 21242
rect 17116 21190 17130 21242
rect 17130 21190 17142 21242
rect 17142 21190 17172 21242
rect 17196 21190 17206 21242
rect 17206 21190 17252 21242
rect 16956 21188 17012 21190
rect 17036 21188 17092 21190
rect 17116 21188 17172 21190
rect 17196 21188 17252 21190
rect 17222 20984 17278 21040
rect 16956 20154 17012 20156
rect 17036 20154 17092 20156
rect 17116 20154 17172 20156
rect 17196 20154 17252 20156
rect 16956 20102 17002 20154
rect 17002 20102 17012 20154
rect 17036 20102 17066 20154
rect 17066 20102 17078 20154
rect 17078 20102 17092 20154
rect 17116 20102 17130 20154
rect 17130 20102 17142 20154
rect 17142 20102 17172 20154
rect 17196 20102 17206 20154
rect 17206 20102 17252 20154
rect 16956 20100 17012 20102
rect 17036 20100 17092 20102
rect 17116 20100 17172 20102
rect 17196 20100 17252 20102
rect 16578 13232 16634 13288
rect 16210 5228 16266 5264
rect 16210 5208 16212 5228
rect 16212 5208 16264 5228
rect 16264 5208 16266 5228
rect 12616 4378 12672 4380
rect 12696 4378 12752 4380
rect 12776 4378 12832 4380
rect 12856 4378 12912 4380
rect 12616 4326 12662 4378
rect 12662 4326 12672 4378
rect 12696 4326 12726 4378
rect 12726 4326 12738 4378
rect 12738 4326 12752 4378
rect 12776 4326 12790 4378
rect 12790 4326 12802 4378
rect 12802 4326 12832 4378
rect 12856 4326 12866 4378
rect 12866 4326 12912 4378
rect 12616 4324 12672 4326
rect 12696 4324 12752 4326
rect 12776 4324 12832 4326
rect 12856 4324 12912 4326
rect 11956 3834 12012 3836
rect 12036 3834 12092 3836
rect 12116 3834 12172 3836
rect 12196 3834 12252 3836
rect 11956 3782 12002 3834
rect 12002 3782 12012 3834
rect 12036 3782 12066 3834
rect 12066 3782 12078 3834
rect 12078 3782 12092 3834
rect 12116 3782 12130 3834
rect 12130 3782 12142 3834
rect 12142 3782 12172 3834
rect 12196 3782 12206 3834
rect 12206 3782 12252 3834
rect 11956 3780 12012 3782
rect 12036 3780 12092 3782
rect 12116 3780 12172 3782
rect 12196 3780 12252 3782
rect 12616 3290 12672 3292
rect 12696 3290 12752 3292
rect 12776 3290 12832 3292
rect 12856 3290 12912 3292
rect 12616 3238 12662 3290
rect 12662 3238 12672 3290
rect 12696 3238 12726 3290
rect 12726 3238 12738 3290
rect 12738 3238 12752 3290
rect 12776 3238 12790 3290
rect 12790 3238 12802 3290
rect 12802 3238 12832 3290
rect 12856 3238 12866 3290
rect 12866 3238 12912 3290
rect 12616 3236 12672 3238
rect 12696 3236 12752 3238
rect 12776 3236 12832 3238
rect 12856 3236 12912 3238
rect 11956 2746 12012 2748
rect 12036 2746 12092 2748
rect 12116 2746 12172 2748
rect 12196 2746 12252 2748
rect 11956 2694 12002 2746
rect 12002 2694 12012 2746
rect 12036 2694 12066 2746
rect 12066 2694 12078 2746
rect 12078 2694 12092 2746
rect 12116 2694 12130 2746
rect 12130 2694 12142 2746
rect 12142 2694 12172 2746
rect 12196 2694 12206 2746
rect 12206 2694 12252 2746
rect 11956 2692 12012 2694
rect 12036 2692 12092 2694
rect 12116 2692 12172 2694
rect 12196 2692 12252 2694
rect 16956 19066 17012 19068
rect 17036 19066 17092 19068
rect 17116 19066 17172 19068
rect 17196 19066 17252 19068
rect 16956 19014 17002 19066
rect 17002 19014 17012 19066
rect 17036 19014 17066 19066
rect 17066 19014 17078 19066
rect 17078 19014 17092 19066
rect 17116 19014 17130 19066
rect 17130 19014 17142 19066
rect 17142 19014 17172 19066
rect 17196 19014 17206 19066
rect 17206 19014 17252 19066
rect 16956 19012 17012 19014
rect 17036 19012 17092 19014
rect 17116 19012 17172 19014
rect 17196 19012 17252 19014
rect 16956 17978 17012 17980
rect 17036 17978 17092 17980
rect 17116 17978 17172 17980
rect 17196 17978 17252 17980
rect 16956 17926 17002 17978
rect 17002 17926 17012 17978
rect 17036 17926 17066 17978
rect 17066 17926 17078 17978
rect 17078 17926 17092 17978
rect 17116 17926 17130 17978
rect 17130 17926 17142 17978
rect 17142 17926 17172 17978
rect 17196 17926 17206 17978
rect 17206 17926 17252 17978
rect 16956 17924 17012 17926
rect 17036 17924 17092 17926
rect 17116 17924 17172 17926
rect 17196 17924 17252 17926
rect 16956 16890 17012 16892
rect 17036 16890 17092 16892
rect 17116 16890 17172 16892
rect 17196 16890 17252 16892
rect 16956 16838 17002 16890
rect 17002 16838 17012 16890
rect 17036 16838 17066 16890
rect 17066 16838 17078 16890
rect 17078 16838 17092 16890
rect 17116 16838 17130 16890
rect 17130 16838 17142 16890
rect 17142 16838 17172 16890
rect 17196 16838 17206 16890
rect 17206 16838 17252 16890
rect 16956 16836 17012 16838
rect 17036 16836 17092 16838
rect 17116 16836 17172 16838
rect 17196 16836 17252 16838
rect 16956 15802 17012 15804
rect 17036 15802 17092 15804
rect 17116 15802 17172 15804
rect 17196 15802 17252 15804
rect 16956 15750 17002 15802
rect 17002 15750 17012 15802
rect 17036 15750 17066 15802
rect 17066 15750 17078 15802
rect 17078 15750 17092 15802
rect 17116 15750 17130 15802
rect 17130 15750 17142 15802
rect 17142 15750 17172 15802
rect 17196 15750 17206 15802
rect 17206 15750 17252 15802
rect 16956 15748 17012 15750
rect 17036 15748 17092 15750
rect 17116 15748 17172 15750
rect 17196 15748 17252 15750
rect 16956 14714 17012 14716
rect 17036 14714 17092 14716
rect 17116 14714 17172 14716
rect 17196 14714 17252 14716
rect 16956 14662 17002 14714
rect 17002 14662 17012 14714
rect 17036 14662 17066 14714
rect 17066 14662 17078 14714
rect 17078 14662 17092 14714
rect 17116 14662 17130 14714
rect 17130 14662 17142 14714
rect 17142 14662 17172 14714
rect 17196 14662 17206 14714
rect 17206 14662 17252 14714
rect 16956 14660 17012 14662
rect 17036 14660 17092 14662
rect 17116 14660 17172 14662
rect 17196 14660 17252 14662
rect 16956 13626 17012 13628
rect 17036 13626 17092 13628
rect 17116 13626 17172 13628
rect 17196 13626 17252 13628
rect 16956 13574 17002 13626
rect 17002 13574 17012 13626
rect 17036 13574 17066 13626
rect 17066 13574 17078 13626
rect 17078 13574 17092 13626
rect 17116 13574 17130 13626
rect 17130 13574 17142 13626
rect 17142 13574 17172 13626
rect 17196 13574 17206 13626
rect 17206 13574 17252 13626
rect 16956 13572 17012 13574
rect 17036 13572 17092 13574
rect 17116 13572 17172 13574
rect 17196 13572 17252 13574
rect 17616 42458 17672 42460
rect 17696 42458 17752 42460
rect 17776 42458 17832 42460
rect 17856 42458 17912 42460
rect 17616 42406 17662 42458
rect 17662 42406 17672 42458
rect 17696 42406 17726 42458
rect 17726 42406 17738 42458
rect 17738 42406 17752 42458
rect 17776 42406 17790 42458
rect 17790 42406 17802 42458
rect 17802 42406 17832 42458
rect 17856 42406 17866 42458
rect 17866 42406 17912 42458
rect 17616 42404 17672 42406
rect 17696 42404 17752 42406
rect 17776 42404 17832 42406
rect 17856 42404 17912 42406
rect 17616 41370 17672 41372
rect 17696 41370 17752 41372
rect 17776 41370 17832 41372
rect 17856 41370 17912 41372
rect 17616 41318 17662 41370
rect 17662 41318 17672 41370
rect 17696 41318 17726 41370
rect 17726 41318 17738 41370
rect 17738 41318 17752 41370
rect 17776 41318 17790 41370
rect 17790 41318 17802 41370
rect 17802 41318 17832 41370
rect 17856 41318 17866 41370
rect 17866 41318 17912 41370
rect 17616 41316 17672 41318
rect 17696 41316 17752 41318
rect 17776 41316 17832 41318
rect 17856 41316 17912 41318
rect 17616 40282 17672 40284
rect 17696 40282 17752 40284
rect 17776 40282 17832 40284
rect 17856 40282 17912 40284
rect 17616 40230 17662 40282
rect 17662 40230 17672 40282
rect 17696 40230 17726 40282
rect 17726 40230 17738 40282
rect 17738 40230 17752 40282
rect 17776 40230 17790 40282
rect 17790 40230 17802 40282
rect 17802 40230 17832 40282
rect 17856 40230 17866 40282
rect 17866 40230 17912 40282
rect 17616 40228 17672 40230
rect 17696 40228 17752 40230
rect 17776 40228 17832 40230
rect 17856 40228 17912 40230
rect 17616 39194 17672 39196
rect 17696 39194 17752 39196
rect 17776 39194 17832 39196
rect 17856 39194 17912 39196
rect 17616 39142 17662 39194
rect 17662 39142 17672 39194
rect 17696 39142 17726 39194
rect 17726 39142 17738 39194
rect 17738 39142 17752 39194
rect 17776 39142 17790 39194
rect 17790 39142 17802 39194
rect 17802 39142 17832 39194
rect 17856 39142 17866 39194
rect 17866 39142 17912 39194
rect 17616 39140 17672 39142
rect 17696 39140 17752 39142
rect 17776 39140 17832 39142
rect 17856 39140 17912 39142
rect 17616 38106 17672 38108
rect 17696 38106 17752 38108
rect 17776 38106 17832 38108
rect 17856 38106 17912 38108
rect 17616 38054 17662 38106
rect 17662 38054 17672 38106
rect 17696 38054 17726 38106
rect 17726 38054 17738 38106
rect 17738 38054 17752 38106
rect 17776 38054 17790 38106
rect 17790 38054 17802 38106
rect 17802 38054 17832 38106
rect 17856 38054 17866 38106
rect 17866 38054 17912 38106
rect 17616 38052 17672 38054
rect 17696 38052 17752 38054
rect 17776 38052 17832 38054
rect 17856 38052 17912 38054
rect 17616 37018 17672 37020
rect 17696 37018 17752 37020
rect 17776 37018 17832 37020
rect 17856 37018 17912 37020
rect 17616 36966 17662 37018
rect 17662 36966 17672 37018
rect 17696 36966 17726 37018
rect 17726 36966 17738 37018
rect 17738 36966 17752 37018
rect 17776 36966 17790 37018
rect 17790 36966 17802 37018
rect 17802 36966 17832 37018
rect 17856 36966 17866 37018
rect 17866 36966 17912 37018
rect 17616 36964 17672 36966
rect 17696 36964 17752 36966
rect 17776 36964 17832 36966
rect 17856 36964 17912 36966
rect 17406 33904 17462 33960
rect 16956 12538 17012 12540
rect 17036 12538 17092 12540
rect 17116 12538 17172 12540
rect 17196 12538 17252 12540
rect 16956 12486 17002 12538
rect 17002 12486 17012 12538
rect 17036 12486 17066 12538
rect 17066 12486 17078 12538
rect 17078 12486 17092 12538
rect 17116 12486 17130 12538
rect 17130 12486 17142 12538
rect 17142 12486 17172 12538
rect 17196 12486 17206 12538
rect 17206 12486 17252 12538
rect 16956 12484 17012 12486
rect 17036 12484 17092 12486
rect 17116 12484 17172 12486
rect 17196 12484 17252 12486
rect 16956 11450 17012 11452
rect 17036 11450 17092 11452
rect 17116 11450 17172 11452
rect 17196 11450 17252 11452
rect 16956 11398 17002 11450
rect 17002 11398 17012 11450
rect 17036 11398 17066 11450
rect 17066 11398 17078 11450
rect 17078 11398 17092 11450
rect 17116 11398 17130 11450
rect 17130 11398 17142 11450
rect 17142 11398 17172 11450
rect 17196 11398 17206 11450
rect 17206 11398 17252 11450
rect 16956 11396 17012 11398
rect 17036 11396 17092 11398
rect 17116 11396 17172 11398
rect 17196 11396 17252 11398
rect 16956 10362 17012 10364
rect 17036 10362 17092 10364
rect 17116 10362 17172 10364
rect 17196 10362 17252 10364
rect 16956 10310 17002 10362
rect 17002 10310 17012 10362
rect 17036 10310 17066 10362
rect 17066 10310 17078 10362
rect 17078 10310 17092 10362
rect 17116 10310 17130 10362
rect 17130 10310 17142 10362
rect 17142 10310 17172 10362
rect 17196 10310 17206 10362
rect 17206 10310 17252 10362
rect 16956 10308 17012 10310
rect 17036 10308 17092 10310
rect 17116 10308 17172 10310
rect 17196 10308 17252 10310
rect 16956 9274 17012 9276
rect 17036 9274 17092 9276
rect 17116 9274 17172 9276
rect 17196 9274 17252 9276
rect 16956 9222 17002 9274
rect 17002 9222 17012 9274
rect 17036 9222 17066 9274
rect 17066 9222 17078 9274
rect 17078 9222 17092 9274
rect 17116 9222 17130 9274
rect 17130 9222 17142 9274
rect 17142 9222 17172 9274
rect 17196 9222 17206 9274
rect 17206 9222 17252 9274
rect 16956 9220 17012 9222
rect 17036 9220 17092 9222
rect 17116 9220 17172 9222
rect 17196 9220 17252 9222
rect 17616 35930 17672 35932
rect 17696 35930 17752 35932
rect 17776 35930 17832 35932
rect 17856 35930 17912 35932
rect 17616 35878 17662 35930
rect 17662 35878 17672 35930
rect 17696 35878 17726 35930
rect 17726 35878 17738 35930
rect 17738 35878 17752 35930
rect 17776 35878 17790 35930
rect 17790 35878 17802 35930
rect 17802 35878 17832 35930
rect 17856 35878 17866 35930
rect 17866 35878 17912 35930
rect 17616 35876 17672 35878
rect 17696 35876 17752 35878
rect 17776 35876 17832 35878
rect 17856 35876 17912 35878
rect 17616 34842 17672 34844
rect 17696 34842 17752 34844
rect 17776 34842 17832 34844
rect 17856 34842 17912 34844
rect 17616 34790 17662 34842
rect 17662 34790 17672 34842
rect 17696 34790 17726 34842
rect 17726 34790 17738 34842
rect 17738 34790 17752 34842
rect 17776 34790 17790 34842
rect 17790 34790 17802 34842
rect 17802 34790 17832 34842
rect 17856 34790 17866 34842
rect 17866 34790 17912 34842
rect 17616 34788 17672 34790
rect 17696 34788 17752 34790
rect 17776 34788 17832 34790
rect 17856 34788 17912 34790
rect 17616 33754 17672 33756
rect 17696 33754 17752 33756
rect 17776 33754 17832 33756
rect 17856 33754 17912 33756
rect 17616 33702 17662 33754
rect 17662 33702 17672 33754
rect 17696 33702 17726 33754
rect 17726 33702 17738 33754
rect 17738 33702 17752 33754
rect 17776 33702 17790 33754
rect 17790 33702 17802 33754
rect 17802 33702 17832 33754
rect 17856 33702 17866 33754
rect 17866 33702 17912 33754
rect 17616 33700 17672 33702
rect 17696 33700 17752 33702
rect 17776 33700 17832 33702
rect 17856 33700 17912 33702
rect 17616 32666 17672 32668
rect 17696 32666 17752 32668
rect 17776 32666 17832 32668
rect 17856 32666 17912 32668
rect 17616 32614 17662 32666
rect 17662 32614 17672 32666
rect 17696 32614 17726 32666
rect 17726 32614 17738 32666
rect 17738 32614 17752 32666
rect 17776 32614 17790 32666
rect 17790 32614 17802 32666
rect 17802 32614 17832 32666
rect 17856 32614 17866 32666
rect 17866 32614 17912 32666
rect 17616 32612 17672 32614
rect 17696 32612 17752 32614
rect 17776 32612 17832 32614
rect 17856 32612 17912 32614
rect 18234 54168 18290 54224
rect 18234 52264 18290 52320
rect 18234 50360 18290 50416
rect 18234 48492 18236 48512
rect 18236 48492 18288 48512
rect 18288 48492 18290 48512
rect 18234 48456 18290 48492
rect 18234 46552 18290 46608
rect 18234 44684 18236 44704
rect 18236 44684 18288 44704
rect 18288 44684 18290 44704
rect 18234 44648 18290 44684
rect 17616 31578 17672 31580
rect 17696 31578 17752 31580
rect 17776 31578 17832 31580
rect 17856 31578 17912 31580
rect 17616 31526 17662 31578
rect 17662 31526 17672 31578
rect 17696 31526 17726 31578
rect 17726 31526 17738 31578
rect 17738 31526 17752 31578
rect 17776 31526 17790 31578
rect 17790 31526 17802 31578
rect 17802 31526 17832 31578
rect 17856 31526 17866 31578
rect 17866 31526 17912 31578
rect 17616 31524 17672 31526
rect 17696 31524 17752 31526
rect 17776 31524 17832 31526
rect 17856 31524 17912 31526
rect 17616 30490 17672 30492
rect 17696 30490 17752 30492
rect 17776 30490 17832 30492
rect 17856 30490 17912 30492
rect 17616 30438 17662 30490
rect 17662 30438 17672 30490
rect 17696 30438 17726 30490
rect 17726 30438 17738 30490
rect 17738 30438 17752 30490
rect 17776 30438 17790 30490
rect 17790 30438 17802 30490
rect 17802 30438 17832 30490
rect 17856 30438 17866 30490
rect 17866 30438 17912 30490
rect 17616 30436 17672 30438
rect 17696 30436 17752 30438
rect 17776 30436 17832 30438
rect 17856 30436 17912 30438
rect 17616 29402 17672 29404
rect 17696 29402 17752 29404
rect 17776 29402 17832 29404
rect 17856 29402 17912 29404
rect 17616 29350 17662 29402
rect 17662 29350 17672 29402
rect 17696 29350 17726 29402
rect 17726 29350 17738 29402
rect 17738 29350 17752 29402
rect 17776 29350 17790 29402
rect 17790 29350 17802 29402
rect 17802 29350 17832 29402
rect 17856 29350 17866 29402
rect 17866 29350 17912 29402
rect 17616 29348 17672 29350
rect 17696 29348 17752 29350
rect 17776 29348 17832 29350
rect 17856 29348 17912 29350
rect 17616 28314 17672 28316
rect 17696 28314 17752 28316
rect 17776 28314 17832 28316
rect 17856 28314 17912 28316
rect 17616 28262 17662 28314
rect 17662 28262 17672 28314
rect 17696 28262 17726 28314
rect 17726 28262 17738 28314
rect 17738 28262 17752 28314
rect 17776 28262 17790 28314
rect 17790 28262 17802 28314
rect 17802 28262 17832 28314
rect 17856 28262 17866 28314
rect 17866 28262 17912 28314
rect 17616 28260 17672 28262
rect 17696 28260 17752 28262
rect 17776 28260 17832 28262
rect 17856 28260 17912 28262
rect 17866 27512 17922 27568
rect 17616 27226 17672 27228
rect 17696 27226 17752 27228
rect 17776 27226 17832 27228
rect 17856 27226 17912 27228
rect 17616 27174 17662 27226
rect 17662 27174 17672 27226
rect 17696 27174 17726 27226
rect 17726 27174 17738 27226
rect 17738 27174 17752 27226
rect 17776 27174 17790 27226
rect 17790 27174 17802 27226
rect 17802 27174 17832 27226
rect 17856 27174 17866 27226
rect 17866 27174 17912 27226
rect 17616 27172 17672 27174
rect 17696 27172 17752 27174
rect 17776 27172 17832 27174
rect 17856 27172 17912 27174
rect 17616 26138 17672 26140
rect 17696 26138 17752 26140
rect 17776 26138 17832 26140
rect 17856 26138 17912 26140
rect 17616 26086 17662 26138
rect 17662 26086 17672 26138
rect 17696 26086 17726 26138
rect 17726 26086 17738 26138
rect 17738 26086 17752 26138
rect 17776 26086 17790 26138
rect 17790 26086 17802 26138
rect 17802 26086 17832 26138
rect 17856 26086 17866 26138
rect 17866 26086 17912 26138
rect 17616 26084 17672 26086
rect 17696 26084 17752 26086
rect 17776 26084 17832 26086
rect 17856 26084 17912 26086
rect 16956 8186 17012 8188
rect 17036 8186 17092 8188
rect 17116 8186 17172 8188
rect 17196 8186 17252 8188
rect 16956 8134 17002 8186
rect 17002 8134 17012 8186
rect 17036 8134 17066 8186
rect 17066 8134 17078 8186
rect 17078 8134 17092 8186
rect 17116 8134 17130 8186
rect 17130 8134 17142 8186
rect 17142 8134 17172 8186
rect 17196 8134 17206 8186
rect 17206 8134 17252 8186
rect 16956 8132 17012 8134
rect 17036 8132 17092 8134
rect 17116 8132 17172 8134
rect 17196 8132 17252 8134
rect 16956 7098 17012 7100
rect 17036 7098 17092 7100
rect 17116 7098 17172 7100
rect 17196 7098 17252 7100
rect 16956 7046 17002 7098
rect 17002 7046 17012 7098
rect 17036 7046 17066 7098
rect 17066 7046 17078 7098
rect 17078 7046 17092 7098
rect 17116 7046 17130 7098
rect 17130 7046 17142 7098
rect 17142 7046 17172 7098
rect 17196 7046 17206 7098
rect 17206 7046 17252 7098
rect 16956 7044 17012 7046
rect 17036 7044 17092 7046
rect 17116 7044 17172 7046
rect 17196 7044 17252 7046
rect 16956 6010 17012 6012
rect 17036 6010 17092 6012
rect 17116 6010 17172 6012
rect 17196 6010 17252 6012
rect 16956 5958 17002 6010
rect 17002 5958 17012 6010
rect 17036 5958 17066 6010
rect 17066 5958 17078 6010
rect 17078 5958 17092 6010
rect 17116 5958 17130 6010
rect 17130 5958 17142 6010
rect 17142 5958 17172 6010
rect 17196 5958 17206 6010
rect 17206 5958 17252 6010
rect 16956 5956 17012 5958
rect 17036 5956 17092 5958
rect 17116 5956 17172 5958
rect 17196 5956 17252 5958
rect 17616 25050 17672 25052
rect 17696 25050 17752 25052
rect 17776 25050 17832 25052
rect 17856 25050 17912 25052
rect 17616 24998 17662 25050
rect 17662 24998 17672 25050
rect 17696 24998 17726 25050
rect 17726 24998 17738 25050
rect 17738 24998 17752 25050
rect 17776 24998 17790 25050
rect 17790 24998 17802 25050
rect 17802 24998 17832 25050
rect 17856 24998 17866 25050
rect 17866 24998 17912 25050
rect 17616 24996 17672 24998
rect 17696 24996 17752 24998
rect 17776 24996 17832 24998
rect 17856 24996 17912 24998
rect 18234 42744 18290 42800
rect 18234 42608 18290 42664
rect 18234 41928 18290 41984
rect 18234 40876 18236 40896
rect 18236 40876 18288 40896
rect 18288 40876 18290 40896
rect 18234 40840 18290 40876
rect 18234 38936 18290 38992
rect 18234 37068 18236 37088
rect 18236 37068 18288 37088
rect 18288 37068 18290 37088
rect 18234 37032 18290 37068
rect 18234 35128 18290 35184
rect 18234 33260 18236 33280
rect 18236 33260 18288 33280
rect 18288 33260 18290 33280
rect 18234 33224 18290 33260
rect 18234 31320 18290 31376
rect 18234 29452 18236 29472
rect 18236 29452 18288 29472
rect 18288 29452 18290 29472
rect 18234 29416 18290 29452
rect 18234 25644 18236 25664
rect 18236 25644 18288 25664
rect 18288 25644 18290 25664
rect 18234 25608 18290 25644
rect 17616 23962 17672 23964
rect 17696 23962 17752 23964
rect 17776 23962 17832 23964
rect 17856 23962 17912 23964
rect 17616 23910 17662 23962
rect 17662 23910 17672 23962
rect 17696 23910 17726 23962
rect 17726 23910 17738 23962
rect 17738 23910 17752 23962
rect 17776 23910 17790 23962
rect 17790 23910 17802 23962
rect 17802 23910 17832 23962
rect 17856 23910 17866 23962
rect 17866 23910 17912 23962
rect 17616 23908 17672 23910
rect 17696 23908 17752 23910
rect 17776 23908 17832 23910
rect 17856 23908 17912 23910
rect 17616 22874 17672 22876
rect 17696 22874 17752 22876
rect 17776 22874 17832 22876
rect 17856 22874 17912 22876
rect 17616 22822 17662 22874
rect 17662 22822 17672 22874
rect 17696 22822 17726 22874
rect 17726 22822 17738 22874
rect 17738 22822 17752 22874
rect 17776 22822 17790 22874
rect 17790 22822 17802 22874
rect 17802 22822 17832 22874
rect 17856 22822 17866 22874
rect 17866 22822 17912 22874
rect 17616 22820 17672 22822
rect 17696 22820 17752 22822
rect 17776 22820 17832 22822
rect 17856 22820 17912 22822
rect 17616 21786 17672 21788
rect 17696 21786 17752 21788
rect 17776 21786 17832 21788
rect 17856 21786 17912 21788
rect 17616 21734 17662 21786
rect 17662 21734 17672 21786
rect 17696 21734 17726 21786
rect 17726 21734 17738 21786
rect 17738 21734 17752 21786
rect 17776 21734 17790 21786
rect 17790 21734 17802 21786
rect 17802 21734 17832 21786
rect 17856 21734 17866 21786
rect 17866 21734 17912 21786
rect 17616 21732 17672 21734
rect 17696 21732 17752 21734
rect 17776 21732 17832 21734
rect 17856 21732 17912 21734
rect 17616 20698 17672 20700
rect 17696 20698 17752 20700
rect 17776 20698 17832 20700
rect 17856 20698 17912 20700
rect 17616 20646 17662 20698
rect 17662 20646 17672 20698
rect 17696 20646 17726 20698
rect 17726 20646 17738 20698
rect 17738 20646 17752 20698
rect 17776 20646 17790 20698
rect 17790 20646 17802 20698
rect 17802 20646 17832 20698
rect 17856 20646 17866 20698
rect 17866 20646 17912 20698
rect 17616 20644 17672 20646
rect 17696 20644 17752 20646
rect 17776 20644 17832 20646
rect 17856 20644 17912 20646
rect 18234 23704 18290 23760
rect 18234 21836 18236 21856
rect 18236 21836 18288 21856
rect 18288 21836 18290 21856
rect 18234 21800 18290 21836
rect 18234 19932 18236 19952
rect 18236 19932 18288 19952
rect 18288 19932 18290 19952
rect 18234 19896 18290 19932
rect 17616 19610 17672 19612
rect 17696 19610 17752 19612
rect 17776 19610 17832 19612
rect 17856 19610 17912 19612
rect 17616 19558 17662 19610
rect 17662 19558 17672 19610
rect 17696 19558 17726 19610
rect 17726 19558 17738 19610
rect 17738 19558 17752 19610
rect 17776 19558 17790 19610
rect 17790 19558 17802 19610
rect 17802 19558 17832 19610
rect 17856 19558 17866 19610
rect 17866 19558 17912 19610
rect 17616 19556 17672 19558
rect 17696 19556 17752 19558
rect 17776 19556 17832 19558
rect 17856 19556 17912 19558
rect 17616 18522 17672 18524
rect 17696 18522 17752 18524
rect 17776 18522 17832 18524
rect 17856 18522 17912 18524
rect 17616 18470 17662 18522
rect 17662 18470 17672 18522
rect 17696 18470 17726 18522
rect 17726 18470 17738 18522
rect 17738 18470 17752 18522
rect 17776 18470 17790 18522
rect 17790 18470 17802 18522
rect 17802 18470 17832 18522
rect 17856 18470 17866 18522
rect 17866 18470 17912 18522
rect 17616 18468 17672 18470
rect 17696 18468 17752 18470
rect 17776 18468 17832 18470
rect 17856 18468 17912 18470
rect 18234 18028 18236 18048
rect 18236 18028 18288 18048
rect 18288 18028 18290 18048
rect 18234 17992 18290 18028
rect 17616 17434 17672 17436
rect 17696 17434 17752 17436
rect 17776 17434 17832 17436
rect 17856 17434 17912 17436
rect 17616 17382 17662 17434
rect 17662 17382 17672 17434
rect 17696 17382 17726 17434
rect 17726 17382 17738 17434
rect 17738 17382 17752 17434
rect 17776 17382 17790 17434
rect 17790 17382 17802 17434
rect 17802 17382 17832 17434
rect 17856 17382 17866 17434
rect 17866 17382 17912 17434
rect 17616 17380 17672 17382
rect 17696 17380 17752 17382
rect 17776 17380 17832 17382
rect 17856 17380 17912 17382
rect 17958 16632 18014 16688
rect 17616 16346 17672 16348
rect 17696 16346 17752 16348
rect 17776 16346 17832 16348
rect 17856 16346 17912 16348
rect 17616 16294 17662 16346
rect 17662 16294 17672 16346
rect 17696 16294 17726 16346
rect 17726 16294 17738 16346
rect 17738 16294 17752 16346
rect 17776 16294 17790 16346
rect 17790 16294 17802 16346
rect 17802 16294 17832 16346
rect 17856 16294 17866 16346
rect 17866 16294 17912 16346
rect 17616 16292 17672 16294
rect 17696 16292 17752 16294
rect 17776 16292 17832 16294
rect 17856 16292 17912 16294
rect 18234 16088 18290 16144
rect 18602 41928 18658 41984
rect 17616 15258 17672 15260
rect 17696 15258 17752 15260
rect 17776 15258 17832 15260
rect 17856 15258 17912 15260
rect 17616 15206 17662 15258
rect 17662 15206 17672 15258
rect 17696 15206 17726 15258
rect 17726 15206 17738 15258
rect 17738 15206 17752 15258
rect 17776 15206 17790 15258
rect 17790 15206 17802 15258
rect 17802 15206 17832 15258
rect 17856 15206 17866 15258
rect 17866 15206 17912 15258
rect 17616 15204 17672 15206
rect 17696 15204 17752 15206
rect 17776 15204 17832 15206
rect 17856 15204 17912 15206
rect 17682 14884 17738 14920
rect 17682 14864 17684 14884
rect 17684 14864 17736 14884
rect 17736 14864 17738 14884
rect 17616 14170 17672 14172
rect 17696 14170 17752 14172
rect 17776 14170 17832 14172
rect 17856 14170 17912 14172
rect 17616 14118 17662 14170
rect 17662 14118 17672 14170
rect 17696 14118 17726 14170
rect 17726 14118 17738 14170
rect 17738 14118 17752 14170
rect 17776 14118 17790 14170
rect 17790 14118 17802 14170
rect 17802 14118 17832 14170
rect 17856 14118 17866 14170
rect 17866 14118 17912 14170
rect 17616 14116 17672 14118
rect 17696 14116 17752 14118
rect 17776 14116 17832 14118
rect 17856 14116 17912 14118
rect 17616 13082 17672 13084
rect 17696 13082 17752 13084
rect 17776 13082 17832 13084
rect 17856 13082 17912 13084
rect 17616 13030 17662 13082
rect 17662 13030 17672 13082
rect 17696 13030 17726 13082
rect 17726 13030 17738 13082
rect 17738 13030 17752 13082
rect 17776 13030 17790 13082
rect 17790 13030 17802 13082
rect 17802 13030 17832 13082
rect 17856 13030 17866 13082
rect 17866 13030 17912 13082
rect 17616 13028 17672 13030
rect 17696 13028 17752 13030
rect 17776 13028 17832 13030
rect 17856 13028 17912 13030
rect 17616 11994 17672 11996
rect 17696 11994 17752 11996
rect 17776 11994 17832 11996
rect 17856 11994 17912 11996
rect 17616 11942 17662 11994
rect 17662 11942 17672 11994
rect 17696 11942 17726 11994
rect 17726 11942 17738 11994
rect 17738 11942 17752 11994
rect 17776 11942 17790 11994
rect 17790 11942 17802 11994
rect 17802 11942 17832 11994
rect 17856 11942 17866 11994
rect 17866 11942 17912 11994
rect 17616 11940 17672 11942
rect 17696 11940 17752 11942
rect 17776 11940 17832 11942
rect 17856 11940 17912 11942
rect 17616 10906 17672 10908
rect 17696 10906 17752 10908
rect 17776 10906 17832 10908
rect 17856 10906 17912 10908
rect 17616 10854 17662 10906
rect 17662 10854 17672 10906
rect 17696 10854 17726 10906
rect 17726 10854 17738 10906
rect 17738 10854 17752 10906
rect 17776 10854 17790 10906
rect 17790 10854 17802 10906
rect 17802 10854 17832 10906
rect 17856 10854 17866 10906
rect 17866 10854 17912 10906
rect 17616 10852 17672 10854
rect 17696 10852 17752 10854
rect 17776 10852 17832 10854
rect 17856 10852 17912 10854
rect 17616 9818 17672 9820
rect 17696 9818 17752 9820
rect 17776 9818 17832 9820
rect 17856 9818 17912 9820
rect 17616 9766 17662 9818
rect 17662 9766 17672 9818
rect 17696 9766 17726 9818
rect 17726 9766 17738 9818
rect 17738 9766 17752 9818
rect 17776 9766 17790 9818
rect 17790 9766 17802 9818
rect 17802 9766 17832 9818
rect 17856 9766 17866 9818
rect 17866 9766 17912 9818
rect 17616 9764 17672 9766
rect 17696 9764 17752 9766
rect 17776 9764 17832 9766
rect 17856 9764 17912 9766
rect 18234 14220 18236 14240
rect 18236 14220 18288 14240
rect 18288 14220 18290 14240
rect 18234 14184 18290 14220
rect 18234 12316 18236 12336
rect 18236 12316 18288 12336
rect 18288 12316 18290 12336
rect 18234 12280 18290 12316
rect 18234 10412 18236 10432
rect 18236 10412 18288 10432
rect 18288 10412 18290 10432
rect 18234 10376 18290 10412
rect 17616 8730 17672 8732
rect 17696 8730 17752 8732
rect 17776 8730 17832 8732
rect 17856 8730 17912 8732
rect 17616 8678 17662 8730
rect 17662 8678 17672 8730
rect 17696 8678 17726 8730
rect 17726 8678 17738 8730
rect 17738 8678 17752 8730
rect 17776 8678 17790 8730
rect 17790 8678 17802 8730
rect 17802 8678 17832 8730
rect 17856 8678 17866 8730
rect 17866 8678 17912 8730
rect 17616 8676 17672 8678
rect 17696 8676 17752 8678
rect 17776 8676 17832 8678
rect 17856 8676 17912 8678
rect 19246 51856 19302 51912
rect 17616 7642 17672 7644
rect 17696 7642 17752 7644
rect 17776 7642 17832 7644
rect 17856 7642 17912 7644
rect 17616 7590 17662 7642
rect 17662 7590 17672 7642
rect 17696 7590 17726 7642
rect 17726 7590 17738 7642
rect 17738 7590 17752 7642
rect 17776 7590 17790 7642
rect 17790 7590 17802 7642
rect 17802 7590 17832 7642
rect 17856 7590 17866 7642
rect 17866 7590 17912 7642
rect 17616 7588 17672 7590
rect 17696 7588 17752 7590
rect 17776 7588 17832 7590
rect 17856 7588 17912 7590
rect 17616 6554 17672 6556
rect 17696 6554 17752 6556
rect 17776 6554 17832 6556
rect 17856 6554 17912 6556
rect 17616 6502 17662 6554
rect 17662 6502 17672 6554
rect 17696 6502 17726 6554
rect 17726 6502 17738 6554
rect 17738 6502 17752 6554
rect 17776 6502 17790 6554
rect 17790 6502 17802 6554
rect 17802 6502 17832 6554
rect 17856 6502 17866 6554
rect 17866 6502 17912 6554
rect 17616 6500 17672 6502
rect 17696 6500 17752 6502
rect 17776 6500 17832 6502
rect 17856 6500 17912 6502
rect 17616 5466 17672 5468
rect 17696 5466 17752 5468
rect 17776 5466 17832 5468
rect 17856 5466 17912 5468
rect 17616 5414 17662 5466
rect 17662 5414 17672 5466
rect 17696 5414 17726 5466
rect 17726 5414 17738 5466
rect 17738 5414 17752 5466
rect 17776 5414 17790 5466
rect 17790 5414 17802 5466
rect 17802 5414 17832 5466
rect 17856 5414 17866 5466
rect 17866 5414 17912 5466
rect 17616 5412 17672 5414
rect 17696 5412 17752 5414
rect 17776 5412 17832 5414
rect 17856 5412 17912 5414
rect 16956 4922 17012 4924
rect 17036 4922 17092 4924
rect 17116 4922 17172 4924
rect 17196 4922 17252 4924
rect 16956 4870 17002 4922
rect 17002 4870 17012 4922
rect 17036 4870 17066 4922
rect 17066 4870 17078 4922
rect 17078 4870 17092 4922
rect 17116 4870 17130 4922
rect 17130 4870 17142 4922
rect 17142 4870 17172 4922
rect 17196 4870 17206 4922
rect 17206 4870 17252 4922
rect 16956 4868 17012 4870
rect 17036 4868 17092 4870
rect 17116 4868 17172 4870
rect 17196 4868 17252 4870
rect 17616 4378 17672 4380
rect 17696 4378 17752 4380
rect 17776 4378 17832 4380
rect 17856 4378 17912 4380
rect 17616 4326 17662 4378
rect 17662 4326 17672 4378
rect 17696 4326 17726 4378
rect 17726 4326 17738 4378
rect 17738 4326 17752 4378
rect 17776 4326 17790 4378
rect 17790 4326 17802 4378
rect 17802 4326 17832 4378
rect 17856 4326 17866 4378
rect 17866 4326 17912 4378
rect 17616 4324 17672 4326
rect 17696 4324 17752 4326
rect 17776 4324 17832 4326
rect 17856 4324 17912 4326
rect 16956 3834 17012 3836
rect 17036 3834 17092 3836
rect 17116 3834 17172 3836
rect 17196 3834 17252 3836
rect 16956 3782 17002 3834
rect 17002 3782 17012 3834
rect 17036 3782 17066 3834
rect 17066 3782 17078 3834
rect 17078 3782 17092 3834
rect 17116 3782 17130 3834
rect 17130 3782 17142 3834
rect 17142 3782 17172 3834
rect 17196 3782 17206 3834
rect 17206 3782 17252 3834
rect 16956 3780 17012 3782
rect 17036 3780 17092 3782
rect 17116 3780 17172 3782
rect 17196 3780 17252 3782
rect 17616 3290 17672 3292
rect 17696 3290 17752 3292
rect 17776 3290 17832 3292
rect 17856 3290 17912 3292
rect 17616 3238 17662 3290
rect 17662 3238 17672 3290
rect 17696 3238 17726 3290
rect 17726 3238 17738 3290
rect 17738 3238 17752 3290
rect 17776 3238 17790 3290
rect 17790 3238 17802 3290
rect 17802 3238 17832 3290
rect 17856 3238 17866 3290
rect 17866 3238 17912 3290
rect 17616 3236 17672 3238
rect 17696 3236 17752 3238
rect 17776 3236 17832 3238
rect 17856 3236 17912 3238
rect 16956 2746 17012 2748
rect 17036 2746 17092 2748
rect 17116 2746 17172 2748
rect 17196 2746 17252 2748
rect 16956 2694 17002 2746
rect 17002 2694 17012 2746
rect 17036 2694 17066 2746
rect 17066 2694 17078 2746
rect 17078 2694 17092 2746
rect 17116 2694 17130 2746
rect 17130 2694 17142 2746
rect 17142 2694 17172 2746
rect 17196 2694 17206 2746
rect 17206 2694 17252 2746
rect 16956 2692 17012 2694
rect 17036 2692 17092 2694
rect 17116 2692 17172 2694
rect 17196 2692 17252 2694
rect 18234 8472 18290 8528
rect 18234 6604 18236 6624
rect 18236 6604 18288 6624
rect 18288 6604 18290 6624
rect 18234 6568 18290 6604
rect 18234 4664 18290 4720
rect 18234 2796 18236 2816
rect 18236 2796 18288 2816
rect 18288 2796 18290 2816
rect 18234 2760 18290 2796
rect 2616 2202 2672 2204
rect 2696 2202 2752 2204
rect 2776 2202 2832 2204
rect 2856 2202 2912 2204
rect 2616 2150 2662 2202
rect 2662 2150 2672 2202
rect 2696 2150 2726 2202
rect 2726 2150 2738 2202
rect 2738 2150 2752 2202
rect 2776 2150 2790 2202
rect 2790 2150 2802 2202
rect 2802 2150 2832 2202
rect 2856 2150 2866 2202
rect 2866 2150 2912 2202
rect 2616 2148 2672 2150
rect 2696 2148 2752 2150
rect 2776 2148 2832 2150
rect 2856 2148 2912 2150
rect 7616 2202 7672 2204
rect 7696 2202 7752 2204
rect 7776 2202 7832 2204
rect 7856 2202 7912 2204
rect 7616 2150 7662 2202
rect 7662 2150 7672 2202
rect 7696 2150 7726 2202
rect 7726 2150 7738 2202
rect 7738 2150 7752 2202
rect 7776 2150 7790 2202
rect 7790 2150 7802 2202
rect 7802 2150 7832 2202
rect 7856 2150 7866 2202
rect 7866 2150 7912 2202
rect 7616 2148 7672 2150
rect 7696 2148 7752 2150
rect 7776 2148 7832 2150
rect 7856 2148 7912 2150
rect 12616 2202 12672 2204
rect 12696 2202 12752 2204
rect 12776 2202 12832 2204
rect 12856 2202 12912 2204
rect 12616 2150 12662 2202
rect 12662 2150 12672 2202
rect 12696 2150 12726 2202
rect 12726 2150 12738 2202
rect 12738 2150 12752 2202
rect 12776 2150 12790 2202
rect 12790 2150 12802 2202
rect 12802 2150 12832 2202
rect 12856 2150 12866 2202
rect 12866 2150 12912 2202
rect 12616 2148 12672 2150
rect 12696 2148 12752 2150
rect 12776 2148 12832 2150
rect 12856 2148 12912 2150
rect 17616 2202 17672 2204
rect 17696 2202 17752 2204
rect 17776 2202 17832 2204
rect 17856 2202 17912 2204
rect 17616 2150 17662 2202
rect 17662 2150 17672 2202
rect 17696 2150 17726 2202
rect 17726 2150 17738 2202
rect 17738 2150 17752 2202
rect 17776 2150 17790 2202
rect 17790 2150 17802 2202
rect 17802 2150 17832 2202
rect 17856 2150 17866 2202
rect 17866 2150 17912 2202
rect 17616 2148 17672 2150
rect 17696 2148 17752 2150
rect 17776 2148 17832 2150
rect 17856 2148 17912 2150
<< metal3 >>
rect 1946 77824 2262 77825
rect 1946 77760 1952 77824
rect 2016 77760 2032 77824
rect 2096 77760 2112 77824
rect 2176 77760 2192 77824
rect 2256 77760 2262 77824
rect 1946 77759 2262 77760
rect 6946 77824 7262 77825
rect 6946 77760 6952 77824
rect 7016 77760 7032 77824
rect 7096 77760 7112 77824
rect 7176 77760 7192 77824
rect 7256 77760 7262 77824
rect 6946 77759 7262 77760
rect 11946 77824 12262 77825
rect 11946 77760 11952 77824
rect 12016 77760 12032 77824
rect 12096 77760 12112 77824
rect 12176 77760 12192 77824
rect 12256 77760 12262 77824
rect 11946 77759 12262 77760
rect 16946 77824 17262 77825
rect 16946 77760 16952 77824
rect 17016 77760 17032 77824
rect 17096 77760 17112 77824
rect 17176 77760 17192 77824
rect 17256 77760 17262 77824
rect 16946 77759 17262 77760
rect 2606 77280 2922 77281
rect 2606 77216 2612 77280
rect 2676 77216 2692 77280
rect 2756 77216 2772 77280
rect 2836 77216 2852 77280
rect 2916 77216 2922 77280
rect 2606 77215 2922 77216
rect 7606 77280 7922 77281
rect 7606 77216 7612 77280
rect 7676 77216 7692 77280
rect 7756 77216 7772 77280
rect 7836 77216 7852 77280
rect 7916 77216 7922 77280
rect 7606 77215 7922 77216
rect 12606 77280 12922 77281
rect 12606 77216 12612 77280
rect 12676 77216 12692 77280
rect 12756 77216 12772 77280
rect 12836 77216 12852 77280
rect 12916 77216 12922 77280
rect 12606 77215 12922 77216
rect 17606 77280 17922 77281
rect 17606 77216 17612 77280
rect 17676 77216 17692 77280
rect 17756 77216 17772 77280
rect 17836 77216 17852 77280
rect 17916 77216 17922 77280
rect 17606 77215 17922 77216
rect 18229 77074 18295 77077
rect 19200 77074 20000 77104
rect 18229 77072 20000 77074
rect 18229 77016 18234 77072
rect 18290 77016 20000 77072
rect 18229 77014 20000 77016
rect 18229 77011 18295 77014
rect 19200 76984 20000 77014
rect 14641 76804 14707 76805
rect 15929 76804 15995 76805
rect 14590 76740 14596 76804
rect 14660 76802 14707 76804
rect 14660 76800 14752 76802
rect 14702 76744 14752 76800
rect 14660 76742 14752 76744
rect 14660 76740 14707 76742
rect 15878 76740 15884 76804
rect 15948 76802 15995 76804
rect 15948 76800 16040 76802
rect 15990 76744 16040 76800
rect 15948 76742 16040 76744
rect 15948 76740 15995 76742
rect 14641 76739 14707 76740
rect 15929 76739 15995 76740
rect 1946 76736 2262 76737
rect 1946 76672 1952 76736
rect 2016 76672 2032 76736
rect 2096 76672 2112 76736
rect 2176 76672 2192 76736
rect 2256 76672 2262 76736
rect 1946 76671 2262 76672
rect 6946 76736 7262 76737
rect 6946 76672 6952 76736
rect 7016 76672 7032 76736
rect 7096 76672 7112 76736
rect 7176 76672 7192 76736
rect 7256 76672 7262 76736
rect 6946 76671 7262 76672
rect 11946 76736 12262 76737
rect 11946 76672 11952 76736
rect 12016 76672 12032 76736
rect 12096 76672 12112 76736
rect 12176 76672 12192 76736
rect 12256 76672 12262 76736
rect 11946 76671 12262 76672
rect 16946 76736 17262 76737
rect 16946 76672 16952 76736
rect 17016 76672 17032 76736
rect 17096 76672 17112 76736
rect 17176 76672 17192 76736
rect 17256 76672 17262 76736
rect 16946 76671 17262 76672
rect 6126 76332 6132 76396
rect 6196 76394 6202 76396
rect 8477 76394 8543 76397
rect 6196 76392 8543 76394
rect 6196 76336 8482 76392
rect 8538 76336 8543 76392
rect 6196 76334 8543 76336
rect 6196 76332 6202 76334
rect 8477 76331 8543 76334
rect 11237 76260 11303 76261
rect 11237 76258 11284 76260
rect 11192 76256 11284 76258
rect 11192 76200 11242 76256
rect 11192 76198 11284 76200
rect 11237 76196 11284 76198
rect 11348 76196 11354 76260
rect 11237 76195 11303 76196
rect 2606 76192 2922 76193
rect 2606 76128 2612 76192
rect 2676 76128 2692 76192
rect 2756 76128 2772 76192
rect 2836 76128 2852 76192
rect 2916 76128 2922 76192
rect 2606 76127 2922 76128
rect 7606 76192 7922 76193
rect 7606 76128 7612 76192
rect 7676 76128 7692 76192
rect 7756 76128 7772 76192
rect 7836 76128 7852 76192
rect 7916 76128 7922 76192
rect 7606 76127 7922 76128
rect 12606 76192 12922 76193
rect 12606 76128 12612 76192
rect 12676 76128 12692 76192
rect 12756 76128 12772 76192
rect 12836 76128 12852 76192
rect 12916 76128 12922 76192
rect 12606 76127 12922 76128
rect 17606 76192 17922 76193
rect 17606 76128 17612 76192
rect 17676 76128 17692 76192
rect 17756 76128 17772 76192
rect 17836 76128 17852 76192
rect 17916 76128 17922 76192
rect 17606 76127 17922 76128
rect 8753 76122 8819 76125
rect 8886 76122 8892 76124
rect 8753 76120 8892 76122
rect 8753 76064 8758 76120
rect 8814 76064 8892 76120
rect 8753 76062 8892 76064
rect 8753 76059 8819 76062
rect 8886 76060 8892 76062
rect 8956 76060 8962 76124
rect 7557 75986 7623 75989
rect 14222 75986 14228 75988
rect 7557 75984 14228 75986
rect 7557 75928 7562 75984
rect 7618 75928 14228 75984
rect 7557 75926 14228 75928
rect 7557 75923 7623 75926
rect 14222 75924 14228 75926
rect 14292 75924 14298 75988
rect 1946 75648 2262 75649
rect 1946 75584 1952 75648
rect 2016 75584 2032 75648
rect 2096 75584 2112 75648
rect 2176 75584 2192 75648
rect 2256 75584 2262 75648
rect 1946 75583 2262 75584
rect 6946 75648 7262 75649
rect 6946 75584 6952 75648
rect 7016 75584 7032 75648
rect 7096 75584 7112 75648
rect 7176 75584 7192 75648
rect 7256 75584 7262 75648
rect 6946 75583 7262 75584
rect 11946 75648 12262 75649
rect 11946 75584 11952 75648
rect 12016 75584 12032 75648
rect 12096 75584 12112 75648
rect 12176 75584 12192 75648
rect 12256 75584 12262 75648
rect 11946 75583 12262 75584
rect 16946 75648 17262 75649
rect 16946 75584 16952 75648
rect 17016 75584 17032 75648
rect 17096 75584 17112 75648
rect 17176 75584 17192 75648
rect 17256 75584 17262 75648
rect 16946 75583 17262 75584
rect 6545 75170 6611 75173
rect 6678 75170 6684 75172
rect 6545 75168 6684 75170
rect 6545 75112 6550 75168
rect 6606 75112 6684 75168
rect 6545 75110 6684 75112
rect 6545 75107 6611 75110
rect 6678 75108 6684 75110
rect 6748 75108 6754 75172
rect 18229 75170 18295 75173
rect 19200 75170 20000 75200
rect 18229 75168 20000 75170
rect 18229 75112 18234 75168
rect 18290 75112 20000 75168
rect 18229 75110 20000 75112
rect 18229 75107 18295 75110
rect 2606 75104 2922 75105
rect 2606 75040 2612 75104
rect 2676 75040 2692 75104
rect 2756 75040 2772 75104
rect 2836 75040 2852 75104
rect 2916 75040 2922 75104
rect 2606 75039 2922 75040
rect 7606 75104 7922 75105
rect 7606 75040 7612 75104
rect 7676 75040 7692 75104
rect 7756 75040 7772 75104
rect 7836 75040 7852 75104
rect 7916 75040 7922 75104
rect 7606 75039 7922 75040
rect 12606 75104 12922 75105
rect 12606 75040 12612 75104
rect 12676 75040 12692 75104
rect 12756 75040 12772 75104
rect 12836 75040 12852 75104
rect 12916 75040 12922 75104
rect 12606 75039 12922 75040
rect 17606 75104 17922 75105
rect 17606 75040 17612 75104
rect 17676 75040 17692 75104
rect 17756 75040 17772 75104
rect 17836 75040 17852 75104
rect 17916 75040 17922 75104
rect 19200 75080 20000 75110
rect 17606 75039 17922 75040
rect 1946 74560 2262 74561
rect 1946 74496 1952 74560
rect 2016 74496 2032 74560
rect 2096 74496 2112 74560
rect 2176 74496 2192 74560
rect 2256 74496 2262 74560
rect 1946 74495 2262 74496
rect 6946 74560 7262 74561
rect 6946 74496 6952 74560
rect 7016 74496 7032 74560
rect 7096 74496 7112 74560
rect 7176 74496 7192 74560
rect 7256 74496 7262 74560
rect 6946 74495 7262 74496
rect 11946 74560 12262 74561
rect 11946 74496 11952 74560
rect 12016 74496 12032 74560
rect 12096 74496 12112 74560
rect 12176 74496 12192 74560
rect 12256 74496 12262 74560
rect 11946 74495 12262 74496
rect 16946 74560 17262 74561
rect 16946 74496 16952 74560
rect 17016 74496 17032 74560
rect 17096 74496 17112 74560
rect 17176 74496 17192 74560
rect 17256 74496 17262 74560
rect 16946 74495 17262 74496
rect 2606 74016 2922 74017
rect 2606 73952 2612 74016
rect 2676 73952 2692 74016
rect 2756 73952 2772 74016
rect 2836 73952 2852 74016
rect 2916 73952 2922 74016
rect 2606 73951 2922 73952
rect 7606 74016 7922 74017
rect 7606 73952 7612 74016
rect 7676 73952 7692 74016
rect 7756 73952 7772 74016
rect 7836 73952 7852 74016
rect 7916 73952 7922 74016
rect 7606 73951 7922 73952
rect 12606 74016 12922 74017
rect 12606 73952 12612 74016
rect 12676 73952 12692 74016
rect 12756 73952 12772 74016
rect 12836 73952 12852 74016
rect 12916 73952 12922 74016
rect 12606 73951 12922 73952
rect 17606 74016 17922 74017
rect 17606 73952 17612 74016
rect 17676 73952 17692 74016
rect 17756 73952 17772 74016
rect 17836 73952 17852 74016
rect 17916 73952 17922 74016
rect 17606 73951 17922 73952
rect 1946 73472 2262 73473
rect 1946 73408 1952 73472
rect 2016 73408 2032 73472
rect 2096 73408 2112 73472
rect 2176 73408 2192 73472
rect 2256 73408 2262 73472
rect 1946 73407 2262 73408
rect 6946 73472 7262 73473
rect 6946 73408 6952 73472
rect 7016 73408 7032 73472
rect 7096 73408 7112 73472
rect 7176 73408 7192 73472
rect 7256 73408 7262 73472
rect 6946 73407 7262 73408
rect 11946 73472 12262 73473
rect 11946 73408 11952 73472
rect 12016 73408 12032 73472
rect 12096 73408 12112 73472
rect 12176 73408 12192 73472
rect 12256 73408 12262 73472
rect 11946 73407 12262 73408
rect 16946 73472 17262 73473
rect 16946 73408 16952 73472
rect 17016 73408 17032 73472
rect 17096 73408 17112 73472
rect 17176 73408 17192 73472
rect 17256 73408 17262 73472
rect 16946 73407 17262 73408
rect 18229 73266 18295 73269
rect 19200 73266 20000 73296
rect 18229 73264 20000 73266
rect 18229 73208 18234 73264
rect 18290 73208 20000 73264
rect 18229 73206 20000 73208
rect 18229 73203 18295 73206
rect 19200 73176 20000 73206
rect 2606 72928 2922 72929
rect 2606 72864 2612 72928
rect 2676 72864 2692 72928
rect 2756 72864 2772 72928
rect 2836 72864 2852 72928
rect 2916 72864 2922 72928
rect 2606 72863 2922 72864
rect 7606 72928 7922 72929
rect 7606 72864 7612 72928
rect 7676 72864 7692 72928
rect 7756 72864 7772 72928
rect 7836 72864 7852 72928
rect 7916 72864 7922 72928
rect 7606 72863 7922 72864
rect 12606 72928 12922 72929
rect 12606 72864 12612 72928
rect 12676 72864 12692 72928
rect 12756 72864 12772 72928
rect 12836 72864 12852 72928
rect 12916 72864 12922 72928
rect 12606 72863 12922 72864
rect 17606 72928 17922 72929
rect 17606 72864 17612 72928
rect 17676 72864 17692 72928
rect 17756 72864 17772 72928
rect 17836 72864 17852 72928
rect 17916 72864 17922 72928
rect 17606 72863 17922 72864
rect 1946 72384 2262 72385
rect 1946 72320 1952 72384
rect 2016 72320 2032 72384
rect 2096 72320 2112 72384
rect 2176 72320 2192 72384
rect 2256 72320 2262 72384
rect 1946 72319 2262 72320
rect 6946 72384 7262 72385
rect 6946 72320 6952 72384
rect 7016 72320 7032 72384
rect 7096 72320 7112 72384
rect 7176 72320 7192 72384
rect 7256 72320 7262 72384
rect 6946 72319 7262 72320
rect 11946 72384 12262 72385
rect 11946 72320 11952 72384
rect 12016 72320 12032 72384
rect 12096 72320 12112 72384
rect 12176 72320 12192 72384
rect 12256 72320 12262 72384
rect 11946 72319 12262 72320
rect 16946 72384 17262 72385
rect 16946 72320 16952 72384
rect 17016 72320 17032 72384
rect 17096 72320 17112 72384
rect 17176 72320 17192 72384
rect 17256 72320 17262 72384
rect 16946 72319 17262 72320
rect 2606 71840 2922 71841
rect 2606 71776 2612 71840
rect 2676 71776 2692 71840
rect 2756 71776 2772 71840
rect 2836 71776 2852 71840
rect 2916 71776 2922 71840
rect 2606 71775 2922 71776
rect 7606 71840 7922 71841
rect 7606 71776 7612 71840
rect 7676 71776 7692 71840
rect 7756 71776 7772 71840
rect 7836 71776 7852 71840
rect 7916 71776 7922 71840
rect 7606 71775 7922 71776
rect 12606 71840 12922 71841
rect 12606 71776 12612 71840
rect 12676 71776 12692 71840
rect 12756 71776 12772 71840
rect 12836 71776 12852 71840
rect 12916 71776 12922 71840
rect 12606 71775 12922 71776
rect 17606 71840 17922 71841
rect 17606 71776 17612 71840
rect 17676 71776 17692 71840
rect 17756 71776 17772 71840
rect 17836 71776 17852 71840
rect 17916 71776 17922 71840
rect 17606 71775 17922 71776
rect 18229 71362 18295 71365
rect 19200 71362 20000 71392
rect 18229 71360 20000 71362
rect 18229 71304 18234 71360
rect 18290 71304 20000 71360
rect 18229 71302 20000 71304
rect 18229 71299 18295 71302
rect 1946 71296 2262 71297
rect 1946 71232 1952 71296
rect 2016 71232 2032 71296
rect 2096 71232 2112 71296
rect 2176 71232 2192 71296
rect 2256 71232 2262 71296
rect 1946 71231 2262 71232
rect 6946 71296 7262 71297
rect 6946 71232 6952 71296
rect 7016 71232 7032 71296
rect 7096 71232 7112 71296
rect 7176 71232 7192 71296
rect 7256 71232 7262 71296
rect 6946 71231 7262 71232
rect 11946 71296 12262 71297
rect 11946 71232 11952 71296
rect 12016 71232 12032 71296
rect 12096 71232 12112 71296
rect 12176 71232 12192 71296
rect 12256 71232 12262 71296
rect 11946 71231 12262 71232
rect 16946 71296 17262 71297
rect 16946 71232 16952 71296
rect 17016 71232 17032 71296
rect 17096 71232 17112 71296
rect 17176 71232 17192 71296
rect 17256 71232 17262 71296
rect 19200 71272 20000 71302
rect 16946 71231 17262 71232
rect 3325 70956 3391 70957
rect 3325 70952 3372 70956
rect 3436 70954 3442 70956
rect 3325 70896 3330 70952
rect 3325 70892 3372 70896
rect 3436 70894 3482 70954
rect 3436 70892 3442 70894
rect 3325 70891 3391 70892
rect 2606 70752 2922 70753
rect 2606 70688 2612 70752
rect 2676 70688 2692 70752
rect 2756 70688 2772 70752
rect 2836 70688 2852 70752
rect 2916 70688 2922 70752
rect 2606 70687 2922 70688
rect 7606 70752 7922 70753
rect 7606 70688 7612 70752
rect 7676 70688 7692 70752
rect 7756 70688 7772 70752
rect 7836 70688 7852 70752
rect 7916 70688 7922 70752
rect 7606 70687 7922 70688
rect 12606 70752 12922 70753
rect 12606 70688 12612 70752
rect 12676 70688 12692 70752
rect 12756 70688 12772 70752
rect 12836 70688 12852 70752
rect 12916 70688 12922 70752
rect 12606 70687 12922 70688
rect 17606 70752 17922 70753
rect 17606 70688 17612 70752
rect 17676 70688 17692 70752
rect 17756 70688 17772 70752
rect 17836 70688 17852 70752
rect 17916 70688 17922 70752
rect 17606 70687 17922 70688
rect 1946 70208 2262 70209
rect 1946 70144 1952 70208
rect 2016 70144 2032 70208
rect 2096 70144 2112 70208
rect 2176 70144 2192 70208
rect 2256 70144 2262 70208
rect 1946 70143 2262 70144
rect 6946 70208 7262 70209
rect 6946 70144 6952 70208
rect 7016 70144 7032 70208
rect 7096 70144 7112 70208
rect 7176 70144 7192 70208
rect 7256 70144 7262 70208
rect 6946 70143 7262 70144
rect 11946 70208 12262 70209
rect 11946 70144 11952 70208
rect 12016 70144 12032 70208
rect 12096 70144 12112 70208
rect 12176 70144 12192 70208
rect 12256 70144 12262 70208
rect 11946 70143 12262 70144
rect 16946 70208 17262 70209
rect 16946 70144 16952 70208
rect 17016 70144 17032 70208
rect 17096 70144 17112 70208
rect 17176 70144 17192 70208
rect 17256 70144 17262 70208
rect 16946 70143 17262 70144
rect 2606 69664 2922 69665
rect 2606 69600 2612 69664
rect 2676 69600 2692 69664
rect 2756 69600 2772 69664
rect 2836 69600 2852 69664
rect 2916 69600 2922 69664
rect 2606 69599 2922 69600
rect 7606 69664 7922 69665
rect 7606 69600 7612 69664
rect 7676 69600 7692 69664
rect 7756 69600 7772 69664
rect 7836 69600 7852 69664
rect 7916 69600 7922 69664
rect 7606 69599 7922 69600
rect 12606 69664 12922 69665
rect 12606 69600 12612 69664
rect 12676 69600 12692 69664
rect 12756 69600 12772 69664
rect 12836 69600 12852 69664
rect 12916 69600 12922 69664
rect 12606 69599 12922 69600
rect 17606 69664 17922 69665
rect 17606 69600 17612 69664
rect 17676 69600 17692 69664
rect 17756 69600 17772 69664
rect 17836 69600 17852 69664
rect 17916 69600 17922 69664
rect 17606 69599 17922 69600
rect 18229 69458 18295 69461
rect 19200 69458 20000 69488
rect 18229 69456 20000 69458
rect 18229 69400 18234 69456
rect 18290 69400 20000 69456
rect 18229 69398 20000 69400
rect 18229 69395 18295 69398
rect 19200 69368 20000 69398
rect 1710 69260 1716 69324
rect 1780 69322 1786 69324
rect 2037 69322 2103 69325
rect 1780 69320 2103 69322
rect 1780 69264 2042 69320
rect 2098 69264 2103 69320
rect 1780 69262 2103 69264
rect 1780 69260 1786 69262
rect 2037 69259 2103 69262
rect 1946 69120 2262 69121
rect 1946 69056 1952 69120
rect 2016 69056 2032 69120
rect 2096 69056 2112 69120
rect 2176 69056 2192 69120
rect 2256 69056 2262 69120
rect 1946 69055 2262 69056
rect 6946 69120 7262 69121
rect 6946 69056 6952 69120
rect 7016 69056 7032 69120
rect 7096 69056 7112 69120
rect 7176 69056 7192 69120
rect 7256 69056 7262 69120
rect 6946 69055 7262 69056
rect 11946 69120 12262 69121
rect 11946 69056 11952 69120
rect 12016 69056 12032 69120
rect 12096 69056 12112 69120
rect 12176 69056 12192 69120
rect 12256 69056 12262 69120
rect 11946 69055 12262 69056
rect 16946 69120 17262 69121
rect 16946 69056 16952 69120
rect 17016 69056 17032 69120
rect 17096 69056 17112 69120
rect 17176 69056 17192 69120
rect 17256 69056 17262 69120
rect 16946 69055 17262 69056
rect 15009 69052 15075 69053
rect 14958 69050 14964 69052
rect 14918 68990 14964 69050
rect 15028 69048 15075 69052
rect 15070 68992 15075 69048
rect 14958 68988 14964 68990
rect 15028 68988 15075 68992
rect 15009 68987 15075 68988
rect 2606 68576 2922 68577
rect 2606 68512 2612 68576
rect 2676 68512 2692 68576
rect 2756 68512 2772 68576
rect 2836 68512 2852 68576
rect 2916 68512 2922 68576
rect 2606 68511 2922 68512
rect 7606 68576 7922 68577
rect 7606 68512 7612 68576
rect 7676 68512 7692 68576
rect 7756 68512 7772 68576
rect 7836 68512 7852 68576
rect 7916 68512 7922 68576
rect 7606 68511 7922 68512
rect 12606 68576 12922 68577
rect 12606 68512 12612 68576
rect 12676 68512 12692 68576
rect 12756 68512 12772 68576
rect 12836 68512 12852 68576
rect 12916 68512 12922 68576
rect 12606 68511 12922 68512
rect 17606 68576 17922 68577
rect 17606 68512 17612 68576
rect 17676 68512 17692 68576
rect 17756 68512 17772 68576
rect 17836 68512 17852 68576
rect 17916 68512 17922 68576
rect 17606 68511 17922 68512
rect 1946 68032 2262 68033
rect 1946 67968 1952 68032
rect 2016 67968 2032 68032
rect 2096 67968 2112 68032
rect 2176 67968 2192 68032
rect 2256 67968 2262 68032
rect 1946 67967 2262 67968
rect 6946 68032 7262 68033
rect 6946 67968 6952 68032
rect 7016 67968 7032 68032
rect 7096 67968 7112 68032
rect 7176 67968 7192 68032
rect 7256 67968 7262 68032
rect 6946 67967 7262 67968
rect 11946 68032 12262 68033
rect 11946 67968 11952 68032
rect 12016 67968 12032 68032
rect 12096 67968 12112 68032
rect 12176 67968 12192 68032
rect 12256 67968 12262 68032
rect 11946 67967 12262 67968
rect 16946 68032 17262 68033
rect 16946 67968 16952 68032
rect 17016 67968 17032 68032
rect 17096 67968 17112 68032
rect 17176 67968 17192 68032
rect 17256 67968 17262 68032
rect 16946 67967 17262 67968
rect 10358 67628 10364 67692
rect 10428 67690 10434 67692
rect 10501 67690 10567 67693
rect 10428 67688 10567 67690
rect 10428 67632 10506 67688
rect 10562 67632 10567 67688
rect 10428 67630 10567 67632
rect 10428 67628 10434 67630
rect 10501 67627 10567 67630
rect 11646 67628 11652 67692
rect 11716 67690 11722 67692
rect 12065 67690 12131 67693
rect 11716 67688 12131 67690
rect 11716 67632 12070 67688
rect 12126 67632 12131 67688
rect 11716 67630 12131 67632
rect 11716 67628 11722 67630
rect 12065 67627 12131 67630
rect 18229 67554 18295 67557
rect 19200 67554 20000 67584
rect 18229 67552 20000 67554
rect 18229 67496 18234 67552
rect 18290 67496 20000 67552
rect 18229 67494 20000 67496
rect 18229 67491 18295 67494
rect 2606 67488 2922 67489
rect 2606 67424 2612 67488
rect 2676 67424 2692 67488
rect 2756 67424 2772 67488
rect 2836 67424 2852 67488
rect 2916 67424 2922 67488
rect 2606 67423 2922 67424
rect 7606 67488 7922 67489
rect 7606 67424 7612 67488
rect 7676 67424 7692 67488
rect 7756 67424 7772 67488
rect 7836 67424 7852 67488
rect 7916 67424 7922 67488
rect 7606 67423 7922 67424
rect 12606 67488 12922 67489
rect 12606 67424 12612 67488
rect 12676 67424 12692 67488
rect 12756 67424 12772 67488
rect 12836 67424 12852 67488
rect 12916 67424 12922 67488
rect 12606 67423 12922 67424
rect 17606 67488 17922 67489
rect 17606 67424 17612 67488
rect 17676 67424 17692 67488
rect 17756 67424 17772 67488
rect 17836 67424 17852 67488
rect 17916 67424 17922 67488
rect 19200 67464 20000 67494
rect 17606 67423 17922 67424
rect 1946 66944 2262 66945
rect 1946 66880 1952 66944
rect 2016 66880 2032 66944
rect 2096 66880 2112 66944
rect 2176 66880 2192 66944
rect 2256 66880 2262 66944
rect 1946 66879 2262 66880
rect 6946 66944 7262 66945
rect 6946 66880 6952 66944
rect 7016 66880 7032 66944
rect 7096 66880 7112 66944
rect 7176 66880 7192 66944
rect 7256 66880 7262 66944
rect 6946 66879 7262 66880
rect 11946 66944 12262 66945
rect 11946 66880 11952 66944
rect 12016 66880 12032 66944
rect 12096 66880 12112 66944
rect 12176 66880 12192 66944
rect 12256 66880 12262 66944
rect 11946 66879 12262 66880
rect 16946 66944 17262 66945
rect 16946 66880 16952 66944
rect 17016 66880 17032 66944
rect 17096 66880 17112 66944
rect 17176 66880 17192 66944
rect 17256 66880 17262 66944
rect 16946 66879 17262 66880
rect 2606 66400 2922 66401
rect 2606 66336 2612 66400
rect 2676 66336 2692 66400
rect 2756 66336 2772 66400
rect 2836 66336 2852 66400
rect 2916 66336 2922 66400
rect 2606 66335 2922 66336
rect 7606 66400 7922 66401
rect 7606 66336 7612 66400
rect 7676 66336 7692 66400
rect 7756 66336 7772 66400
rect 7836 66336 7852 66400
rect 7916 66336 7922 66400
rect 7606 66335 7922 66336
rect 12606 66400 12922 66401
rect 12606 66336 12612 66400
rect 12676 66336 12692 66400
rect 12756 66336 12772 66400
rect 12836 66336 12852 66400
rect 12916 66336 12922 66400
rect 12606 66335 12922 66336
rect 17606 66400 17922 66401
rect 17606 66336 17612 66400
rect 17676 66336 17692 66400
rect 17756 66336 17772 66400
rect 17836 66336 17852 66400
rect 17916 66336 17922 66400
rect 17606 66335 17922 66336
rect 1946 65856 2262 65857
rect 1946 65792 1952 65856
rect 2016 65792 2032 65856
rect 2096 65792 2112 65856
rect 2176 65792 2192 65856
rect 2256 65792 2262 65856
rect 1946 65791 2262 65792
rect 6946 65856 7262 65857
rect 6946 65792 6952 65856
rect 7016 65792 7032 65856
rect 7096 65792 7112 65856
rect 7176 65792 7192 65856
rect 7256 65792 7262 65856
rect 6946 65791 7262 65792
rect 11946 65856 12262 65857
rect 11946 65792 11952 65856
rect 12016 65792 12032 65856
rect 12096 65792 12112 65856
rect 12176 65792 12192 65856
rect 12256 65792 12262 65856
rect 11946 65791 12262 65792
rect 16946 65856 17262 65857
rect 16946 65792 16952 65856
rect 17016 65792 17032 65856
rect 17096 65792 17112 65856
rect 17176 65792 17192 65856
rect 17256 65792 17262 65856
rect 16946 65791 17262 65792
rect 18229 65650 18295 65653
rect 19200 65650 20000 65680
rect 18229 65648 20000 65650
rect 18229 65592 18234 65648
rect 18290 65592 20000 65648
rect 18229 65590 20000 65592
rect 18229 65587 18295 65590
rect 19200 65560 20000 65590
rect 2606 65312 2922 65313
rect 2606 65248 2612 65312
rect 2676 65248 2692 65312
rect 2756 65248 2772 65312
rect 2836 65248 2852 65312
rect 2916 65248 2922 65312
rect 2606 65247 2922 65248
rect 7606 65312 7922 65313
rect 7606 65248 7612 65312
rect 7676 65248 7692 65312
rect 7756 65248 7772 65312
rect 7836 65248 7852 65312
rect 7916 65248 7922 65312
rect 7606 65247 7922 65248
rect 12606 65312 12922 65313
rect 12606 65248 12612 65312
rect 12676 65248 12692 65312
rect 12756 65248 12772 65312
rect 12836 65248 12852 65312
rect 12916 65248 12922 65312
rect 12606 65247 12922 65248
rect 17606 65312 17922 65313
rect 17606 65248 17612 65312
rect 17676 65248 17692 65312
rect 17756 65248 17772 65312
rect 17836 65248 17852 65312
rect 17916 65248 17922 65312
rect 17606 65247 17922 65248
rect 3918 65180 3924 65244
rect 3988 65242 3994 65244
rect 4061 65242 4127 65245
rect 3988 65240 4127 65242
rect 3988 65184 4066 65240
rect 4122 65184 4127 65240
rect 3988 65182 4127 65184
rect 3988 65180 3994 65182
rect 4061 65179 4127 65182
rect 15694 65044 15700 65108
rect 15764 65106 15770 65108
rect 17493 65106 17559 65109
rect 15764 65104 17559 65106
rect 15764 65048 17498 65104
rect 17554 65048 17559 65104
rect 15764 65046 17559 65048
rect 15764 65044 15770 65046
rect 17493 65043 17559 65046
rect 1946 64768 2262 64769
rect 1946 64704 1952 64768
rect 2016 64704 2032 64768
rect 2096 64704 2112 64768
rect 2176 64704 2192 64768
rect 2256 64704 2262 64768
rect 1946 64703 2262 64704
rect 6946 64768 7262 64769
rect 6946 64704 6952 64768
rect 7016 64704 7032 64768
rect 7096 64704 7112 64768
rect 7176 64704 7192 64768
rect 7256 64704 7262 64768
rect 6946 64703 7262 64704
rect 11946 64768 12262 64769
rect 11946 64704 11952 64768
rect 12016 64704 12032 64768
rect 12096 64704 12112 64768
rect 12176 64704 12192 64768
rect 12256 64704 12262 64768
rect 11946 64703 12262 64704
rect 16946 64768 17262 64769
rect 16946 64704 16952 64768
rect 17016 64704 17032 64768
rect 17096 64704 17112 64768
rect 17176 64704 17192 64768
rect 17256 64704 17262 64768
rect 16946 64703 17262 64704
rect 2606 64224 2922 64225
rect 2606 64160 2612 64224
rect 2676 64160 2692 64224
rect 2756 64160 2772 64224
rect 2836 64160 2852 64224
rect 2916 64160 2922 64224
rect 2606 64159 2922 64160
rect 7606 64224 7922 64225
rect 7606 64160 7612 64224
rect 7676 64160 7692 64224
rect 7756 64160 7772 64224
rect 7836 64160 7852 64224
rect 7916 64160 7922 64224
rect 7606 64159 7922 64160
rect 12606 64224 12922 64225
rect 12606 64160 12612 64224
rect 12676 64160 12692 64224
rect 12756 64160 12772 64224
rect 12836 64160 12852 64224
rect 12916 64160 12922 64224
rect 12606 64159 12922 64160
rect 17606 64224 17922 64225
rect 17606 64160 17612 64224
rect 17676 64160 17692 64224
rect 17756 64160 17772 64224
rect 17836 64160 17852 64224
rect 17916 64160 17922 64224
rect 17606 64159 17922 64160
rect 18229 63746 18295 63749
rect 19200 63746 20000 63776
rect 18229 63744 20000 63746
rect 18229 63688 18234 63744
rect 18290 63688 20000 63744
rect 18229 63686 20000 63688
rect 18229 63683 18295 63686
rect 1946 63680 2262 63681
rect 1946 63616 1952 63680
rect 2016 63616 2032 63680
rect 2096 63616 2112 63680
rect 2176 63616 2192 63680
rect 2256 63616 2262 63680
rect 1946 63615 2262 63616
rect 6946 63680 7262 63681
rect 6946 63616 6952 63680
rect 7016 63616 7032 63680
rect 7096 63616 7112 63680
rect 7176 63616 7192 63680
rect 7256 63616 7262 63680
rect 6946 63615 7262 63616
rect 11946 63680 12262 63681
rect 11946 63616 11952 63680
rect 12016 63616 12032 63680
rect 12096 63616 12112 63680
rect 12176 63616 12192 63680
rect 12256 63616 12262 63680
rect 11946 63615 12262 63616
rect 16946 63680 17262 63681
rect 16946 63616 16952 63680
rect 17016 63616 17032 63680
rect 17096 63616 17112 63680
rect 17176 63616 17192 63680
rect 17256 63616 17262 63680
rect 19200 63656 20000 63686
rect 16946 63615 17262 63616
rect 4838 63276 4844 63340
rect 4908 63338 4914 63340
rect 14457 63338 14523 63341
rect 4908 63336 14523 63338
rect 4908 63280 14462 63336
rect 14518 63280 14523 63336
rect 4908 63278 14523 63280
rect 4908 63276 4914 63278
rect 14457 63275 14523 63278
rect 2606 63136 2922 63137
rect 2606 63072 2612 63136
rect 2676 63072 2692 63136
rect 2756 63072 2772 63136
rect 2836 63072 2852 63136
rect 2916 63072 2922 63136
rect 2606 63071 2922 63072
rect 7606 63136 7922 63137
rect 7606 63072 7612 63136
rect 7676 63072 7692 63136
rect 7756 63072 7772 63136
rect 7836 63072 7852 63136
rect 7916 63072 7922 63136
rect 7606 63071 7922 63072
rect 12606 63136 12922 63137
rect 12606 63072 12612 63136
rect 12676 63072 12692 63136
rect 12756 63072 12772 63136
rect 12836 63072 12852 63136
rect 12916 63072 12922 63136
rect 12606 63071 12922 63072
rect 17606 63136 17922 63137
rect 17606 63072 17612 63136
rect 17676 63072 17692 63136
rect 17756 63072 17772 63136
rect 17836 63072 17852 63136
rect 17916 63072 17922 63136
rect 17606 63071 17922 63072
rect 8753 62660 8819 62661
rect 8702 62596 8708 62660
rect 8772 62658 8819 62660
rect 8772 62656 8864 62658
rect 8814 62600 8864 62656
rect 8772 62598 8864 62600
rect 8772 62596 8819 62598
rect 8753 62595 8819 62596
rect 1946 62592 2262 62593
rect 1946 62528 1952 62592
rect 2016 62528 2032 62592
rect 2096 62528 2112 62592
rect 2176 62528 2192 62592
rect 2256 62528 2262 62592
rect 1946 62527 2262 62528
rect 6946 62592 7262 62593
rect 6946 62528 6952 62592
rect 7016 62528 7032 62592
rect 7096 62528 7112 62592
rect 7176 62528 7192 62592
rect 7256 62528 7262 62592
rect 6946 62527 7262 62528
rect 11946 62592 12262 62593
rect 11946 62528 11952 62592
rect 12016 62528 12032 62592
rect 12096 62528 12112 62592
rect 12176 62528 12192 62592
rect 12256 62528 12262 62592
rect 11946 62527 12262 62528
rect 16946 62592 17262 62593
rect 16946 62528 16952 62592
rect 17016 62528 17032 62592
rect 17096 62528 17112 62592
rect 17176 62528 17192 62592
rect 17256 62528 17262 62592
rect 16946 62527 17262 62528
rect 4245 62252 4311 62253
rect 4245 62248 4292 62252
rect 4356 62250 4362 62252
rect 4245 62192 4250 62248
rect 4245 62188 4292 62192
rect 4356 62190 4402 62250
rect 4356 62188 4362 62190
rect 4245 62187 4311 62188
rect 2606 62048 2922 62049
rect 2606 61984 2612 62048
rect 2676 61984 2692 62048
rect 2756 61984 2772 62048
rect 2836 61984 2852 62048
rect 2916 61984 2922 62048
rect 2606 61983 2922 61984
rect 7606 62048 7922 62049
rect 7606 61984 7612 62048
rect 7676 61984 7692 62048
rect 7756 61984 7772 62048
rect 7836 61984 7852 62048
rect 7916 61984 7922 62048
rect 7606 61983 7922 61984
rect 12606 62048 12922 62049
rect 12606 61984 12612 62048
rect 12676 61984 12692 62048
rect 12756 61984 12772 62048
rect 12836 61984 12852 62048
rect 12916 61984 12922 62048
rect 12606 61983 12922 61984
rect 17606 62048 17922 62049
rect 17606 61984 17612 62048
rect 17676 61984 17692 62048
rect 17756 61984 17772 62048
rect 17836 61984 17852 62048
rect 17916 61984 17922 62048
rect 17606 61983 17922 61984
rect 18229 61842 18295 61845
rect 19200 61842 20000 61872
rect 18229 61840 20000 61842
rect 18229 61784 18234 61840
rect 18290 61784 20000 61840
rect 18229 61782 20000 61784
rect 18229 61779 18295 61782
rect 19200 61752 20000 61782
rect 1946 61504 2262 61505
rect 1946 61440 1952 61504
rect 2016 61440 2032 61504
rect 2096 61440 2112 61504
rect 2176 61440 2192 61504
rect 2256 61440 2262 61504
rect 1946 61439 2262 61440
rect 6946 61504 7262 61505
rect 6946 61440 6952 61504
rect 7016 61440 7032 61504
rect 7096 61440 7112 61504
rect 7176 61440 7192 61504
rect 7256 61440 7262 61504
rect 6946 61439 7262 61440
rect 11946 61504 12262 61505
rect 11946 61440 11952 61504
rect 12016 61440 12032 61504
rect 12096 61440 12112 61504
rect 12176 61440 12192 61504
rect 12256 61440 12262 61504
rect 11946 61439 12262 61440
rect 16946 61504 17262 61505
rect 16946 61440 16952 61504
rect 17016 61440 17032 61504
rect 17096 61440 17112 61504
rect 17176 61440 17192 61504
rect 17256 61440 17262 61504
rect 16946 61439 17262 61440
rect 2606 60960 2922 60961
rect 2606 60896 2612 60960
rect 2676 60896 2692 60960
rect 2756 60896 2772 60960
rect 2836 60896 2852 60960
rect 2916 60896 2922 60960
rect 2606 60895 2922 60896
rect 7606 60960 7922 60961
rect 7606 60896 7612 60960
rect 7676 60896 7692 60960
rect 7756 60896 7772 60960
rect 7836 60896 7852 60960
rect 7916 60896 7922 60960
rect 7606 60895 7922 60896
rect 12606 60960 12922 60961
rect 12606 60896 12612 60960
rect 12676 60896 12692 60960
rect 12756 60896 12772 60960
rect 12836 60896 12852 60960
rect 12916 60896 12922 60960
rect 12606 60895 12922 60896
rect 17606 60960 17922 60961
rect 17606 60896 17612 60960
rect 17676 60896 17692 60960
rect 17756 60896 17772 60960
rect 17836 60896 17852 60960
rect 17916 60896 17922 60960
rect 17606 60895 17922 60896
rect 1946 60416 2262 60417
rect 1946 60352 1952 60416
rect 2016 60352 2032 60416
rect 2096 60352 2112 60416
rect 2176 60352 2192 60416
rect 2256 60352 2262 60416
rect 1946 60351 2262 60352
rect 6946 60416 7262 60417
rect 6946 60352 6952 60416
rect 7016 60352 7032 60416
rect 7096 60352 7112 60416
rect 7176 60352 7192 60416
rect 7256 60352 7262 60416
rect 6946 60351 7262 60352
rect 11946 60416 12262 60417
rect 11946 60352 11952 60416
rect 12016 60352 12032 60416
rect 12096 60352 12112 60416
rect 12176 60352 12192 60416
rect 12256 60352 12262 60416
rect 11946 60351 12262 60352
rect 16946 60416 17262 60417
rect 16946 60352 16952 60416
rect 17016 60352 17032 60416
rect 17096 60352 17112 60416
rect 17176 60352 17192 60416
rect 17256 60352 17262 60416
rect 16946 60351 17262 60352
rect 16389 60076 16455 60077
rect 16389 60074 16436 60076
rect 16344 60072 16436 60074
rect 16344 60016 16394 60072
rect 16344 60014 16436 60016
rect 16389 60012 16436 60014
rect 16500 60012 16506 60076
rect 16389 60011 16455 60012
rect 8109 59938 8175 59941
rect 9070 59938 9076 59940
rect 8109 59936 9076 59938
rect 8109 59880 8114 59936
rect 8170 59880 9076 59936
rect 8109 59878 9076 59880
rect 8109 59875 8175 59878
rect 9070 59876 9076 59878
rect 9140 59876 9146 59940
rect 18229 59938 18295 59941
rect 19200 59938 20000 59968
rect 18229 59936 20000 59938
rect 18229 59880 18234 59936
rect 18290 59880 20000 59936
rect 18229 59878 20000 59880
rect 18229 59875 18295 59878
rect 2606 59872 2922 59873
rect 2606 59808 2612 59872
rect 2676 59808 2692 59872
rect 2756 59808 2772 59872
rect 2836 59808 2852 59872
rect 2916 59808 2922 59872
rect 2606 59807 2922 59808
rect 7606 59872 7922 59873
rect 7606 59808 7612 59872
rect 7676 59808 7692 59872
rect 7756 59808 7772 59872
rect 7836 59808 7852 59872
rect 7916 59808 7922 59872
rect 7606 59807 7922 59808
rect 12606 59872 12922 59873
rect 12606 59808 12612 59872
rect 12676 59808 12692 59872
rect 12756 59808 12772 59872
rect 12836 59808 12852 59872
rect 12916 59808 12922 59872
rect 12606 59807 12922 59808
rect 17606 59872 17922 59873
rect 17606 59808 17612 59872
rect 17676 59808 17692 59872
rect 17756 59808 17772 59872
rect 17836 59808 17852 59872
rect 17916 59808 17922 59872
rect 19200 59848 20000 59878
rect 17606 59807 17922 59808
rect 1946 59328 2262 59329
rect 1946 59264 1952 59328
rect 2016 59264 2032 59328
rect 2096 59264 2112 59328
rect 2176 59264 2192 59328
rect 2256 59264 2262 59328
rect 1946 59263 2262 59264
rect 6946 59328 7262 59329
rect 6946 59264 6952 59328
rect 7016 59264 7032 59328
rect 7096 59264 7112 59328
rect 7176 59264 7192 59328
rect 7256 59264 7262 59328
rect 6946 59263 7262 59264
rect 11946 59328 12262 59329
rect 11946 59264 11952 59328
rect 12016 59264 12032 59328
rect 12096 59264 12112 59328
rect 12176 59264 12192 59328
rect 12256 59264 12262 59328
rect 11946 59263 12262 59264
rect 16946 59328 17262 59329
rect 16946 59264 16952 59328
rect 17016 59264 17032 59328
rect 17096 59264 17112 59328
rect 17176 59264 17192 59328
rect 17256 59264 17262 59328
rect 16946 59263 17262 59264
rect 13721 58852 13787 58853
rect 13670 58788 13676 58852
rect 13740 58850 13787 58852
rect 13740 58848 13832 58850
rect 13782 58792 13832 58848
rect 13740 58790 13832 58792
rect 13740 58788 13787 58790
rect 13721 58787 13787 58788
rect 2606 58784 2922 58785
rect 2606 58720 2612 58784
rect 2676 58720 2692 58784
rect 2756 58720 2772 58784
rect 2836 58720 2852 58784
rect 2916 58720 2922 58784
rect 2606 58719 2922 58720
rect 7606 58784 7922 58785
rect 7606 58720 7612 58784
rect 7676 58720 7692 58784
rect 7756 58720 7772 58784
rect 7836 58720 7852 58784
rect 7916 58720 7922 58784
rect 7606 58719 7922 58720
rect 12606 58784 12922 58785
rect 12606 58720 12612 58784
rect 12676 58720 12692 58784
rect 12756 58720 12772 58784
rect 12836 58720 12852 58784
rect 12916 58720 12922 58784
rect 12606 58719 12922 58720
rect 17606 58784 17922 58785
rect 17606 58720 17612 58784
rect 17676 58720 17692 58784
rect 17756 58720 17772 58784
rect 17836 58720 17852 58784
rect 17916 58720 17922 58784
rect 17606 58719 17922 58720
rect 1946 58240 2262 58241
rect 1946 58176 1952 58240
rect 2016 58176 2032 58240
rect 2096 58176 2112 58240
rect 2176 58176 2192 58240
rect 2256 58176 2262 58240
rect 1946 58175 2262 58176
rect 6946 58240 7262 58241
rect 6946 58176 6952 58240
rect 7016 58176 7032 58240
rect 7096 58176 7112 58240
rect 7176 58176 7192 58240
rect 7256 58176 7262 58240
rect 6946 58175 7262 58176
rect 11946 58240 12262 58241
rect 11946 58176 11952 58240
rect 12016 58176 12032 58240
rect 12096 58176 12112 58240
rect 12176 58176 12192 58240
rect 12256 58176 12262 58240
rect 11946 58175 12262 58176
rect 16946 58240 17262 58241
rect 16946 58176 16952 58240
rect 17016 58176 17032 58240
rect 17096 58176 17112 58240
rect 17176 58176 17192 58240
rect 17256 58176 17262 58240
rect 16946 58175 17262 58176
rect 18229 58034 18295 58037
rect 19200 58034 20000 58064
rect 18229 58032 20000 58034
rect 18229 57976 18234 58032
rect 18290 57976 20000 58032
rect 18229 57974 20000 57976
rect 18229 57971 18295 57974
rect 19200 57944 20000 57974
rect 2606 57696 2922 57697
rect 2606 57632 2612 57696
rect 2676 57632 2692 57696
rect 2756 57632 2772 57696
rect 2836 57632 2852 57696
rect 2916 57632 2922 57696
rect 2606 57631 2922 57632
rect 7606 57696 7922 57697
rect 7606 57632 7612 57696
rect 7676 57632 7692 57696
rect 7756 57632 7772 57696
rect 7836 57632 7852 57696
rect 7916 57632 7922 57696
rect 7606 57631 7922 57632
rect 12606 57696 12922 57697
rect 12606 57632 12612 57696
rect 12676 57632 12692 57696
rect 12756 57632 12772 57696
rect 12836 57632 12852 57696
rect 12916 57632 12922 57696
rect 12606 57631 12922 57632
rect 17606 57696 17922 57697
rect 17606 57632 17612 57696
rect 17676 57632 17692 57696
rect 17756 57632 17772 57696
rect 17836 57632 17852 57696
rect 17916 57632 17922 57696
rect 17606 57631 17922 57632
rect 1946 57152 2262 57153
rect 1946 57088 1952 57152
rect 2016 57088 2032 57152
rect 2096 57088 2112 57152
rect 2176 57088 2192 57152
rect 2256 57088 2262 57152
rect 1946 57087 2262 57088
rect 6946 57152 7262 57153
rect 6946 57088 6952 57152
rect 7016 57088 7032 57152
rect 7096 57088 7112 57152
rect 7176 57088 7192 57152
rect 7256 57088 7262 57152
rect 6946 57087 7262 57088
rect 11946 57152 12262 57153
rect 11946 57088 11952 57152
rect 12016 57088 12032 57152
rect 12096 57088 12112 57152
rect 12176 57088 12192 57152
rect 12256 57088 12262 57152
rect 11946 57087 12262 57088
rect 16946 57152 17262 57153
rect 16946 57088 16952 57152
rect 17016 57088 17032 57152
rect 17096 57088 17112 57152
rect 17176 57088 17192 57152
rect 17256 57088 17262 57152
rect 16946 57087 17262 57088
rect 3049 56674 3115 56677
rect 6310 56674 6316 56676
rect 3049 56672 6316 56674
rect 3049 56616 3054 56672
rect 3110 56616 6316 56672
rect 3049 56614 6316 56616
rect 3049 56611 3115 56614
rect 6310 56612 6316 56614
rect 6380 56612 6386 56676
rect 2606 56608 2922 56609
rect 2606 56544 2612 56608
rect 2676 56544 2692 56608
rect 2756 56544 2772 56608
rect 2836 56544 2852 56608
rect 2916 56544 2922 56608
rect 2606 56543 2922 56544
rect 7606 56608 7922 56609
rect 7606 56544 7612 56608
rect 7676 56544 7692 56608
rect 7756 56544 7772 56608
rect 7836 56544 7852 56608
rect 7916 56544 7922 56608
rect 7606 56543 7922 56544
rect 12606 56608 12922 56609
rect 12606 56544 12612 56608
rect 12676 56544 12692 56608
rect 12756 56544 12772 56608
rect 12836 56544 12852 56608
rect 12916 56544 12922 56608
rect 12606 56543 12922 56544
rect 17606 56608 17922 56609
rect 17606 56544 17612 56608
rect 17676 56544 17692 56608
rect 17756 56544 17772 56608
rect 17836 56544 17852 56608
rect 17916 56544 17922 56608
rect 17606 56543 17922 56544
rect 18229 56130 18295 56133
rect 19200 56130 20000 56160
rect 18229 56128 20000 56130
rect 18229 56072 18234 56128
rect 18290 56072 20000 56128
rect 18229 56070 20000 56072
rect 18229 56067 18295 56070
rect 1946 56064 2262 56065
rect 1946 56000 1952 56064
rect 2016 56000 2032 56064
rect 2096 56000 2112 56064
rect 2176 56000 2192 56064
rect 2256 56000 2262 56064
rect 1946 55999 2262 56000
rect 6946 56064 7262 56065
rect 6946 56000 6952 56064
rect 7016 56000 7032 56064
rect 7096 56000 7112 56064
rect 7176 56000 7192 56064
rect 7256 56000 7262 56064
rect 6946 55999 7262 56000
rect 11946 56064 12262 56065
rect 11946 56000 11952 56064
rect 12016 56000 12032 56064
rect 12096 56000 12112 56064
rect 12176 56000 12192 56064
rect 12256 56000 12262 56064
rect 11946 55999 12262 56000
rect 16946 56064 17262 56065
rect 16946 56000 16952 56064
rect 17016 56000 17032 56064
rect 17096 56000 17112 56064
rect 17176 56000 17192 56064
rect 17256 56000 17262 56064
rect 19200 56040 20000 56070
rect 16946 55999 17262 56000
rect 11421 55858 11487 55861
rect 11421 55856 14658 55858
rect 11421 55800 11426 55856
rect 11482 55800 14658 55856
rect 11421 55798 14658 55800
rect 11421 55795 11487 55798
rect 1526 55660 1532 55724
rect 1596 55722 1602 55724
rect 1669 55722 1735 55725
rect 1596 55720 1735 55722
rect 1596 55664 1674 55720
rect 1730 55664 1735 55720
rect 1596 55662 1735 55664
rect 1596 55660 1602 55662
rect 1669 55659 1735 55662
rect 12433 55722 12499 55725
rect 14406 55722 14412 55724
rect 12433 55720 14412 55722
rect 12433 55664 12438 55720
rect 12494 55664 14412 55720
rect 12433 55662 14412 55664
rect 12433 55659 12499 55662
rect 14406 55660 14412 55662
rect 14476 55660 14482 55724
rect 14598 55722 14658 55798
rect 16614 55722 16620 55724
rect 14598 55662 16620 55722
rect 16614 55660 16620 55662
rect 16684 55660 16690 55724
rect 2606 55520 2922 55521
rect 2606 55456 2612 55520
rect 2676 55456 2692 55520
rect 2756 55456 2772 55520
rect 2836 55456 2852 55520
rect 2916 55456 2922 55520
rect 2606 55455 2922 55456
rect 7606 55520 7922 55521
rect 7606 55456 7612 55520
rect 7676 55456 7692 55520
rect 7756 55456 7772 55520
rect 7836 55456 7852 55520
rect 7916 55456 7922 55520
rect 7606 55455 7922 55456
rect 12606 55520 12922 55521
rect 12606 55456 12612 55520
rect 12676 55456 12692 55520
rect 12756 55456 12772 55520
rect 12836 55456 12852 55520
rect 12916 55456 12922 55520
rect 12606 55455 12922 55456
rect 17606 55520 17922 55521
rect 17606 55456 17612 55520
rect 17676 55456 17692 55520
rect 17756 55456 17772 55520
rect 17836 55456 17852 55520
rect 17916 55456 17922 55520
rect 17606 55455 17922 55456
rect 1946 54976 2262 54977
rect 1946 54912 1952 54976
rect 2016 54912 2032 54976
rect 2096 54912 2112 54976
rect 2176 54912 2192 54976
rect 2256 54912 2262 54976
rect 1946 54911 2262 54912
rect 6946 54976 7262 54977
rect 6946 54912 6952 54976
rect 7016 54912 7032 54976
rect 7096 54912 7112 54976
rect 7176 54912 7192 54976
rect 7256 54912 7262 54976
rect 6946 54911 7262 54912
rect 11946 54976 12262 54977
rect 11946 54912 11952 54976
rect 12016 54912 12032 54976
rect 12096 54912 12112 54976
rect 12176 54912 12192 54976
rect 12256 54912 12262 54976
rect 11946 54911 12262 54912
rect 16946 54976 17262 54977
rect 16946 54912 16952 54976
rect 17016 54912 17032 54976
rect 17096 54912 17112 54976
rect 17176 54912 17192 54976
rect 17256 54912 17262 54976
rect 16946 54911 17262 54912
rect 2606 54432 2922 54433
rect 2606 54368 2612 54432
rect 2676 54368 2692 54432
rect 2756 54368 2772 54432
rect 2836 54368 2852 54432
rect 2916 54368 2922 54432
rect 2606 54367 2922 54368
rect 7606 54432 7922 54433
rect 7606 54368 7612 54432
rect 7676 54368 7692 54432
rect 7756 54368 7772 54432
rect 7836 54368 7852 54432
rect 7916 54368 7922 54432
rect 7606 54367 7922 54368
rect 12606 54432 12922 54433
rect 12606 54368 12612 54432
rect 12676 54368 12692 54432
rect 12756 54368 12772 54432
rect 12836 54368 12852 54432
rect 12916 54368 12922 54432
rect 12606 54367 12922 54368
rect 17606 54432 17922 54433
rect 17606 54368 17612 54432
rect 17676 54368 17692 54432
rect 17756 54368 17772 54432
rect 17836 54368 17852 54432
rect 17916 54368 17922 54432
rect 17606 54367 17922 54368
rect 18229 54226 18295 54229
rect 19200 54226 20000 54256
rect 18229 54224 20000 54226
rect 18229 54168 18234 54224
rect 18290 54168 20000 54224
rect 18229 54166 20000 54168
rect 18229 54163 18295 54166
rect 19200 54136 20000 54166
rect 10174 54028 10180 54092
rect 10244 54090 10250 54092
rect 12433 54090 12499 54093
rect 10244 54088 12499 54090
rect 10244 54032 12438 54088
rect 12494 54032 12499 54088
rect 10244 54030 12499 54032
rect 10244 54028 10250 54030
rect 12433 54027 12499 54030
rect 1946 53888 2262 53889
rect 1946 53824 1952 53888
rect 2016 53824 2032 53888
rect 2096 53824 2112 53888
rect 2176 53824 2192 53888
rect 2256 53824 2262 53888
rect 1946 53823 2262 53824
rect 6946 53888 7262 53889
rect 6946 53824 6952 53888
rect 7016 53824 7032 53888
rect 7096 53824 7112 53888
rect 7176 53824 7192 53888
rect 7256 53824 7262 53888
rect 6946 53823 7262 53824
rect 11946 53888 12262 53889
rect 11946 53824 11952 53888
rect 12016 53824 12032 53888
rect 12096 53824 12112 53888
rect 12176 53824 12192 53888
rect 12256 53824 12262 53888
rect 11946 53823 12262 53824
rect 16946 53888 17262 53889
rect 16946 53824 16952 53888
rect 17016 53824 17032 53888
rect 17096 53824 17112 53888
rect 17176 53824 17192 53888
rect 17256 53824 17262 53888
rect 16946 53823 17262 53824
rect 2606 53344 2922 53345
rect 2606 53280 2612 53344
rect 2676 53280 2692 53344
rect 2756 53280 2772 53344
rect 2836 53280 2852 53344
rect 2916 53280 2922 53344
rect 2606 53279 2922 53280
rect 7606 53344 7922 53345
rect 7606 53280 7612 53344
rect 7676 53280 7692 53344
rect 7756 53280 7772 53344
rect 7836 53280 7852 53344
rect 7916 53280 7922 53344
rect 7606 53279 7922 53280
rect 12606 53344 12922 53345
rect 12606 53280 12612 53344
rect 12676 53280 12692 53344
rect 12756 53280 12772 53344
rect 12836 53280 12852 53344
rect 12916 53280 12922 53344
rect 12606 53279 12922 53280
rect 17606 53344 17922 53345
rect 17606 53280 17612 53344
rect 17676 53280 17692 53344
rect 17756 53280 17772 53344
rect 17836 53280 17852 53344
rect 17916 53280 17922 53344
rect 17606 53279 17922 53280
rect 1946 52800 2262 52801
rect 1946 52736 1952 52800
rect 2016 52736 2032 52800
rect 2096 52736 2112 52800
rect 2176 52736 2192 52800
rect 2256 52736 2262 52800
rect 1946 52735 2262 52736
rect 6946 52800 7262 52801
rect 6946 52736 6952 52800
rect 7016 52736 7032 52800
rect 7096 52736 7112 52800
rect 7176 52736 7192 52800
rect 7256 52736 7262 52800
rect 6946 52735 7262 52736
rect 11946 52800 12262 52801
rect 11946 52736 11952 52800
rect 12016 52736 12032 52800
rect 12096 52736 12112 52800
rect 12176 52736 12192 52800
rect 12256 52736 12262 52800
rect 11946 52735 12262 52736
rect 16946 52800 17262 52801
rect 16946 52736 16952 52800
rect 17016 52736 17032 52800
rect 17096 52736 17112 52800
rect 17176 52736 17192 52800
rect 17256 52736 17262 52800
rect 16946 52735 17262 52736
rect 8518 52532 8524 52596
rect 8588 52594 8594 52596
rect 9489 52594 9555 52597
rect 8588 52592 9555 52594
rect 8588 52536 9494 52592
rect 9550 52536 9555 52592
rect 8588 52534 9555 52536
rect 8588 52532 8594 52534
rect 9489 52531 9555 52534
rect 10593 52458 10659 52461
rect 10910 52458 10916 52460
rect 10593 52456 10916 52458
rect 10593 52400 10598 52456
rect 10654 52400 10916 52456
rect 10593 52398 10916 52400
rect 10593 52395 10659 52398
rect 10910 52396 10916 52398
rect 10980 52396 10986 52460
rect 18229 52322 18295 52325
rect 19200 52322 20000 52352
rect 18229 52320 20000 52322
rect 18229 52264 18234 52320
rect 18290 52264 20000 52320
rect 18229 52262 20000 52264
rect 18229 52259 18295 52262
rect 2606 52256 2922 52257
rect 2606 52192 2612 52256
rect 2676 52192 2692 52256
rect 2756 52192 2772 52256
rect 2836 52192 2852 52256
rect 2916 52192 2922 52256
rect 2606 52191 2922 52192
rect 7606 52256 7922 52257
rect 7606 52192 7612 52256
rect 7676 52192 7692 52256
rect 7756 52192 7772 52256
rect 7836 52192 7852 52256
rect 7916 52192 7922 52256
rect 7606 52191 7922 52192
rect 12606 52256 12922 52257
rect 12606 52192 12612 52256
rect 12676 52192 12692 52256
rect 12756 52192 12772 52256
rect 12836 52192 12852 52256
rect 12916 52192 12922 52256
rect 12606 52191 12922 52192
rect 17606 52256 17922 52257
rect 17606 52192 17612 52256
rect 17676 52192 17692 52256
rect 17756 52192 17772 52256
rect 17836 52192 17852 52256
rect 17916 52192 17922 52256
rect 19200 52232 20000 52262
rect 17606 52191 17922 52192
rect 7833 51914 7899 51917
rect 8150 51914 8156 51916
rect 7833 51912 8156 51914
rect 7833 51856 7838 51912
rect 7894 51856 8156 51912
rect 7833 51854 8156 51856
rect 7833 51851 7899 51854
rect 8150 51852 8156 51854
rect 8220 51914 8226 51916
rect 19241 51914 19307 51917
rect 8220 51912 19307 51914
rect 8220 51856 19246 51912
rect 19302 51856 19307 51912
rect 8220 51854 19307 51856
rect 8220 51852 8226 51854
rect 19241 51851 19307 51854
rect 1946 51712 2262 51713
rect 1946 51648 1952 51712
rect 2016 51648 2032 51712
rect 2096 51648 2112 51712
rect 2176 51648 2192 51712
rect 2256 51648 2262 51712
rect 1946 51647 2262 51648
rect 6946 51712 7262 51713
rect 6946 51648 6952 51712
rect 7016 51648 7032 51712
rect 7096 51648 7112 51712
rect 7176 51648 7192 51712
rect 7256 51648 7262 51712
rect 6946 51647 7262 51648
rect 11946 51712 12262 51713
rect 11946 51648 11952 51712
rect 12016 51648 12032 51712
rect 12096 51648 12112 51712
rect 12176 51648 12192 51712
rect 12256 51648 12262 51712
rect 11946 51647 12262 51648
rect 16946 51712 17262 51713
rect 16946 51648 16952 51712
rect 17016 51648 17032 51712
rect 17096 51648 17112 51712
rect 17176 51648 17192 51712
rect 17256 51648 17262 51712
rect 16946 51647 17262 51648
rect 11421 51370 11487 51373
rect 13118 51370 13124 51372
rect 11421 51368 13124 51370
rect 11421 51312 11426 51368
rect 11482 51312 13124 51368
rect 11421 51310 13124 51312
rect 11421 51307 11487 51310
rect 13118 51308 13124 51310
rect 13188 51308 13194 51372
rect 2606 51168 2922 51169
rect 2606 51104 2612 51168
rect 2676 51104 2692 51168
rect 2756 51104 2772 51168
rect 2836 51104 2852 51168
rect 2916 51104 2922 51168
rect 2606 51103 2922 51104
rect 7606 51168 7922 51169
rect 7606 51104 7612 51168
rect 7676 51104 7692 51168
rect 7756 51104 7772 51168
rect 7836 51104 7852 51168
rect 7916 51104 7922 51168
rect 7606 51103 7922 51104
rect 12606 51168 12922 51169
rect 12606 51104 12612 51168
rect 12676 51104 12692 51168
rect 12756 51104 12772 51168
rect 12836 51104 12852 51168
rect 12916 51104 12922 51168
rect 12606 51103 12922 51104
rect 17606 51168 17922 51169
rect 17606 51104 17612 51168
rect 17676 51104 17692 51168
rect 17756 51104 17772 51168
rect 17836 51104 17852 51168
rect 17916 51104 17922 51168
rect 17606 51103 17922 51104
rect 6913 50826 6979 50829
rect 7414 50826 7420 50828
rect 6913 50824 7420 50826
rect 6913 50768 6918 50824
rect 6974 50768 7420 50824
rect 6913 50766 7420 50768
rect 6913 50763 6979 50766
rect 7414 50764 7420 50766
rect 7484 50826 7490 50828
rect 7557 50826 7623 50829
rect 7484 50824 7623 50826
rect 7484 50768 7562 50824
rect 7618 50768 7623 50824
rect 7484 50766 7623 50768
rect 7484 50764 7490 50766
rect 7557 50763 7623 50766
rect 10685 50692 10751 50693
rect 10685 50690 10732 50692
rect 10640 50688 10732 50690
rect 10640 50632 10690 50688
rect 10640 50630 10732 50632
rect 10685 50628 10732 50630
rect 10796 50628 10802 50692
rect 10685 50627 10751 50628
rect 1946 50624 2262 50625
rect 1946 50560 1952 50624
rect 2016 50560 2032 50624
rect 2096 50560 2112 50624
rect 2176 50560 2192 50624
rect 2256 50560 2262 50624
rect 1946 50559 2262 50560
rect 6946 50624 7262 50625
rect 6946 50560 6952 50624
rect 7016 50560 7032 50624
rect 7096 50560 7112 50624
rect 7176 50560 7192 50624
rect 7256 50560 7262 50624
rect 6946 50559 7262 50560
rect 11946 50624 12262 50625
rect 11946 50560 11952 50624
rect 12016 50560 12032 50624
rect 12096 50560 12112 50624
rect 12176 50560 12192 50624
rect 12256 50560 12262 50624
rect 11946 50559 12262 50560
rect 16946 50624 17262 50625
rect 16946 50560 16952 50624
rect 17016 50560 17032 50624
rect 17096 50560 17112 50624
rect 17176 50560 17192 50624
rect 17256 50560 17262 50624
rect 16946 50559 17262 50560
rect 18229 50418 18295 50421
rect 19200 50418 20000 50448
rect 18229 50416 20000 50418
rect 18229 50360 18234 50416
rect 18290 50360 20000 50416
rect 18229 50358 20000 50360
rect 18229 50355 18295 50358
rect 19200 50328 20000 50358
rect 2606 50080 2922 50081
rect 2606 50016 2612 50080
rect 2676 50016 2692 50080
rect 2756 50016 2772 50080
rect 2836 50016 2852 50080
rect 2916 50016 2922 50080
rect 2606 50015 2922 50016
rect 7606 50080 7922 50081
rect 7606 50016 7612 50080
rect 7676 50016 7692 50080
rect 7756 50016 7772 50080
rect 7836 50016 7852 50080
rect 7916 50016 7922 50080
rect 7606 50015 7922 50016
rect 12606 50080 12922 50081
rect 12606 50016 12612 50080
rect 12676 50016 12692 50080
rect 12756 50016 12772 50080
rect 12836 50016 12852 50080
rect 12916 50016 12922 50080
rect 12606 50015 12922 50016
rect 17606 50080 17922 50081
rect 17606 50016 17612 50080
rect 17676 50016 17692 50080
rect 17756 50016 17772 50080
rect 17836 50016 17852 50080
rect 17916 50016 17922 50080
rect 17606 50015 17922 50016
rect 4429 49740 4495 49741
rect 4429 49736 4476 49740
rect 4540 49738 4546 49740
rect 4429 49680 4434 49736
rect 4429 49676 4476 49680
rect 4540 49678 4586 49738
rect 4540 49676 4546 49678
rect 4429 49675 4495 49676
rect 15878 49540 15884 49604
rect 15948 49602 15954 49604
rect 16297 49602 16363 49605
rect 15948 49600 16363 49602
rect 15948 49544 16302 49600
rect 16358 49544 16363 49600
rect 15948 49542 16363 49544
rect 15948 49540 15954 49542
rect 16297 49539 16363 49542
rect 1946 49536 2262 49537
rect 1946 49472 1952 49536
rect 2016 49472 2032 49536
rect 2096 49472 2112 49536
rect 2176 49472 2192 49536
rect 2256 49472 2262 49536
rect 1946 49471 2262 49472
rect 6946 49536 7262 49537
rect 6946 49472 6952 49536
rect 7016 49472 7032 49536
rect 7096 49472 7112 49536
rect 7176 49472 7192 49536
rect 7256 49472 7262 49536
rect 6946 49471 7262 49472
rect 11946 49536 12262 49537
rect 11946 49472 11952 49536
rect 12016 49472 12032 49536
rect 12096 49472 12112 49536
rect 12176 49472 12192 49536
rect 12256 49472 12262 49536
rect 11946 49471 12262 49472
rect 16946 49536 17262 49537
rect 16946 49472 16952 49536
rect 17016 49472 17032 49536
rect 17096 49472 17112 49536
rect 17176 49472 17192 49536
rect 17256 49472 17262 49536
rect 16946 49471 17262 49472
rect 2606 48992 2922 48993
rect 2606 48928 2612 48992
rect 2676 48928 2692 48992
rect 2756 48928 2772 48992
rect 2836 48928 2852 48992
rect 2916 48928 2922 48992
rect 2606 48927 2922 48928
rect 7606 48992 7922 48993
rect 7606 48928 7612 48992
rect 7676 48928 7692 48992
rect 7756 48928 7772 48992
rect 7836 48928 7852 48992
rect 7916 48928 7922 48992
rect 7606 48927 7922 48928
rect 12606 48992 12922 48993
rect 12606 48928 12612 48992
rect 12676 48928 12692 48992
rect 12756 48928 12772 48992
rect 12836 48928 12852 48992
rect 12916 48928 12922 48992
rect 12606 48927 12922 48928
rect 17606 48992 17922 48993
rect 17606 48928 17612 48992
rect 17676 48928 17692 48992
rect 17756 48928 17772 48992
rect 17836 48928 17852 48992
rect 17916 48928 17922 48992
rect 17606 48927 17922 48928
rect 16757 48650 16823 48653
rect 16757 48648 16866 48650
rect 16757 48592 16762 48648
rect 16818 48592 16866 48648
rect 16757 48587 16866 48592
rect 1946 48448 2262 48449
rect 1946 48384 1952 48448
rect 2016 48384 2032 48448
rect 2096 48384 2112 48448
rect 2176 48384 2192 48448
rect 2256 48384 2262 48448
rect 1946 48383 2262 48384
rect 6946 48448 7262 48449
rect 6946 48384 6952 48448
rect 7016 48384 7032 48448
rect 7096 48384 7112 48448
rect 7176 48384 7192 48448
rect 7256 48384 7262 48448
rect 6946 48383 7262 48384
rect 11946 48448 12262 48449
rect 11946 48384 11952 48448
rect 12016 48384 12032 48448
rect 12096 48384 12112 48448
rect 12176 48384 12192 48448
rect 12256 48384 12262 48448
rect 11946 48383 12262 48384
rect 16021 48380 16087 48381
rect 16021 48376 16068 48380
rect 16132 48378 16138 48380
rect 16021 48320 16026 48376
rect 16021 48316 16068 48320
rect 16132 48318 16178 48378
rect 16132 48316 16138 48318
rect 16021 48315 16087 48316
rect 16806 48245 16866 48587
rect 18229 48514 18295 48517
rect 19200 48514 20000 48544
rect 18229 48512 20000 48514
rect 18229 48456 18234 48512
rect 18290 48456 20000 48512
rect 18229 48454 20000 48456
rect 18229 48451 18295 48454
rect 16946 48448 17262 48449
rect 16946 48384 16952 48448
rect 17016 48384 17032 48448
rect 17096 48384 17112 48448
rect 17176 48384 17192 48448
rect 17256 48384 17262 48448
rect 19200 48424 20000 48454
rect 16946 48383 17262 48384
rect 3693 48242 3759 48245
rect 4654 48242 4660 48244
rect 3693 48240 4660 48242
rect 3693 48184 3698 48240
rect 3754 48184 4660 48240
rect 3693 48182 4660 48184
rect 3693 48179 3759 48182
rect 4654 48180 4660 48182
rect 4724 48180 4730 48244
rect 16757 48240 16866 48245
rect 16757 48184 16762 48240
rect 16818 48184 16866 48240
rect 16757 48182 16866 48184
rect 16757 48179 16823 48182
rect 2606 47904 2922 47905
rect 2606 47840 2612 47904
rect 2676 47840 2692 47904
rect 2756 47840 2772 47904
rect 2836 47840 2852 47904
rect 2916 47840 2922 47904
rect 2606 47839 2922 47840
rect 7606 47904 7922 47905
rect 7606 47840 7612 47904
rect 7676 47840 7692 47904
rect 7756 47840 7772 47904
rect 7836 47840 7852 47904
rect 7916 47840 7922 47904
rect 7606 47839 7922 47840
rect 12606 47904 12922 47905
rect 12606 47840 12612 47904
rect 12676 47840 12692 47904
rect 12756 47840 12772 47904
rect 12836 47840 12852 47904
rect 12916 47840 12922 47904
rect 12606 47839 12922 47840
rect 17606 47904 17922 47905
rect 17606 47840 17612 47904
rect 17676 47840 17692 47904
rect 17756 47840 17772 47904
rect 17836 47840 17852 47904
rect 17916 47840 17922 47904
rect 17606 47839 17922 47840
rect 1946 47360 2262 47361
rect 1946 47296 1952 47360
rect 2016 47296 2032 47360
rect 2096 47296 2112 47360
rect 2176 47296 2192 47360
rect 2256 47296 2262 47360
rect 1946 47295 2262 47296
rect 6946 47360 7262 47361
rect 6946 47296 6952 47360
rect 7016 47296 7032 47360
rect 7096 47296 7112 47360
rect 7176 47296 7192 47360
rect 7256 47296 7262 47360
rect 6946 47295 7262 47296
rect 11946 47360 12262 47361
rect 11946 47296 11952 47360
rect 12016 47296 12032 47360
rect 12096 47296 12112 47360
rect 12176 47296 12192 47360
rect 12256 47296 12262 47360
rect 11946 47295 12262 47296
rect 16946 47360 17262 47361
rect 16946 47296 16952 47360
rect 17016 47296 17032 47360
rect 17096 47296 17112 47360
rect 17176 47296 17192 47360
rect 17256 47296 17262 47360
rect 16946 47295 17262 47296
rect 3049 47290 3115 47293
rect 3182 47290 3188 47292
rect 3049 47288 3188 47290
rect 3049 47232 3054 47288
rect 3110 47232 3188 47288
rect 3049 47230 3188 47232
rect 3049 47227 3115 47230
rect 3182 47228 3188 47230
rect 3252 47228 3258 47292
rect 2606 46816 2922 46817
rect 2606 46752 2612 46816
rect 2676 46752 2692 46816
rect 2756 46752 2772 46816
rect 2836 46752 2852 46816
rect 2916 46752 2922 46816
rect 2606 46751 2922 46752
rect 7606 46816 7922 46817
rect 7606 46752 7612 46816
rect 7676 46752 7692 46816
rect 7756 46752 7772 46816
rect 7836 46752 7852 46816
rect 7916 46752 7922 46816
rect 7606 46751 7922 46752
rect 12606 46816 12922 46817
rect 12606 46752 12612 46816
rect 12676 46752 12692 46816
rect 12756 46752 12772 46816
rect 12836 46752 12852 46816
rect 12916 46752 12922 46816
rect 12606 46751 12922 46752
rect 17606 46816 17922 46817
rect 17606 46752 17612 46816
rect 17676 46752 17692 46816
rect 17756 46752 17772 46816
rect 17836 46752 17852 46816
rect 17916 46752 17922 46816
rect 17606 46751 17922 46752
rect 18229 46610 18295 46613
rect 19200 46610 20000 46640
rect 18229 46608 20000 46610
rect 18229 46552 18234 46608
rect 18290 46552 20000 46608
rect 18229 46550 20000 46552
rect 18229 46547 18295 46550
rect 19200 46520 20000 46550
rect 1946 46272 2262 46273
rect 1946 46208 1952 46272
rect 2016 46208 2032 46272
rect 2096 46208 2112 46272
rect 2176 46208 2192 46272
rect 2256 46208 2262 46272
rect 1946 46207 2262 46208
rect 6946 46272 7262 46273
rect 6946 46208 6952 46272
rect 7016 46208 7032 46272
rect 7096 46208 7112 46272
rect 7176 46208 7192 46272
rect 7256 46208 7262 46272
rect 6946 46207 7262 46208
rect 11946 46272 12262 46273
rect 11946 46208 11952 46272
rect 12016 46208 12032 46272
rect 12096 46208 12112 46272
rect 12176 46208 12192 46272
rect 12256 46208 12262 46272
rect 11946 46207 12262 46208
rect 16946 46272 17262 46273
rect 16946 46208 16952 46272
rect 17016 46208 17032 46272
rect 17096 46208 17112 46272
rect 17176 46208 17192 46272
rect 17256 46208 17262 46272
rect 16946 46207 17262 46208
rect 2606 45728 2922 45729
rect 2606 45664 2612 45728
rect 2676 45664 2692 45728
rect 2756 45664 2772 45728
rect 2836 45664 2852 45728
rect 2916 45664 2922 45728
rect 2606 45663 2922 45664
rect 7606 45728 7922 45729
rect 7606 45664 7612 45728
rect 7676 45664 7692 45728
rect 7756 45664 7772 45728
rect 7836 45664 7852 45728
rect 7916 45664 7922 45728
rect 7606 45663 7922 45664
rect 12606 45728 12922 45729
rect 12606 45664 12612 45728
rect 12676 45664 12692 45728
rect 12756 45664 12772 45728
rect 12836 45664 12852 45728
rect 12916 45664 12922 45728
rect 12606 45663 12922 45664
rect 17606 45728 17922 45729
rect 17606 45664 17612 45728
rect 17676 45664 17692 45728
rect 17756 45664 17772 45728
rect 17836 45664 17852 45728
rect 17916 45664 17922 45728
rect 17606 45663 17922 45664
rect 1946 45184 2262 45185
rect 1946 45120 1952 45184
rect 2016 45120 2032 45184
rect 2096 45120 2112 45184
rect 2176 45120 2192 45184
rect 2256 45120 2262 45184
rect 1946 45119 2262 45120
rect 6946 45184 7262 45185
rect 6946 45120 6952 45184
rect 7016 45120 7032 45184
rect 7096 45120 7112 45184
rect 7176 45120 7192 45184
rect 7256 45120 7262 45184
rect 6946 45119 7262 45120
rect 11946 45184 12262 45185
rect 11946 45120 11952 45184
rect 12016 45120 12032 45184
rect 12096 45120 12112 45184
rect 12176 45120 12192 45184
rect 12256 45120 12262 45184
rect 11946 45119 12262 45120
rect 16946 45184 17262 45185
rect 16946 45120 16952 45184
rect 17016 45120 17032 45184
rect 17096 45120 17112 45184
rect 17176 45120 17192 45184
rect 17256 45120 17262 45184
rect 16946 45119 17262 45120
rect 18229 44706 18295 44709
rect 19200 44706 20000 44736
rect 18229 44704 20000 44706
rect 18229 44648 18234 44704
rect 18290 44648 20000 44704
rect 18229 44646 20000 44648
rect 18229 44643 18295 44646
rect 2606 44640 2922 44641
rect 2606 44576 2612 44640
rect 2676 44576 2692 44640
rect 2756 44576 2772 44640
rect 2836 44576 2852 44640
rect 2916 44576 2922 44640
rect 2606 44575 2922 44576
rect 7606 44640 7922 44641
rect 7606 44576 7612 44640
rect 7676 44576 7692 44640
rect 7756 44576 7772 44640
rect 7836 44576 7852 44640
rect 7916 44576 7922 44640
rect 7606 44575 7922 44576
rect 12606 44640 12922 44641
rect 12606 44576 12612 44640
rect 12676 44576 12692 44640
rect 12756 44576 12772 44640
rect 12836 44576 12852 44640
rect 12916 44576 12922 44640
rect 12606 44575 12922 44576
rect 17606 44640 17922 44641
rect 17606 44576 17612 44640
rect 17676 44576 17692 44640
rect 17756 44576 17772 44640
rect 17836 44576 17852 44640
rect 17916 44576 17922 44640
rect 19200 44616 20000 44646
rect 17606 44575 17922 44576
rect 1946 44096 2262 44097
rect 1946 44032 1952 44096
rect 2016 44032 2032 44096
rect 2096 44032 2112 44096
rect 2176 44032 2192 44096
rect 2256 44032 2262 44096
rect 1946 44031 2262 44032
rect 6946 44096 7262 44097
rect 6946 44032 6952 44096
rect 7016 44032 7032 44096
rect 7096 44032 7112 44096
rect 7176 44032 7192 44096
rect 7256 44032 7262 44096
rect 6946 44031 7262 44032
rect 11946 44096 12262 44097
rect 11946 44032 11952 44096
rect 12016 44032 12032 44096
rect 12096 44032 12112 44096
rect 12176 44032 12192 44096
rect 12256 44032 12262 44096
rect 11946 44031 12262 44032
rect 16946 44096 17262 44097
rect 16946 44032 16952 44096
rect 17016 44032 17032 44096
rect 17096 44032 17112 44096
rect 17176 44032 17192 44096
rect 17256 44032 17262 44096
rect 16946 44031 17262 44032
rect 2606 43552 2922 43553
rect 2606 43488 2612 43552
rect 2676 43488 2692 43552
rect 2756 43488 2772 43552
rect 2836 43488 2852 43552
rect 2916 43488 2922 43552
rect 2606 43487 2922 43488
rect 7606 43552 7922 43553
rect 7606 43488 7612 43552
rect 7676 43488 7692 43552
rect 7756 43488 7772 43552
rect 7836 43488 7852 43552
rect 7916 43488 7922 43552
rect 7606 43487 7922 43488
rect 12606 43552 12922 43553
rect 12606 43488 12612 43552
rect 12676 43488 12692 43552
rect 12756 43488 12772 43552
rect 12836 43488 12852 43552
rect 12916 43488 12922 43552
rect 12606 43487 12922 43488
rect 17606 43552 17922 43553
rect 17606 43488 17612 43552
rect 17676 43488 17692 43552
rect 17756 43488 17772 43552
rect 17836 43488 17852 43552
rect 17916 43488 17922 43552
rect 17606 43487 17922 43488
rect 7414 43284 7420 43348
rect 7484 43346 7490 43348
rect 7557 43346 7623 43349
rect 7484 43344 7623 43346
rect 7484 43288 7562 43344
rect 7618 43288 7623 43344
rect 7484 43286 7623 43288
rect 7484 43284 7490 43286
rect 7557 43283 7623 43286
rect 1946 43008 2262 43009
rect 1946 42944 1952 43008
rect 2016 42944 2032 43008
rect 2096 42944 2112 43008
rect 2176 42944 2192 43008
rect 2256 42944 2262 43008
rect 1946 42943 2262 42944
rect 6946 43008 7262 43009
rect 6946 42944 6952 43008
rect 7016 42944 7032 43008
rect 7096 42944 7112 43008
rect 7176 42944 7192 43008
rect 7256 42944 7262 43008
rect 6946 42943 7262 42944
rect 11946 43008 12262 43009
rect 11946 42944 11952 43008
rect 12016 42944 12032 43008
rect 12096 42944 12112 43008
rect 12176 42944 12192 43008
rect 12256 42944 12262 43008
rect 11946 42943 12262 42944
rect 16946 43008 17262 43009
rect 16946 42944 16952 43008
rect 17016 42944 17032 43008
rect 17096 42944 17112 43008
rect 17176 42944 17192 43008
rect 17256 42944 17262 43008
rect 16946 42943 17262 42944
rect 6494 42876 6500 42940
rect 6564 42938 6570 42940
rect 6729 42938 6795 42941
rect 6564 42936 6795 42938
rect 6564 42880 6734 42936
rect 6790 42880 6795 42936
rect 6564 42878 6795 42880
rect 6564 42876 6570 42878
rect 6729 42875 6795 42878
rect 11053 42802 11119 42805
rect 11278 42802 11284 42804
rect 11053 42800 11284 42802
rect 11053 42744 11058 42800
rect 11114 42744 11284 42800
rect 11053 42742 11284 42744
rect 11053 42739 11119 42742
rect 11278 42740 11284 42742
rect 11348 42740 11354 42804
rect 11462 42740 11468 42804
rect 11532 42802 11538 42804
rect 11605 42802 11671 42805
rect 11532 42800 11671 42802
rect 11532 42744 11610 42800
rect 11666 42744 11671 42800
rect 11532 42742 11671 42744
rect 11532 42740 11538 42742
rect 11605 42739 11671 42742
rect 18229 42802 18295 42805
rect 19200 42802 20000 42832
rect 18229 42800 20000 42802
rect 18229 42744 18234 42800
rect 18290 42744 20000 42800
rect 18229 42742 20000 42744
rect 18229 42739 18295 42742
rect 19200 42712 20000 42742
rect 10409 42666 10475 42669
rect 18229 42666 18295 42669
rect 10409 42664 18295 42666
rect 10409 42608 10414 42664
rect 10470 42608 18234 42664
rect 18290 42608 18295 42664
rect 10409 42606 18295 42608
rect 10409 42603 10475 42606
rect 18229 42603 18295 42606
rect 2606 42464 2922 42465
rect 2606 42400 2612 42464
rect 2676 42400 2692 42464
rect 2756 42400 2772 42464
rect 2836 42400 2852 42464
rect 2916 42400 2922 42464
rect 2606 42399 2922 42400
rect 7606 42464 7922 42465
rect 7606 42400 7612 42464
rect 7676 42400 7692 42464
rect 7756 42400 7772 42464
rect 7836 42400 7852 42464
rect 7916 42400 7922 42464
rect 7606 42399 7922 42400
rect 12606 42464 12922 42465
rect 12606 42400 12612 42464
rect 12676 42400 12692 42464
rect 12756 42400 12772 42464
rect 12836 42400 12852 42464
rect 12916 42400 12922 42464
rect 12606 42399 12922 42400
rect 17606 42464 17922 42465
rect 17606 42400 17612 42464
rect 17676 42400 17692 42464
rect 17756 42400 17772 42464
rect 17836 42400 17852 42464
rect 17916 42400 17922 42464
rect 17606 42399 17922 42400
rect 18229 41986 18295 41989
rect 18597 41986 18663 41989
rect 18229 41984 18663 41986
rect 18229 41928 18234 41984
rect 18290 41928 18602 41984
rect 18658 41928 18663 41984
rect 18229 41926 18663 41928
rect 18229 41923 18295 41926
rect 18597 41923 18663 41926
rect 1946 41920 2262 41921
rect 1946 41856 1952 41920
rect 2016 41856 2032 41920
rect 2096 41856 2112 41920
rect 2176 41856 2192 41920
rect 2256 41856 2262 41920
rect 1946 41855 2262 41856
rect 6946 41920 7262 41921
rect 6946 41856 6952 41920
rect 7016 41856 7032 41920
rect 7096 41856 7112 41920
rect 7176 41856 7192 41920
rect 7256 41856 7262 41920
rect 6946 41855 7262 41856
rect 11946 41920 12262 41921
rect 11946 41856 11952 41920
rect 12016 41856 12032 41920
rect 12096 41856 12112 41920
rect 12176 41856 12192 41920
rect 12256 41856 12262 41920
rect 11946 41855 12262 41856
rect 16946 41920 17262 41921
rect 16946 41856 16952 41920
rect 17016 41856 17032 41920
rect 17096 41856 17112 41920
rect 17176 41856 17192 41920
rect 17256 41856 17262 41920
rect 16946 41855 17262 41856
rect 2606 41376 2922 41377
rect 2606 41312 2612 41376
rect 2676 41312 2692 41376
rect 2756 41312 2772 41376
rect 2836 41312 2852 41376
rect 2916 41312 2922 41376
rect 2606 41311 2922 41312
rect 7606 41376 7922 41377
rect 7606 41312 7612 41376
rect 7676 41312 7692 41376
rect 7756 41312 7772 41376
rect 7836 41312 7852 41376
rect 7916 41312 7922 41376
rect 7606 41311 7922 41312
rect 12606 41376 12922 41377
rect 12606 41312 12612 41376
rect 12676 41312 12692 41376
rect 12756 41312 12772 41376
rect 12836 41312 12852 41376
rect 12916 41312 12922 41376
rect 12606 41311 12922 41312
rect 17606 41376 17922 41377
rect 17606 41312 17612 41376
rect 17676 41312 17692 41376
rect 17756 41312 17772 41376
rect 17836 41312 17852 41376
rect 17916 41312 17922 41376
rect 17606 41311 17922 41312
rect 1761 40898 1827 40901
rect 1718 40896 1827 40898
rect 1718 40840 1766 40896
rect 1822 40840 1827 40896
rect 1718 40835 1827 40840
rect 18229 40898 18295 40901
rect 19200 40898 20000 40928
rect 18229 40896 20000 40898
rect 18229 40840 18234 40896
rect 18290 40840 20000 40896
rect 18229 40838 20000 40840
rect 18229 40835 18295 40838
rect 1577 40626 1643 40629
rect 1718 40626 1778 40835
rect 1946 40832 2262 40833
rect 1946 40768 1952 40832
rect 2016 40768 2032 40832
rect 2096 40768 2112 40832
rect 2176 40768 2192 40832
rect 2256 40768 2262 40832
rect 1946 40767 2262 40768
rect 6946 40832 7262 40833
rect 6946 40768 6952 40832
rect 7016 40768 7032 40832
rect 7096 40768 7112 40832
rect 7176 40768 7192 40832
rect 7256 40768 7262 40832
rect 6946 40767 7262 40768
rect 11946 40832 12262 40833
rect 11946 40768 11952 40832
rect 12016 40768 12032 40832
rect 12096 40768 12112 40832
rect 12176 40768 12192 40832
rect 12256 40768 12262 40832
rect 11946 40767 12262 40768
rect 16946 40832 17262 40833
rect 16946 40768 16952 40832
rect 17016 40768 17032 40832
rect 17096 40768 17112 40832
rect 17176 40768 17192 40832
rect 17256 40768 17262 40832
rect 19200 40808 20000 40838
rect 16946 40767 17262 40768
rect 1577 40624 1778 40626
rect 1577 40568 1582 40624
rect 1638 40568 1778 40624
rect 1577 40566 1778 40568
rect 1577 40563 1643 40566
rect 9070 40564 9076 40628
rect 9140 40626 9146 40628
rect 16941 40626 17007 40629
rect 9140 40624 17007 40626
rect 9140 40568 16946 40624
rect 17002 40568 17007 40624
rect 9140 40566 17007 40568
rect 9140 40564 9146 40566
rect 16941 40563 17007 40566
rect 9254 40428 9260 40492
rect 9324 40490 9330 40492
rect 9489 40490 9555 40493
rect 9324 40488 9555 40490
rect 9324 40432 9494 40488
rect 9550 40432 9555 40488
rect 9324 40430 9555 40432
rect 9324 40428 9330 40430
rect 9489 40427 9555 40430
rect 2606 40288 2922 40289
rect 2606 40224 2612 40288
rect 2676 40224 2692 40288
rect 2756 40224 2772 40288
rect 2836 40224 2852 40288
rect 2916 40224 2922 40288
rect 2606 40223 2922 40224
rect 7606 40288 7922 40289
rect 7606 40224 7612 40288
rect 7676 40224 7692 40288
rect 7756 40224 7772 40288
rect 7836 40224 7852 40288
rect 7916 40224 7922 40288
rect 7606 40223 7922 40224
rect 12606 40288 12922 40289
rect 12606 40224 12612 40288
rect 12676 40224 12692 40288
rect 12756 40224 12772 40288
rect 12836 40224 12852 40288
rect 12916 40224 12922 40288
rect 12606 40223 12922 40224
rect 17606 40288 17922 40289
rect 17606 40224 17612 40288
rect 17676 40224 17692 40288
rect 17756 40224 17772 40288
rect 17836 40224 17852 40288
rect 17916 40224 17922 40288
rect 17606 40223 17922 40224
rect 1946 39744 2262 39745
rect 1946 39680 1952 39744
rect 2016 39680 2032 39744
rect 2096 39680 2112 39744
rect 2176 39680 2192 39744
rect 2256 39680 2262 39744
rect 1946 39679 2262 39680
rect 6946 39744 7262 39745
rect 6946 39680 6952 39744
rect 7016 39680 7032 39744
rect 7096 39680 7112 39744
rect 7176 39680 7192 39744
rect 7256 39680 7262 39744
rect 6946 39679 7262 39680
rect 11946 39744 12262 39745
rect 11946 39680 11952 39744
rect 12016 39680 12032 39744
rect 12096 39680 12112 39744
rect 12176 39680 12192 39744
rect 12256 39680 12262 39744
rect 11946 39679 12262 39680
rect 16946 39744 17262 39745
rect 16946 39680 16952 39744
rect 17016 39680 17032 39744
rect 17096 39680 17112 39744
rect 17176 39680 17192 39744
rect 17256 39680 17262 39744
rect 16946 39679 17262 39680
rect 2606 39200 2922 39201
rect 2606 39136 2612 39200
rect 2676 39136 2692 39200
rect 2756 39136 2772 39200
rect 2836 39136 2852 39200
rect 2916 39136 2922 39200
rect 2606 39135 2922 39136
rect 7606 39200 7922 39201
rect 7606 39136 7612 39200
rect 7676 39136 7692 39200
rect 7756 39136 7772 39200
rect 7836 39136 7852 39200
rect 7916 39136 7922 39200
rect 7606 39135 7922 39136
rect 12606 39200 12922 39201
rect 12606 39136 12612 39200
rect 12676 39136 12692 39200
rect 12756 39136 12772 39200
rect 12836 39136 12852 39200
rect 12916 39136 12922 39200
rect 12606 39135 12922 39136
rect 17606 39200 17922 39201
rect 17606 39136 17612 39200
rect 17676 39136 17692 39200
rect 17756 39136 17772 39200
rect 17836 39136 17852 39200
rect 17916 39136 17922 39200
rect 17606 39135 17922 39136
rect 18229 38994 18295 38997
rect 19200 38994 20000 39024
rect 18229 38992 20000 38994
rect 18229 38936 18234 38992
rect 18290 38936 20000 38992
rect 18229 38934 20000 38936
rect 18229 38931 18295 38934
rect 19200 38904 20000 38934
rect 1946 38656 2262 38657
rect 1946 38592 1952 38656
rect 2016 38592 2032 38656
rect 2096 38592 2112 38656
rect 2176 38592 2192 38656
rect 2256 38592 2262 38656
rect 1946 38591 2262 38592
rect 6946 38656 7262 38657
rect 6946 38592 6952 38656
rect 7016 38592 7032 38656
rect 7096 38592 7112 38656
rect 7176 38592 7192 38656
rect 7256 38592 7262 38656
rect 6946 38591 7262 38592
rect 11946 38656 12262 38657
rect 11946 38592 11952 38656
rect 12016 38592 12032 38656
rect 12096 38592 12112 38656
rect 12176 38592 12192 38656
rect 12256 38592 12262 38656
rect 11946 38591 12262 38592
rect 16946 38656 17262 38657
rect 16946 38592 16952 38656
rect 17016 38592 17032 38656
rect 17096 38592 17112 38656
rect 17176 38592 17192 38656
rect 17256 38592 17262 38656
rect 16946 38591 17262 38592
rect 2606 38112 2922 38113
rect 2606 38048 2612 38112
rect 2676 38048 2692 38112
rect 2756 38048 2772 38112
rect 2836 38048 2852 38112
rect 2916 38048 2922 38112
rect 2606 38047 2922 38048
rect 7606 38112 7922 38113
rect 7606 38048 7612 38112
rect 7676 38048 7692 38112
rect 7756 38048 7772 38112
rect 7836 38048 7852 38112
rect 7916 38048 7922 38112
rect 7606 38047 7922 38048
rect 12606 38112 12922 38113
rect 12606 38048 12612 38112
rect 12676 38048 12692 38112
rect 12756 38048 12772 38112
rect 12836 38048 12852 38112
rect 12916 38048 12922 38112
rect 12606 38047 12922 38048
rect 17606 38112 17922 38113
rect 17606 38048 17612 38112
rect 17676 38048 17692 38112
rect 17756 38048 17772 38112
rect 17836 38048 17852 38112
rect 17916 38048 17922 38112
rect 17606 38047 17922 38048
rect 1946 37568 2262 37569
rect 1946 37504 1952 37568
rect 2016 37504 2032 37568
rect 2096 37504 2112 37568
rect 2176 37504 2192 37568
rect 2256 37504 2262 37568
rect 1946 37503 2262 37504
rect 6946 37568 7262 37569
rect 6946 37504 6952 37568
rect 7016 37504 7032 37568
rect 7096 37504 7112 37568
rect 7176 37504 7192 37568
rect 7256 37504 7262 37568
rect 6946 37503 7262 37504
rect 11946 37568 12262 37569
rect 11946 37504 11952 37568
rect 12016 37504 12032 37568
rect 12096 37504 12112 37568
rect 12176 37504 12192 37568
rect 12256 37504 12262 37568
rect 11946 37503 12262 37504
rect 16946 37568 17262 37569
rect 16946 37504 16952 37568
rect 17016 37504 17032 37568
rect 17096 37504 17112 37568
rect 17176 37504 17192 37568
rect 17256 37504 17262 37568
rect 16946 37503 17262 37504
rect 15142 37300 15148 37364
rect 15212 37362 15218 37364
rect 16297 37362 16363 37365
rect 15212 37360 16363 37362
rect 15212 37304 16302 37360
rect 16358 37304 16363 37360
rect 15212 37302 16363 37304
rect 15212 37300 15218 37302
rect 16297 37299 16363 37302
rect 18229 37090 18295 37093
rect 19200 37090 20000 37120
rect 18229 37088 20000 37090
rect 18229 37032 18234 37088
rect 18290 37032 20000 37088
rect 18229 37030 20000 37032
rect 18229 37027 18295 37030
rect 2606 37024 2922 37025
rect 2606 36960 2612 37024
rect 2676 36960 2692 37024
rect 2756 36960 2772 37024
rect 2836 36960 2852 37024
rect 2916 36960 2922 37024
rect 2606 36959 2922 36960
rect 7606 37024 7922 37025
rect 7606 36960 7612 37024
rect 7676 36960 7692 37024
rect 7756 36960 7772 37024
rect 7836 36960 7852 37024
rect 7916 36960 7922 37024
rect 7606 36959 7922 36960
rect 12606 37024 12922 37025
rect 12606 36960 12612 37024
rect 12676 36960 12692 37024
rect 12756 36960 12772 37024
rect 12836 36960 12852 37024
rect 12916 36960 12922 37024
rect 12606 36959 12922 36960
rect 17606 37024 17922 37025
rect 17606 36960 17612 37024
rect 17676 36960 17692 37024
rect 17756 36960 17772 37024
rect 17836 36960 17852 37024
rect 17916 36960 17922 37024
rect 19200 37000 20000 37030
rect 17606 36959 17922 36960
rect 1946 36480 2262 36481
rect 1946 36416 1952 36480
rect 2016 36416 2032 36480
rect 2096 36416 2112 36480
rect 2176 36416 2192 36480
rect 2256 36416 2262 36480
rect 1946 36415 2262 36416
rect 6946 36480 7262 36481
rect 6946 36416 6952 36480
rect 7016 36416 7032 36480
rect 7096 36416 7112 36480
rect 7176 36416 7192 36480
rect 7256 36416 7262 36480
rect 6946 36415 7262 36416
rect 11946 36480 12262 36481
rect 11946 36416 11952 36480
rect 12016 36416 12032 36480
rect 12096 36416 12112 36480
rect 12176 36416 12192 36480
rect 12256 36416 12262 36480
rect 11946 36415 12262 36416
rect 16946 36480 17262 36481
rect 16946 36416 16952 36480
rect 17016 36416 17032 36480
rect 17096 36416 17112 36480
rect 17176 36416 17192 36480
rect 17256 36416 17262 36480
rect 16946 36415 17262 36416
rect 9806 36348 9812 36412
rect 9876 36410 9882 36412
rect 10041 36410 10107 36413
rect 9876 36408 10107 36410
rect 9876 36352 10046 36408
rect 10102 36352 10107 36408
rect 9876 36350 10107 36352
rect 9876 36348 9882 36350
rect 10041 36347 10107 36350
rect 2606 35936 2922 35937
rect 2606 35872 2612 35936
rect 2676 35872 2692 35936
rect 2756 35872 2772 35936
rect 2836 35872 2852 35936
rect 2916 35872 2922 35936
rect 2606 35871 2922 35872
rect 7606 35936 7922 35937
rect 7606 35872 7612 35936
rect 7676 35872 7692 35936
rect 7756 35872 7772 35936
rect 7836 35872 7852 35936
rect 7916 35872 7922 35936
rect 7606 35871 7922 35872
rect 12606 35936 12922 35937
rect 12606 35872 12612 35936
rect 12676 35872 12692 35936
rect 12756 35872 12772 35936
rect 12836 35872 12852 35936
rect 12916 35872 12922 35936
rect 12606 35871 12922 35872
rect 17606 35936 17922 35937
rect 17606 35872 17612 35936
rect 17676 35872 17692 35936
rect 17756 35872 17772 35936
rect 17836 35872 17852 35936
rect 17916 35872 17922 35936
rect 17606 35871 17922 35872
rect 10910 35668 10916 35732
rect 10980 35730 10986 35732
rect 14089 35730 14155 35733
rect 10980 35728 14155 35730
rect 10980 35672 14094 35728
rect 14150 35672 14155 35728
rect 10980 35670 14155 35672
rect 10980 35668 10986 35670
rect 14089 35667 14155 35670
rect 3366 35532 3372 35596
rect 3436 35594 3442 35596
rect 12433 35594 12499 35597
rect 3436 35592 12499 35594
rect 3436 35536 12438 35592
rect 12494 35536 12499 35592
rect 3436 35534 12499 35536
rect 3436 35532 3442 35534
rect 12433 35531 12499 35534
rect 1946 35392 2262 35393
rect 1946 35328 1952 35392
rect 2016 35328 2032 35392
rect 2096 35328 2112 35392
rect 2176 35328 2192 35392
rect 2256 35328 2262 35392
rect 1946 35327 2262 35328
rect 6946 35392 7262 35393
rect 6946 35328 6952 35392
rect 7016 35328 7032 35392
rect 7096 35328 7112 35392
rect 7176 35328 7192 35392
rect 7256 35328 7262 35392
rect 6946 35327 7262 35328
rect 11946 35392 12262 35393
rect 11946 35328 11952 35392
rect 12016 35328 12032 35392
rect 12096 35328 12112 35392
rect 12176 35328 12192 35392
rect 12256 35328 12262 35392
rect 11946 35327 12262 35328
rect 16946 35392 17262 35393
rect 16946 35328 16952 35392
rect 17016 35328 17032 35392
rect 17096 35328 17112 35392
rect 17176 35328 17192 35392
rect 17256 35328 17262 35392
rect 16946 35327 17262 35328
rect 18229 35186 18295 35189
rect 19200 35186 20000 35216
rect 18229 35184 20000 35186
rect 18229 35128 18234 35184
rect 18290 35128 20000 35184
rect 18229 35126 20000 35128
rect 18229 35123 18295 35126
rect 19200 35096 20000 35126
rect 2606 34848 2922 34849
rect 2606 34784 2612 34848
rect 2676 34784 2692 34848
rect 2756 34784 2772 34848
rect 2836 34784 2852 34848
rect 2916 34784 2922 34848
rect 2606 34783 2922 34784
rect 7606 34848 7922 34849
rect 7606 34784 7612 34848
rect 7676 34784 7692 34848
rect 7756 34784 7772 34848
rect 7836 34784 7852 34848
rect 7916 34784 7922 34848
rect 7606 34783 7922 34784
rect 12606 34848 12922 34849
rect 12606 34784 12612 34848
rect 12676 34784 12692 34848
rect 12756 34784 12772 34848
rect 12836 34784 12852 34848
rect 12916 34784 12922 34848
rect 12606 34783 12922 34784
rect 17606 34848 17922 34849
rect 17606 34784 17612 34848
rect 17676 34784 17692 34848
rect 17756 34784 17772 34848
rect 17836 34784 17852 34848
rect 17916 34784 17922 34848
rect 17606 34783 17922 34784
rect 1946 34304 2262 34305
rect 1946 34240 1952 34304
rect 2016 34240 2032 34304
rect 2096 34240 2112 34304
rect 2176 34240 2192 34304
rect 2256 34240 2262 34304
rect 1946 34239 2262 34240
rect 6946 34304 7262 34305
rect 6946 34240 6952 34304
rect 7016 34240 7032 34304
rect 7096 34240 7112 34304
rect 7176 34240 7192 34304
rect 7256 34240 7262 34304
rect 6946 34239 7262 34240
rect 11946 34304 12262 34305
rect 11946 34240 11952 34304
rect 12016 34240 12032 34304
rect 12096 34240 12112 34304
rect 12176 34240 12192 34304
rect 12256 34240 12262 34304
rect 11946 34239 12262 34240
rect 16946 34304 17262 34305
rect 16946 34240 16952 34304
rect 17016 34240 17032 34304
rect 17096 34240 17112 34304
rect 17176 34240 17192 34304
rect 17256 34240 17262 34304
rect 16946 34239 17262 34240
rect 16757 34234 16823 34237
rect 16757 34232 16866 34234
rect 16757 34176 16762 34232
rect 16818 34176 16866 34232
rect 16757 34171 16866 34176
rect 16806 33962 16866 34171
rect 17401 33962 17467 33965
rect 16806 33960 17467 33962
rect 16806 33904 17406 33960
rect 17462 33904 17467 33960
rect 16806 33902 17467 33904
rect 17401 33899 17467 33902
rect 2606 33760 2922 33761
rect 2606 33696 2612 33760
rect 2676 33696 2692 33760
rect 2756 33696 2772 33760
rect 2836 33696 2852 33760
rect 2916 33696 2922 33760
rect 2606 33695 2922 33696
rect 7606 33760 7922 33761
rect 7606 33696 7612 33760
rect 7676 33696 7692 33760
rect 7756 33696 7772 33760
rect 7836 33696 7852 33760
rect 7916 33696 7922 33760
rect 7606 33695 7922 33696
rect 12606 33760 12922 33761
rect 12606 33696 12612 33760
rect 12676 33696 12692 33760
rect 12756 33696 12772 33760
rect 12836 33696 12852 33760
rect 12916 33696 12922 33760
rect 12606 33695 12922 33696
rect 17606 33760 17922 33761
rect 17606 33696 17612 33760
rect 17676 33696 17692 33760
rect 17756 33696 17772 33760
rect 17836 33696 17852 33760
rect 17916 33696 17922 33760
rect 17606 33695 17922 33696
rect 18229 33282 18295 33285
rect 19200 33282 20000 33312
rect 18229 33280 20000 33282
rect 18229 33224 18234 33280
rect 18290 33224 20000 33280
rect 18229 33222 20000 33224
rect 18229 33219 18295 33222
rect 1946 33216 2262 33217
rect 1946 33152 1952 33216
rect 2016 33152 2032 33216
rect 2096 33152 2112 33216
rect 2176 33152 2192 33216
rect 2256 33152 2262 33216
rect 1946 33151 2262 33152
rect 6946 33216 7262 33217
rect 6946 33152 6952 33216
rect 7016 33152 7032 33216
rect 7096 33152 7112 33216
rect 7176 33152 7192 33216
rect 7256 33152 7262 33216
rect 6946 33151 7262 33152
rect 11946 33216 12262 33217
rect 11946 33152 11952 33216
rect 12016 33152 12032 33216
rect 12096 33152 12112 33216
rect 12176 33152 12192 33216
rect 12256 33152 12262 33216
rect 11946 33151 12262 33152
rect 16946 33216 17262 33217
rect 16946 33152 16952 33216
rect 17016 33152 17032 33216
rect 17096 33152 17112 33216
rect 17176 33152 17192 33216
rect 17256 33152 17262 33216
rect 19200 33192 20000 33222
rect 16946 33151 17262 33152
rect 8702 33084 8708 33148
rect 8772 33146 8778 33148
rect 8937 33146 9003 33149
rect 8772 33144 9003 33146
rect 8772 33088 8942 33144
rect 8998 33088 9003 33144
rect 8772 33086 9003 33088
rect 8772 33084 8778 33086
rect 8937 33083 9003 33086
rect 8477 33010 8543 33013
rect 9070 33010 9076 33012
rect 8477 33008 9076 33010
rect 8477 32952 8482 33008
rect 8538 32952 9076 33008
rect 8477 32950 9076 32952
rect 8477 32947 8543 32950
rect 9070 32948 9076 32950
rect 9140 32948 9146 33012
rect 2606 32672 2922 32673
rect 2606 32608 2612 32672
rect 2676 32608 2692 32672
rect 2756 32608 2772 32672
rect 2836 32608 2852 32672
rect 2916 32608 2922 32672
rect 2606 32607 2922 32608
rect 7606 32672 7922 32673
rect 7606 32608 7612 32672
rect 7676 32608 7692 32672
rect 7756 32608 7772 32672
rect 7836 32608 7852 32672
rect 7916 32608 7922 32672
rect 7606 32607 7922 32608
rect 12606 32672 12922 32673
rect 12606 32608 12612 32672
rect 12676 32608 12692 32672
rect 12756 32608 12772 32672
rect 12836 32608 12852 32672
rect 12916 32608 12922 32672
rect 12606 32607 12922 32608
rect 17606 32672 17922 32673
rect 17606 32608 17612 32672
rect 17676 32608 17692 32672
rect 17756 32608 17772 32672
rect 17836 32608 17852 32672
rect 17916 32608 17922 32672
rect 17606 32607 17922 32608
rect 16941 32330 17007 32333
rect 16806 32328 17007 32330
rect 16806 32272 16946 32328
rect 17002 32272 17007 32328
rect 16806 32270 17007 32272
rect 1946 32128 2262 32129
rect 1946 32064 1952 32128
rect 2016 32064 2032 32128
rect 2096 32064 2112 32128
rect 2176 32064 2192 32128
rect 2256 32064 2262 32128
rect 1946 32063 2262 32064
rect 6946 32128 7262 32129
rect 6946 32064 6952 32128
rect 7016 32064 7032 32128
rect 7096 32064 7112 32128
rect 7176 32064 7192 32128
rect 7256 32064 7262 32128
rect 6946 32063 7262 32064
rect 11946 32128 12262 32129
rect 11946 32064 11952 32128
rect 12016 32064 12032 32128
rect 12096 32064 12112 32128
rect 12176 32064 12192 32128
rect 12256 32064 12262 32128
rect 11946 32063 12262 32064
rect 16806 31789 16866 32270
rect 16941 32267 17007 32270
rect 16946 32128 17262 32129
rect 16946 32064 16952 32128
rect 17016 32064 17032 32128
rect 17096 32064 17112 32128
rect 17176 32064 17192 32128
rect 17256 32064 17262 32128
rect 16946 32063 17262 32064
rect 2497 31786 2563 31789
rect 4838 31786 4844 31788
rect 2497 31784 4844 31786
rect 2497 31728 2502 31784
rect 2558 31728 4844 31784
rect 2497 31726 4844 31728
rect 2497 31723 2563 31726
rect 4838 31724 4844 31726
rect 4908 31724 4914 31788
rect 16757 31784 16866 31789
rect 16757 31728 16762 31784
rect 16818 31728 16866 31784
rect 16757 31726 16866 31728
rect 16757 31723 16823 31726
rect 2606 31584 2922 31585
rect 2606 31520 2612 31584
rect 2676 31520 2692 31584
rect 2756 31520 2772 31584
rect 2836 31520 2852 31584
rect 2916 31520 2922 31584
rect 2606 31519 2922 31520
rect 7606 31584 7922 31585
rect 7606 31520 7612 31584
rect 7676 31520 7692 31584
rect 7756 31520 7772 31584
rect 7836 31520 7852 31584
rect 7916 31520 7922 31584
rect 7606 31519 7922 31520
rect 12606 31584 12922 31585
rect 12606 31520 12612 31584
rect 12676 31520 12692 31584
rect 12756 31520 12772 31584
rect 12836 31520 12852 31584
rect 12916 31520 12922 31584
rect 12606 31519 12922 31520
rect 17606 31584 17922 31585
rect 17606 31520 17612 31584
rect 17676 31520 17692 31584
rect 17756 31520 17772 31584
rect 17836 31520 17852 31584
rect 17916 31520 17922 31584
rect 17606 31519 17922 31520
rect 18229 31378 18295 31381
rect 19200 31378 20000 31408
rect 18229 31376 20000 31378
rect 18229 31320 18234 31376
rect 18290 31320 20000 31376
rect 18229 31318 20000 31320
rect 18229 31315 18295 31318
rect 19200 31288 20000 31318
rect 1946 31040 2262 31041
rect 1946 30976 1952 31040
rect 2016 30976 2032 31040
rect 2096 30976 2112 31040
rect 2176 30976 2192 31040
rect 2256 30976 2262 31040
rect 1946 30975 2262 30976
rect 6946 31040 7262 31041
rect 6946 30976 6952 31040
rect 7016 30976 7032 31040
rect 7096 30976 7112 31040
rect 7176 30976 7192 31040
rect 7256 30976 7262 31040
rect 6946 30975 7262 30976
rect 11946 31040 12262 31041
rect 11946 30976 11952 31040
rect 12016 30976 12032 31040
rect 12096 30976 12112 31040
rect 12176 30976 12192 31040
rect 12256 30976 12262 31040
rect 11946 30975 12262 30976
rect 16946 31040 17262 31041
rect 16946 30976 16952 31040
rect 17016 30976 17032 31040
rect 17096 30976 17112 31040
rect 17176 30976 17192 31040
rect 17256 30976 17262 31040
rect 16946 30975 17262 30976
rect 2606 30496 2922 30497
rect 2606 30432 2612 30496
rect 2676 30432 2692 30496
rect 2756 30432 2772 30496
rect 2836 30432 2852 30496
rect 2916 30432 2922 30496
rect 2606 30431 2922 30432
rect 7606 30496 7922 30497
rect 7606 30432 7612 30496
rect 7676 30432 7692 30496
rect 7756 30432 7772 30496
rect 7836 30432 7852 30496
rect 7916 30432 7922 30496
rect 7606 30431 7922 30432
rect 12606 30496 12922 30497
rect 12606 30432 12612 30496
rect 12676 30432 12692 30496
rect 12756 30432 12772 30496
rect 12836 30432 12852 30496
rect 12916 30432 12922 30496
rect 12606 30431 12922 30432
rect 17606 30496 17922 30497
rect 17606 30432 17612 30496
rect 17676 30432 17692 30496
rect 17756 30432 17772 30496
rect 17836 30432 17852 30496
rect 17916 30432 17922 30496
rect 17606 30431 17922 30432
rect 1946 29952 2262 29953
rect 1946 29888 1952 29952
rect 2016 29888 2032 29952
rect 2096 29888 2112 29952
rect 2176 29888 2192 29952
rect 2256 29888 2262 29952
rect 1946 29887 2262 29888
rect 6946 29952 7262 29953
rect 6946 29888 6952 29952
rect 7016 29888 7032 29952
rect 7096 29888 7112 29952
rect 7176 29888 7192 29952
rect 7256 29888 7262 29952
rect 6946 29887 7262 29888
rect 11946 29952 12262 29953
rect 11946 29888 11952 29952
rect 12016 29888 12032 29952
rect 12096 29888 12112 29952
rect 12176 29888 12192 29952
rect 12256 29888 12262 29952
rect 11946 29887 12262 29888
rect 16946 29952 17262 29953
rect 16946 29888 16952 29952
rect 17016 29888 17032 29952
rect 17096 29888 17112 29952
rect 17176 29888 17192 29952
rect 17256 29888 17262 29952
rect 16946 29887 17262 29888
rect 14181 29882 14247 29885
rect 14958 29882 14964 29884
rect 14181 29880 14964 29882
rect 14181 29824 14186 29880
rect 14242 29824 14964 29880
rect 14181 29822 14964 29824
rect 14181 29819 14247 29822
rect 14958 29820 14964 29822
rect 15028 29820 15034 29884
rect 18229 29474 18295 29477
rect 19200 29474 20000 29504
rect 18229 29472 20000 29474
rect 18229 29416 18234 29472
rect 18290 29416 20000 29472
rect 18229 29414 20000 29416
rect 18229 29411 18295 29414
rect 2606 29408 2922 29409
rect 2606 29344 2612 29408
rect 2676 29344 2692 29408
rect 2756 29344 2772 29408
rect 2836 29344 2852 29408
rect 2916 29344 2922 29408
rect 2606 29343 2922 29344
rect 7606 29408 7922 29409
rect 7606 29344 7612 29408
rect 7676 29344 7692 29408
rect 7756 29344 7772 29408
rect 7836 29344 7852 29408
rect 7916 29344 7922 29408
rect 7606 29343 7922 29344
rect 12606 29408 12922 29409
rect 12606 29344 12612 29408
rect 12676 29344 12692 29408
rect 12756 29344 12772 29408
rect 12836 29344 12852 29408
rect 12916 29344 12922 29408
rect 12606 29343 12922 29344
rect 17606 29408 17922 29409
rect 17606 29344 17612 29408
rect 17676 29344 17692 29408
rect 17756 29344 17772 29408
rect 17836 29344 17852 29408
rect 17916 29344 17922 29408
rect 19200 29384 20000 29414
rect 17606 29343 17922 29344
rect 1946 28864 2262 28865
rect 1946 28800 1952 28864
rect 2016 28800 2032 28864
rect 2096 28800 2112 28864
rect 2176 28800 2192 28864
rect 2256 28800 2262 28864
rect 1946 28799 2262 28800
rect 6946 28864 7262 28865
rect 6946 28800 6952 28864
rect 7016 28800 7032 28864
rect 7096 28800 7112 28864
rect 7176 28800 7192 28864
rect 7256 28800 7262 28864
rect 6946 28799 7262 28800
rect 11946 28864 12262 28865
rect 11946 28800 11952 28864
rect 12016 28800 12032 28864
rect 12096 28800 12112 28864
rect 12176 28800 12192 28864
rect 12256 28800 12262 28864
rect 11946 28799 12262 28800
rect 16946 28864 17262 28865
rect 16946 28800 16952 28864
rect 17016 28800 17032 28864
rect 17096 28800 17112 28864
rect 17176 28800 17192 28864
rect 17256 28800 17262 28864
rect 16946 28799 17262 28800
rect 7925 28522 7991 28525
rect 8334 28522 8340 28524
rect 7925 28520 8340 28522
rect 7925 28464 7930 28520
rect 7986 28464 8340 28520
rect 7925 28462 8340 28464
rect 7925 28459 7991 28462
rect 8334 28460 8340 28462
rect 8404 28460 8410 28524
rect 2606 28320 2922 28321
rect 2606 28256 2612 28320
rect 2676 28256 2692 28320
rect 2756 28256 2772 28320
rect 2836 28256 2852 28320
rect 2916 28256 2922 28320
rect 2606 28255 2922 28256
rect 7606 28320 7922 28321
rect 7606 28256 7612 28320
rect 7676 28256 7692 28320
rect 7756 28256 7772 28320
rect 7836 28256 7852 28320
rect 7916 28256 7922 28320
rect 7606 28255 7922 28256
rect 12606 28320 12922 28321
rect 12606 28256 12612 28320
rect 12676 28256 12692 28320
rect 12756 28256 12772 28320
rect 12836 28256 12852 28320
rect 12916 28256 12922 28320
rect 12606 28255 12922 28256
rect 17606 28320 17922 28321
rect 17606 28256 17612 28320
rect 17676 28256 17692 28320
rect 17756 28256 17772 28320
rect 17836 28256 17852 28320
rect 17916 28256 17922 28320
rect 17606 28255 17922 28256
rect 1946 27776 2262 27777
rect 1946 27712 1952 27776
rect 2016 27712 2032 27776
rect 2096 27712 2112 27776
rect 2176 27712 2192 27776
rect 2256 27712 2262 27776
rect 1946 27711 2262 27712
rect 6946 27776 7262 27777
rect 6946 27712 6952 27776
rect 7016 27712 7032 27776
rect 7096 27712 7112 27776
rect 7176 27712 7192 27776
rect 7256 27712 7262 27776
rect 6946 27711 7262 27712
rect 11946 27776 12262 27777
rect 11946 27712 11952 27776
rect 12016 27712 12032 27776
rect 12096 27712 12112 27776
rect 12176 27712 12192 27776
rect 12256 27712 12262 27776
rect 11946 27711 12262 27712
rect 16946 27776 17262 27777
rect 16946 27712 16952 27776
rect 17016 27712 17032 27776
rect 17096 27712 17112 27776
rect 17176 27712 17192 27776
rect 17256 27712 17262 27776
rect 16946 27711 17262 27712
rect 17861 27570 17927 27573
rect 19200 27570 20000 27600
rect 17861 27568 20000 27570
rect 17861 27512 17866 27568
rect 17922 27512 20000 27568
rect 17861 27510 20000 27512
rect 17861 27507 17927 27510
rect 19200 27480 20000 27510
rect 2606 27232 2922 27233
rect 2606 27168 2612 27232
rect 2676 27168 2692 27232
rect 2756 27168 2772 27232
rect 2836 27168 2852 27232
rect 2916 27168 2922 27232
rect 2606 27167 2922 27168
rect 7606 27232 7922 27233
rect 7606 27168 7612 27232
rect 7676 27168 7692 27232
rect 7756 27168 7772 27232
rect 7836 27168 7852 27232
rect 7916 27168 7922 27232
rect 7606 27167 7922 27168
rect 12606 27232 12922 27233
rect 12606 27168 12612 27232
rect 12676 27168 12692 27232
rect 12756 27168 12772 27232
rect 12836 27168 12852 27232
rect 12916 27168 12922 27232
rect 12606 27167 12922 27168
rect 17606 27232 17922 27233
rect 17606 27168 17612 27232
rect 17676 27168 17692 27232
rect 17756 27168 17772 27232
rect 17836 27168 17852 27232
rect 17916 27168 17922 27232
rect 17606 27167 17922 27168
rect 8937 27026 9003 27029
rect 9438 27026 9444 27028
rect 8937 27024 9444 27026
rect 8937 26968 8942 27024
rect 8998 26968 9444 27024
rect 8937 26966 9444 26968
rect 8937 26963 9003 26966
rect 9438 26964 9444 26966
rect 9508 26964 9514 27028
rect 8477 26890 8543 26893
rect 9254 26890 9260 26892
rect 8477 26888 9260 26890
rect 8477 26832 8482 26888
rect 8538 26832 9260 26888
rect 8477 26830 9260 26832
rect 8477 26827 8543 26830
rect 9254 26828 9260 26830
rect 9324 26828 9330 26892
rect 1946 26688 2262 26689
rect 1946 26624 1952 26688
rect 2016 26624 2032 26688
rect 2096 26624 2112 26688
rect 2176 26624 2192 26688
rect 2256 26624 2262 26688
rect 1946 26623 2262 26624
rect 6946 26688 7262 26689
rect 6946 26624 6952 26688
rect 7016 26624 7032 26688
rect 7096 26624 7112 26688
rect 7176 26624 7192 26688
rect 7256 26624 7262 26688
rect 6946 26623 7262 26624
rect 11946 26688 12262 26689
rect 11946 26624 11952 26688
rect 12016 26624 12032 26688
rect 12096 26624 12112 26688
rect 12176 26624 12192 26688
rect 12256 26624 12262 26688
rect 11946 26623 12262 26624
rect 16946 26688 17262 26689
rect 16946 26624 16952 26688
rect 17016 26624 17032 26688
rect 17096 26624 17112 26688
rect 17176 26624 17192 26688
rect 17256 26624 17262 26688
rect 16946 26623 17262 26624
rect 8109 26346 8175 26349
rect 8109 26344 8218 26346
rect 8109 26288 8114 26344
rect 8170 26288 8218 26344
rect 8109 26283 8218 26288
rect 2606 26144 2922 26145
rect 2606 26080 2612 26144
rect 2676 26080 2692 26144
rect 2756 26080 2772 26144
rect 2836 26080 2852 26144
rect 2916 26080 2922 26144
rect 2606 26079 2922 26080
rect 7606 26144 7922 26145
rect 7606 26080 7612 26144
rect 7676 26080 7692 26144
rect 7756 26080 7772 26144
rect 7836 26080 7852 26144
rect 7916 26080 7922 26144
rect 7606 26079 7922 26080
rect 8017 26074 8083 26077
rect 8158 26074 8218 26283
rect 11145 26210 11211 26213
rect 11278 26210 11284 26212
rect 11145 26208 11284 26210
rect 11145 26152 11150 26208
rect 11206 26152 11284 26208
rect 11145 26150 11284 26152
rect 11145 26147 11211 26150
rect 11278 26148 11284 26150
rect 11348 26148 11354 26212
rect 12606 26144 12922 26145
rect 12606 26080 12612 26144
rect 12676 26080 12692 26144
rect 12756 26080 12772 26144
rect 12836 26080 12852 26144
rect 12916 26080 12922 26144
rect 12606 26079 12922 26080
rect 17606 26144 17922 26145
rect 17606 26080 17612 26144
rect 17676 26080 17692 26144
rect 17756 26080 17772 26144
rect 17836 26080 17852 26144
rect 17916 26080 17922 26144
rect 17606 26079 17922 26080
rect 8017 26072 8218 26074
rect 8017 26016 8022 26072
rect 8078 26016 8218 26072
rect 8017 26014 8218 26016
rect 8293 26076 8359 26077
rect 10133 26076 10199 26077
rect 8293 26072 8340 26076
rect 8404 26074 8410 26076
rect 10133 26074 10180 26076
rect 8293 26016 8298 26072
rect 8017 26011 8083 26014
rect 8293 26012 8340 26016
rect 8404 26014 8450 26074
rect 10088 26072 10180 26074
rect 10088 26016 10138 26072
rect 10088 26014 10180 26016
rect 8404 26012 8410 26014
rect 10133 26012 10180 26014
rect 10244 26012 10250 26076
rect 11053 26074 11119 26077
rect 11646 26074 11652 26076
rect 11053 26072 11652 26074
rect 11053 26016 11058 26072
rect 11114 26016 11652 26072
rect 11053 26014 11652 26016
rect 8293 26011 8359 26012
rect 10133 26011 10199 26012
rect 11053 26011 11119 26014
rect 11646 26012 11652 26014
rect 11716 26012 11722 26076
rect 18229 25666 18295 25669
rect 19200 25666 20000 25696
rect 18229 25664 20000 25666
rect 18229 25608 18234 25664
rect 18290 25608 20000 25664
rect 18229 25606 20000 25608
rect 18229 25603 18295 25606
rect 1946 25600 2262 25601
rect 1946 25536 1952 25600
rect 2016 25536 2032 25600
rect 2096 25536 2112 25600
rect 2176 25536 2192 25600
rect 2256 25536 2262 25600
rect 1946 25535 2262 25536
rect 6946 25600 7262 25601
rect 6946 25536 6952 25600
rect 7016 25536 7032 25600
rect 7096 25536 7112 25600
rect 7176 25536 7192 25600
rect 7256 25536 7262 25600
rect 6946 25535 7262 25536
rect 11946 25600 12262 25601
rect 11946 25536 11952 25600
rect 12016 25536 12032 25600
rect 12096 25536 12112 25600
rect 12176 25536 12192 25600
rect 12256 25536 12262 25600
rect 11946 25535 12262 25536
rect 16946 25600 17262 25601
rect 16946 25536 16952 25600
rect 17016 25536 17032 25600
rect 17096 25536 17112 25600
rect 17176 25536 17192 25600
rect 17256 25536 17262 25600
rect 19200 25576 20000 25606
rect 16946 25535 17262 25536
rect 10317 25396 10383 25397
rect 10317 25394 10364 25396
rect 10272 25392 10364 25394
rect 10272 25336 10322 25392
rect 10272 25334 10364 25336
rect 10317 25332 10364 25334
rect 10428 25332 10434 25396
rect 10317 25331 10383 25332
rect 2606 25056 2922 25057
rect 2606 24992 2612 25056
rect 2676 24992 2692 25056
rect 2756 24992 2772 25056
rect 2836 24992 2852 25056
rect 2916 24992 2922 25056
rect 2606 24991 2922 24992
rect 7606 25056 7922 25057
rect 7606 24992 7612 25056
rect 7676 24992 7692 25056
rect 7756 24992 7772 25056
rect 7836 24992 7852 25056
rect 7916 24992 7922 25056
rect 7606 24991 7922 24992
rect 12606 25056 12922 25057
rect 12606 24992 12612 25056
rect 12676 24992 12692 25056
rect 12756 24992 12772 25056
rect 12836 24992 12852 25056
rect 12916 24992 12922 25056
rect 12606 24991 12922 24992
rect 17606 25056 17922 25057
rect 17606 24992 17612 25056
rect 17676 24992 17692 25056
rect 17756 24992 17772 25056
rect 17836 24992 17852 25056
rect 17916 24992 17922 25056
rect 17606 24991 17922 24992
rect 1710 24788 1716 24852
rect 1780 24850 1786 24852
rect 9765 24850 9831 24853
rect 1780 24848 9831 24850
rect 1780 24792 9770 24848
rect 9826 24792 9831 24848
rect 1780 24790 9831 24792
rect 1780 24788 1786 24790
rect 9765 24787 9831 24790
rect 13302 24788 13308 24852
rect 13372 24850 13378 24852
rect 13537 24850 13603 24853
rect 13372 24848 13603 24850
rect 13372 24792 13542 24848
rect 13598 24792 13603 24848
rect 13372 24790 13603 24792
rect 13372 24788 13378 24790
rect 13537 24787 13603 24790
rect 13118 24652 13124 24716
rect 13188 24714 13194 24716
rect 16389 24714 16455 24717
rect 13188 24712 16455 24714
rect 13188 24656 16394 24712
rect 16450 24656 16455 24712
rect 13188 24654 16455 24656
rect 13188 24652 13194 24654
rect 16389 24651 16455 24654
rect 1946 24512 2262 24513
rect 1946 24448 1952 24512
rect 2016 24448 2032 24512
rect 2096 24448 2112 24512
rect 2176 24448 2192 24512
rect 2256 24448 2262 24512
rect 1946 24447 2262 24448
rect 6946 24512 7262 24513
rect 6946 24448 6952 24512
rect 7016 24448 7032 24512
rect 7096 24448 7112 24512
rect 7176 24448 7192 24512
rect 7256 24448 7262 24512
rect 6946 24447 7262 24448
rect 11946 24512 12262 24513
rect 11946 24448 11952 24512
rect 12016 24448 12032 24512
rect 12096 24448 12112 24512
rect 12176 24448 12192 24512
rect 12256 24448 12262 24512
rect 11946 24447 12262 24448
rect 16946 24512 17262 24513
rect 16946 24448 16952 24512
rect 17016 24448 17032 24512
rect 17096 24448 17112 24512
rect 17176 24448 17192 24512
rect 17256 24448 17262 24512
rect 16946 24447 17262 24448
rect 2606 23968 2922 23969
rect 2606 23904 2612 23968
rect 2676 23904 2692 23968
rect 2756 23904 2772 23968
rect 2836 23904 2852 23968
rect 2916 23904 2922 23968
rect 2606 23903 2922 23904
rect 7606 23968 7922 23969
rect 7606 23904 7612 23968
rect 7676 23904 7692 23968
rect 7756 23904 7772 23968
rect 7836 23904 7852 23968
rect 7916 23904 7922 23968
rect 7606 23903 7922 23904
rect 12606 23968 12922 23969
rect 12606 23904 12612 23968
rect 12676 23904 12692 23968
rect 12756 23904 12772 23968
rect 12836 23904 12852 23968
rect 12916 23904 12922 23968
rect 12606 23903 12922 23904
rect 17606 23968 17922 23969
rect 17606 23904 17612 23968
rect 17676 23904 17692 23968
rect 17756 23904 17772 23968
rect 17836 23904 17852 23968
rect 17916 23904 17922 23968
rect 17606 23903 17922 23904
rect 18229 23762 18295 23765
rect 19200 23762 20000 23792
rect 18229 23760 20000 23762
rect 18229 23704 18234 23760
rect 18290 23704 20000 23760
rect 18229 23702 20000 23704
rect 18229 23699 18295 23702
rect 19200 23672 20000 23702
rect 4286 23564 4292 23628
rect 4356 23626 4362 23628
rect 16941 23626 17007 23629
rect 4356 23624 17007 23626
rect 4356 23568 16946 23624
rect 17002 23568 17007 23624
rect 4356 23566 17007 23568
rect 4356 23564 4362 23566
rect 16941 23563 17007 23566
rect 1946 23424 2262 23425
rect 1946 23360 1952 23424
rect 2016 23360 2032 23424
rect 2096 23360 2112 23424
rect 2176 23360 2192 23424
rect 2256 23360 2262 23424
rect 1946 23359 2262 23360
rect 6946 23424 7262 23425
rect 6946 23360 6952 23424
rect 7016 23360 7032 23424
rect 7096 23360 7112 23424
rect 7176 23360 7192 23424
rect 7256 23360 7262 23424
rect 6946 23359 7262 23360
rect 11946 23424 12262 23425
rect 11946 23360 11952 23424
rect 12016 23360 12032 23424
rect 12096 23360 12112 23424
rect 12176 23360 12192 23424
rect 12256 23360 12262 23424
rect 11946 23359 12262 23360
rect 16946 23424 17262 23425
rect 16946 23360 16952 23424
rect 17016 23360 17032 23424
rect 17096 23360 17112 23424
rect 17176 23360 17192 23424
rect 17256 23360 17262 23424
rect 16946 23359 17262 23360
rect 2606 22880 2922 22881
rect 2606 22816 2612 22880
rect 2676 22816 2692 22880
rect 2756 22816 2772 22880
rect 2836 22816 2852 22880
rect 2916 22816 2922 22880
rect 2606 22815 2922 22816
rect 7606 22880 7922 22881
rect 7606 22816 7612 22880
rect 7676 22816 7692 22880
rect 7756 22816 7772 22880
rect 7836 22816 7852 22880
rect 7916 22816 7922 22880
rect 7606 22815 7922 22816
rect 12606 22880 12922 22881
rect 12606 22816 12612 22880
rect 12676 22816 12692 22880
rect 12756 22816 12772 22880
rect 12836 22816 12852 22880
rect 12916 22816 12922 22880
rect 12606 22815 12922 22816
rect 17606 22880 17922 22881
rect 17606 22816 17612 22880
rect 17676 22816 17692 22880
rect 17756 22816 17772 22880
rect 17836 22816 17852 22880
rect 17916 22816 17922 22880
rect 17606 22815 17922 22816
rect 14406 22476 14412 22540
rect 14476 22538 14482 22540
rect 17217 22538 17283 22541
rect 14476 22536 17283 22538
rect 14476 22480 17222 22536
rect 17278 22480 17283 22536
rect 14476 22478 17283 22480
rect 14476 22476 14482 22478
rect 17217 22475 17283 22478
rect 1946 22336 2262 22337
rect 1946 22272 1952 22336
rect 2016 22272 2032 22336
rect 2096 22272 2112 22336
rect 2176 22272 2192 22336
rect 2256 22272 2262 22336
rect 1946 22271 2262 22272
rect 6946 22336 7262 22337
rect 6946 22272 6952 22336
rect 7016 22272 7032 22336
rect 7096 22272 7112 22336
rect 7176 22272 7192 22336
rect 7256 22272 7262 22336
rect 6946 22271 7262 22272
rect 11946 22336 12262 22337
rect 11946 22272 11952 22336
rect 12016 22272 12032 22336
rect 12096 22272 12112 22336
rect 12176 22272 12192 22336
rect 12256 22272 12262 22336
rect 11946 22271 12262 22272
rect 16946 22336 17262 22337
rect 16946 22272 16952 22336
rect 17016 22272 17032 22336
rect 17096 22272 17112 22336
rect 17176 22272 17192 22336
rect 17256 22272 17262 22336
rect 16946 22271 17262 22272
rect 4153 21994 4219 21997
rect 4470 21994 4476 21996
rect 4153 21992 4476 21994
rect 4153 21936 4158 21992
rect 4214 21936 4476 21992
rect 4153 21934 4476 21936
rect 4153 21931 4219 21934
rect 4470 21932 4476 21934
rect 4540 21932 4546 21996
rect 18229 21858 18295 21861
rect 19200 21858 20000 21888
rect 18229 21856 20000 21858
rect 18229 21800 18234 21856
rect 18290 21800 20000 21856
rect 18229 21798 20000 21800
rect 18229 21795 18295 21798
rect 2606 21792 2922 21793
rect 2606 21728 2612 21792
rect 2676 21728 2692 21792
rect 2756 21728 2772 21792
rect 2836 21728 2852 21792
rect 2916 21728 2922 21792
rect 2606 21727 2922 21728
rect 7606 21792 7922 21793
rect 7606 21728 7612 21792
rect 7676 21728 7692 21792
rect 7756 21728 7772 21792
rect 7836 21728 7852 21792
rect 7916 21728 7922 21792
rect 7606 21727 7922 21728
rect 12606 21792 12922 21793
rect 12606 21728 12612 21792
rect 12676 21728 12692 21792
rect 12756 21728 12772 21792
rect 12836 21728 12852 21792
rect 12916 21728 12922 21792
rect 12606 21727 12922 21728
rect 17606 21792 17922 21793
rect 17606 21728 17612 21792
rect 17676 21728 17692 21792
rect 17756 21728 17772 21792
rect 17836 21728 17852 21792
rect 17916 21728 17922 21792
rect 19200 21768 20000 21798
rect 17606 21727 17922 21728
rect 1946 21248 2262 21249
rect 1946 21184 1952 21248
rect 2016 21184 2032 21248
rect 2096 21184 2112 21248
rect 2176 21184 2192 21248
rect 2256 21184 2262 21248
rect 1946 21183 2262 21184
rect 6946 21248 7262 21249
rect 6946 21184 6952 21248
rect 7016 21184 7032 21248
rect 7096 21184 7112 21248
rect 7176 21184 7192 21248
rect 7256 21184 7262 21248
rect 6946 21183 7262 21184
rect 11946 21248 12262 21249
rect 11946 21184 11952 21248
rect 12016 21184 12032 21248
rect 12096 21184 12112 21248
rect 12176 21184 12192 21248
rect 12256 21184 12262 21248
rect 11946 21183 12262 21184
rect 16946 21248 17262 21249
rect 16946 21184 16952 21248
rect 17016 21184 17032 21248
rect 17096 21184 17112 21248
rect 17176 21184 17192 21248
rect 17256 21184 17262 21248
rect 16946 21183 17262 21184
rect 11421 21042 11487 21045
rect 16430 21042 16436 21044
rect 11421 21040 16436 21042
rect 11421 20984 11426 21040
rect 11482 20984 16436 21040
rect 11421 20982 16436 20984
rect 11421 20979 11487 20982
rect 16430 20980 16436 20982
rect 16500 21042 16506 21044
rect 17217 21042 17283 21045
rect 16500 21040 17283 21042
rect 16500 20984 17222 21040
rect 17278 20984 17283 21040
rect 16500 20982 17283 20984
rect 16500 20980 16506 20982
rect 17217 20979 17283 20982
rect 4470 20708 4476 20772
rect 4540 20770 4546 20772
rect 4797 20770 4863 20773
rect 4540 20768 4863 20770
rect 4540 20712 4802 20768
rect 4858 20712 4863 20768
rect 4540 20710 4863 20712
rect 4540 20708 4546 20710
rect 4797 20707 4863 20710
rect 2606 20704 2922 20705
rect 2606 20640 2612 20704
rect 2676 20640 2692 20704
rect 2756 20640 2772 20704
rect 2836 20640 2852 20704
rect 2916 20640 2922 20704
rect 2606 20639 2922 20640
rect 7606 20704 7922 20705
rect 7606 20640 7612 20704
rect 7676 20640 7692 20704
rect 7756 20640 7772 20704
rect 7836 20640 7852 20704
rect 7916 20640 7922 20704
rect 7606 20639 7922 20640
rect 12606 20704 12922 20705
rect 12606 20640 12612 20704
rect 12676 20640 12692 20704
rect 12756 20640 12772 20704
rect 12836 20640 12852 20704
rect 12916 20640 12922 20704
rect 12606 20639 12922 20640
rect 17606 20704 17922 20705
rect 17606 20640 17612 20704
rect 17676 20640 17692 20704
rect 17756 20640 17772 20704
rect 17836 20640 17852 20704
rect 17916 20640 17922 20704
rect 17606 20639 17922 20640
rect 1946 20160 2262 20161
rect 1946 20096 1952 20160
rect 2016 20096 2032 20160
rect 2096 20096 2112 20160
rect 2176 20096 2192 20160
rect 2256 20096 2262 20160
rect 1946 20095 2262 20096
rect 6946 20160 7262 20161
rect 6946 20096 6952 20160
rect 7016 20096 7032 20160
rect 7096 20096 7112 20160
rect 7176 20096 7192 20160
rect 7256 20096 7262 20160
rect 6946 20095 7262 20096
rect 11946 20160 12262 20161
rect 11946 20096 11952 20160
rect 12016 20096 12032 20160
rect 12096 20096 12112 20160
rect 12176 20096 12192 20160
rect 12256 20096 12262 20160
rect 11946 20095 12262 20096
rect 16946 20160 17262 20161
rect 16946 20096 16952 20160
rect 17016 20096 17032 20160
rect 17096 20096 17112 20160
rect 17176 20096 17192 20160
rect 17256 20096 17262 20160
rect 16946 20095 17262 20096
rect 6494 19892 6500 19956
rect 6564 19954 6570 19956
rect 12157 19954 12223 19957
rect 6564 19952 12223 19954
rect 6564 19896 12162 19952
rect 12218 19896 12223 19952
rect 6564 19894 12223 19896
rect 6564 19892 6570 19894
rect 12157 19891 12223 19894
rect 18229 19954 18295 19957
rect 19200 19954 20000 19984
rect 18229 19952 20000 19954
rect 18229 19896 18234 19952
rect 18290 19896 20000 19952
rect 18229 19894 20000 19896
rect 18229 19891 18295 19894
rect 19200 19864 20000 19894
rect 2606 19616 2922 19617
rect 2606 19552 2612 19616
rect 2676 19552 2692 19616
rect 2756 19552 2772 19616
rect 2836 19552 2852 19616
rect 2916 19552 2922 19616
rect 2606 19551 2922 19552
rect 7606 19616 7922 19617
rect 7606 19552 7612 19616
rect 7676 19552 7692 19616
rect 7756 19552 7772 19616
rect 7836 19552 7852 19616
rect 7916 19552 7922 19616
rect 7606 19551 7922 19552
rect 12606 19616 12922 19617
rect 12606 19552 12612 19616
rect 12676 19552 12692 19616
rect 12756 19552 12772 19616
rect 12836 19552 12852 19616
rect 12916 19552 12922 19616
rect 12606 19551 12922 19552
rect 17606 19616 17922 19617
rect 17606 19552 17612 19616
rect 17676 19552 17692 19616
rect 17756 19552 17772 19616
rect 17836 19552 17852 19616
rect 17916 19552 17922 19616
rect 17606 19551 17922 19552
rect 1946 19072 2262 19073
rect 1946 19008 1952 19072
rect 2016 19008 2032 19072
rect 2096 19008 2112 19072
rect 2176 19008 2192 19072
rect 2256 19008 2262 19072
rect 1946 19007 2262 19008
rect 6946 19072 7262 19073
rect 6946 19008 6952 19072
rect 7016 19008 7032 19072
rect 7096 19008 7112 19072
rect 7176 19008 7192 19072
rect 7256 19008 7262 19072
rect 6946 19007 7262 19008
rect 11946 19072 12262 19073
rect 11946 19008 11952 19072
rect 12016 19008 12032 19072
rect 12096 19008 12112 19072
rect 12176 19008 12192 19072
rect 12256 19008 12262 19072
rect 11946 19007 12262 19008
rect 16946 19072 17262 19073
rect 16946 19008 16952 19072
rect 17016 19008 17032 19072
rect 17096 19008 17112 19072
rect 17176 19008 17192 19072
rect 17256 19008 17262 19072
rect 16946 19007 17262 19008
rect 2606 18528 2922 18529
rect 2606 18464 2612 18528
rect 2676 18464 2692 18528
rect 2756 18464 2772 18528
rect 2836 18464 2852 18528
rect 2916 18464 2922 18528
rect 2606 18463 2922 18464
rect 7606 18528 7922 18529
rect 7606 18464 7612 18528
rect 7676 18464 7692 18528
rect 7756 18464 7772 18528
rect 7836 18464 7852 18528
rect 7916 18464 7922 18528
rect 7606 18463 7922 18464
rect 12606 18528 12922 18529
rect 12606 18464 12612 18528
rect 12676 18464 12692 18528
rect 12756 18464 12772 18528
rect 12836 18464 12852 18528
rect 12916 18464 12922 18528
rect 12606 18463 12922 18464
rect 17606 18528 17922 18529
rect 17606 18464 17612 18528
rect 17676 18464 17692 18528
rect 17756 18464 17772 18528
rect 17836 18464 17852 18528
rect 17916 18464 17922 18528
rect 17606 18463 17922 18464
rect 18229 18050 18295 18053
rect 19200 18050 20000 18080
rect 18229 18048 20000 18050
rect 18229 17992 18234 18048
rect 18290 17992 20000 18048
rect 18229 17990 20000 17992
rect 18229 17987 18295 17990
rect 1946 17984 2262 17985
rect 1946 17920 1952 17984
rect 2016 17920 2032 17984
rect 2096 17920 2112 17984
rect 2176 17920 2192 17984
rect 2256 17920 2262 17984
rect 1946 17919 2262 17920
rect 6946 17984 7262 17985
rect 6946 17920 6952 17984
rect 7016 17920 7032 17984
rect 7096 17920 7112 17984
rect 7176 17920 7192 17984
rect 7256 17920 7262 17984
rect 6946 17919 7262 17920
rect 11946 17984 12262 17985
rect 11946 17920 11952 17984
rect 12016 17920 12032 17984
rect 12096 17920 12112 17984
rect 12176 17920 12192 17984
rect 12256 17920 12262 17984
rect 11946 17919 12262 17920
rect 16946 17984 17262 17985
rect 16946 17920 16952 17984
rect 17016 17920 17032 17984
rect 17096 17920 17112 17984
rect 17176 17920 17192 17984
rect 17256 17920 17262 17984
rect 19200 17960 20000 17990
rect 16946 17919 17262 17920
rect 2606 17440 2922 17441
rect 2606 17376 2612 17440
rect 2676 17376 2692 17440
rect 2756 17376 2772 17440
rect 2836 17376 2852 17440
rect 2916 17376 2922 17440
rect 2606 17375 2922 17376
rect 7606 17440 7922 17441
rect 7606 17376 7612 17440
rect 7676 17376 7692 17440
rect 7756 17376 7772 17440
rect 7836 17376 7852 17440
rect 7916 17376 7922 17440
rect 7606 17375 7922 17376
rect 12606 17440 12922 17441
rect 12606 17376 12612 17440
rect 12676 17376 12692 17440
rect 12756 17376 12772 17440
rect 12836 17376 12852 17440
rect 12916 17376 12922 17440
rect 12606 17375 12922 17376
rect 17606 17440 17922 17441
rect 17606 17376 17612 17440
rect 17676 17376 17692 17440
rect 17756 17376 17772 17440
rect 17836 17376 17852 17440
rect 17916 17376 17922 17440
rect 17606 17375 17922 17376
rect 1946 16896 2262 16897
rect 1946 16832 1952 16896
rect 2016 16832 2032 16896
rect 2096 16832 2112 16896
rect 2176 16832 2192 16896
rect 2256 16832 2262 16896
rect 1946 16831 2262 16832
rect 6946 16896 7262 16897
rect 6946 16832 6952 16896
rect 7016 16832 7032 16896
rect 7096 16832 7112 16896
rect 7176 16832 7192 16896
rect 7256 16832 7262 16896
rect 6946 16831 7262 16832
rect 11946 16896 12262 16897
rect 11946 16832 11952 16896
rect 12016 16832 12032 16896
rect 12096 16832 12112 16896
rect 12176 16832 12192 16896
rect 12256 16832 12262 16896
rect 11946 16831 12262 16832
rect 16946 16896 17262 16897
rect 16946 16832 16952 16896
rect 17016 16832 17032 16896
rect 17096 16832 17112 16896
rect 17176 16832 17192 16896
rect 17256 16832 17262 16896
rect 16946 16831 17262 16832
rect 6310 16628 6316 16692
rect 6380 16690 6386 16692
rect 17953 16690 18019 16693
rect 6380 16688 18019 16690
rect 6380 16632 17958 16688
rect 18014 16632 18019 16688
rect 6380 16630 18019 16632
rect 6380 16628 6386 16630
rect 17953 16627 18019 16630
rect 9029 16554 9095 16557
rect 14590 16554 14596 16556
rect 9029 16552 14596 16554
rect 9029 16496 9034 16552
rect 9090 16496 14596 16552
rect 9029 16494 14596 16496
rect 9029 16491 9095 16494
rect 14590 16492 14596 16494
rect 14660 16492 14666 16556
rect 2606 16352 2922 16353
rect 2606 16288 2612 16352
rect 2676 16288 2692 16352
rect 2756 16288 2772 16352
rect 2836 16288 2852 16352
rect 2916 16288 2922 16352
rect 2606 16287 2922 16288
rect 7606 16352 7922 16353
rect 7606 16288 7612 16352
rect 7676 16288 7692 16352
rect 7756 16288 7772 16352
rect 7836 16288 7852 16352
rect 7916 16288 7922 16352
rect 7606 16287 7922 16288
rect 12606 16352 12922 16353
rect 12606 16288 12612 16352
rect 12676 16288 12692 16352
rect 12756 16288 12772 16352
rect 12836 16288 12852 16352
rect 12916 16288 12922 16352
rect 12606 16287 12922 16288
rect 17606 16352 17922 16353
rect 17606 16288 17612 16352
rect 17676 16288 17692 16352
rect 17756 16288 17772 16352
rect 17836 16288 17852 16352
rect 17916 16288 17922 16352
rect 17606 16287 17922 16288
rect 18229 16146 18295 16149
rect 19200 16146 20000 16176
rect 18229 16144 20000 16146
rect 18229 16088 18234 16144
rect 18290 16088 20000 16144
rect 18229 16086 20000 16088
rect 18229 16083 18295 16086
rect 19200 16056 20000 16086
rect 1946 15808 2262 15809
rect 1946 15744 1952 15808
rect 2016 15744 2032 15808
rect 2096 15744 2112 15808
rect 2176 15744 2192 15808
rect 2256 15744 2262 15808
rect 1946 15743 2262 15744
rect 6946 15808 7262 15809
rect 6946 15744 6952 15808
rect 7016 15744 7032 15808
rect 7096 15744 7112 15808
rect 7176 15744 7192 15808
rect 7256 15744 7262 15808
rect 6946 15743 7262 15744
rect 11946 15808 12262 15809
rect 11946 15744 11952 15808
rect 12016 15744 12032 15808
rect 12096 15744 12112 15808
rect 12176 15744 12192 15808
rect 12256 15744 12262 15808
rect 11946 15743 12262 15744
rect 16946 15808 17262 15809
rect 16946 15744 16952 15808
rect 17016 15744 17032 15808
rect 17096 15744 17112 15808
rect 17176 15744 17192 15808
rect 17256 15744 17262 15808
rect 16946 15743 17262 15744
rect 11278 15540 11284 15604
rect 11348 15602 11354 15604
rect 12985 15602 13051 15605
rect 11348 15600 13051 15602
rect 11348 15544 12990 15600
rect 13046 15544 13051 15600
rect 11348 15542 13051 15544
rect 11348 15540 11354 15542
rect 12985 15539 13051 15542
rect 2606 15264 2922 15265
rect 2606 15200 2612 15264
rect 2676 15200 2692 15264
rect 2756 15200 2772 15264
rect 2836 15200 2852 15264
rect 2916 15200 2922 15264
rect 2606 15199 2922 15200
rect 7606 15264 7922 15265
rect 7606 15200 7612 15264
rect 7676 15200 7692 15264
rect 7756 15200 7772 15264
rect 7836 15200 7852 15264
rect 7916 15200 7922 15264
rect 7606 15199 7922 15200
rect 12606 15264 12922 15265
rect 12606 15200 12612 15264
rect 12676 15200 12692 15264
rect 12756 15200 12772 15264
rect 12836 15200 12852 15264
rect 12916 15200 12922 15264
rect 12606 15199 12922 15200
rect 17606 15264 17922 15265
rect 17606 15200 17612 15264
rect 17676 15200 17692 15264
rect 17756 15200 17772 15264
rect 17836 15200 17852 15264
rect 17916 15200 17922 15264
rect 17606 15199 17922 15200
rect 8385 15194 8451 15197
rect 8518 15194 8524 15196
rect 8385 15192 8524 15194
rect 8385 15136 8390 15192
rect 8446 15136 8524 15192
rect 8385 15134 8524 15136
rect 8385 15131 8451 15134
rect 8518 15132 8524 15134
rect 8588 15132 8594 15196
rect 3918 14996 3924 15060
rect 3988 15058 3994 15060
rect 7833 15058 7899 15061
rect 3988 15056 7899 15058
rect 3988 15000 7838 15056
rect 7894 15000 7899 15056
rect 3988 14998 7899 15000
rect 3988 14996 3994 14998
rect 7833 14995 7899 14998
rect 1526 14860 1532 14924
rect 1596 14922 1602 14924
rect 17677 14922 17743 14925
rect 1596 14920 17743 14922
rect 1596 14864 17682 14920
rect 17738 14864 17743 14920
rect 1596 14862 17743 14864
rect 1596 14860 1602 14862
rect 17677 14859 17743 14862
rect 1946 14720 2262 14721
rect 1946 14656 1952 14720
rect 2016 14656 2032 14720
rect 2096 14656 2112 14720
rect 2176 14656 2192 14720
rect 2256 14656 2262 14720
rect 1946 14655 2262 14656
rect 6946 14720 7262 14721
rect 6946 14656 6952 14720
rect 7016 14656 7032 14720
rect 7096 14656 7112 14720
rect 7176 14656 7192 14720
rect 7256 14656 7262 14720
rect 6946 14655 7262 14656
rect 11946 14720 12262 14721
rect 11946 14656 11952 14720
rect 12016 14656 12032 14720
rect 12096 14656 12112 14720
rect 12176 14656 12192 14720
rect 12256 14656 12262 14720
rect 11946 14655 12262 14656
rect 16946 14720 17262 14721
rect 16946 14656 16952 14720
rect 17016 14656 17032 14720
rect 17096 14656 17112 14720
rect 17176 14656 17192 14720
rect 17256 14656 17262 14720
rect 16946 14655 17262 14656
rect 18229 14242 18295 14245
rect 19200 14242 20000 14272
rect 18229 14240 20000 14242
rect 18229 14184 18234 14240
rect 18290 14184 20000 14240
rect 18229 14182 20000 14184
rect 18229 14179 18295 14182
rect 2606 14176 2922 14177
rect 2606 14112 2612 14176
rect 2676 14112 2692 14176
rect 2756 14112 2772 14176
rect 2836 14112 2852 14176
rect 2916 14112 2922 14176
rect 2606 14111 2922 14112
rect 7606 14176 7922 14177
rect 7606 14112 7612 14176
rect 7676 14112 7692 14176
rect 7756 14112 7772 14176
rect 7836 14112 7852 14176
rect 7916 14112 7922 14176
rect 7606 14111 7922 14112
rect 12606 14176 12922 14177
rect 12606 14112 12612 14176
rect 12676 14112 12692 14176
rect 12756 14112 12772 14176
rect 12836 14112 12852 14176
rect 12916 14112 12922 14176
rect 12606 14111 12922 14112
rect 17606 14176 17922 14177
rect 17606 14112 17612 14176
rect 17676 14112 17692 14176
rect 17756 14112 17772 14176
rect 17836 14112 17852 14176
rect 17916 14112 17922 14176
rect 19200 14152 20000 14182
rect 17606 14111 17922 14112
rect 1946 13632 2262 13633
rect 1946 13568 1952 13632
rect 2016 13568 2032 13632
rect 2096 13568 2112 13632
rect 2176 13568 2192 13632
rect 2256 13568 2262 13632
rect 1946 13567 2262 13568
rect 6946 13632 7262 13633
rect 6946 13568 6952 13632
rect 7016 13568 7032 13632
rect 7096 13568 7112 13632
rect 7176 13568 7192 13632
rect 7256 13568 7262 13632
rect 6946 13567 7262 13568
rect 11946 13632 12262 13633
rect 11946 13568 11952 13632
rect 12016 13568 12032 13632
rect 12096 13568 12112 13632
rect 12176 13568 12192 13632
rect 12256 13568 12262 13632
rect 11946 13567 12262 13568
rect 16946 13632 17262 13633
rect 16946 13568 16952 13632
rect 17016 13568 17032 13632
rect 17096 13568 17112 13632
rect 17176 13568 17192 13632
rect 17256 13568 17262 13632
rect 16946 13567 17262 13568
rect 11462 13228 11468 13292
rect 11532 13290 11538 13292
rect 16573 13290 16639 13293
rect 11532 13288 16639 13290
rect 11532 13232 16578 13288
rect 16634 13232 16639 13288
rect 11532 13230 16639 13232
rect 11532 13228 11538 13230
rect 16573 13227 16639 13230
rect 2606 13088 2922 13089
rect 2606 13024 2612 13088
rect 2676 13024 2692 13088
rect 2756 13024 2772 13088
rect 2836 13024 2852 13088
rect 2916 13024 2922 13088
rect 2606 13023 2922 13024
rect 7606 13088 7922 13089
rect 7606 13024 7612 13088
rect 7676 13024 7692 13088
rect 7756 13024 7772 13088
rect 7836 13024 7852 13088
rect 7916 13024 7922 13088
rect 7606 13023 7922 13024
rect 12606 13088 12922 13089
rect 12606 13024 12612 13088
rect 12676 13024 12692 13088
rect 12756 13024 12772 13088
rect 12836 13024 12852 13088
rect 12916 13024 12922 13088
rect 12606 13023 12922 13024
rect 17606 13088 17922 13089
rect 17606 13024 17612 13088
rect 17676 13024 17692 13088
rect 17756 13024 17772 13088
rect 17836 13024 17852 13088
rect 17916 13024 17922 13088
rect 17606 13023 17922 13024
rect 1946 12544 2262 12545
rect 1946 12480 1952 12544
rect 2016 12480 2032 12544
rect 2096 12480 2112 12544
rect 2176 12480 2192 12544
rect 2256 12480 2262 12544
rect 1946 12479 2262 12480
rect 6946 12544 7262 12545
rect 6946 12480 6952 12544
rect 7016 12480 7032 12544
rect 7096 12480 7112 12544
rect 7176 12480 7192 12544
rect 7256 12480 7262 12544
rect 6946 12479 7262 12480
rect 11946 12544 12262 12545
rect 11946 12480 11952 12544
rect 12016 12480 12032 12544
rect 12096 12480 12112 12544
rect 12176 12480 12192 12544
rect 12256 12480 12262 12544
rect 11946 12479 12262 12480
rect 16946 12544 17262 12545
rect 16946 12480 16952 12544
rect 17016 12480 17032 12544
rect 17096 12480 17112 12544
rect 17176 12480 17192 12544
rect 17256 12480 17262 12544
rect 16946 12479 17262 12480
rect 9070 12276 9076 12340
rect 9140 12338 9146 12340
rect 12157 12338 12223 12341
rect 9140 12336 12223 12338
rect 9140 12280 12162 12336
rect 12218 12280 12223 12336
rect 9140 12278 12223 12280
rect 9140 12276 9146 12278
rect 12157 12275 12223 12278
rect 18229 12338 18295 12341
rect 19200 12338 20000 12368
rect 18229 12336 20000 12338
rect 18229 12280 18234 12336
rect 18290 12280 20000 12336
rect 18229 12278 20000 12280
rect 18229 12275 18295 12278
rect 19200 12248 20000 12278
rect 10685 12202 10751 12205
rect 13670 12202 13676 12204
rect 10685 12200 13676 12202
rect 10685 12144 10690 12200
rect 10746 12144 13676 12200
rect 10685 12142 13676 12144
rect 10685 12139 10751 12142
rect 13670 12140 13676 12142
rect 13740 12140 13746 12204
rect 2606 12000 2922 12001
rect 2606 11936 2612 12000
rect 2676 11936 2692 12000
rect 2756 11936 2772 12000
rect 2836 11936 2852 12000
rect 2916 11936 2922 12000
rect 2606 11935 2922 11936
rect 7606 12000 7922 12001
rect 7606 11936 7612 12000
rect 7676 11936 7692 12000
rect 7756 11936 7772 12000
rect 7836 11936 7852 12000
rect 7916 11936 7922 12000
rect 7606 11935 7922 11936
rect 12606 12000 12922 12001
rect 12606 11936 12612 12000
rect 12676 11936 12692 12000
rect 12756 11936 12772 12000
rect 12836 11936 12852 12000
rect 12916 11936 12922 12000
rect 12606 11935 12922 11936
rect 17606 12000 17922 12001
rect 17606 11936 17612 12000
rect 17676 11936 17692 12000
rect 17756 11936 17772 12000
rect 17836 11936 17852 12000
rect 17916 11936 17922 12000
rect 17606 11935 17922 11936
rect 1946 11456 2262 11457
rect 1946 11392 1952 11456
rect 2016 11392 2032 11456
rect 2096 11392 2112 11456
rect 2176 11392 2192 11456
rect 2256 11392 2262 11456
rect 1946 11391 2262 11392
rect 6946 11456 7262 11457
rect 6946 11392 6952 11456
rect 7016 11392 7032 11456
rect 7096 11392 7112 11456
rect 7176 11392 7192 11456
rect 7256 11392 7262 11456
rect 6946 11391 7262 11392
rect 11946 11456 12262 11457
rect 11946 11392 11952 11456
rect 12016 11392 12032 11456
rect 12096 11392 12112 11456
rect 12176 11392 12192 11456
rect 12256 11392 12262 11456
rect 11946 11391 12262 11392
rect 16946 11456 17262 11457
rect 16946 11392 16952 11456
rect 17016 11392 17032 11456
rect 17096 11392 17112 11456
rect 17176 11392 17192 11456
rect 17256 11392 17262 11456
rect 16946 11391 17262 11392
rect 8886 11188 8892 11252
rect 8956 11250 8962 11252
rect 15285 11250 15351 11253
rect 8956 11248 15351 11250
rect 8956 11192 15290 11248
rect 15346 11192 15351 11248
rect 8956 11190 15351 11192
rect 8956 11188 8962 11190
rect 15285 11187 15351 11190
rect 8293 11114 8359 11117
rect 15694 11114 15700 11116
rect 8293 11112 15700 11114
rect 8293 11056 8298 11112
rect 8354 11056 15700 11112
rect 8293 11054 15700 11056
rect 8293 11051 8359 11054
rect 15694 11052 15700 11054
rect 15764 11052 15770 11116
rect 2606 10912 2922 10913
rect 2606 10848 2612 10912
rect 2676 10848 2692 10912
rect 2756 10848 2772 10912
rect 2836 10848 2852 10912
rect 2916 10848 2922 10912
rect 2606 10847 2922 10848
rect 7606 10912 7922 10913
rect 7606 10848 7612 10912
rect 7676 10848 7692 10912
rect 7756 10848 7772 10912
rect 7836 10848 7852 10912
rect 7916 10848 7922 10912
rect 7606 10847 7922 10848
rect 12606 10912 12922 10913
rect 12606 10848 12612 10912
rect 12676 10848 12692 10912
rect 12756 10848 12772 10912
rect 12836 10848 12852 10912
rect 12916 10848 12922 10912
rect 12606 10847 12922 10848
rect 17606 10912 17922 10913
rect 17606 10848 17612 10912
rect 17676 10848 17692 10912
rect 17756 10848 17772 10912
rect 17836 10848 17852 10912
rect 17916 10848 17922 10912
rect 17606 10847 17922 10848
rect 2589 10706 2655 10709
rect 6126 10706 6132 10708
rect 2589 10704 6132 10706
rect 2589 10648 2594 10704
rect 2650 10648 6132 10704
rect 2589 10646 6132 10648
rect 2589 10643 2655 10646
rect 6126 10644 6132 10646
rect 6196 10644 6202 10708
rect 7925 10570 7991 10573
rect 15142 10570 15148 10572
rect 7925 10568 15148 10570
rect 7925 10512 7930 10568
rect 7986 10512 15148 10568
rect 7925 10510 15148 10512
rect 7925 10507 7991 10510
rect 15142 10508 15148 10510
rect 15212 10508 15218 10572
rect 18229 10434 18295 10437
rect 19200 10434 20000 10464
rect 18229 10432 20000 10434
rect 18229 10376 18234 10432
rect 18290 10376 20000 10432
rect 18229 10374 20000 10376
rect 18229 10371 18295 10374
rect 1946 10368 2262 10369
rect 1946 10304 1952 10368
rect 2016 10304 2032 10368
rect 2096 10304 2112 10368
rect 2176 10304 2192 10368
rect 2256 10304 2262 10368
rect 1946 10303 2262 10304
rect 6946 10368 7262 10369
rect 6946 10304 6952 10368
rect 7016 10304 7032 10368
rect 7096 10304 7112 10368
rect 7176 10304 7192 10368
rect 7256 10304 7262 10368
rect 6946 10303 7262 10304
rect 11946 10368 12262 10369
rect 11946 10304 11952 10368
rect 12016 10304 12032 10368
rect 12096 10304 12112 10368
rect 12176 10304 12192 10368
rect 12256 10304 12262 10368
rect 11946 10303 12262 10304
rect 16946 10368 17262 10369
rect 16946 10304 16952 10368
rect 17016 10304 17032 10368
rect 17096 10304 17112 10368
rect 17176 10304 17192 10368
rect 17256 10304 17262 10368
rect 19200 10344 20000 10374
rect 16946 10303 17262 10304
rect 3182 9964 3188 10028
rect 3252 10026 3258 10028
rect 7005 10026 7071 10029
rect 3252 10024 7071 10026
rect 3252 9968 7010 10024
rect 7066 9968 7071 10024
rect 3252 9966 7071 9968
rect 3252 9964 3258 9966
rect 7005 9963 7071 9966
rect 2606 9824 2922 9825
rect 2606 9760 2612 9824
rect 2676 9760 2692 9824
rect 2756 9760 2772 9824
rect 2836 9760 2852 9824
rect 2916 9760 2922 9824
rect 2606 9759 2922 9760
rect 7606 9824 7922 9825
rect 7606 9760 7612 9824
rect 7676 9760 7692 9824
rect 7756 9760 7772 9824
rect 7836 9760 7852 9824
rect 7916 9760 7922 9824
rect 7606 9759 7922 9760
rect 12606 9824 12922 9825
rect 12606 9760 12612 9824
rect 12676 9760 12692 9824
rect 12756 9760 12772 9824
rect 12836 9760 12852 9824
rect 12916 9760 12922 9824
rect 12606 9759 12922 9760
rect 17606 9824 17922 9825
rect 17606 9760 17612 9824
rect 17676 9760 17692 9824
rect 17756 9760 17772 9824
rect 17836 9760 17852 9824
rect 17916 9760 17922 9824
rect 17606 9759 17922 9760
rect 6637 9620 6703 9621
rect 6637 9618 6684 9620
rect 6592 9616 6684 9618
rect 6592 9560 6642 9616
rect 6592 9558 6684 9560
rect 6637 9556 6684 9558
rect 6748 9556 6754 9620
rect 6637 9555 6703 9556
rect 1946 9280 2262 9281
rect 1946 9216 1952 9280
rect 2016 9216 2032 9280
rect 2096 9216 2112 9280
rect 2176 9216 2192 9280
rect 2256 9216 2262 9280
rect 1946 9215 2262 9216
rect 6946 9280 7262 9281
rect 6946 9216 6952 9280
rect 7016 9216 7032 9280
rect 7096 9216 7112 9280
rect 7176 9216 7192 9280
rect 7256 9216 7262 9280
rect 6946 9215 7262 9216
rect 11946 9280 12262 9281
rect 11946 9216 11952 9280
rect 12016 9216 12032 9280
rect 12096 9216 12112 9280
rect 12176 9216 12192 9280
rect 12256 9216 12262 9280
rect 11946 9215 12262 9216
rect 16946 9280 17262 9281
rect 16946 9216 16952 9280
rect 17016 9216 17032 9280
rect 17096 9216 17112 9280
rect 17176 9216 17192 9280
rect 17256 9216 17262 9280
rect 16946 9215 17262 9216
rect 2606 8736 2922 8737
rect 2606 8672 2612 8736
rect 2676 8672 2692 8736
rect 2756 8672 2772 8736
rect 2836 8672 2852 8736
rect 2916 8672 2922 8736
rect 2606 8671 2922 8672
rect 7606 8736 7922 8737
rect 7606 8672 7612 8736
rect 7676 8672 7692 8736
rect 7756 8672 7772 8736
rect 7836 8672 7852 8736
rect 7916 8672 7922 8736
rect 7606 8671 7922 8672
rect 12606 8736 12922 8737
rect 12606 8672 12612 8736
rect 12676 8672 12692 8736
rect 12756 8672 12772 8736
rect 12836 8672 12852 8736
rect 12916 8672 12922 8736
rect 12606 8671 12922 8672
rect 17606 8736 17922 8737
rect 17606 8672 17612 8736
rect 17676 8672 17692 8736
rect 17756 8672 17772 8736
rect 17836 8672 17852 8736
rect 17916 8672 17922 8736
rect 17606 8671 17922 8672
rect 18229 8530 18295 8533
rect 19200 8530 20000 8560
rect 18229 8528 20000 8530
rect 18229 8472 18234 8528
rect 18290 8472 20000 8528
rect 18229 8470 20000 8472
rect 18229 8467 18295 8470
rect 19200 8440 20000 8470
rect 14181 8260 14247 8261
rect 14181 8256 14228 8260
rect 14292 8258 14298 8260
rect 14181 8200 14186 8256
rect 14181 8196 14228 8200
rect 14292 8198 14338 8258
rect 14292 8196 14298 8198
rect 14181 8195 14247 8196
rect 1946 8192 2262 8193
rect 1946 8128 1952 8192
rect 2016 8128 2032 8192
rect 2096 8128 2112 8192
rect 2176 8128 2192 8192
rect 2256 8128 2262 8192
rect 1946 8127 2262 8128
rect 6946 8192 7262 8193
rect 6946 8128 6952 8192
rect 7016 8128 7032 8192
rect 7096 8128 7112 8192
rect 7176 8128 7192 8192
rect 7256 8128 7262 8192
rect 6946 8127 7262 8128
rect 11946 8192 12262 8193
rect 11946 8128 11952 8192
rect 12016 8128 12032 8192
rect 12096 8128 12112 8192
rect 12176 8128 12192 8192
rect 12256 8128 12262 8192
rect 11946 8127 12262 8128
rect 16946 8192 17262 8193
rect 16946 8128 16952 8192
rect 17016 8128 17032 8192
rect 17096 8128 17112 8192
rect 17176 8128 17192 8192
rect 17256 8128 17262 8192
rect 16946 8127 17262 8128
rect 9438 8060 9444 8124
rect 9508 8122 9514 8124
rect 11513 8122 11579 8125
rect 9508 8120 11579 8122
rect 9508 8064 11518 8120
rect 11574 8064 11579 8120
rect 9508 8062 11579 8064
rect 9508 8060 9514 8062
rect 11513 8059 11579 8062
rect 12249 7986 12315 7989
rect 16614 7986 16620 7988
rect 12249 7984 16620 7986
rect 12249 7928 12254 7984
rect 12310 7928 16620 7984
rect 12249 7926 16620 7928
rect 12249 7923 12315 7926
rect 16614 7924 16620 7926
rect 16684 7924 16690 7988
rect 2606 7648 2922 7649
rect 2606 7584 2612 7648
rect 2676 7584 2692 7648
rect 2756 7584 2772 7648
rect 2836 7584 2852 7648
rect 2916 7584 2922 7648
rect 2606 7583 2922 7584
rect 7606 7648 7922 7649
rect 7606 7584 7612 7648
rect 7676 7584 7692 7648
rect 7756 7584 7772 7648
rect 7836 7584 7852 7648
rect 7916 7584 7922 7648
rect 7606 7583 7922 7584
rect 12606 7648 12922 7649
rect 12606 7584 12612 7648
rect 12676 7584 12692 7648
rect 12756 7584 12772 7648
rect 12836 7584 12852 7648
rect 12916 7584 12922 7648
rect 12606 7583 12922 7584
rect 17606 7648 17922 7649
rect 17606 7584 17612 7648
rect 17676 7584 17692 7648
rect 17756 7584 17772 7648
rect 17836 7584 17852 7648
rect 17916 7584 17922 7648
rect 17606 7583 17922 7584
rect 4654 7244 4660 7308
rect 4724 7306 4730 7308
rect 13813 7306 13879 7309
rect 4724 7304 13879 7306
rect 4724 7248 13818 7304
rect 13874 7248 13879 7304
rect 4724 7246 13879 7248
rect 4724 7244 4730 7246
rect 13813 7243 13879 7246
rect 1946 7104 2262 7105
rect 1946 7040 1952 7104
rect 2016 7040 2032 7104
rect 2096 7040 2112 7104
rect 2176 7040 2192 7104
rect 2256 7040 2262 7104
rect 1946 7039 2262 7040
rect 6946 7104 7262 7105
rect 6946 7040 6952 7104
rect 7016 7040 7032 7104
rect 7096 7040 7112 7104
rect 7176 7040 7192 7104
rect 7256 7040 7262 7104
rect 6946 7039 7262 7040
rect 11946 7104 12262 7105
rect 11946 7040 11952 7104
rect 12016 7040 12032 7104
rect 12096 7040 12112 7104
rect 12176 7040 12192 7104
rect 12256 7040 12262 7104
rect 11946 7039 12262 7040
rect 16946 7104 17262 7105
rect 16946 7040 16952 7104
rect 17016 7040 17032 7104
rect 17096 7040 17112 7104
rect 17176 7040 17192 7104
rect 17256 7040 17262 7104
rect 16946 7039 17262 7040
rect 7373 6898 7439 6901
rect 8150 6898 8156 6900
rect 7373 6896 8156 6898
rect 7373 6840 7378 6896
rect 7434 6840 8156 6896
rect 7373 6838 8156 6840
rect 7373 6835 7439 6838
rect 8150 6836 8156 6838
rect 8220 6836 8226 6900
rect 12709 6898 12775 6901
rect 13353 6900 13419 6901
rect 13302 6898 13308 6900
rect 8342 6838 12450 6898
rect 6913 6762 6979 6765
rect 8342 6762 8402 6838
rect 6913 6760 8402 6762
rect 6913 6704 6918 6760
rect 6974 6704 8402 6760
rect 6913 6702 8402 6704
rect 9673 6762 9739 6765
rect 9806 6762 9812 6764
rect 9673 6760 9812 6762
rect 9673 6704 9678 6760
rect 9734 6704 9812 6760
rect 9673 6702 9812 6704
rect 6913 6699 6979 6702
rect 9673 6699 9739 6702
rect 9806 6700 9812 6702
rect 9876 6700 9882 6764
rect 12390 6762 12450 6838
rect 12709 6896 13308 6898
rect 13372 6898 13419 6900
rect 13372 6896 13500 6898
rect 12709 6840 12714 6896
rect 12770 6840 13308 6896
rect 13414 6840 13500 6896
rect 12709 6838 13308 6840
rect 12709 6835 12775 6838
rect 13302 6836 13308 6838
rect 13372 6838 13500 6840
rect 13372 6836 13419 6838
rect 13353 6835 13419 6836
rect 16062 6762 16068 6764
rect 12390 6702 16068 6762
rect 16062 6700 16068 6702
rect 16132 6700 16138 6764
rect 18229 6626 18295 6629
rect 19200 6626 20000 6656
rect 18229 6624 20000 6626
rect 18229 6568 18234 6624
rect 18290 6568 20000 6624
rect 18229 6566 20000 6568
rect 18229 6563 18295 6566
rect 2606 6560 2922 6561
rect 2606 6496 2612 6560
rect 2676 6496 2692 6560
rect 2756 6496 2772 6560
rect 2836 6496 2852 6560
rect 2916 6496 2922 6560
rect 2606 6495 2922 6496
rect 7606 6560 7922 6561
rect 7606 6496 7612 6560
rect 7676 6496 7692 6560
rect 7756 6496 7772 6560
rect 7836 6496 7852 6560
rect 7916 6496 7922 6560
rect 7606 6495 7922 6496
rect 12606 6560 12922 6561
rect 12606 6496 12612 6560
rect 12676 6496 12692 6560
rect 12756 6496 12772 6560
rect 12836 6496 12852 6560
rect 12916 6496 12922 6560
rect 12606 6495 12922 6496
rect 17606 6560 17922 6561
rect 17606 6496 17612 6560
rect 17676 6496 17692 6560
rect 17756 6496 17772 6560
rect 17836 6496 17852 6560
rect 17916 6496 17922 6560
rect 19200 6536 20000 6566
rect 17606 6495 17922 6496
rect 1946 6016 2262 6017
rect 1946 5952 1952 6016
rect 2016 5952 2032 6016
rect 2096 5952 2112 6016
rect 2176 5952 2192 6016
rect 2256 5952 2262 6016
rect 1946 5951 2262 5952
rect 6946 6016 7262 6017
rect 6946 5952 6952 6016
rect 7016 5952 7032 6016
rect 7096 5952 7112 6016
rect 7176 5952 7192 6016
rect 7256 5952 7262 6016
rect 6946 5951 7262 5952
rect 11946 6016 12262 6017
rect 11946 5952 11952 6016
rect 12016 5952 12032 6016
rect 12096 5952 12112 6016
rect 12176 5952 12192 6016
rect 12256 5952 12262 6016
rect 11946 5951 12262 5952
rect 16946 6016 17262 6017
rect 16946 5952 16952 6016
rect 17016 5952 17032 6016
rect 17096 5952 17112 6016
rect 17176 5952 17192 6016
rect 17256 5952 17262 6016
rect 16946 5951 17262 5952
rect 2606 5472 2922 5473
rect 2606 5408 2612 5472
rect 2676 5408 2692 5472
rect 2756 5408 2772 5472
rect 2836 5408 2852 5472
rect 2916 5408 2922 5472
rect 2606 5407 2922 5408
rect 7606 5472 7922 5473
rect 7606 5408 7612 5472
rect 7676 5408 7692 5472
rect 7756 5408 7772 5472
rect 7836 5408 7852 5472
rect 7916 5408 7922 5472
rect 7606 5407 7922 5408
rect 12606 5472 12922 5473
rect 12606 5408 12612 5472
rect 12676 5408 12692 5472
rect 12756 5408 12772 5472
rect 12836 5408 12852 5472
rect 12916 5408 12922 5472
rect 12606 5407 12922 5408
rect 17606 5472 17922 5473
rect 17606 5408 17612 5472
rect 17676 5408 17692 5472
rect 17756 5408 17772 5472
rect 17836 5408 17852 5472
rect 17916 5408 17922 5472
rect 17606 5407 17922 5408
rect 10910 5204 10916 5268
rect 10980 5266 10986 5268
rect 16205 5266 16271 5269
rect 10980 5264 16271 5266
rect 10980 5208 16210 5264
rect 16266 5208 16271 5264
rect 10980 5206 16271 5208
rect 10980 5204 10986 5206
rect 16205 5203 16271 5206
rect 1946 4928 2262 4929
rect 1946 4864 1952 4928
rect 2016 4864 2032 4928
rect 2096 4864 2112 4928
rect 2176 4864 2192 4928
rect 2256 4864 2262 4928
rect 1946 4863 2262 4864
rect 6946 4928 7262 4929
rect 6946 4864 6952 4928
rect 7016 4864 7032 4928
rect 7096 4864 7112 4928
rect 7176 4864 7192 4928
rect 7256 4864 7262 4928
rect 6946 4863 7262 4864
rect 11946 4928 12262 4929
rect 11946 4864 11952 4928
rect 12016 4864 12032 4928
rect 12096 4864 12112 4928
rect 12176 4864 12192 4928
rect 12256 4864 12262 4928
rect 11946 4863 12262 4864
rect 16946 4928 17262 4929
rect 16946 4864 16952 4928
rect 17016 4864 17032 4928
rect 17096 4864 17112 4928
rect 17176 4864 17192 4928
rect 17256 4864 17262 4928
rect 16946 4863 17262 4864
rect 18229 4722 18295 4725
rect 19200 4722 20000 4752
rect 18229 4720 20000 4722
rect 18229 4664 18234 4720
rect 18290 4664 20000 4720
rect 18229 4662 20000 4664
rect 18229 4659 18295 4662
rect 19200 4632 20000 4662
rect 2606 4384 2922 4385
rect 2606 4320 2612 4384
rect 2676 4320 2692 4384
rect 2756 4320 2772 4384
rect 2836 4320 2852 4384
rect 2916 4320 2922 4384
rect 2606 4319 2922 4320
rect 7606 4384 7922 4385
rect 7606 4320 7612 4384
rect 7676 4320 7692 4384
rect 7756 4320 7772 4384
rect 7836 4320 7852 4384
rect 7916 4320 7922 4384
rect 7606 4319 7922 4320
rect 12606 4384 12922 4385
rect 12606 4320 12612 4384
rect 12676 4320 12692 4384
rect 12756 4320 12772 4384
rect 12836 4320 12852 4384
rect 12916 4320 12922 4384
rect 12606 4319 12922 4320
rect 17606 4384 17922 4385
rect 17606 4320 17612 4384
rect 17676 4320 17692 4384
rect 17756 4320 17772 4384
rect 17836 4320 17852 4384
rect 17916 4320 17922 4384
rect 17606 4319 17922 4320
rect 1946 3840 2262 3841
rect 1946 3776 1952 3840
rect 2016 3776 2032 3840
rect 2096 3776 2112 3840
rect 2176 3776 2192 3840
rect 2256 3776 2262 3840
rect 1946 3775 2262 3776
rect 6946 3840 7262 3841
rect 6946 3776 6952 3840
rect 7016 3776 7032 3840
rect 7096 3776 7112 3840
rect 7176 3776 7192 3840
rect 7256 3776 7262 3840
rect 6946 3775 7262 3776
rect 11946 3840 12262 3841
rect 11946 3776 11952 3840
rect 12016 3776 12032 3840
rect 12096 3776 12112 3840
rect 12176 3776 12192 3840
rect 12256 3776 12262 3840
rect 11946 3775 12262 3776
rect 16946 3840 17262 3841
rect 16946 3776 16952 3840
rect 17016 3776 17032 3840
rect 17096 3776 17112 3840
rect 17176 3776 17192 3840
rect 17256 3776 17262 3840
rect 16946 3775 17262 3776
rect 2606 3296 2922 3297
rect 2606 3232 2612 3296
rect 2676 3232 2692 3296
rect 2756 3232 2772 3296
rect 2836 3232 2852 3296
rect 2916 3232 2922 3296
rect 2606 3231 2922 3232
rect 7606 3296 7922 3297
rect 7606 3232 7612 3296
rect 7676 3232 7692 3296
rect 7756 3232 7772 3296
rect 7836 3232 7852 3296
rect 7916 3232 7922 3296
rect 7606 3231 7922 3232
rect 12606 3296 12922 3297
rect 12606 3232 12612 3296
rect 12676 3232 12692 3296
rect 12756 3232 12772 3296
rect 12836 3232 12852 3296
rect 12916 3232 12922 3296
rect 12606 3231 12922 3232
rect 17606 3296 17922 3297
rect 17606 3232 17612 3296
rect 17676 3232 17692 3296
rect 17756 3232 17772 3296
rect 17836 3232 17852 3296
rect 17916 3232 17922 3296
rect 17606 3231 17922 3232
rect 18229 2818 18295 2821
rect 19200 2818 20000 2848
rect 18229 2816 20000 2818
rect 18229 2760 18234 2816
rect 18290 2760 20000 2816
rect 18229 2758 20000 2760
rect 18229 2755 18295 2758
rect 1946 2752 2262 2753
rect 1946 2688 1952 2752
rect 2016 2688 2032 2752
rect 2096 2688 2112 2752
rect 2176 2688 2192 2752
rect 2256 2688 2262 2752
rect 1946 2687 2262 2688
rect 6946 2752 7262 2753
rect 6946 2688 6952 2752
rect 7016 2688 7032 2752
rect 7096 2688 7112 2752
rect 7176 2688 7192 2752
rect 7256 2688 7262 2752
rect 6946 2687 7262 2688
rect 11946 2752 12262 2753
rect 11946 2688 11952 2752
rect 12016 2688 12032 2752
rect 12096 2688 12112 2752
rect 12176 2688 12192 2752
rect 12256 2688 12262 2752
rect 11946 2687 12262 2688
rect 16946 2752 17262 2753
rect 16946 2688 16952 2752
rect 17016 2688 17032 2752
rect 17096 2688 17112 2752
rect 17176 2688 17192 2752
rect 17256 2688 17262 2752
rect 19200 2728 20000 2758
rect 16946 2687 17262 2688
rect 2606 2208 2922 2209
rect 2606 2144 2612 2208
rect 2676 2144 2692 2208
rect 2756 2144 2772 2208
rect 2836 2144 2852 2208
rect 2916 2144 2922 2208
rect 2606 2143 2922 2144
rect 7606 2208 7922 2209
rect 7606 2144 7612 2208
rect 7676 2144 7692 2208
rect 7756 2144 7772 2208
rect 7836 2144 7852 2208
rect 7916 2144 7922 2208
rect 7606 2143 7922 2144
rect 12606 2208 12922 2209
rect 12606 2144 12612 2208
rect 12676 2144 12692 2208
rect 12756 2144 12772 2208
rect 12836 2144 12852 2208
rect 12916 2144 12922 2208
rect 12606 2143 12922 2144
rect 17606 2208 17922 2209
rect 17606 2144 17612 2208
rect 17676 2144 17692 2208
rect 17756 2144 17772 2208
rect 17836 2144 17852 2208
rect 17916 2144 17922 2208
rect 17606 2143 17922 2144
<< via3 >>
rect 1952 77820 2016 77824
rect 1952 77764 1956 77820
rect 1956 77764 2012 77820
rect 2012 77764 2016 77820
rect 1952 77760 2016 77764
rect 2032 77820 2096 77824
rect 2032 77764 2036 77820
rect 2036 77764 2092 77820
rect 2092 77764 2096 77820
rect 2032 77760 2096 77764
rect 2112 77820 2176 77824
rect 2112 77764 2116 77820
rect 2116 77764 2172 77820
rect 2172 77764 2176 77820
rect 2112 77760 2176 77764
rect 2192 77820 2256 77824
rect 2192 77764 2196 77820
rect 2196 77764 2252 77820
rect 2252 77764 2256 77820
rect 2192 77760 2256 77764
rect 6952 77820 7016 77824
rect 6952 77764 6956 77820
rect 6956 77764 7012 77820
rect 7012 77764 7016 77820
rect 6952 77760 7016 77764
rect 7032 77820 7096 77824
rect 7032 77764 7036 77820
rect 7036 77764 7092 77820
rect 7092 77764 7096 77820
rect 7032 77760 7096 77764
rect 7112 77820 7176 77824
rect 7112 77764 7116 77820
rect 7116 77764 7172 77820
rect 7172 77764 7176 77820
rect 7112 77760 7176 77764
rect 7192 77820 7256 77824
rect 7192 77764 7196 77820
rect 7196 77764 7252 77820
rect 7252 77764 7256 77820
rect 7192 77760 7256 77764
rect 11952 77820 12016 77824
rect 11952 77764 11956 77820
rect 11956 77764 12012 77820
rect 12012 77764 12016 77820
rect 11952 77760 12016 77764
rect 12032 77820 12096 77824
rect 12032 77764 12036 77820
rect 12036 77764 12092 77820
rect 12092 77764 12096 77820
rect 12032 77760 12096 77764
rect 12112 77820 12176 77824
rect 12112 77764 12116 77820
rect 12116 77764 12172 77820
rect 12172 77764 12176 77820
rect 12112 77760 12176 77764
rect 12192 77820 12256 77824
rect 12192 77764 12196 77820
rect 12196 77764 12252 77820
rect 12252 77764 12256 77820
rect 12192 77760 12256 77764
rect 16952 77820 17016 77824
rect 16952 77764 16956 77820
rect 16956 77764 17012 77820
rect 17012 77764 17016 77820
rect 16952 77760 17016 77764
rect 17032 77820 17096 77824
rect 17032 77764 17036 77820
rect 17036 77764 17092 77820
rect 17092 77764 17096 77820
rect 17032 77760 17096 77764
rect 17112 77820 17176 77824
rect 17112 77764 17116 77820
rect 17116 77764 17172 77820
rect 17172 77764 17176 77820
rect 17112 77760 17176 77764
rect 17192 77820 17256 77824
rect 17192 77764 17196 77820
rect 17196 77764 17252 77820
rect 17252 77764 17256 77820
rect 17192 77760 17256 77764
rect 2612 77276 2676 77280
rect 2612 77220 2616 77276
rect 2616 77220 2672 77276
rect 2672 77220 2676 77276
rect 2612 77216 2676 77220
rect 2692 77276 2756 77280
rect 2692 77220 2696 77276
rect 2696 77220 2752 77276
rect 2752 77220 2756 77276
rect 2692 77216 2756 77220
rect 2772 77276 2836 77280
rect 2772 77220 2776 77276
rect 2776 77220 2832 77276
rect 2832 77220 2836 77276
rect 2772 77216 2836 77220
rect 2852 77276 2916 77280
rect 2852 77220 2856 77276
rect 2856 77220 2912 77276
rect 2912 77220 2916 77276
rect 2852 77216 2916 77220
rect 7612 77276 7676 77280
rect 7612 77220 7616 77276
rect 7616 77220 7672 77276
rect 7672 77220 7676 77276
rect 7612 77216 7676 77220
rect 7692 77276 7756 77280
rect 7692 77220 7696 77276
rect 7696 77220 7752 77276
rect 7752 77220 7756 77276
rect 7692 77216 7756 77220
rect 7772 77276 7836 77280
rect 7772 77220 7776 77276
rect 7776 77220 7832 77276
rect 7832 77220 7836 77276
rect 7772 77216 7836 77220
rect 7852 77276 7916 77280
rect 7852 77220 7856 77276
rect 7856 77220 7912 77276
rect 7912 77220 7916 77276
rect 7852 77216 7916 77220
rect 12612 77276 12676 77280
rect 12612 77220 12616 77276
rect 12616 77220 12672 77276
rect 12672 77220 12676 77276
rect 12612 77216 12676 77220
rect 12692 77276 12756 77280
rect 12692 77220 12696 77276
rect 12696 77220 12752 77276
rect 12752 77220 12756 77276
rect 12692 77216 12756 77220
rect 12772 77276 12836 77280
rect 12772 77220 12776 77276
rect 12776 77220 12832 77276
rect 12832 77220 12836 77276
rect 12772 77216 12836 77220
rect 12852 77276 12916 77280
rect 12852 77220 12856 77276
rect 12856 77220 12912 77276
rect 12912 77220 12916 77276
rect 12852 77216 12916 77220
rect 17612 77276 17676 77280
rect 17612 77220 17616 77276
rect 17616 77220 17672 77276
rect 17672 77220 17676 77276
rect 17612 77216 17676 77220
rect 17692 77276 17756 77280
rect 17692 77220 17696 77276
rect 17696 77220 17752 77276
rect 17752 77220 17756 77276
rect 17692 77216 17756 77220
rect 17772 77276 17836 77280
rect 17772 77220 17776 77276
rect 17776 77220 17832 77276
rect 17832 77220 17836 77276
rect 17772 77216 17836 77220
rect 17852 77276 17916 77280
rect 17852 77220 17856 77276
rect 17856 77220 17912 77276
rect 17912 77220 17916 77276
rect 17852 77216 17916 77220
rect 14596 76800 14660 76804
rect 14596 76744 14646 76800
rect 14646 76744 14660 76800
rect 14596 76740 14660 76744
rect 15884 76800 15948 76804
rect 15884 76744 15934 76800
rect 15934 76744 15948 76800
rect 15884 76740 15948 76744
rect 1952 76732 2016 76736
rect 1952 76676 1956 76732
rect 1956 76676 2012 76732
rect 2012 76676 2016 76732
rect 1952 76672 2016 76676
rect 2032 76732 2096 76736
rect 2032 76676 2036 76732
rect 2036 76676 2092 76732
rect 2092 76676 2096 76732
rect 2032 76672 2096 76676
rect 2112 76732 2176 76736
rect 2112 76676 2116 76732
rect 2116 76676 2172 76732
rect 2172 76676 2176 76732
rect 2112 76672 2176 76676
rect 2192 76732 2256 76736
rect 2192 76676 2196 76732
rect 2196 76676 2252 76732
rect 2252 76676 2256 76732
rect 2192 76672 2256 76676
rect 6952 76732 7016 76736
rect 6952 76676 6956 76732
rect 6956 76676 7012 76732
rect 7012 76676 7016 76732
rect 6952 76672 7016 76676
rect 7032 76732 7096 76736
rect 7032 76676 7036 76732
rect 7036 76676 7092 76732
rect 7092 76676 7096 76732
rect 7032 76672 7096 76676
rect 7112 76732 7176 76736
rect 7112 76676 7116 76732
rect 7116 76676 7172 76732
rect 7172 76676 7176 76732
rect 7112 76672 7176 76676
rect 7192 76732 7256 76736
rect 7192 76676 7196 76732
rect 7196 76676 7252 76732
rect 7252 76676 7256 76732
rect 7192 76672 7256 76676
rect 11952 76732 12016 76736
rect 11952 76676 11956 76732
rect 11956 76676 12012 76732
rect 12012 76676 12016 76732
rect 11952 76672 12016 76676
rect 12032 76732 12096 76736
rect 12032 76676 12036 76732
rect 12036 76676 12092 76732
rect 12092 76676 12096 76732
rect 12032 76672 12096 76676
rect 12112 76732 12176 76736
rect 12112 76676 12116 76732
rect 12116 76676 12172 76732
rect 12172 76676 12176 76732
rect 12112 76672 12176 76676
rect 12192 76732 12256 76736
rect 12192 76676 12196 76732
rect 12196 76676 12252 76732
rect 12252 76676 12256 76732
rect 12192 76672 12256 76676
rect 16952 76732 17016 76736
rect 16952 76676 16956 76732
rect 16956 76676 17012 76732
rect 17012 76676 17016 76732
rect 16952 76672 17016 76676
rect 17032 76732 17096 76736
rect 17032 76676 17036 76732
rect 17036 76676 17092 76732
rect 17092 76676 17096 76732
rect 17032 76672 17096 76676
rect 17112 76732 17176 76736
rect 17112 76676 17116 76732
rect 17116 76676 17172 76732
rect 17172 76676 17176 76732
rect 17112 76672 17176 76676
rect 17192 76732 17256 76736
rect 17192 76676 17196 76732
rect 17196 76676 17252 76732
rect 17252 76676 17256 76732
rect 17192 76672 17256 76676
rect 6132 76332 6196 76396
rect 11284 76256 11348 76260
rect 11284 76200 11298 76256
rect 11298 76200 11348 76256
rect 11284 76196 11348 76200
rect 2612 76188 2676 76192
rect 2612 76132 2616 76188
rect 2616 76132 2672 76188
rect 2672 76132 2676 76188
rect 2612 76128 2676 76132
rect 2692 76188 2756 76192
rect 2692 76132 2696 76188
rect 2696 76132 2752 76188
rect 2752 76132 2756 76188
rect 2692 76128 2756 76132
rect 2772 76188 2836 76192
rect 2772 76132 2776 76188
rect 2776 76132 2832 76188
rect 2832 76132 2836 76188
rect 2772 76128 2836 76132
rect 2852 76188 2916 76192
rect 2852 76132 2856 76188
rect 2856 76132 2912 76188
rect 2912 76132 2916 76188
rect 2852 76128 2916 76132
rect 7612 76188 7676 76192
rect 7612 76132 7616 76188
rect 7616 76132 7672 76188
rect 7672 76132 7676 76188
rect 7612 76128 7676 76132
rect 7692 76188 7756 76192
rect 7692 76132 7696 76188
rect 7696 76132 7752 76188
rect 7752 76132 7756 76188
rect 7692 76128 7756 76132
rect 7772 76188 7836 76192
rect 7772 76132 7776 76188
rect 7776 76132 7832 76188
rect 7832 76132 7836 76188
rect 7772 76128 7836 76132
rect 7852 76188 7916 76192
rect 7852 76132 7856 76188
rect 7856 76132 7912 76188
rect 7912 76132 7916 76188
rect 7852 76128 7916 76132
rect 12612 76188 12676 76192
rect 12612 76132 12616 76188
rect 12616 76132 12672 76188
rect 12672 76132 12676 76188
rect 12612 76128 12676 76132
rect 12692 76188 12756 76192
rect 12692 76132 12696 76188
rect 12696 76132 12752 76188
rect 12752 76132 12756 76188
rect 12692 76128 12756 76132
rect 12772 76188 12836 76192
rect 12772 76132 12776 76188
rect 12776 76132 12832 76188
rect 12832 76132 12836 76188
rect 12772 76128 12836 76132
rect 12852 76188 12916 76192
rect 12852 76132 12856 76188
rect 12856 76132 12912 76188
rect 12912 76132 12916 76188
rect 12852 76128 12916 76132
rect 17612 76188 17676 76192
rect 17612 76132 17616 76188
rect 17616 76132 17672 76188
rect 17672 76132 17676 76188
rect 17612 76128 17676 76132
rect 17692 76188 17756 76192
rect 17692 76132 17696 76188
rect 17696 76132 17752 76188
rect 17752 76132 17756 76188
rect 17692 76128 17756 76132
rect 17772 76188 17836 76192
rect 17772 76132 17776 76188
rect 17776 76132 17832 76188
rect 17832 76132 17836 76188
rect 17772 76128 17836 76132
rect 17852 76188 17916 76192
rect 17852 76132 17856 76188
rect 17856 76132 17912 76188
rect 17912 76132 17916 76188
rect 17852 76128 17916 76132
rect 8892 76060 8956 76124
rect 14228 75924 14292 75988
rect 1952 75644 2016 75648
rect 1952 75588 1956 75644
rect 1956 75588 2012 75644
rect 2012 75588 2016 75644
rect 1952 75584 2016 75588
rect 2032 75644 2096 75648
rect 2032 75588 2036 75644
rect 2036 75588 2092 75644
rect 2092 75588 2096 75644
rect 2032 75584 2096 75588
rect 2112 75644 2176 75648
rect 2112 75588 2116 75644
rect 2116 75588 2172 75644
rect 2172 75588 2176 75644
rect 2112 75584 2176 75588
rect 2192 75644 2256 75648
rect 2192 75588 2196 75644
rect 2196 75588 2252 75644
rect 2252 75588 2256 75644
rect 2192 75584 2256 75588
rect 6952 75644 7016 75648
rect 6952 75588 6956 75644
rect 6956 75588 7012 75644
rect 7012 75588 7016 75644
rect 6952 75584 7016 75588
rect 7032 75644 7096 75648
rect 7032 75588 7036 75644
rect 7036 75588 7092 75644
rect 7092 75588 7096 75644
rect 7032 75584 7096 75588
rect 7112 75644 7176 75648
rect 7112 75588 7116 75644
rect 7116 75588 7172 75644
rect 7172 75588 7176 75644
rect 7112 75584 7176 75588
rect 7192 75644 7256 75648
rect 7192 75588 7196 75644
rect 7196 75588 7252 75644
rect 7252 75588 7256 75644
rect 7192 75584 7256 75588
rect 11952 75644 12016 75648
rect 11952 75588 11956 75644
rect 11956 75588 12012 75644
rect 12012 75588 12016 75644
rect 11952 75584 12016 75588
rect 12032 75644 12096 75648
rect 12032 75588 12036 75644
rect 12036 75588 12092 75644
rect 12092 75588 12096 75644
rect 12032 75584 12096 75588
rect 12112 75644 12176 75648
rect 12112 75588 12116 75644
rect 12116 75588 12172 75644
rect 12172 75588 12176 75644
rect 12112 75584 12176 75588
rect 12192 75644 12256 75648
rect 12192 75588 12196 75644
rect 12196 75588 12252 75644
rect 12252 75588 12256 75644
rect 12192 75584 12256 75588
rect 16952 75644 17016 75648
rect 16952 75588 16956 75644
rect 16956 75588 17012 75644
rect 17012 75588 17016 75644
rect 16952 75584 17016 75588
rect 17032 75644 17096 75648
rect 17032 75588 17036 75644
rect 17036 75588 17092 75644
rect 17092 75588 17096 75644
rect 17032 75584 17096 75588
rect 17112 75644 17176 75648
rect 17112 75588 17116 75644
rect 17116 75588 17172 75644
rect 17172 75588 17176 75644
rect 17112 75584 17176 75588
rect 17192 75644 17256 75648
rect 17192 75588 17196 75644
rect 17196 75588 17252 75644
rect 17252 75588 17256 75644
rect 17192 75584 17256 75588
rect 6684 75108 6748 75172
rect 2612 75100 2676 75104
rect 2612 75044 2616 75100
rect 2616 75044 2672 75100
rect 2672 75044 2676 75100
rect 2612 75040 2676 75044
rect 2692 75100 2756 75104
rect 2692 75044 2696 75100
rect 2696 75044 2752 75100
rect 2752 75044 2756 75100
rect 2692 75040 2756 75044
rect 2772 75100 2836 75104
rect 2772 75044 2776 75100
rect 2776 75044 2832 75100
rect 2832 75044 2836 75100
rect 2772 75040 2836 75044
rect 2852 75100 2916 75104
rect 2852 75044 2856 75100
rect 2856 75044 2912 75100
rect 2912 75044 2916 75100
rect 2852 75040 2916 75044
rect 7612 75100 7676 75104
rect 7612 75044 7616 75100
rect 7616 75044 7672 75100
rect 7672 75044 7676 75100
rect 7612 75040 7676 75044
rect 7692 75100 7756 75104
rect 7692 75044 7696 75100
rect 7696 75044 7752 75100
rect 7752 75044 7756 75100
rect 7692 75040 7756 75044
rect 7772 75100 7836 75104
rect 7772 75044 7776 75100
rect 7776 75044 7832 75100
rect 7832 75044 7836 75100
rect 7772 75040 7836 75044
rect 7852 75100 7916 75104
rect 7852 75044 7856 75100
rect 7856 75044 7912 75100
rect 7912 75044 7916 75100
rect 7852 75040 7916 75044
rect 12612 75100 12676 75104
rect 12612 75044 12616 75100
rect 12616 75044 12672 75100
rect 12672 75044 12676 75100
rect 12612 75040 12676 75044
rect 12692 75100 12756 75104
rect 12692 75044 12696 75100
rect 12696 75044 12752 75100
rect 12752 75044 12756 75100
rect 12692 75040 12756 75044
rect 12772 75100 12836 75104
rect 12772 75044 12776 75100
rect 12776 75044 12832 75100
rect 12832 75044 12836 75100
rect 12772 75040 12836 75044
rect 12852 75100 12916 75104
rect 12852 75044 12856 75100
rect 12856 75044 12912 75100
rect 12912 75044 12916 75100
rect 12852 75040 12916 75044
rect 17612 75100 17676 75104
rect 17612 75044 17616 75100
rect 17616 75044 17672 75100
rect 17672 75044 17676 75100
rect 17612 75040 17676 75044
rect 17692 75100 17756 75104
rect 17692 75044 17696 75100
rect 17696 75044 17752 75100
rect 17752 75044 17756 75100
rect 17692 75040 17756 75044
rect 17772 75100 17836 75104
rect 17772 75044 17776 75100
rect 17776 75044 17832 75100
rect 17832 75044 17836 75100
rect 17772 75040 17836 75044
rect 17852 75100 17916 75104
rect 17852 75044 17856 75100
rect 17856 75044 17912 75100
rect 17912 75044 17916 75100
rect 17852 75040 17916 75044
rect 1952 74556 2016 74560
rect 1952 74500 1956 74556
rect 1956 74500 2012 74556
rect 2012 74500 2016 74556
rect 1952 74496 2016 74500
rect 2032 74556 2096 74560
rect 2032 74500 2036 74556
rect 2036 74500 2092 74556
rect 2092 74500 2096 74556
rect 2032 74496 2096 74500
rect 2112 74556 2176 74560
rect 2112 74500 2116 74556
rect 2116 74500 2172 74556
rect 2172 74500 2176 74556
rect 2112 74496 2176 74500
rect 2192 74556 2256 74560
rect 2192 74500 2196 74556
rect 2196 74500 2252 74556
rect 2252 74500 2256 74556
rect 2192 74496 2256 74500
rect 6952 74556 7016 74560
rect 6952 74500 6956 74556
rect 6956 74500 7012 74556
rect 7012 74500 7016 74556
rect 6952 74496 7016 74500
rect 7032 74556 7096 74560
rect 7032 74500 7036 74556
rect 7036 74500 7092 74556
rect 7092 74500 7096 74556
rect 7032 74496 7096 74500
rect 7112 74556 7176 74560
rect 7112 74500 7116 74556
rect 7116 74500 7172 74556
rect 7172 74500 7176 74556
rect 7112 74496 7176 74500
rect 7192 74556 7256 74560
rect 7192 74500 7196 74556
rect 7196 74500 7252 74556
rect 7252 74500 7256 74556
rect 7192 74496 7256 74500
rect 11952 74556 12016 74560
rect 11952 74500 11956 74556
rect 11956 74500 12012 74556
rect 12012 74500 12016 74556
rect 11952 74496 12016 74500
rect 12032 74556 12096 74560
rect 12032 74500 12036 74556
rect 12036 74500 12092 74556
rect 12092 74500 12096 74556
rect 12032 74496 12096 74500
rect 12112 74556 12176 74560
rect 12112 74500 12116 74556
rect 12116 74500 12172 74556
rect 12172 74500 12176 74556
rect 12112 74496 12176 74500
rect 12192 74556 12256 74560
rect 12192 74500 12196 74556
rect 12196 74500 12252 74556
rect 12252 74500 12256 74556
rect 12192 74496 12256 74500
rect 16952 74556 17016 74560
rect 16952 74500 16956 74556
rect 16956 74500 17012 74556
rect 17012 74500 17016 74556
rect 16952 74496 17016 74500
rect 17032 74556 17096 74560
rect 17032 74500 17036 74556
rect 17036 74500 17092 74556
rect 17092 74500 17096 74556
rect 17032 74496 17096 74500
rect 17112 74556 17176 74560
rect 17112 74500 17116 74556
rect 17116 74500 17172 74556
rect 17172 74500 17176 74556
rect 17112 74496 17176 74500
rect 17192 74556 17256 74560
rect 17192 74500 17196 74556
rect 17196 74500 17252 74556
rect 17252 74500 17256 74556
rect 17192 74496 17256 74500
rect 2612 74012 2676 74016
rect 2612 73956 2616 74012
rect 2616 73956 2672 74012
rect 2672 73956 2676 74012
rect 2612 73952 2676 73956
rect 2692 74012 2756 74016
rect 2692 73956 2696 74012
rect 2696 73956 2752 74012
rect 2752 73956 2756 74012
rect 2692 73952 2756 73956
rect 2772 74012 2836 74016
rect 2772 73956 2776 74012
rect 2776 73956 2832 74012
rect 2832 73956 2836 74012
rect 2772 73952 2836 73956
rect 2852 74012 2916 74016
rect 2852 73956 2856 74012
rect 2856 73956 2912 74012
rect 2912 73956 2916 74012
rect 2852 73952 2916 73956
rect 7612 74012 7676 74016
rect 7612 73956 7616 74012
rect 7616 73956 7672 74012
rect 7672 73956 7676 74012
rect 7612 73952 7676 73956
rect 7692 74012 7756 74016
rect 7692 73956 7696 74012
rect 7696 73956 7752 74012
rect 7752 73956 7756 74012
rect 7692 73952 7756 73956
rect 7772 74012 7836 74016
rect 7772 73956 7776 74012
rect 7776 73956 7832 74012
rect 7832 73956 7836 74012
rect 7772 73952 7836 73956
rect 7852 74012 7916 74016
rect 7852 73956 7856 74012
rect 7856 73956 7912 74012
rect 7912 73956 7916 74012
rect 7852 73952 7916 73956
rect 12612 74012 12676 74016
rect 12612 73956 12616 74012
rect 12616 73956 12672 74012
rect 12672 73956 12676 74012
rect 12612 73952 12676 73956
rect 12692 74012 12756 74016
rect 12692 73956 12696 74012
rect 12696 73956 12752 74012
rect 12752 73956 12756 74012
rect 12692 73952 12756 73956
rect 12772 74012 12836 74016
rect 12772 73956 12776 74012
rect 12776 73956 12832 74012
rect 12832 73956 12836 74012
rect 12772 73952 12836 73956
rect 12852 74012 12916 74016
rect 12852 73956 12856 74012
rect 12856 73956 12912 74012
rect 12912 73956 12916 74012
rect 12852 73952 12916 73956
rect 17612 74012 17676 74016
rect 17612 73956 17616 74012
rect 17616 73956 17672 74012
rect 17672 73956 17676 74012
rect 17612 73952 17676 73956
rect 17692 74012 17756 74016
rect 17692 73956 17696 74012
rect 17696 73956 17752 74012
rect 17752 73956 17756 74012
rect 17692 73952 17756 73956
rect 17772 74012 17836 74016
rect 17772 73956 17776 74012
rect 17776 73956 17832 74012
rect 17832 73956 17836 74012
rect 17772 73952 17836 73956
rect 17852 74012 17916 74016
rect 17852 73956 17856 74012
rect 17856 73956 17912 74012
rect 17912 73956 17916 74012
rect 17852 73952 17916 73956
rect 1952 73468 2016 73472
rect 1952 73412 1956 73468
rect 1956 73412 2012 73468
rect 2012 73412 2016 73468
rect 1952 73408 2016 73412
rect 2032 73468 2096 73472
rect 2032 73412 2036 73468
rect 2036 73412 2092 73468
rect 2092 73412 2096 73468
rect 2032 73408 2096 73412
rect 2112 73468 2176 73472
rect 2112 73412 2116 73468
rect 2116 73412 2172 73468
rect 2172 73412 2176 73468
rect 2112 73408 2176 73412
rect 2192 73468 2256 73472
rect 2192 73412 2196 73468
rect 2196 73412 2252 73468
rect 2252 73412 2256 73468
rect 2192 73408 2256 73412
rect 6952 73468 7016 73472
rect 6952 73412 6956 73468
rect 6956 73412 7012 73468
rect 7012 73412 7016 73468
rect 6952 73408 7016 73412
rect 7032 73468 7096 73472
rect 7032 73412 7036 73468
rect 7036 73412 7092 73468
rect 7092 73412 7096 73468
rect 7032 73408 7096 73412
rect 7112 73468 7176 73472
rect 7112 73412 7116 73468
rect 7116 73412 7172 73468
rect 7172 73412 7176 73468
rect 7112 73408 7176 73412
rect 7192 73468 7256 73472
rect 7192 73412 7196 73468
rect 7196 73412 7252 73468
rect 7252 73412 7256 73468
rect 7192 73408 7256 73412
rect 11952 73468 12016 73472
rect 11952 73412 11956 73468
rect 11956 73412 12012 73468
rect 12012 73412 12016 73468
rect 11952 73408 12016 73412
rect 12032 73468 12096 73472
rect 12032 73412 12036 73468
rect 12036 73412 12092 73468
rect 12092 73412 12096 73468
rect 12032 73408 12096 73412
rect 12112 73468 12176 73472
rect 12112 73412 12116 73468
rect 12116 73412 12172 73468
rect 12172 73412 12176 73468
rect 12112 73408 12176 73412
rect 12192 73468 12256 73472
rect 12192 73412 12196 73468
rect 12196 73412 12252 73468
rect 12252 73412 12256 73468
rect 12192 73408 12256 73412
rect 16952 73468 17016 73472
rect 16952 73412 16956 73468
rect 16956 73412 17012 73468
rect 17012 73412 17016 73468
rect 16952 73408 17016 73412
rect 17032 73468 17096 73472
rect 17032 73412 17036 73468
rect 17036 73412 17092 73468
rect 17092 73412 17096 73468
rect 17032 73408 17096 73412
rect 17112 73468 17176 73472
rect 17112 73412 17116 73468
rect 17116 73412 17172 73468
rect 17172 73412 17176 73468
rect 17112 73408 17176 73412
rect 17192 73468 17256 73472
rect 17192 73412 17196 73468
rect 17196 73412 17252 73468
rect 17252 73412 17256 73468
rect 17192 73408 17256 73412
rect 2612 72924 2676 72928
rect 2612 72868 2616 72924
rect 2616 72868 2672 72924
rect 2672 72868 2676 72924
rect 2612 72864 2676 72868
rect 2692 72924 2756 72928
rect 2692 72868 2696 72924
rect 2696 72868 2752 72924
rect 2752 72868 2756 72924
rect 2692 72864 2756 72868
rect 2772 72924 2836 72928
rect 2772 72868 2776 72924
rect 2776 72868 2832 72924
rect 2832 72868 2836 72924
rect 2772 72864 2836 72868
rect 2852 72924 2916 72928
rect 2852 72868 2856 72924
rect 2856 72868 2912 72924
rect 2912 72868 2916 72924
rect 2852 72864 2916 72868
rect 7612 72924 7676 72928
rect 7612 72868 7616 72924
rect 7616 72868 7672 72924
rect 7672 72868 7676 72924
rect 7612 72864 7676 72868
rect 7692 72924 7756 72928
rect 7692 72868 7696 72924
rect 7696 72868 7752 72924
rect 7752 72868 7756 72924
rect 7692 72864 7756 72868
rect 7772 72924 7836 72928
rect 7772 72868 7776 72924
rect 7776 72868 7832 72924
rect 7832 72868 7836 72924
rect 7772 72864 7836 72868
rect 7852 72924 7916 72928
rect 7852 72868 7856 72924
rect 7856 72868 7912 72924
rect 7912 72868 7916 72924
rect 7852 72864 7916 72868
rect 12612 72924 12676 72928
rect 12612 72868 12616 72924
rect 12616 72868 12672 72924
rect 12672 72868 12676 72924
rect 12612 72864 12676 72868
rect 12692 72924 12756 72928
rect 12692 72868 12696 72924
rect 12696 72868 12752 72924
rect 12752 72868 12756 72924
rect 12692 72864 12756 72868
rect 12772 72924 12836 72928
rect 12772 72868 12776 72924
rect 12776 72868 12832 72924
rect 12832 72868 12836 72924
rect 12772 72864 12836 72868
rect 12852 72924 12916 72928
rect 12852 72868 12856 72924
rect 12856 72868 12912 72924
rect 12912 72868 12916 72924
rect 12852 72864 12916 72868
rect 17612 72924 17676 72928
rect 17612 72868 17616 72924
rect 17616 72868 17672 72924
rect 17672 72868 17676 72924
rect 17612 72864 17676 72868
rect 17692 72924 17756 72928
rect 17692 72868 17696 72924
rect 17696 72868 17752 72924
rect 17752 72868 17756 72924
rect 17692 72864 17756 72868
rect 17772 72924 17836 72928
rect 17772 72868 17776 72924
rect 17776 72868 17832 72924
rect 17832 72868 17836 72924
rect 17772 72864 17836 72868
rect 17852 72924 17916 72928
rect 17852 72868 17856 72924
rect 17856 72868 17912 72924
rect 17912 72868 17916 72924
rect 17852 72864 17916 72868
rect 1952 72380 2016 72384
rect 1952 72324 1956 72380
rect 1956 72324 2012 72380
rect 2012 72324 2016 72380
rect 1952 72320 2016 72324
rect 2032 72380 2096 72384
rect 2032 72324 2036 72380
rect 2036 72324 2092 72380
rect 2092 72324 2096 72380
rect 2032 72320 2096 72324
rect 2112 72380 2176 72384
rect 2112 72324 2116 72380
rect 2116 72324 2172 72380
rect 2172 72324 2176 72380
rect 2112 72320 2176 72324
rect 2192 72380 2256 72384
rect 2192 72324 2196 72380
rect 2196 72324 2252 72380
rect 2252 72324 2256 72380
rect 2192 72320 2256 72324
rect 6952 72380 7016 72384
rect 6952 72324 6956 72380
rect 6956 72324 7012 72380
rect 7012 72324 7016 72380
rect 6952 72320 7016 72324
rect 7032 72380 7096 72384
rect 7032 72324 7036 72380
rect 7036 72324 7092 72380
rect 7092 72324 7096 72380
rect 7032 72320 7096 72324
rect 7112 72380 7176 72384
rect 7112 72324 7116 72380
rect 7116 72324 7172 72380
rect 7172 72324 7176 72380
rect 7112 72320 7176 72324
rect 7192 72380 7256 72384
rect 7192 72324 7196 72380
rect 7196 72324 7252 72380
rect 7252 72324 7256 72380
rect 7192 72320 7256 72324
rect 11952 72380 12016 72384
rect 11952 72324 11956 72380
rect 11956 72324 12012 72380
rect 12012 72324 12016 72380
rect 11952 72320 12016 72324
rect 12032 72380 12096 72384
rect 12032 72324 12036 72380
rect 12036 72324 12092 72380
rect 12092 72324 12096 72380
rect 12032 72320 12096 72324
rect 12112 72380 12176 72384
rect 12112 72324 12116 72380
rect 12116 72324 12172 72380
rect 12172 72324 12176 72380
rect 12112 72320 12176 72324
rect 12192 72380 12256 72384
rect 12192 72324 12196 72380
rect 12196 72324 12252 72380
rect 12252 72324 12256 72380
rect 12192 72320 12256 72324
rect 16952 72380 17016 72384
rect 16952 72324 16956 72380
rect 16956 72324 17012 72380
rect 17012 72324 17016 72380
rect 16952 72320 17016 72324
rect 17032 72380 17096 72384
rect 17032 72324 17036 72380
rect 17036 72324 17092 72380
rect 17092 72324 17096 72380
rect 17032 72320 17096 72324
rect 17112 72380 17176 72384
rect 17112 72324 17116 72380
rect 17116 72324 17172 72380
rect 17172 72324 17176 72380
rect 17112 72320 17176 72324
rect 17192 72380 17256 72384
rect 17192 72324 17196 72380
rect 17196 72324 17252 72380
rect 17252 72324 17256 72380
rect 17192 72320 17256 72324
rect 2612 71836 2676 71840
rect 2612 71780 2616 71836
rect 2616 71780 2672 71836
rect 2672 71780 2676 71836
rect 2612 71776 2676 71780
rect 2692 71836 2756 71840
rect 2692 71780 2696 71836
rect 2696 71780 2752 71836
rect 2752 71780 2756 71836
rect 2692 71776 2756 71780
rect 2772 71836 2836 71840
rect 2772 71780 2776 71836
rect 2776 71780 2832 71836
rect 2832 71780 2836 71836
rect 2772 71776 2836 71780
rect 2852 71836 2916 71840
rect 2852 71780 2856 71836
rect 2856 71780 2912 71836
rect 2912 71780 2916 71836
rect 2852 71776 2916 71780
rect 7612 71836 7676 71840
rect 7612 71780 7616 71836
rect 7616 71780 7672 71836
rect 7672 71780 7676 71836
rect 7612 71776 7676 71780
rect 7692 71836 7756 71840
rect 7692 71780 7696 71836
rect 7696 71780 7752 71836
rect 7752 71780 7756 71836
rect 7692 71776 7756 71780
rect 7772 71836 7836 71840
rect 7772 71780 7776 71836
rect 7776 71780 7832 71836
rect 7832 71780 7836 71836
rect 7772 71776 7836 71780
rect 7852 71836 7916 71840
rect 7852 71780 7856 71836
rect 7856 71780 7912 71836
rect 7912 71780 7916 71836
rect 7852 71776 7916 71780
rect 12612 71836 12676 71840
rect 12612 71780 12616 71836
rect 12616 71780 12672 71836
rect 12672 71780 12676 71836
rect 12612 71776 12676 71780
rect 12692 71836 12756 71840
rect 12692 71780 12696 71836
rect 12696 71780 12752 71836
rect 12752 71780 12756 71836
rect 12692 71776 12756 71780
rect 12772 71836 12836 71840
rect 12772 71780 12776 71836
rect 12776 71780 12832 71836
rect 12832 71780 12836 71836
rect 12772 71776 12836 71780
rect 12852 71836 12916 71840
rect 12852 71780 12856 71836
rect 12856 71780 12912 71836
rect 12912 71780 12916 71836
rect 12852 71776 12916 71780
rect 17612 71836 17676 71840
rect 17612 71780 17616 71836
rect 17616 71780 17672 71836
rect 17672 71780 17676 71836
rect 17612 71776 17676 71780
rect 17692 71836 17756 71840
rect 17692 71780 17696 71836
rect 17696 71780 17752 71836
rect 17752 71780 17756 71836
rect 17692 71776 17756 71780
rect 17772 71836 17836 71840
rect 17772 71780 17776 71836
rect 17776 71780 17832 71836
rect 17832 71780 17836 71836
rect 17772 71776 17836 71780
rect 17852 71836 17916 71840
rect 17852 71780 17856 71836
rect 17856 71780 17912 71836
rect 17912 71780 17916 71836
rect 17852 71776 17916 71780
rect 1952 71292 2016 71296
rect 1952 71236 1956 71292
rect 1956 71236 2012 71292
rect 2012 71236 2016 71292
rect 1952 71232 2016 71236
rect 2032 71292 2096 71296
rect 2032 71236 2036 71292
rect 2036 71236 2092 71292
rect 2092 71236 2096 71292
rect 2032 71232 2096 71236
rect 2112 71292 2176 71296
rect 2112 71236 2116 71292
rect 2116 71236 2172 71292
rect 2172 71236 2176 71292
rect 2112 71232 2176 71236
rect 2192 71292 2256 71296
rect 2192 71236 2196 71292
rect 2196 71236 2252 71292
rect 2252 71236 2256 71292
rect 2192 71232 2256 71236
rect 6952 71292 7016 71296
rect 6952 71236 6956 71292
rect 6956 71236 7012 71292
rect 7012 71236 7016 71292
rect 6952 71232 7016 71236
rect 7032 71292 7096 71296
rect 7032 71236 7036 71292
rect 7036 71236 7092 71292
rect 7092 71236 7096 71292
rect 7032 71232 7096 71236
rect 7112 71292 7176 71296
rect 7112 71236 7116 71292
rect 7116 71236 7172 71292
rect 7172 71236 7176 71292
rect 7112 71232 7176 71236
rect 7192 71292 7256 71296
rect 7192 71236 7196 71292
rect 7196 71236 7252 71292
rect 7252 71236 7256 71292
rect 7192 71232 7256 71236
rect 11952 71292 12016 71296
rect 11952 71236 11956 71292
rect 11956 71236 12012 71292
rect 12012 71236 12016 71292
rect 11952 71232 12016 71236
rect 12032 71292 12096 71296
rect 12032 71236 12036 71292
rect 12036 71236 12092 71292
rect 12092 71236 12096 71292
rect 12032 71232 12096 71236
rect 12112 71292 12176 71296
rect 12112 71236 12116 71292
rect 12116 71236 12172 71292
rect 12172 71236 12176 71292
rect 12112 71232 12176 71236
rect 12192 71292 12256 71296
rect 12192 71236 12196 71292
rect 12196 71236 12252 71292
rect 12252 71236 12256 71292
rect 12192 71232 12256 71236
rect 16952 71292 17016 71296
rect 16952 71236 16956 71292
rect 16956 71236 17012 71292
rect 17012 71236 17016 71292
rect 16952 71232 17016 71236
rect 17032 71292 17096 71296
rect 17032 71236 17036 71292
rect 17036 71236 17092 71292
rect 17092 71236 17096 71292
rect 17032 71232 17096 71236
rect 17112 71292 17176 71296
rect 17112 71236 17116 71292
rect 17116 71236 17172 71292
rect 17172 71236 17176 71292
rect 17112 71232 17176 71236
rect 17192 71292 17256 71296
rect 17192 71236 17196 71292
rect 17196 71236 17252 71292
rect 17252 71236 17256 71292
rect 17192 71232 17256 71236
rect 3372 70952 3436 70956
rect 3372 70896 3386 70952
rect 3386 70896 3436 70952
rect 3372 70892 3436 70896
rect 2612 70748 2676 70752
rect 2612 70692 2616 70748
rect 2616 70692 2672 70748
rect 2672 70692 2676 70748
rect 2612 70688 2676 70692
rect 2692 70748 2756 70752
rect 2692 70692 2696 70748
rect 2696 70692 2752 70748
rect 2752 70692 2756 70748
rect 2692 70688 2756 70692
rect 2772 70748 2836 70752
rect 2772 70692 2776 70748
rect 2776 70692 2832 70748
rect 2832 70692 2836 70748
rect 2772 70688 2836 70692
rect 2852 70748 2916 70752
rect 2852 70692 2856 70748
rect 2856 70692 2912 70748
rect 2912 70692 2916 70748
rect 2852 70688 2916 70692
rect 7612 70748 7676 70752
rect 7612 70692 7616 70748
rect 7616 70692 7672 70748
rect 7672 70692 7676 70748
rect 7612 70688 7676 70692
rect 7692 70748 7756 70752
rect 7692 70692 7696 70748
rect 7696 70692 7752 70748
rect 7752 70692 7756 70748
rect 7692 70688 7756 70692
rect 7772 70748 7836 70752
rect 7772 70692 7776 70748
rect 7776 70692 7832 70748
rect 7832 70692 7836 70748
rect 7772 70688 7836 70692
rect 7852 70748 7916 70752
rect 7852 70692 7856 70748
rect 7856 70692 7912 70748
rect 7912 70692 7916 70748
rect 7852 70688 7916 70692
rect 12612 70748 12676 70752
rect 12612 70692 12616 70748
rect 12616 70692 12672 70748
rect 12672 70692 12676 70748
rect 12612 70688 12676 70692
rect 12692 70748 12756 70752
rect 12692 70692 12696 70748
rect 12696 70692 12752 70748
rect 12752 70692 12756 70748
rect 12692 70688 12756 70692
rect 12772 70748 12836 70752
rect 12772 70692 12776 70748
rect 12776 70692 12832 70748
rect 12832 70692 12836 70748
rect 12772 70688 12836 70692
rect 12852 70748 12916 70752
rect 12852 70692 12856 70748
rect 12856 70692 12912 70748
rect 12912 70692 12916 70748
rect 12852 70688 12916 70692
rect 17612 70748 17676 70752
rect 17612 70692 17616 70748
rect 17616 70692 17672 70748
rect 17672 70692 17676 70748
rect 17612 70688 17676 70692
rect 17692 70748 17756 70752
rect 17692 70692 17696 70748
rect 17696 70692 17752 70748
rect 17752 70692 17756 70748
rect 17692 70688 17756 70692
rect 17772 70748 17836 70752
rect 17772 70692 17776 70748
rect 17776 70692 17832 70748
rect 17832 70692 17836 70748
rect 17772 70688 17836 70692
rect 17852 70748 17916 70752
rect 17852 70692 17856 70748
rect 17856 70692 17912 70748
rect 17912 70692 17916 70748
rect 17852 70688 17916 70692
rect 1952 70204 2016 70208
rect 1952 70148 1956 70204
rect 1956 70148 2012 70204
rect 2012 70148 2016 70204
rect 1952 70144 2016 70148
rect 2032 70204 2096 70208
rect 2032 70148 2036 70204
rect 2036 70148 2092 70204
rect 2092 70148 2096 70204
rect 2032 70144 2096 70148
rect 2112 70204 2176 70208
rect 2112 70148 2116 70204
rect 2116 70148 2172 70204
rect 2172 70148 2176 70204
rect 2112 70144 2176 70148
rect 2192 70204 2256 70208
rect 2192 70148 2196 70204
rect 2196 70148 2252 70204
rect 2252 70148 2256 70204
rect 2192 70144 2256 70148
rect 6952 70204 7016 70208
rect 6952 70148 6956 70204
rect 6956 70148 7012 70204
rect 7012 70148 7016 70204
rect 6952 70144 7016 70148
rect 7032 70204 7096 70208
rect 7032 70148 7036 70204
rect 7036 70148 7092 70204
rect 7092 70148 7096 70204
rect 7032 70144 7096 70148
rect 7112 70204 7176 70208
rect 7112 70148 7116 70204
rect 7116 70148 7172 70204
rect 7172 70148 7176 70204
rect 7112 70144 7176 70148
rect 7192 70204 7256 70208
rect 7192 70148 7196 70204
rect 7196 70148 7252 70204
rect 7252 70148 7256 70204
rect 7192 70144 7256 70148
rect 11952 70204 12016 70208
rect 11952 70148 11956 70204
rect 11956 70148 12012 70204
rect 12012 70148 12016 70204
rect 11952 70144 12016 70148
rect 12032 70204 12096 70208
rect 12032 70148 12036 70204
rect 12036 70148 12092 70204
rect 12092 70148 12096 70204
rect 12032 70144 12096 70148
rect 12112 70204 12176 70208
rect 12112 70148 12116 70204
rect 12116 70148 12172 70204
rect 12172 70148 12176 70204
rect 12112 70144 12176 70148
rect 12192 70204 12256 70208
rect 12192 70148 12196 70204
rect 12196 70148 12252 70204
rect 12252 70148 12256 70204
rect 12192 70144 12256 70148
rect 16952 70204 17016 70208
rect 16952 70148 16956 70204
rect 16956 70148 17012 70204
rect 17012 70148 17016 70204
rect 16952 70144 17016 70148
rect 17032 70204 17096 70208
rect 17032 70148 17036 70204
rect 17036 70148 17092 70204
rect 17092 70148 17096 70204
rect 17032 70144 17096 70148
rect 17112 70204 17176 70208
rect 17112 70148 17116 70204
rect 17116 70148 17172 70204
rect 17172 70148 17176 70204
rect 17112 70144 17176 70148
rect 17192 70204 17256 70208
rect 17192 70148 17196 70204
rect 17196 70148 17252 70204
rect 17252 70148 17256 70204
rect 17192 70144 17256 70148
rect 2612 69660 2676 69664
rect 2612 69604 2616 69660
rect 2616 69604 2672 69660
rect 2672 69604 2676 69660
rect 2612 69600 2676 69604
rect 2692 69660 2756 69664
rect 2692 69604 2696 69660
rect 2696 69604 2752 69660
rect 2752 69604 2756 69660
rect 2692 69600 2756 69604
rect 2772 69660 2836 69664
rect 2772 69604 2776 69660
rect 2776 69604 2832 69660
rect 2832 69604 2836 69660
rect 2772 69600 2836 69604
rect 2852 69660 2916 69664
rect 2852 69604 2856 69660
rect 2856 69604 2912 69660
rect 2912 69604 2916 69660
rect 2852 69600 2916 69604
rect 7612 69660 7676 69664
rect 7612 69604 7616 69660
rect 7616 69604 7672 69660
rect 7672 69604 7676 69660
rect 7612 69600 7676 69604
rect 7692 69660 7756 69664
rect 7692 69604 7696 69660
rect 7696 69604 7752 69660
rect 7752 69604 7756 69660
rect 7692 69600 7756 69604
rect 7772 69660 7836 69664
rect 7772 69604 7776 69660
rect 7776 69604 7832 69660
rect 7832 69604 7836 69660
rect 7772 69600 7836 69604
rect 7852 69660 7916 69664
rect 7852 69604 7856 69660
rect 7856 69604 7912 69660
rect 7912 69604 7916 69660
rect 7852 69600 7916 69604
rect 12612 69660 12676 69664
rect 12612 69604 12616 69660
rect 12616 69604 12672 69660
rect 12672 69604 12676 69660
rect 12612 69600 12676 69604
rect 12692 69660 12756 69664
rect 12692 69604 12696 69660
rect 12696 69604 12752 69660
rect 12752 69604 12756 69660
rect 12692 69600 12756 69604
rect 12772 69660 12836 69664
rect 12772 69604 12776 69660
rect 12776 69604 12832 69660
rect 12832 69604 12836 69660
rect 12772 69600 12836 69604
rect 12852 69660 12916 69664
rect 12852 69604 12856 69660
rect 12856 69604 12912 69660
rect 12912 69604 12916 69660
rect 12852 69600 12916 69604
rect 17612 69660 17676 69664
rect 17612 69604 17616 69660
rect 17616 69604 17672 69660
rect 17672 69604 17676 69660
rect 17612 69600 17676 69604
rect 17692 69660 17756 69664
rect 17692 69604 17696 69660
rect 17696 69604 17752 69660
rect 17752 69604 17756 69660
rect 17692 69600 17756 69604
rect 17772 69660 17836 69664
rect 17772 69604 17776 69660
rect 17776 69604 17832 69660
rect 17832 69604 17836 69660
rect 17772 69600 17836 69604
rect 17852 69660 17916 69664
rect 17852 69604 17856 69660
rect 17856 69604 17912 69660
rect 17912 69604 17916 69660
rect 17852 69600 17916 69604
rect 1716 69260 1780 69324
rect 1952 69116 2016 69120
rect 1952 69060 1956 69116
rect 1956 69060 2012 69116
rect 2012 69060 2016 69116
rect 1952 69056 2016 69060
rect 2032 69116 2096 69120
rect 2032 69060 2036 69116
rect 2036 69060 2092 69116
rect 2092 69060 2096 69116
rect 2032 69056 2096 69060
rect 2112 69116 2176 69120
rect 2112 69060 2116 69116
rect 2116 69060 2172 69116
rect 2172 69060 2176 69116
rect 2112 69056 2176 69060
rect 2192 69116 2256 69120
rect 2192 69060 2196 69116
rect 2196 69060 2252 69116
rect 2252 69060 2256 69116
rect 2192 69056 2256 69060
rect 6952 69116 7016 69120
rect 6952 69060 6956 69116
rect 6956 69060 7012 69116
rect 7012 69060 7016 69116
rect 6952 69056 7016 69060
rect 7032 69116 7096 69120
rect 7032 69060 7036 69116
rect 7036 69060 7092 69116
rect 7092 69060 7096 69116
rect 7032 69056 7096 69060
rect 7112 69116 7176 69120
rect 7112 69060 7116 69116
rect 7116 69060 7172 69116
rect 7172 69060 7176 69116
rect 7112 69056 7176 69060
rect 7192 69116 7256 69120
rect 7192 69060 7196 69116
rect 7196 69060 7252 69116
rect 7252 69060 7256 69116
rect 7192 69056 7256 69060
rect 11952 69116 12016 69120
rect 11952 69060 11956 69116
rect 11956 69060 12012 69116
rect 12012 69060 12016 69116
rect 11952 69056 12016 69060
rect 12032 69116 12096 69120
rect 12032 69060 12036 69116
rect 12036 69060 12092 69116
rect 12092 69060 12096 69116
rect 12032 69056 12096 69060
rect 12112 69116 12176 69120
rect 12112 69060 12116 69116
rect 12116 69060 12172 69116
rect 12172 69060 12176 69116
rect 12112 69056 12176 69060
rect 12192 69116 12256 69120
rect 12192 69060 12196 69116
rect 12196 69060 12252 69116
rect 12252 69060 12256 69116
rect 12192 69056 12256 69060
rect 16952 69116 17016 69120
rect 16952 69060 16956 69116
rect 16956 69060 17012 69116
rect 17012 69060 17016 69116
rect 16952 69056 17016 69060
rect 17032 69116 17096 69120
rect 17032 69060 17036 69116
rect 17036 69060 17092 69116
rect 17092 69060 17096 69116
rect 17032 69056 17096 69060
rect 17112 69116 17176 69120
rect 17112 69060 17116 69116
rect 17116 69060 17172 69116
rect 17172 69060 17176 69116
rect 17112 69056 17176 69060
rect 17192 69116 17256 69120
rect 17192 69060 17196 69116
rect 17196 69060 17252 69116
rect 17252 69060 17256 69116
rect 17192 69056 17256 69060
rect 14964 69048 15028 69052
rect 14964 68992 15014 69048
rect 15014 68992 15028 69048
rect 14964 68988 15028 68992
rect 2612 68572 2676 68576
rect 2612 68516 2616 68572
rect 2616 68516 2672 68572
rect 2672 68516 2676 68572
rect 2612 68512 2676 68516
rect 2692 68572 2756 68576
rect 2692 68516 2696 68572
rect 2696 68516 2752 68572
rect 2752 68516 2756 68572
rect 2692 68512 2756 68516
rect 2772 68572 2836 68576
rect 2772 68516 2776 68572
rect 2776 68516 2832 68572
rect 2832 68516 2836 68572
rect 2772 68512 2836 68516
rect 2852 68572 2916 68576
rect 2852 68516 2856 68572
rect 2856 68516 2912 68572
rect 2912 68516 2916 68572
rect 2852 68512 2916 68516
rect 7612 68572 7676 68576
rect 7612 68516 7616 68572
rect 7616 68516 7672 68572
rect 7672 68516 7676 68572
rect 7612 68512 7676 68516
rect 7692 68572 7756 68576
rect 7692 68516 7696 68572
rect 7696 68516 7752 68572
rect 7752 68516 7756 68572
rect 7692 68512 7756 68516
rect 7772 68572 7836 68576
rect 7772 68516 7776 68572
rect 7776 68516 7832 68572
rect 7832 68516 7836 68572
rect 7772 68512 7836 68516
rect 7852 68572 7916 68576
rect 7852 68516 7856 68572
rect 7856 68516 7912 68572
rect 7912 68516 7916 68572
rect 7852 68512 7916 68516
rect 12612 68572 12676 68576
rect 12612 68516 12616 68572
rect 12616 68516 12672 68572
rect 12672 68516 12676 68572
rect 12612 68512 12676 68516
rect 12692 68572 12756 68576
rect 12692 68516 12696 68572
rect 12696 68516 12752 68572
rect 12752 68516 12756 68572
rect 12692 68512 12756 68516
rect 12772 68572 12836 68576
rect 12772 68516 12776 68572
rect 12776 68516 12832 68572
rect 12832 68516 12836 68572
rect 12772 68512 12836 68516
rect 12852 68572 12916 68576
rect 12852 68516 12856 68572
rect 12856 68516 12912 68572
rect 12912 68516 12916 68572
rect 12852 68512 12916 68516
rect 17612 68572 17676 68576
rect 17612 68516 17616 68572
rect 17616 68516 17672 68572
rect 17672 68516 17676 68572
rect 17612 68512 17676 68516
rect 17692 68572 17756 68576
rect 17692 68516 17696 68572
rect 17696 68516 17752 68572
rect 17752 68516 17756 68572
rect 17692 68512 17756 68516
rect 17772 68572 17836 68576
rect 17772 68516 17776 68572
rect 17776 68516 17832 68572
rect 17832 68516 17836 68572
rect 17772 68512 17836 68516
rect 17852 68572 17916 68576
rect 17852 68516 17856 68572
rect 17856 68516 17912 68572
rect 17912 68516 17916 68572
rect 17852 68512 17916 68516
rect 1952 68028 2016 68032
rect 1952 67972 1956 68028
rect 1956 67972 2012 68028
rect 2012 67972 2016 68028
rect 1952 67968 2016 67972
rect 2032 68028 2096 68032
rect 2032 67972 2036 68028
rect 2036 67972 2092 68028
rect 2092 67972 2096 68028
rect 2032 67968 2096 67972
rect 2112 68028 2176 68032
rect 2112 67972 2116 68028
rect 2116 67972 2172 68028
rect 2172 67972 2176 68028
rect 2112 67968 2176 67972
rect 2192 68028 2256 68032
rect 2192 67972 2196 68028
rect 2196 67972 2252 68028
rect 2252 67972 2256 68028
rect 2192 67968 2256 67972
rect 6952 68028 7016 68032
rect 6952 67972 6956 68028
rect 6956 67972 7012 68028
rect 7012 67972 7016 68028
rect 6952 67968 7016 67972
rect 7032 68028 7096 68032
rect 7032 67972 7036 68028
rect 7036 67972 7092 68028
rect 7092 67972 7096 68028
rect 7032 67968 7096 67972
rect 7112 68028 7176 68032
rect 7112 67972 7116 68028
rect 7116 67972 7172 68028
rect 7172 67972 7176 68028
rect 7112 67968 7176 67972
rect 7192 68028 7256 68032
rect 7192 67972 7196 68028
rect 7196 67972 7252 68028
rect 7252 67972 7256 68028
rect 7192 67968 7256 67972
rect 11952 68028 12016 68032
rect 11952 67972 11956 68028
rect 11956 67972 12012 68028
rect 12012 67972 12016 68028
rect 11952 67968 12016 67972
rect 12032 68028 12096 68032
rect 12032 67972 12036 68028
rect 12036 67972 12092 68028
rect 12092 67972 12096 68028
rect 12032 67968 12096 67972
rect 12112 68028 12176 68032
rect 12112 67972 12116 68028
rect 12116 67972 12172 68028
rect 12172 67972 12176 68028
rect 12112 67968 12176 67972
rect 12192 68028 12256 68032
rect 12192 67972 12196 68028
rect 12196 67972 12252 68028
rect 12252 67972 12256 68028
rect 12192 67968 12256 67972
rect 16952 68028 17016 68032
rect 16952 67972 16956 68028
rect 16956 67972 17012 68028
rect 17012 67972 17016 68028
rect 16952 67968 17016 67972
rect 17032 68028 17096 68032
rect 17032 67972 17036 68028
rect 17036 67972 17092 68028
rect 17092 67972 17096 68028
rect 17032 67968 17096 67972
rect 17112 68028 17176 68032
rect 17112 67972 17116 68028
rect 17116 67972 17172 68028
rect 17172 67972 17176 68028
rect 17112 67968 17176 67972
rect 17192 68028 17256 68032
rect 17192 67972 17196 68028
rect 17196 67972 17252 68028
rect 17252 67972 17256 68028
rect 17192 67968 17256 67972
rect 10364 67628 10428 67692
rect 11652 67628 11716 67692
rect 2612 67484 2676 67488
rect 2612 67428 2616 67484
rect 2616 67428 2672 67484
rect 2672 67428 2676 67484
rect 2612 67424 2676 67428
rect 2692 67484 2756 67488
rect 2692 67428 2696 67484
rect 2696 67428 2752 67484
rect 2752 67428 2756 67484
rect 2692 67424 2756 67428
rect 2772 67484 2836 67488
rect 2772 67428 2776 67484
rect 2776 67428 2832 67484
rect 2832 67428 2836 67484
rect 2772 67424 2836 67428
rect 2852 67484 2916 67488
rect 2852 67428 2856 67484
rect 2856 67428 2912 67484
rect 2912 67428 2916 67484
rect 2852 67424 2916 67428
rect 7612 67484 7676 67488
rect 7612 67428 7616 67484
rect 7616 67428 7672 67484
rect 7672 67428 7676 67484
rect 7612 67424 7676 67428
rect 7692 67484 7756 67488
rect 7692 67428 7696 67484
rect 7696 67428 7752 67484
rect 7752 67428 7756 67484
rect 7692 67424 7756 67428
rect 7772 67484 7836 67488
rect 7772 67428 7776 67484
rect 7776 67428 7832 67484
rect 7832 67428 7836 67484
rect 7772 67424 7836 67428
rect 7852 67484 7916 67488
rect 7852 67428 7856 67484
rect 7856 67428 7912 67484
rect 7912 67428 7916 67484
rect 7852 67424 7916 67428
rect 12612 67484 12676 67488
rect 12612 67428 12616 67484
rect 12616 67428 12672 67484
rect 12672 67428 12676 67484
rect 12612 67424 12676 67428
rect 12692 67484 12756 67488
rect 12692 67428 12696 67484
rect 12696 67428 12752 67484
rect 12752 67428 12756 67484
rect 12692 67424 12756 67428
rect 12772 67484 12836 67488
rect 12772 67428 12776 67484
rect 12776 67428 12832 67484
rect 12832 67428 12836 67484
rect 12772 67424 12836 67428
rect 12852 67484 12916 67488
rect 12852 67428 12856 67484
rect 12856 67428 12912 67484
rect 12912 67428 12916 67484
rect 12852 67424 12916 67428
rect 17612 67484 17676 67488
rect 17612 67428 17616 67484
rect 17616 67428 17672 67484
rect 17672 67428 17676 67484
rect 17612 67424 17676 67428
rect 17692 67484 17756 67488
rect 17692 67428 17696 67484
rect 17696 67428 17752 67484
rect 17752 67428 17756 67484
rect 17692 67424 17756 67428
rect 17772 67484 17836 67488
rect 17772 67428 17776 67484
rect 17776 67428 17832 67484
rect 17832 67428 17836 67484
rect 17772 67424 17836 67428
rect 17852 67484 17916 67488
rect 17852 67428 17856 67484
rect 17856 67428 17912 67484
rect 17912 67428 17916 67484
rect 17852 67424 17916 67428
rect 1952 66940 2016 66944
rect 1952 66884 1956 66940
rect 1956 66884 2012 66940
rect 2012 66884 2016 66940
rect 1952 66880 2016 66884
rect 2032 66940 2096 66944
rect 2032 66884 2036 66940
rect 2036 66884 2092 66940
rect 2092 66884 2096 66940
rect 2032 66880 2096 66884
rect 2112 66940 2176 66944
rect 2112 66884 2116 66940
rect 2116 66884 2172 66940
rect 2172 66884 2176 66940
rect 2112 66880 2176 66884
rect 2192 66940 2256 66944
rect 2192 66884 2196 66940
rect 2196 66884 2252 66940
rect 2252 66884 2256 66940
rect 2192 66880 2256 66884
rect 6952 66940 7016 66944
rect 6952 66884 6956 66940
rect 6956 66884 7012 66940
rect 7012 66884 7016 66940
rect 6952 66880 7016 66884
rect 7032 66940 7096 66944
rect 7032 66884 7036 66940
rect 7036 66884 7092 66940
rect 7092 66884 7096 66940
rect 7032 66880 7096 66884
rect 7112 66940 7176 66944
rect 7112 66884 7116 66940
rect 7116 66884 7172 66940
rect 7172 66884 7176 66940
rect 7112 66880 7176 66884
rect 7192 66940 7256 66944
rect 7192 66884 7196 66940
rect 7196 66884 7252 66940
rect 7252 66884 7256 66940
rect 7192 66880 7256 66884
rect 11952 66940 12016 66944
rect 11952 66884 11956 66940
rect 11956 66884 12012 66940
rect 12012 66884 12016 66940
rect 11952 66880 12016 66884
rect 12032 66940 12096 66944
rect 12032 66884 12036 66940
rect 12036 66884 12092 66940
rect 12092 66884 12096 66940
rect 12032 66880 12096 66884
rect 12112 66940 12176 66944
rect 12112 66884 12116 66940
rect 12116 66884 12172 66940
rect 12172 66884 12176 66940
rect 12112 66880 12176 66884
rect 12192 66940 12256 66944
rect 12192 66884 12196 66940
rect 12196 66884 12252 66940
rect 12252 66884 12256 66940
rect 12192 66880 12256 66884
rect 16952 66940 17016 66944
rect 16952 66884 16956 66940
rect 16956 66884 17012 66940
rect 17012 66884 17016 66940
rect 16952 66880 17016 66884
rect 17032 66940 17096 66944
rect 17032 66884 17036 66940
rect 17036 66884 17092 66940
rect 17092 66884 17096 66940
rect 17032 66880 17096 66884
rect 17112 66940 17176 66944
rect 17112 66884 17116 66940
rect 17116 66884 17172 66940
rect 17172 66884 17176 66940
rect 17112 66880 17176 66884
rect 17192 66940 17256 66944
rect 17192 66884 17196 66940
rect 17196 66884 17252 66940
rect 17252 66884 17256 66940
rect 17192 66880 17256 66884
rect 2612 66396 2676 66400
rect 2612 66340 2616 66396
rect 2616 66340 2672 66396
rect 2672 66340 2676 66396
rect 2612 66336 2676 66340
rect 2692 66396 2756 66400
rect 2692 66340 2696 66396
rect 2696 66340 2752 66396
rect 2752 66340 2756 66396
rect 2692 66336 2756 66340
rect 2772 66396 2836 66400
rect 2772 66340 2776 66396
rect 2776 66340 2832 66396
rect 2832 66340 2836 66396
rect 2772 66336 2836 66340
rect 2852 66396 2916 66400
rect 2852 66340 2856 66396
rect 2856 66340 2912 66396
rect 2912 66340 2916 66396
rect 2852 66336 2916 66340
rect 7612 66396 7676 66400
rect 7612 66340 7616 66396
rect 7616 66340 7672 66396
rect 7672 66340 7676 66396
rect 7612 66336 7676 66340
rect 7692 66396 7756 66400
rect 7692 66340 7696 66396
rect 7696 66340 7752 66396
rect 7752 66340 7756 66396
rect 7692 66336 7756 66340
rect 7772 66396 7836 66400
rect 7772 66340 7776 66396
rect 7776 66340 7832 66396
rect 7832 66340 7836 66396
rect 7772 66336 7836 66340
rect 7852 66396 7916 66400
rect 7852 66340 7856 66396
rect 7856 66340 7912 66396
rect 7912 66340 7916 66396
rect 7852 66336 7916 66340
rect 12612 66396 12676 66400
rect 12612 66340 12616 66396
rect 12616 66340 12672 66396
rect 12672 66340 12676 66396
rect 12612 66336 12676 66340
rect 12692 66396 12756 66400
rect 12692 66340 12696 66396
rect 12696 66340 12752 66396
rect 12752 66340 12756 66396
rect 12692 66336 12756 66340
rect 12772 66396 12836 66400
rect 12772 66340 12776 66396
rect 12776 66340 12832 66396
rect 12832 66340 12836 66396
rect 12772 66336 12836 66340
rect 12852 66396 12916 66400
rect 12852 66340 12856 66396
rect 12856 66340 12912 66396
rect 12912 66340 12916 66396
rect 12852 66336 12916 66340
rect 17612 66396 17676 66400
rect 17612 66340 17616 66396
rect 17616 66340 17672 66396
rect 17672 66340 17676 66396
rect 17612 66336 17676 66340
rect 17692 66396 17756 66400
rect 17692 66340 17696 66396
rect 17696 66340 17752 66396
rect 17752 66340 17756 66396
rect 17692 66336 17756 66340
rect 17772 66396 17836 66400
rect 17772 66340 17776 66396
rect 17776 66340 17832 66396
rect 17832 66340 17836 66396
rect 17772 66336 17836 66340
rect 17852 66396 17916 66400
rect 17852 66340 17856 66396
rect 17856 66340 17912 66396
rect 17912 66340 17916 66396
rect 17852 66336 17916 66340
rect 1952 65852 2016 65856
rect 1952 65796 1956 65852
rect 1956 65796 2012 65852
rect 2012 65796 2016 65852
rect 1952 65792 2016 65796
rect 2032 65852 2096 65856
rect 2032 65796 2036 65852
rect 2036 65796 2092 65852
rect 2092 65796 2096 65852
rect 2032 65792 2096 65796
rect 2112 65852 2176 65856
rect 2112 65796 2116 65852
rect 2116 65796 2172 65852
rect 2172 65796 2176 65852
rect 2112 65792 2176 65796
rect 2192 65852 2256 65856
rect 2192 65796 2196 65852
rect 2196 65796 2252 65852
rect 2252 65796 2256 65852
rect 2192 65792 2256 65796
rect 6952 65852 7016 65856
rect 6952 65796 6956 65852
rect 6956 65796 7012 65852
rect 7012 65796 7016 65852
rect 6952 65792 7016 65796
rect 7032 65852 7096 65856
rect 7032 65796 7036 65852
rect 7036 65796 7092 65852
rect 7092 65796 7096 65852
rect 7032 65792 7096 65796
rect 7112 65852 7176 65856
rect 7112 65796 7116 65852
rect 7116 65796 7172 65852
rect 7172 65796 7176 65852
rect 7112 65792 7176 65796
rect 7192 65852 7256 65856
rect 7192 65796 7196 65852
rect 7196 65796 7252 65852
rect 7252 65796 7256 65852
rect 7192 65792 7256 65796
rect 11952 65852 12016 65856
rect 11952 65796 11956 65852
rect 11956 65796 12012 65852
rect 12012 65796 12016 65852
rect 11952 65792 12016 65796
rect 12032 65852 12096 65856
rect 12032 65796 12036 65852
rect 12036 65796 12092 65852
rect 12092 65796 12096 65852
rect 12032 65792 12096 65796
rect 12112 65852 12176 65856
rect 12112 65796 12116 65852
rect 12116 65796 12172 65852
rect 12172 65796 12176 65852
rect 12112 65792 12176 65796
rect 12192 65852 12256 65856
rect 12192 65796 12196 65852
rect 12196 65796 12252 65852
rect 12252 65796 12256 65852
rect 12192 65792 12256 65796
rect 16952 65852 17016 65856
rect 16952 65796 16956 65852
rect 16956 65796 17012 65852
rect 17012 65796 17016 65852
rect 16952 65792 17016 65796
rect 17032 65852 17096 65856
rect 17032 65796 17036 65852
rect 17036 65796 17092 65852
rect 17092 65796 17096 65852
rect 17032 65792 17096 65796
rect 17112 65852 17176 65856
rect 17112 65796 17116 65852
rect 17116 65796 17172 65852
rect 17172 65796 17176 65852
rect 17112 65792 17176 65796
rect 17192 65852 17256 65856
rect 17192 65796 17196 65852
rect 17196 65796 17252 65852
rect 17252 65796 17256 65852
rect 17192 65792 17256 65796
rect 2612 65308 2676 65312
rect 2612 65252 2616 65308
rect 2616 65252 2672 65308
rect 2672 65252 2676 65308
rect 2612 65248 2676 65252
rect 2692 65308 2756 65312
rect 2692 65252 2696 65308
rect 2696 65252 2752 65308
rect 2752 65252 2756 65308
rect 2692 65248 2756 65252
rect 2772 65308 2836 65312
rect 2772 65252 2776 65308
rect 2776 65252 2832 65308
rect 2832 65252 2836 65308
rect 2772 65248 2836 65252
rect 2852 65308 2916 65312
rect 2852 65252 2856 65308
rect 2856 65252 2912 65308
rect 2912 65252 2916 65308
rect 2852 65248 2916 65252
rect 7612 65308 7676 65312
rect 7612 65252 7616 65308
rect 7616 65252 7672 65308
rect 7672 65252 7676 65308
rect 7612 65248 7676 65252
rect 7692 65308 7756 65312
rect 7692 65252 7696 65308
rect 7696 65252 7752 65308
rect 7752 65252 7756 65308
rect 7692 65248 7756 65252
rect 7772 65308 7836 65312
rect 7772 65252 7776 65308
rect 7776 65252 7832 65308
rect 7832 65252 7836 65308
rect 7772 65248 7836 65252
rect 7852 65308 7916 65312
rect 7852 65252 7856 65308
rect 7856 65252 7912 65308
rect 7912 65252 7916 65308
rect 7852 65248 7916 65252
rect 12612 65308 12676 65312
rect 12612 65252 12616 65308
rect 12616 65252 12672 65308
rect 12672 65252 12676 65308
rect 12612 65248 12676 65252
rect 12692 65308 12756 65312
rect 12692 65252 12696 65308
rect 12696 65252 12752 65308
rect 12752 65252 12756 65308
rect 12692 65248 12756 65252
rect 12772 65308 12836 65312
rect 12772 65252 12776 65308
rect 12776 65252 12832 65308
rect 12832 65252 12836 65308
rect 12772 65248 12836 65252
rect 12852 65308 12916 65312
rect 12852 65252 12856 65308
rect 12856 65252 12912 65308
rect 12912 65252 12916 65308
rect 12852 65248 12916 65252
rect 17612 65308 17676 65312
rect 17612 65252 17616 65308
rect 17616 65252 17672 65308
rect 17672 65252 17676 65308
rect 17612 65248 17676 65252
rect 17692 65308 17756 65312
rect 17692 65252 17696 65308
rect 17696 65252 17752 65308
rect 17752 65252 17756 65308
rect 17692 65248 17756 65252
rect 17772 65308 17836 65312
rect 17772 65252 17776 65308
rect 17776 65252 17832 65308
rect 17832 65252 17836 65308
rect 17772 65248 17836 65252
rect 17852 65308 17916 65312
rect 17852 65252 17856 65308
rect 17856 65252 17912 65308
rect 17912 65252 17916 65308
rect 17852 65248 17916 65252
rect 3924 65180 3988 65244
rect 15700 65044 15764 65108
rect 1952 64764 2016 64768
rect 1952 64708 1956 64764
rect 1956 64708 2012 64764
rect 2012 64708 2016 64764
rect 1952 64704 2016 64708
rect 2032 64764 2096 64768
rect 2032 64708 2036 64764
rect 2036 64708 2092 64764
rect 2092 64708 2096 64764
rect 2032 64704 2096 64708
rect 2112 64764 2176 64768
rect 2112 64708 2116 64764
rect 2116 64708 2172 64764
rect 2172 64708 2176 64764
rect 2112 64704 2176 64708
rect 2192 64764 2256 64768
rect 2192 64708 2196 64764
rect 2196 64708 2252 64764
rect 2252 64708 2256 64764
rect 2192 64704 2256 64708
rect 6952 64764 7016 64768
rect 6952 64708 6956 64764
rect 6956 64708 7012 64764
rect 7012 64708 7016 64764
rect 6952 64704 7016 64708
rect 7032 64764 7096 64768
rect 7032 64708 7036 64764
rect 7036 64708 7092 64764
rect 7092 64708 7096 64764
rect 7032 64704 7096 64708
rect 7112 64764 7176 64768
rect 7112 64708 7116 64764
rect 7116 64708 7172 64764
rect 7172 64708 7176 64764
rect 7112 64704 7176 64708
rect 7192 64764 7256 64768
rect 7192 64708 7196 64764
rect 7196 64708 7252 64764
rect 7252 64708 7256 64764
rect 7192 64704 7256 64708
rect 11952 64764 12016 64768
rect 11952 64708 11956 64764
rect 11956 64708 12012 64764
rect 12012 64708 12016 64764
rect 11952 64704 12016 64708
rect 12032 64764 12096 64768
rect 12032 64708 12036 64764
rect 12036 64708 12092 64764
rect 12092 64708 12096 64764
rect 12032 64704 12096 64708
rect 12112 64764 12176 64768
rect 12112 64708 12116 64764
rect 12116 64708 12172 64764
rect 12172 64708 12176 64764
rect 12112 64704 12176 64708
rect 12192 64764 12256 64768
rect 12192 64708 12196 64764
rect 12196 64708 12252 64764
rect 12252 64708 12256 64764
rect 12192 64704 12256 64708
rect 16952 64764 17016 64768
rect 16952 64708 16956 64764
rect 16956 64708 17012 64764
rect 17012 64708 17016 64764
rect 16952 64704 17016 64708
rect 17032 64764 17096 64768
rect 17032 64708 17036 64764
rect 17036 64708 17092 64764
rect 17092 64708 17096 64764
rect 17032 64704 17096 64708
rect 17112 64764 17176 64768
rect 17112 64708 17116 64764
rect 17116 64708 17172 64764
rect 17172 64708 17176 64764
rect 17112 64704 17176 64708
rect 17192 64764 17256 64768
rect 17192 64708 17196 64764
rect 17196 64708 17252 64764
rect 17252 64708 17256 64764
rect 17192 64704 17256 64708
rect 2612 64220 2676 64224
rect 2612 64164 2616 64220
rect 2616 64164 2672 64220
rect 2672 64164 2676 64220
rect 2612 64160 2676 64164
rect 2692 64220 2756 64224
rect 2692 64164 2696 64220
rect 2696 64164 2752 64220
rect 2752 64164 2756 64220
rect 2692 64160 2756 64164
rect 2772 64220 2836 64224
rect 2772 64164 2776 64220
rect 2776 64164 2832 64220
rect 2832 64164 2836 64220
rect 2772 64160 2836 64164
rect 2852 64220 2916 64224
rect 2852 64164 2856 64220
rect 2856 64164 2912 64220
rect 2912 64164 2916 64220
rect 2852 64160 2916 64164
rect 7612 64220 7676 64224
rect 7612 64164 7616 64220
rect 7616 64164 7672 64220
rect 7672 64164 7676 64220
rect 7612 64160 7676 64164
rect 7692 64220 7756 64224
rect 7692 64164 7696 64220
rect 7696 64164 7752 64220
rect 7752 64164 7756 64220
rect 7692 64160 7756 64164
rect 7772 64220 7836 64224
rect 7772 64164 7776 64220
rect 7776 64164 7832 64220
rect 7832 64164 7836 64220
rect 7772 64160 7836 64164
rect 7852 64220 7916 64224
rect 7852 64164 7856 64220
rect 7856 64164 7912 64220
rect 7912 64164 7916 64220
rect 7852 64160 7916 64164
rect 12612 64220 12676 64224
rect 12612 64164 12616 64220
rect 12616 64164 12672 64220
rect 12672 64164 12676 64220
rect 12612 64160 12676 64164
rect 12692 64220 12756 64224
rect 12692 64164 12696 64220
rect 12696 64164 12752 64220
rect 12752 64164 12756 64220
rect 12692 64160 12756 64164
rect 12772 64220 12836 64224
rect 12772 64164 12776 64220
rect 12776 64164 12832 64220
rect 12832 64164 12836 64220
rect 12772 64160 12836 64164
rect 12852 64220 12916 64224
rect 12852 64164 12856 64220
rect 12856 64164 12912 64220
rect 12912 64164 12916 64220
rect 12852 64160 12916 64164
rect 17612 64220 17676 64224
rect 17612 64164 17616 64220
rect 17616 64164 17672 64220
rect 17672 64164 17676 64220
rect 17612 64160 17676 64164
rect 17692 64220 17756 64224
rect 17692 64164 17696 64220
rect 17696 64164 17752 64220
rect 17752 64164 17756 64220
rect 17692 64160 17756 64164
rect 17772 64220 17836 64224
rect 17772 64164 17776 64220
rect 17776 64164 17832 64220
rect 17832 64164 17836 64220
rect 17772 64160 17836 64164
rect 17852 64220 17916 64224
rect 17852 64164 17856 64220
rect 17856 64164 17912 64220
rect 17912 64164 17916 64220
rect 17852 64160 17916 64164
rect 1952 63676 2016 63680
rect 1952 63620 1956 63676
rect 1956 63620 2012 63676
rect 2012 63620 2016 63676
rect 1952 63616 2016 63620
rect 2032 63676 2096 63680
rect 2032 63620 2036 63676
rect 2036 63620 2092 63676
rect 2092 63620 2096 63676
rect 2032 63616 2096 63620
rect 2112 63676 2176 63680
rect 2112 63620 2116 63676
rect 2116 63620 2172 63676
rect 2172 63620 2176 63676
rect 2112 63616 2176 63620
rect 2192 63676 2256 63680
rect 2192 63620 2196 63676
rect 2196 63620 2252 63676
rect 2252 63620 2256 63676
rect 2192 63616 2256 63620
rect 6952 63676 7016 63680
rect 6952 63620 6956 63676
rect 6956 63620 7012 63676
rect 7012 63620 7016 63676
rect 6952 63616 7016 63620
rect 7032 63676 7096 63680
rect 7032 63620 7036 63676
rect 7036 63620 7092 63676
rect 7092 63620 7096 63676
rect 7032 63616 7096 63620
rect 7112 63676 7176 63680
rect 7112 63620 7116 63676
rect 7116 63620 7172 63676
rect 7172 63620 7176 63676
rect 7112 63616 7176 63620
rect 7192 63676 7256 63680
rect 7192 63620 7196 63676
rect 7196 63620 7252 63676
rect 7252 63620 7256 63676
rect 7192 63616 7256 63620
rect 11952 63676 12016 63680
rect 11952 63620 11956 63676
rect 11956 63620 12012 63676
rect 12012 63620 12016 63676
rect 11952 63616 12016 63620
rect 12032 63676 12096 63680
rect 12032 63620 12036 63676
rect 12036 63620 12092 63676
rect 12092 63620 12096 63676
rect 12032 63616 12096 63620
rect 12112 63676 12176 63680
rect 12112 63620 12116 63676
rect 12116 63620 12172 63676
rect 12172 63620 12176 63676
rect 12112 63616 12176 63620
rect 12192 63676 12256 63680
rect 12192 63620 12196 63676
rect 12196 63620 12252 63676
rect 12252 63620 12256 63676
rect 12192 63616 12256 63620
rect 16952 63676 17016 63680
rect 16952 63620 16956 63676
rect 16956 63620 17012 63676
rect 17012 63620 17016 63676
rect 16952 63616 17016 63620
rect 17032 63676 17096 63680
rect 17032 63620 17036 63676
rect 17036 63620 17092 63676
rect 17092 63620 17096 63676
rect 17032 63616 17096 63620
rect 17112 63676 17176 63680
rect 17112 63620 17116 63676
rect 17116 63620 17172 63676
rect 17172 63620 17176 63676
rect 17112 63616 17176 63620
rect 17192 63676 17256 63680
rect 17192 63620 17196 63676
rect 17196 63620 17252 63676
rect 17252 63620 17256 63676
rect 17192 63616 17256 63620
rect 4844 63276 4908 63340
rect 2612 63132 2676 63136
rect 2612 63076 2616 63132
rect 2616 63076 2672 63132
rect 2672 63076 2676 63132
rect 2612 63072 2676 63076
rect 2692 63132 2756 63136
rect 2692 63076 2696 63132
rect 2696 63076 2752 63132
rect 2752 63076 2756 63132
rect 2692 63072 2756 63076
rect 2772 63132 2836 63136
rect 2772 63076 2776 63132
rect 2776 63076 2832 63132
rect 2832 63076 2836 63132
rect 2772 63072 2836 63076
rect 2852 63132 2916 63136
rect 2852 63076 2856 63132
rect 2856 63076 2912 63132
rect 2912 63076 2916 63132
rect 2852 63072 2916 63076
rect 7612 63132 7676 63136
rect 7612 63076 7616 63132
rect 7616 63076 7672 63132
rect 7672 63076 7676 63132
rect 7612 63072 7676 63076
rect 7692 63132 7756 63136
rect 7692 63076 7696 63132
rect 7696 63076 7752 63132
rect 7752 63076 7756 63132
rect 7692 63072 7756 63076
rect 7772 63132 7836 63136
rect 7772 63076 7776 63132
rect 7776 63076 7832 63132
rect 7832 63076 7836 63132
rect 7772 63072 7836 63076
rect 7852 63132 7916 63136
rect 7852 63076 7856 63132
rect 7856 63076 7912 63132
rect 7912 63076 7916 63132
rect 7852 63072 7916 63076
rect 12612 63132 12676 63136
rect 12612 63076 12616 63132
rect 12616 63076 12672 63132
rect 12672 63076 12676 63132
rect 12612 63072 12676 63076
rect 12692 63132 12756 63136
rect 12692 63076 12696 63132
rect 12696 63076 12752 63132
rect 12752 63076 12756 63132
rect 12692 63072 12756 63076
rect 12772 63132 12836 63136
rect 12772 63076 12776 63132
rect 12776 63076 12832 63132
rect 12832 63076 12836 63132
rect 12772 63072 12836 63076
rect 12852 63132 12916 63136
rect 12852 63076 12856 63132
rect 12856 63076 12912 63132
rect 12912 63076 12916 63132
rect 12852 63072 12916 63076
rect 17612 63132 17676 63136
rect 17612 63076 17616 63132
rect 17616 63076 17672 63132
rect 17672 63076 17676 63132
rect 17612 63072 17676 63076
rect 17692 63132 17756 63136
rect 17692 63076 17696 63132
rect 17696 63076 17752 63132
rect 17752 63076 17756 63132
rect 17692 63072 17756 63076
rect 17772 63132 17836 63136
rect 17772 63076 17776 63132
rect 17776 63076 17832 63132
rect 17832 63076 17836 63132
rect 17772 63072 17836 63076
rect 17852 63132 17916 63136
rect 17852 63076 17856 63132
rect 17856 63076 17912 63132
rect 17912 63076 17916 63132
rect 17852 63072 17916 63076
rect 8708 62656 8772 62660
rect 8708 62600 8758 62656
rect 8758 62600 8772 62656
rect 8708 62596 8772 62600
rect 1952 62588 2016 62592
rect 1952 62532 1956 62588
rect 1956 62532 2012 62588
rect 2012 62532 2016 62588
rect 1952 62528 2016 62532
rect 2032 62588 2096 62592
rect 2032 62532 2036 62588
rect 2036 62532 2092 62588
rect 2092 62532 2096 62588
rect 2032 62528 2096 62532
rect 2112 62588 2176 62592
rect 2112 62532 2116 62588
rect 2116 62532 2172 62588
rect 2172 62532 2176 62588
rect 2112 62528 2176 62532
rect 2192 62588 2256 62592
rect 2192 62532 2196 62588
rect 2196 62532 2252 62588
rect 2252 62532 2256 62588
rect 2192 62528 2256 62532
rect 6952 62588 7016 62592
rect 6952 62532 6956 62588
rect 6956 62532 7012 62588
rect 7012 62532 7016 62588
rect 6952 62528 7016 62532
rect 7032 62588 7096 62592
rect 7032 62532 7036 62588
rect 7036 62532 7092 62588
rect 7092 62532 7096 62588
rect 7032 62528 7096 62532
rect 7112 62588 7176 62592
rect 7112 62532 7116 62588
rect 7116 62532 7172 62588
rect 7172 62532 7176 62588
rect 7112 62528 7176 62532
rect 7192 62588 7256 62592
rect 7192 62532 7196 62588
rect 7196 62532 7252 62588
rect 7252 62532 7256 62588
rect 7192 62528 7256 62532
rect 11952 62588 12016 62592
rect 11952 62532 11956 62588
rect 11956 62532 12012 62588
rect 12012 62532 12016 62588
rect 11952 62528 12016 62532
rect 12032 62588 12096 62592
rect 12032 62532 12036 62588
rect 12036 62532 12092 62588
rect 12092 62532 12096 62588
rect 12032 62528 12096 62532
rect 12112 62588 12176 62592
rect 12112 62532 12116 62588
rect 12116 62532 12172 62588
rect 12172 62532 12176 62588
rect 12112 62528 12176 62532
rect 12192 62588 12256 62592
rect 12192 62532 12196 62588
rect 12196 62532 12252 62588
rect 12252 62532 12256 62588
rect 12192 62528 12256 62532
rect 16952 62588 17016 62592
rect 16952 62532 16956 62588
rect 16956 62532 17012 62588
rect 17012 62532 17016 62588
rect 16952 62528 17016 62532
rect 17032 62588 17096 62592
rect 17032 62532 17036 62588
rect 17036 62532 17092 62588
rect 17092 62532 17096 62588
rect 17032 62528 17096 62532
rect 17112 62588 17176 62592
rect 17112 62532 17116 62588
rect 17116 62532 17172 62588
rect 17172 62532 17176 62588
rect 17112 62528 17176 62532
rect 17192 62588 17256 62592
rect 17192 62532 17196 62588
rect 17196 62532 17252 62588
rect 17252 62532 17256 62588
rect 17192 62528 17256 62532
rect 4292 62248 4356 62252
rect 4292 62192 4306 62248
rect 4306 62192 4356 62248
rect 4292 62188 4356 62192
rect 2612 62044 2676 62048
rect 2612 61988 2616 62044
rect 2616 61988 2672 62044
rect 2672 61988 2676 62044
rect 2612 61984 2676 61988
rect 2692 62044 2756 62048
rect 2692 61988 2696 62044
rect 2696 61988 2752 62044
rect 2752 61988 2756 62044
rect 2692 61984 2756 61988
rect 2772 62044 2836 62048
rect 2772 61988 2776 62044
rect 2776 61988 2832 62044
rect 2832 61988 2836 62044
rect 2772 61984 2836 61988
rect 2852 62044 2916 62048
rect 2852 61988 2856 62044
rect 2856 61988 2912 62044
rect 2912 61988 2916 62044
rect 2852 61984 2916 61988
rect 7612 62044 7676 62048
rect 7612 61988 7616 62044
rect 7616 61988 7672 62044
rect 7672 61988 7676 62044
rect 7612 61984 7676 61988
rect 7692 62044 7756 62048
rect 7692 61988 7696 62044
rect 7696 61988 7752 62044
rect 7752 61988 7756 62044
rect 7692 61984 7756 61988
rect 7772 62044 7836 62048
rect 7772 61988 7776 62044
rect 7776 61988 7832 62044
rect 7832 61988 7836 62044
rect 7772 61984 7836 61988
rect 7852 62044 7916 62048
rect 7852 61988 7856 62044
rect 7856 61988 7912 62044
rect 7912 61988 7916 62044
rect 7852 61984 7916 61988
rect 12612 62044 12676 62048
rect 12612 61988 12616 62044
rect 12616 61988 12672 62044
rect 12672 61988 12676 62044
rect 12612 61984 12676 61988
rect 12692 62044 12756 62048
rect 12692 61988 12696 62044
rect 12696 61988 12752 62044
rect 12752 61988 12756 62044
rect 12692 61984 12756 61988
rect 12772 62044 12836 62048
rect 12772 61988 12776 62044
rect 12776 61988 12832 62044
rect 12832 61988 12836 62044
rect 12772 61984 12836 61988
rect 12852 62044 12916 62048
rect 12852 61988 12856 62044
rect 12856 61988 12912 62044
rect 12912 61988 12916 62044
rect 12852 61984 12916 61988
rect 17612 62044 17676 62048
rect 17612 61988 17616 62044
rect 17616 61988 17672 62044
rect 17672 61988 17676 62044
rect 17612 61984 17676 61988
rect 17692 62044 17756 62048
rect 17692 61988 17696 62044
rect 17696 61988 17752 62044
rect 17752 61988 17756 62044
rect 17692 61984 17756 61988
rect 17772 62044 17836 62048
rect 17772 61988 17776 62044
rect 17776 61988 17832 62044
rect 17832 61988 17836 62044
rect 17772 61984 17836 61988
rect 17852 62044 17916 62048
rect 17852 61988 17856 62044
rect 17856 61988 17912 62044
rect 17912 61988 17916 62044
rect 17852 61984 17916 61988
rect 1952 61500 2016 61504
rect 1952 61444 1956 61500
rect 1956 61444 2012 61500
rect 2012 61444 2016 61500
rect 1952 61440 2016 61444
rect 2032 61500 2096 61504
rect 2032 61444 2036 61500
rect 2036 61444 2092 61500
rect 2092 61444 2096 61500
rect 2032 61440 2096 61444
rect 2112 61500 2176 61504
rect 2112 61444 2116 61500
rect 2116 61444 2172 61500
rect 2172 61444 2176 61500
rect 2112 61440 2176 61444
rect 2192 61500 2256 61504
rect 2192 61444 2196 61500
rect 2196 61444 2252 61500
rect 2252 61444 2256 61500
rect 2192 61440 2256 61444
rect 6952 61500 7016 61504
rect 6952 61444 6956 61500
rect 6956 61444 7012 61500
rect 7012 61444 7016 61500
rect 6952 61440 7016 61444
rect 7032 61500 7096 61504
rect 7032 61444 7036 61500
rect 7036 61444 7092 61500
rect 7092 61444 7096 61500
rect 7032 61440 7096 61444
rect 7112 61500 7176 61504
rect 7112 61444 7116 61500
rect 7116 61444 7172 61500
rect 7172 61444 7176 61500
rect 7112 61440 7176 61444
rect 7192 61500 7256 61504
rect 7192 61444 7196 61500
rect 7196 61444 7252 61500
rect 7252 61444 7256 61500
rect 7192 61440 7256 61444
rect 11952 61500 12016 61504
rect 11952 61444 11956 61500
rect 11956 61444 12012 61500
rect 12012 61444 12016 61500
rect 11952 61440 12016 61444
rect 12032 61500 12096 61504
rect 12032 61444 12036 61500
rect 12036 61444 12092 61500
rect 12092 61444 12096 61500
rect 12032 61440 12096 61444
rect 12112 61500 12176 61504
rect 12112 61444 12116 61500
rect 12116 61444 12172 61500
rect 12172 61444 12176 61500
rect 12112 61440 12176 61444
rect 12192 61500 12256 61504
rect 12192 61444 12196 61500
rect 12196 61444 12252 61500
rect 12252 61444 12256 61500
rect 12192 61440 12256 61444
rect 16952 61500 17016 61504
rect 16952 61444 16956 61500
rect 16956 61444 17012 61500
rect 17012 61444 17016 61500
rect 16952 61440 17016 61444
rect 17032 61500 17096 61504
rect 17032 61444 17036 61500
rect 17036 61444 17092 61500
rect 17092 61444 17096 61500
rect 17032 61440 17096 61444
rect 17112 61500 17176 61504
rect 17112 61444 17116 61500
rect 17116 61444 17172 61500
rect 17172 61444 17176 61500
rect 17112 61440 17176 61444
rect 17192 61500 17256 61504
rect 17192 61444 17196 61500
rect 17196 61444 17252 61500
rect 17252 61444 17256 61500
rect 17192 61440 17256 61444
rect 2612 60956 2676 60960
rect 2612 60900 2616 60956
rect 2616 60900 2672 60956
rect 2672 60900 2676 60956
rect 2612 60896 2676 60900
rect 2692 60956 2756 60960
rect 2692 60900 2696 60956
rect 2696 60900 2752 60956
rect 2752 60900 2756 60956
rect 2692 60896 2756 60900
rect 2772 60956 2836 60960
rect 2772 60900 2776 60956
rect 2776 60900 2832 60956
rect 2832 60900 2836 60956
rect 2772 60896 2836 60900
rect 2852 60956 2916 60960
rect 2852 60900 2856 60956
rect 2856 60900 2912 60956
rect 2912 60900 2916 60956
rect 2852 60896 2916 60900
rect 7612 60956 7676 60960
rect 7612 60900 7616 60956
rect 7616 60900 7672 60956
rect 7672 60900 7676 60956
rect 7612 60896 7676 60900
rect 7692 60956 7756 60960
rect 7692 60900 7696 60956
rect 7696 60900 7752 60956
rect 7752 60900 7756 60956
rect 7692 60896 7756 60900
rect 7772 60956 7836 60960
rect 7772 60900 7776 60956
rect 7776 60900 7832 60956
rect 7832 60900 7836 60956
rect 7772 60896 7836 60900
rect 7852 60956 7916 60960
rect 7852 60900 7856 60956
rect 7856 60900 7912 60956
rect 7912 60900 7916 60956
rect 7852 60896 7916 60900
rect 12612 60956 12676 60960
rect 12612 60900 12616 60956
rect 12616 60900 12672 60956
rect 12672 60900 12676 60956
rect 12612 60896 12676 60900
rect 12692 60956 12756 60960
rect 12692 60900 12696 60956
rect 12696 60900 12752 60956
rect 12752 60900 12756 60956
rect 12692 60896 12756 60900
rect 12772 60956 12836 60960
rect 12772 60900 12776 60956
rect 12776 60900 12832 60956
rect 12832 60900 12836 60956
rect 12772 60896 12836 60900
rect 12852 60956 12916 60960
rect 12852 60900 12856 60956
rect 12856 60900 12912 60956
rect 12912 60900 12916 60956
rect 12852 60896 12916 60900
rect 17612 60956 17676 60960
rect 17612 60900 17616 60956
rect 17616 60900 17672 60956
rect 17672 60900 17676 60956
rect 17612 60896 17676 60900
rect 17692 60956 17756 60960
rect 17692 60900 17696 60956
rect 17696 60900 17752 60956
rect 17752 60900 17756 60956
rect 17692 60896 17756 60900
rect 17772 60956 17836 60960
rect 17772 60900 17776 60956
rect 17776 60900 17832 60956
rect 17832 60900 17836 60956
rect 17772 60896 17836 60900
rect 17852 60956 17916 60960
rect 17852 60900 17856 60956
rect 17856 60900 17912 60956
rect 17912 60900 17916 60956
rect 17852 60896 17916 60900
rect 1952 60412 2016 60416
rect 1952 60356 1956 60412
rect 1956 60356 2012 60412
rect 2012 60356 2016 60412
rect 1952 60352 2016 60356
rect 2032 60412 2096 60416
rect 2032 60356 2036 60412
rect 2036 60356 2092 60412
rect 2092 60356 2096 60412
rect 2032 60352 2096 60356
rect 2112 60412 2176 60416
rect 2112 60356 2116 60412
rect 2116 60356 2172 60412
rect 2172 60356 2176 60412
rect 2112 60352 2176 60356
rect 2192 60412 2256 60416
rect 2192 60356 2196 60412
rect 2196 60356 2252 60412
rect 2252 60356 2256 60412
rect 2192 60352 2256 60356
rect 6952 60412 7016 60416
rect 6952 60356 6956 60412
rect 6956 60356 7012 60412
rect 7012 60356 7016 60412
rect 6952 60352 7016 60356
rect 7032 60412 7096 60416
rect 7032 60356 7036 60412
rect 7036 60356 7092 60412
rect 7092 60356 7096 60412
rect 7032 60352 7096 60356
rect 7112 60412 7176 60416
rect 7112 60356 7116 60412
rect 7116 60356 7172 60412
rect 7172 60356 7176 60412
rect 7112 60352 7176 60356
rect 7192 60412 7256 60416
rect 7192 60356 7196 60412
rect 7196 60356 7252 60412
rect 7252 60356 7256 60412
rect 7192 60352 7256 60356
rect 11952 60412 12016 60416
rect 11952 60356 11956 60412
rect 11956 60356 12012 60412
rect 12012 60356 12016 60412
rect 11952 60352 12016 60356
rect 12032 60412 12096 60416
rect 12032 60356 12036 60412
rect 12036 60356 12092 60412
rect 12092 60356 12096 60412
rect 12032 60352 12096 60356
rect 12112 60412 12176 60416
rect 12112 60356 12116 60412
rect 12116 60356 12172 60412
rect 12172 60356 12176 60412
rect 12112 60352 12176 60356
rect 12192 60412 12256 60416
rect 12192 60356 12196 60412
rect 12196 60356 12252 60412
rect 12252 60356 12256 60412
rect 12192 60352 12256 60356
rect 16952 60412 17016 60416
rect 16952 60356 16956 60412
rect 16956 60356 17012 60412
rect 17012 60356 17016 60412
rect 16952 60352 17016 60356
rect 17032 60412 17096 60416
rect 17032 60356 17036 60412
rect 17036 60356 17092 60412
rect 17092 60356 17096 60412
rect 17032 60352 17096 60356
rect 17112 60412 17176 60416
rect 17112 60356 17116 60412
rect 17116 60356 17172 60412
rect 17172 60356 17176 60412
rect 17112 60352 17176 60356
rect 17192 60412 17256 60416
rect 17192 60356 17196 60412
rect 17196 60356 17252 60412
rect 17252 60356 17256 60412
rect 17192 60352 17256 60356
rect 16436 60072 16500 60076
rect 16436 60016 16450 60072
rect 16450 60016 16500 60072
rect 16436 60012 16500 60016
rect 9076 59876 9140 59940
rect 2612 59868 2676 59872
rect 2612 59812 2616 59868
rect 2616 59812 2672 59868
rect 2672 59812 2676 59868
rect 2612 59808 2676 59812
rect 2692 59868 2756 59872
rect 2692 59812 2696 59868
rect 2696 59812 2752 59868
rect 2752 59812 2756 59868
rect 2692 59808 2756 59812
rect 2772 59868 2836 59872
rect 2772 59812 2776 59868
rect 2776 59812 2832 59868
rect 2832 59812 2836 59868
rect 2772 59808 2836 59812
rect 2852 59868 2916 59872
rect 2852 59812 2856 59868
rect 2856 59812 2912 59868
rect 2912 59812 2916 59868
rect 2852 59808 2916 59812
rect 7612 59868 7676 59872
rect 7612 59812 7616 59868
rect 7616 59812 7672 59868
rect 7672 59812 7676 59868
rect 7612 59808 7676 59812
rect 7692 59868 7756 59872
rect 7692 59812 7696 59868
rect 7696 59812 7752 59868
rect 7752 59812 7756 59868
rect 7692 59808 7756 59812
rect 7772 59868 7836 59872
rect 7772 59812 7776 59868
rect 7776 59812 7832 59868
rect 7832 59812 7836 59868
rect 7772 59808 7836 59812
rect 7852 59868 7916 59872
rect 7852 59812 7856 59868
rect 7856 59812 7912 59868
rect 7912 59812 7916 59868
rect 7852 59808 7916 59812
rect 12612 59868 12676 59872
rect 12612 59812 12616 59868
rect 12616 59812 12672 59868
rect 12672 59812 12676 59868
rect 12612 59808 12676 59812
rect 12692 59868 12756 59872
rect 12692 59812 12696 59868
rect 12696 59812 12752 59868
rect 12752 59812 12756 59868
rect 12692 59808 12756 59812
rect 12772 59868 12836 59872
rect 12772 59812 12776 59868
rect 12776 59812 12832 59868
rect 12832 59812 12836 59868
rect 12772 59808 12836 59812
rect 12852 59868 12916 59872
rect 12852 59812 12856 59868
rect 12856 59812 12912 59868
rect 12912 59812 12916 59868
rect 12852 59808 12916 59812
rect 17612 59868 17676 59872
rect 17612 59812 17616 59868
rect 17616 59812 17672 59868
rect 17672 59812 17676 59868
rect 17612 59808 17676 59812
rect 17692 59868 17756 59872
rect 17692 59812 17696 59868
rect 17696 59812 17752 59868
rect 17752 59812 17756 59868
rect 17692 59808 17756 59812
rect 17772 59868 17836 59872
rect 17772 59812 17776 59868
rect 17776 59812 17832 59868
rect 17832 59812 17836 59868
rect 17772 59808 17836 59812
rect 17852 59868 17916 59872
rect 17852 59812 17856 59868
rect 17856 59812 17912 59868
rect 17912 59812 17916 59868
rect 17852 59808 17916 59812
rect 1952 59324 2016 59328
rect 1952 59268 1956 59324
rect 1956 59268 2012 59324
rect 2012 59268 2016 59324
rect 1952 59264 2016 59268
rect 2032 59324 2096 59328
rect 2032 59268 2036 59324
rect 2036 59268 2092 59324
rect 2092 59268 2096 59324
rect 2032 59264 2096 59268
rect 2112 59324 2176 59328
rect 2112 59268 2116 59324
rect 2116 59268 2172 59324
rect 2172 59268 2176 59324
rect 2112 59264 2176 59268
rect 2192 59324 2256 59328
rect 2192 59268 2196 59324
rect 2196 59268 2252 59324
rect 2252 59268 2256 59324
rect 2192 59264 2256 59268
rect 6952 59324 7016 59328
rect 6952 59268 6956 59324
rect 6956 59268 7012 59324
rect 7012 59268 7016 59324
rect 6952 59264 7016 59268
rect 7032 59324 7096 59328
rect 7032 59268 7036 59324
rect 7036 59268 7092 59324
rect 7092 59268 7096 59324
rect 7032 59264 7096 59268
rect 7112 59324 7176 59328
rect 7112 59268 7116 59324
rect 7116 59268 7172 59324
rect 7172 59268 7176 59324
rect 7112 59264 7176 59268
rect 7192 59324 7256 59328
rect 7192 59268 7196 59324
rect 7196 59268 7252 59324
rect 7252 59268 7256 59324
rect 7192 59264 7256 59268
rect 11952 59324 12016 59328
rect 11952 59268 11956 59324
rect 11956 59268 12012 59324
rect 12012 59268 12016 59324
rect 11952 59264 12016 59268
rect 12032 59324 12096 59328
rect 12032 59268 12036 59324
rect 12036 59268 12092 59324
rect 12092 59268 12096 59324
rect 12032 59264 12096 59268
rect 12112 59324 12176 59328
rect 12112 59268 12116 59324
rect 12116 59268 12172 59324
rect 12172 59268 12176 59324
rect 12112 59264 12176 59268
rect 12192 59324 12256 59328
rect 12192 59268 12196 59324
rect 12196 59268 12252 59324
rect 12252 59268 12256 59324
rect 12192 59264 12256 59268
rect 16952 59324 17016 59328
rect 16952 59268 16956 59324
rect 16956 59268 17012 59324
rect 17012 59268 17016 59324
rect 16952 59264 17016 59268
rect 17032 59324 17096 59328
rect 17032 59268 17036 59324
rect 17036 59268 17092 59324
rect 17092 59268 17096 59324
rect 17032 59264 17096 59268
rect 17112 59324 17176 59328
rect 17112 59268 17116 59324
rect 17116 59268 17172 59324
rect 17172 59268 17176 59324
rect 17112 59264 17176 59268
rect 17192 59324 17256 59328
rect 17192 59268 17196 59324
rect 17196 59268 17252 59324
rect 17252 59268 17256 59324
rect 17192 59264 17256 59268
rect 13676 58848 13740 58852
rect 13676 58792 13726 58848
rect 13726 58792 13740 58848
rect 13676 58788 13740 58792
rect 2612 58780 2676 58784
rect 2612 58724 2616 58780
rect 2616 58724 2672 58780
rect 2672 58724 2676 58780
rect 2612 58720 2676 58724
rect 2692 58780 2756 58784
rect 2692 58724 2696 58780
rect 2696 58724 2752 58780
rect 2752 58724 2756 58780
rect 2692 58720 2756 58724
rect 2772 58780 2836 58784
rect 2772 58724 2776 58780
rect 2776 58724 2832 58780
rect 2832 58724 2836 58780
rect 2772 58720 2836 58724
rect 2852 58780 2916 58784
rect 2852 58724 2856 58780
rect 2856 58724 2912 58780
rect 2912 58724 2916 58780
rect 2852 58720 2916 58724
rect 7612 58780 7676 58784
rect 7612 58724 7616 58780
rect 7616 58724 7672 58780
rect 7672 58724 7676 58780
rect 7612 58720 7676 58724
rect 7692 58780 7756 58784
rect 7692 58724 7696 58780
rect 7696 58724 7752 58780
rect 7752 58724 7756 58780
rect 7692 58720 7756 58724
rect 7772 58780 7836 58784
rect 7772 58724 7776 58780
rect 7776 58724 7832 58780
rect 7832 58724 7836 58780
rect 7772 58720 7836 58724
rect 7852 58780 7916 58784
rect 7852 58724 7856 58780
rect 7856 58724 7912 58780
rect 7912 58724 7916 58780
rect 7852 58720 7916 58724
rect 12612 58780 12676 58784
rect 12612 58724 12616 58780
rect 12616 58724 12672 58780
rect 12672 58724 12676 58780
rect 12612 58720 12676 58724
rect 12692 58780 12756 58784
rect 12692 58724 12696 58780
rect 12696 58724 12752 58780
rect 12752 58724 12756 58780
rect 12692 58720 12756 58724
rect 12772 58780 12836 58784
rect 12772 58724 12776 58780
rect 12776 58724 12832 58780
rect 12832 58724 12836 58780
rect 12772 58720 12836 58724
rect 12852 58780 12916 58784
rect 12852 58724 12856 58780
rect 12856 58724 12912 58780
rect 12912 58724 12916 58780
rect 12852 58720 12916 58724
rect 17612 58780 17676 58784
rect 17612 58724 17616 58780
rect 17616 58724 17672 58780
rect 17672 58724 17676 58780
rect 17612 58720 17676 58724
rect 17692 58780 17756 58784
rect 17692 58724 17696 58780
rect 17696 58724 17752 58780
rect 17752 58724 17756 58780
rect 17692 58720 17756 58724
rect 17772 58780 17836 58784
rect 17772 58724 17776 58780
rect 17776 58724 17832 58780
rect 17832 58724 17836 58780
rect 17772 58720 17836 58724
rect 17852 58780 17916 58784
rect 17852 58724 17856 58780
rect 17856 58724 17912 58780
rect 17912 58724 17916 58780
rect 17852 58720 17916 58724
rect 1952 58236 2016 58240
rect 1952 58180 1956 58236
rect 1956 58180 2012 58236
rect 2012 58180 2016 58236
rect 1952 58176 2016 58180
rect 2032 58236 2096 58240
rect 2032 58180 2036 58236
rect 2036 58180 2092 58236
rect 2092 58180 2096 58236
rect 2032 58176 2096 58180
rect 2112 58236 2176 58240
rect 2112 58180 2116 58236
rect 2116 58180 2172 58236
rect 2172 58180 2176 58236
rect 2112 58176 2176 58180
rect 2192 58236 2256 58240
rect 2192 58180 2196 58236
rect 2196 58180 2252 58236
rect 2252 58180 2256 58236
rect 2192 58176 2256 58180
rect 6952 58236 7016 58240
rect 6952 58180 6956 58236
rect 6956 58180 7012 58236
rect 7012 58180 7016 58236
rect 6952 58176 7016 58180
rect 7032 58236 7096 58240
rect 7032 58180 7036 58236
rect 7036 58180 7092 58236
rect 7092 58180 7096 58236
rect 7032 58176 7096 58180
rect 7112 58236 7176 58240
rect 7112 58180 7116 58236
rect 7116 58180 7172 58236
rect 7172 58180 7176 58236
rect 7112 58176 7176 58180
rect 7192 58236 7256 58240
rect 7192 58180 7196 58236
rect 7196 58180 7252 58236
rect 7252 58180 7256 58236
rect 7192 58176 7256 58180
rect 11952 58236 12016 58240
rect 11952 58180 11956 58236
rect 11956 58180 12012 58236
rect 12012 58180 12016 58236
rect 11952 58176 12016 58180
rect 12032 58236 12096 58240
rect 12032 58180 12036 58236
rect 12036 58180 12092 58236
rect 12092 58180 12096 58236
rect 12032 58176 12096 58180
rect 12112 58236 12176 58240
rect 12112 58180 12116 58236
rect 12116 58180 12172 58236
rect 12172 58180 12176 58236
rect 12112 58176 12176 58180
rect 12192 58236 12256 58240
rect 12192 58180 12196 58236
rect 12196 58180 12252 58236
rect 12252 58180 12256 58236
rect 12192 58176 12256 58180
rect 16952 58236 17016 58240
rect 16952 58180 16956 58236
rect 16956 58180 17012 58236
rect 17012 58180 17016 58236
rect 16952 58176 17016 58180
rect 17032 58236 17096 58240
rect 17032 58180 17036 58236
rect 17036 58180 17092 58236
rect 17092 58180 17096 58236
rect 17032 58176 17096 58180
rect 17112 58236 17176 58240
rect 17112 58180 17116 58236
rect 17116 58180 17172 58236
rect 17172 58180 17176 58236
rect 17112 58176 17176 58180
rect 17192 58236 17256 58240
rect 17192 58180 17196 58236
rect 17196 58180 17252 58236
rect 17252 58180 17256 58236
rect 17192 58176 17256 58180
rect 2612 57692 2676 57696
rect 2612 57636 2616 57692
rect 2616 57636 2672 57692
rect 2672 57636 2676 57692
rect 2612 57632 2676 57636
rect 2692 57692 2756 57696
rect 2692 57636 2696 57692
rect 2696 57636 2752 57692
rect 2752 57636 2756 57692
rect 2692 57632 2756 57636
rect 2772 57692 2836 57696
rect 2772 57636 2776 57692
rect 2776 57636 2832 57692
rect 2832 57636 2836 57692
rect 2772 57632 2836 57636
rect 2852 57692 2916 57696
rect 2852 57636 2856 57692
rect 2856 57636 2912 57692
rect 2912 57636 2916 57692
rect 2852 57632 2916 57636
rect 7612 57692 7676 57696
rect 7612 57636 7616 57692
rect 7616 57636 7672 57692
rect 7672 57636 7676 57692
rect 7612 57632 7676 57636
rect 7692 57692 7756 57696
rect 7692 57636 7696 57692
rect 7696 57636 7752 57692
rect 7752 57636 7756 57692
rect 7692 57632 7756 57636
rect 7772 57692 7836 57696
rect 7772 57636 7776 57692
rect 7776 57636 7832 57692
rect 7832 57636 7836 57692
rect 7772 57632 7836 57636
rect 7852 57692 7916 57696
rect 7852 57636 7856 57692
rect 7856 57636 7912 57692
rect 7912 57636 7916 57692
rect 7852 57632 7916 57636
rect 12612 57692 12676 57696
rect 12612 57636 12616 57692
rect 12616 57636 12672 57692
rect 12672 57636 12676 57692
rect 12612 57632 12676 57636
rect 12692 57692 12756 57696
rect 12692 57636 12696 57692
rect 12696 57636 12752 57692
rect 12752 57636 12756 57692
rect 12692 57632 12756 57636
rect 12772 57692 12836 57696
rect 12772 57636 12776 57692
rect 12776 57636 12832 57692
rect 12832 57636 12836 57692
rect 12772 57632 12836 57636
rect 12852 57692 12916 57696
rect 12852 57636 12856 57692
rect 12856 57636 12912 57692
rect 12912 57636 12916 57692
rect 12852 57632 12916 57636
rect 17612 57692 17676 57696
rect 17612 57636 17616 57692
rect 17616 57636 17672 57692
rect 17672 57636 17676 57692
rect 17612 57632 17676 57636
rect 17692 57692 17756 57696
rect 17692 57636 17696 57692
rect 17696 57636 17752 57692
rect 17752 57636 17756 57692
rect 17692 57632 17756 57636
rect 17772 57692 17836 57696
rect 17772 57636 17776 57692
rect 17776 57636 17832 57692
rect 17832 57636 17836 57692
rect 17772 57632 17836 57636
rect 17852 57692 17916 57696
rect 17852 57636 17856 57692
rect 17856 57636 17912 57692
rect 17912 57636 17916 57692
rect 17852 57632 17916 57636
rect 1952 57148 2016 57152
rect 1952 57092 1956 57148
rect 1956 57092 2012 57148
rect 2012 57092 2016 57148
rect 1952 57088 2016 57092
rect 2032 57148 2096 57152
rect 2032 57092 2036 57148
rect 2036 57092 2092 57148
rect 2092 57092 2096 57148
rect 2032 57088 2096 57092
rect 2112 57148 2176 57152
rect 2112 57092 2116 57148
rect 2116 57092 2172 57148
rect 2172 57092 2176 57148
rect 2112 57088 2176 57092
rect 2192 57148 2256 57152
rect 2192 57092 2196 57148
rect 2196 57092 2252 57148
rect 2252 57092 2256 57148
rect 2192 57088 2256 57092
rect 6952 57148 7016 57152
rect 6952 57092 6956 57148
rect 6956 57092 7012 57148
rect 7012 57092 7016 57148
rect 6952 57088 7016 57092
rect 7032 57148 7096 57152
rect 7032 57092 7036 57148
rect 7036 57092 7092 57148
rect 7092 57092 7096 57148
rect 7032 57088 7096 57092
rect 7112 57148 7176 57152
rect 7112 57092 7116 57148
rect 7116 57092 7172 57148
rect 7172 57092 7176 57148
rect 7112 57088 7176 57092
rect 7192 57148 7256 57152
rect 7192 57092 7196 57148
rect 7196 57092 7252 57148
rect 7252 57092 7256 57148
rect 7192 57088 7256 57092
rect 11952 57148 12016 57152
rect 11952 57092 11956 57148
rect 11956 57092 12012 57148
rect 12012 57092 12016 57148
rect 11952 57088 12016 57092
rect 12032 57148 12096 57152
rect 12032 57092 12036 57148
rect 12036 57092 12092 57148
rect 12092 57092 12096 57148
rect 12032 57088 12096 57092
rect 12112 57148 12176 57152
rect 12112 57092 12116 57148
rect 12116 57092 12172 57148
rect 12172 57092 12176 57148
rect 12112 57088 12176 57092
rect 12192 57148 12256 57152
rect 12192 57092 12196 57148
rect 12196 57092 12252 57148
rect 12252 57092 12256 57148
rect 12192 57088 12256 57092
rect 16952 57148 17016 57152
rect 16952 57092 16956 57148
rect 16956 57092 17012 57148
rect 17012 57092 17016 57148
rect 16952 57088 17016 57092
rect 17032 57148 17096 57152
rect 17032 57092 17036 57148
rect 17036 57092 17092 57148
rect 17092 57092 17096 57148
rect 17032 57088 17096 57092
rect 17112 57148 17176 57152
rect 17112 57092 17116 57148
rect 17116 57092 17172 57148
rect 17172 57092 17176 57148
rect 17112 57088 17176 57092
rect 17192 57148 17256 57152
rect 17192 57092 17196 57148
rect 17196 57092 17252 57148
rect 17252 57092 17256 57148
rect 17192 57088 17256 57092
rect 6316 56612 6380 56676
rect 2612 56604 2676 56608
rect 2612 56548 2616 56604
rect 2616 56548 2672 56604
rect 2672 56548 2676 56604
rect 2612 56544 2676 56548
rect 2692 56604 2756 56608
rect 2692 56548 2696 56604
rect 2696 56548 2752 56604
rect 2752 56548 2756 56604
rect 2692 56544 2756 56548
rect 2772 56604 2836 56608
rect 2772 56548 2776 56604
rect 2776 56548 2832 56604
rect 2832 56548 2836 56604
rect 2772 56544 2836 56548
rect 2852 56604 2916 56608
rect 2852 56548 2856 56604
rect 2856 56548 2912 56604
rect 2912 56548 2916 56604
rect 2852 56544 2916 56548
rect 7612 56604 7676 56608
rect 7612 56548 7616 56604
rect 7616 56548 7672 56604
rect 7672 56548 7676 56604
rect 7612 56544 7676 56548
rect 7692 56604 7756 56608
rect 7692 56548 7696 56604
rect 7696 56548 7752 56604
rect 7752 56548 7756 56604
rect 7692 56544 7756 56548
rect 7772 56604 7836 56608
rect 7772 56548 7776 56604
rect 7776 56548 7832 56604
rect 7832 56548 7836 56604
rect 7772 56544 7836 56548
rect 7852 56604 7916 56608
rect 7852 56548 7856 56604
rect 7856 56548 7912 56604
rect 7912 56548 7916 56604
rect 7852 56544 7916 56548
rect 12612 56604 12676 56608
rect 12612 56548 12616 56604
rect 12616 56548 12672 56604
rect 12672 56548 12676 56604
rect 12612 56544 12676 56548
rect 12692 56604 12756 56608
rect 12692 56548 12696 56604
rect 12696 56548 12752 56604
rect 12752 56548 12756 56604
rect 12692 56544 12756 56548
rect 12772 56604 12836 56608
rect 12772 56548 12776 56604
rect 12776 56548 12832 56604
rect 12832 56548 12836 56604
rect 12772 56544 12836 56548
rect 12852 56604 12916 56608
rect 12852 56548 12856 56604
rect 12856 56548 12912 56604
rect 12912 56548 12916 56604
rect 12852 56544 12916 56548
rect 17612 56604 17676 56608
rect 17612 56548 17616 56604
rect 17616 56548 17672 56604
rect 17672 56548 17676 56604
rect 17612 56544 17676 56548
rect 17692 56604 17756 56608
rect 17692 56548 17696 56604
rect 17696 56548 17752 56604
rect 17752 56548 17756 56604
rect 17692 56544 17756 56548
rect 17772 56604 17836 56608
rect 17772 56548 17776 56604
rect 17776 56548 17832 56604
rect 17832 56548 17836 56604
rect 17772 56544 17836 56548
rect 17852 56604 17916 56608
rect 17852 56548 17856 56604
rect 17856 56548 17912 56604
rect 17912 56548 17916 56604
rect 17852 56544 17916 56548
rect 1952 56060 2016 56064
rect 1952 56004 1956 56060
rect 1956 56004 2012 56060
rect 2012 56004 2016 56060
rect 1952 56000 2016 56004
rect 2032 56060 2096 56064
rect 2032 56004 2036 56060
rect 2036 56004 2092 56060
rect 2092 56004 2096 56060
rect 2032 56000 2096 56004
rect 2112 56060 2176 56064
rect 2112 56004 2116 56060
rect 2116 56004 2172 56060
rect 2172 56004 2176 56060
rect 2112 56000 2176 56004
rect 2192 56060 2256 56064
rect 2192 56004 2196 56060
rect 2196 56004 2252 56060
rect 2252 56004 2256 56060
rect 2192 56000 2256 56004
rect 6952 56060 7016 56064
rect 6952 56004 6956 56060
rect 6956 56004 7012 56060
rect 7012 56004 7016 56060
rect 6952 56000 7016 56004
rect 7032 56060 7096 56064
rect 7032 56004 7036 56060
rect 7036 56004 7092 56060
rect 7092 56004 7096 56060
rect 7032 56000 7096 56004
rect 7112 56060 7176 56064
rect 7112 56004 7116 56060
rect 7116 56004 7172 56060
rect 7172 56004 7176 56060
rect 7112 56000 7176 56004
rect 7192 56060 7256 56064
rect 7192 56004 7196 56060
rect 7196 56004 7252 56060
rect 7252 56004 7256 56060
rect 7192 56000 7256 56004
rect 11952 56060 12016 56064
rect 11952 56004 11956 56060
rect 11956 56004 12012 56060
rect 12012 56004 12016 56060
rect 11952 56000 12016 56004
rect 12032 56060 12096 56064
rect 12032 56004 12036 56060
rect 12036 56004 12092 56060
rect 12092 56004 12096 56060
rect 12032 56000 12096 56004
rect 12112 56060 12176 56064
rect 12112 56004 12116 56060
rect 12116 56004 12172 56060
rect 12172 56004 12176 56060
rect 12112 56000 12176 56004
rect 12192 56060 12256 56064
rect 12192 56004 12196 56060
rect 12196 56004 12252 56060
rect 12252 56004 12256 56060
rect 12192 56000 12256 56004
rect 16952 56060 17016 56064
rect 16952 56004 16956 56060
rect 16956 56004 17012 56060
rect 17012 56004 17016 56060
rect 16952 56000 17016 56004
rect 17032 56060 17096 56064
rect 17032 56004 17036 56060
rect 17036 56004 17092 56060
rect 17092 56004 17096 56060
rect 17032 56000 17096 56004
rect 17112 56060 17176 56064
rect 17112 56004 17116 56060
rect 17116 56004 17172 56060
rect 17172 56004 17176 56060
rect 17112 56000 17176 56004
rect 17192 56060 17256 56064
rect 17192 56004 17196 56060
rect 17196 56004 17252 56060
rect 17252 56004 17256 56060
rect 17192 56000 17256 56004
rect 1532 55660 1596 55724
rect 14412 55660 14476 55724
rect 16620 55660 16684 55724
rect 2612 55516 2676 55520
rect 2612 55460 2616 55516
rect 2616 55460 2672 55516
rect 2672 55460 2676 55516
rect 2612 55456 2676 55460
rect 2692 55516 2756 55520
rect 2692 55460 2696 55516
rect 2696 55460 2752 55516
rect 2752 55460 2756 55516
rect 2692 55456 2756 55460
rect 2772 55516 2836 55520
rect 2772 55460 2776 55516
rect 2776 55460 2832 55516
rect 2832 55460 2836 55516
rect 2772 55456 2836 55460
rect 2852 55516 2916 55520
rect 2852 55460 2856 55516
rect 2856 55460 2912 55516
rect 2912 55460 2916 55516
rect 2852 55456 2916 55460
rect 7612 55516 7676 55520
rect 7612 55460 7616 55516
rect 7616 55460 7672 55516
rect 7672 55460 7676 55516
rect 7612 55456 7676 55460
rect 7692 55516 7756 55520
rect 7692 55460 7696 55516
rect 7696 55460 7752 55516
rect 7752 55460 7756 55516
rect 7692 55456 7756 55460
rect 7772 55516 7836 55520
rect 7772 55460 7776 55516
rect 7776 55460 7832 55516
rect 7832 55460 7836 55516
rect 7772 55456 7836 55460
rect 7852 55516 7916 55520
rect 7852 55460 7856 55516
rect 7856 55460 7912 55516
rect 7912 55460 7916 55516
rect 7852 55456 7916 55460
rect 12612 55516 12676 55520
rect 12612 55460 12616 55516
rect 12616 55460 12672 55516
rect 12672 55460 12676 55516
rect 12612 55456 12676 55460
rect 12692 55516 12756 55520
rect 12692 55460 12696 55516
rect 12696 55460 12752 55516
rect 12752 55460 12756 55516
rect 12692 55456 12756 55460
rect 12772 55516 12836 55520
rect 12772 55460 12776 55516
rect 12776 55460 12832 55516
rect 12832 55460 12836 55516
rect 12772 55456 12836 55460
rect 12852 55516 12916 55520
rect 12852 55460 12856 55516
rect 12856 55460 12912 55516
rect 12912 55460 12916 55516
rect 12852 55456 12916 55460
rect 17612 55516 17676 55520
rect 17612 55460 17616 55516
rect 17616 55460 17672 55516
rect 17672 55460 17676 55516
rect 17612 55456 17676 55460
rect 17692 55516 17756 55520
rect 17692 55460 17696 55516
rect 17696 55460 17752 55516
rect 17752 55460 17756 55516
rect 17692 55456 17756 55460
rect 17772 55516 17836 55520
rect 17772 55460 17776 55516
rect 17776 55460 17832 55516
rect 17832 55460 17836 55516
rect 17772 55456 17836 55460
rect 17852 55516 17916 55520
rect 17852 55460 17856 55516
rect 17856 55460 17912 55516
rect 17912 55460 17916 55516
rect 17852 55456 17916 55460
rect 1952 54972 2016 54976
rect 1952 54916 1956 54972
rect 1956 54916 2012 54972
rect 2012 54916 2016 54972
rect 1952 54912 2016 54916
rect 2032 54972 2096 54976
rect 2032 54916 2036 54972
rect 2036 54916 2092 54972
rect 2092 54916 2096 54972
rect 2032 54912 2096 54916
rect 2112 54972 2176 54976
rect 2112 54916 2116 54972
rect 2116 54916 2172 54972
rect 2172 54916 2176 54972
rect 2112 54912 2176 54916
rect 2192 54972 2256 54976
rect 2192 54916 2196 54972
rect 2196 54916 2252 54972
rect 2252 54916 2256 54972
rect 2192 54912 2256 54916
rect 6952 54972 7016 54976
rect 6952 54916 6956 54972
rect 6956 54916 7012 54972
rect 7012 54916 7016 54972
rect 6952 54912 7016 54916
rect 7032 54972 7096 54976
rect 7032 54916 7036 54972
rect 7036 54916 7092 54972
rect 7092 54916 7096 54972
rect 7032 54912 7096 54916
rect 7112 54972 7176 54976
rect 7112 54916 7116 54972
rect 7116 54916 7172 54972
rect 7172 54916 7176 54972
rect 7112 54912 7176 54916
rect 7192 54972 7256 54976
rect 7192 54916 7196 54972
rect 7196 54916 7252 54972
rect 7252 54916 7256 54972
rect 7192 54912 7256 54916
rect 11952 54972 12016 54976
rect 11952 54916 11956 54972
rect 11956 54916 12012 54972
rect 12012 54916 12016 54972
rect 11952 54912 12016 54916
rect 12032 54972 12096 54976
rect 12032 54916 12036 54972
rect 12036 54916 12092 54972
rect 12092 54916 12096 54972
rect 12032 54912 12096 54916
rect 12112 54972 12176 54976
rect 12112 54916 12116 54972
rect 12116 54916 12172 54972
rect 12172 54916 12176 54972
rect 12112 54912 12176 54916
rect 12192 54972 12256 54976
rect 12192 54916 12196 54972
rect 12196 54916 12252 54972
rect 12252 54916 12256 54972
rect 12192 54912 12256 54916
rect 16952 54972 17016 54976
rect 16952 54916 16956 54972
rect 16956 54916 17012 54972
rect 17012 54916 17016 54972
rect 16952 54912 17016 54916
rect 17032 54972 17096 54976
rect 17032 54916 17036 54972
rect 17036 54916 17092 54972
rect 17092 54916 17096 54972
rect 17032 54912 17096 54916
rect 17112 54972 17176 54976
rect 17112 54916 17116 54972
rect 17116 54916 17172 54972
rect 17172 54916 17176 54972
rect 17112 54912 17176 54916
rect 17192 54972 17256 54976
rect 17192 54916 17196 54972
rect 17196 54916 17252 54972
rect 17252 54916 17256 54972
rect 17192 54912 17256 54916
rect 2612 54428 2676 54432
rect 2612 54372 2616 54428
rect 2616 54372 2672 54428
rect 2672 54372 2676 54428
rect 2612 54368 2676 54372
rect 2692 54428 2756 54432
rect 2692 54372 2696 54428
rect 2696 54372 2752 54428
rect 2752 54372 2756 54428
rect 2692 54368 2756 54372
rect 2772 54428 2836 54432
rect 2772 54372 2776 54428
rect 2776 54372 2832 54428
rect 2832 54372 2836 54428
rect 2772 54368 2836 54372
rect 2852 54428 2916 54432
rect 2852 54372 2856 54428
rect 2856 54372 2912 54428
rect 2912 54372 2916 54428
rect 2852 54368 2916 54372
rect 7612 54428 7676 54432
rect 7612 54372 7616 54428
rect 7616 54372 7672 54428
rect 7672 54372 7676 54428
rect 7612 54368 7676 54372
rect 7692 54428 7756 54432
rect 7692 54372 7696 54428
rect 7696 54372 7752 54428
rect 7752 54372 7756 54428
rect 7692 54368 7756 54372
rect 7772 54428 7836 54432
rect 7772 54372 7776 54428
rect 7776 54372 7832 54428
rect 7832 54372 7836 54428
rect 7772 54368 7836 54372
rect 7852 54428 7916 54432
rect 7852 54372 7856 54428
rect 7856 54372 7912 54428
rect 7912 54372 7916 54428
rect 7852 54368 7916 54372
rect 12612 54428 12676 54432
rect 12612 54372 12616 54428
rect 12616 54372 12672 54428
rect 12672 54372 12676 54428
rect 12612 54368 12676 54372
rect 12692 54428 12756 54432
rect 12692 54372 12696 54428
rect 12696 54372 12752 54428
rect 12752 54372 12756 54428
rect 12692 54368 12756 54372
rect 12772 54428 12836 54432
rect 12772 54372 12776 54428
rect 12776 54372 12832 54428
rect 12832 54372 12836 54428
rect 12772 54368 12836 54372
rect 12852 54428 12916 54432
rect 12852 54372 12856 54428
rect 12856 54372 12912 54428
rect 12912 54372 12916 54428
rect 12852 54368 12916 54372
rect 17612 54428 17676 54432
rect 17612 54372 17616 54428
rect 17616 54372 17672 54428
rect 17672 54372 17676 54428
rect 17612 54368 17676 54372
rect 17692 54428 17756 54432
rect 17692 54372 17696 54428
rect 17696 54372 17752 54428
rect 17752 54372 17756 54428
rect 17692 54368 17756 54372
rect 17772 54428 17836 54432
rect 17772 54372 17776 54428
rect 17776 54372 17832 54428
rect 17832 54372 17836 54428
rect 17772 54368 17836 54372
rect 17852 54428 17916 54432
rect 17852 54372 17856 54428
rect 17856 54372 17912 54428
rect 17912 54372 17916 54428
rect 17852 54368 17916 54372
rect 10180 54028 10244 54092
rect 1952 53884 2016 53888
rect 1952 53828 1956 53884
rect 1956 53828 2012 53884
rect 2012 53828 2016 53884
rect 1952 53824 2016 53828
rect 2032 53884 2096 53888
rect 2032 53828 2036 53884
rect 2036 53828 2092 53884
rect 2092 53828 2096 53884
rect 2032 53824 2096 53828
rect 2112 53884 2176 53888
rect 2112 53828 2116 53884
rect 2116 53828 2172 53884
rect 2172 53828 2176 53884
rect 2112 53824 2176 53828
rect 2192 53884 2256 53888
rect 2192 53828 2196 53884
rect 2196 53828 2252 53884
rect 2252 53828 2256 53884
rect 2192 53824 2256 53828
rect 6952 53884 7016 53888
rect 6952 53828 6956 53884
rect 6956 53828 7012 53884
rect 7012 53828 7016 53884
rect 6952 53824 7016 53828
rect 7032 53884 7096 53888
rect 7032 53828 7036 53884
rect 7036 53828 7092 53884
rect 7092 53828 7096 53884
rect 7032 53824 7096 53828
rect 7112 53884 7176 53888
rect 7112 53828 7116 53884
rect 7116 53828 7172 53884
rect 7172 53828 7176 53884
rect 7112 53824 7176 53828
rect 7192 53884 7256 53888
rect 7192 53828 7196 53884
rect 7196 53828 7252 53884
rect 7252 53828 7256 53884
rect 7192 53824 7256 53828
rect 11952 53884 12016 53888
rect 11952 53828 11956 53884
rect 11956 53828 12012 53884
rect 12012 53828 12016 53884
rect 11952 53824 12016 53828
rect 12032 53884 12096 53888
rect 12032 53828 12036 53884
rect 12036 53828 12092 53884
rect 12092 53828 12096 53884
rect 12032 53824 12096 53828
rect 12112 53884 12176 53888
rect 12112 53828 12116 53884
rect 12116 53828 12172 53884
rect 12172 53828 12176 53884
rect 12112 53824 12176 53828
rect 12192 53884 12256 53888
rect 12192 53828 12196 53884
rect 12196 53828 12252 53884
rect 12252 53828 12256 53884
rect 12192 53824 12256 53828
rect 16952 53884 17016 53888
rect 16952 53828 16956 53884
rect 16956 53828 17012 53884
rect 17012 53828 17016 53884
rect 16952 53824 17016 53828
rect 17032 53884 17096 53888
rect 17032 53828 17036 53884
rect 17036 53828 17092 53884
rect 17092 53828 17096 53884
rect 17032 53824 17096 53828
rect 17112 53884 17176 53888
rect 17112 53828 17116 53884
rect 17116 53828 17172 53884
rect 17172 53828 17176 53884
rect 17112 53824 17176 53828
rect 17192 53884 17256 53888
rect 17192 53828 17196 53884
rect 17196 53828 17252 53884
rect 17252 53828 17256 53884
rect 17192 53824 17256 53828
rect 2612 53340 2676 53344
rect 2612 53284 2616 53340
rect 2616 53284 2672 53340
rect 2672 53284 2676 53340
rect 2612 53280 2676 53284
rect 2692 53340 2756 53344
rect 2692 53284 2696 53340
rect 2696 53284 2752 53340
rect 2752 53284 2756 53340
rect 2692 53280 2756 53284
rect 2772 53340 2836 53344
rect 2772 53284 2776 53340
rect 2776 53284 2832 53340
rect 2832 53284 2836 53340
rect 2772 53280 2836 53284
rect 2852 53340 2916 53344
rect 2852 53284 2856 53340
rect 2856 53284 2912 53340
rect 2912 53284 2916 53340
rect 2852 53280 2916 53284
rect 7612 53340 7676 53344
rect 7612 53284 7616 53340
rect 7616 53284 7672 53340
rect 7672 53284 7676 53340
rect 7612 53280 7676 53284
rect 7692 53340 7756 53344
rect 7692 53284 7696 53340
rect 7696 53284 7752 53340
rect 7752 53284 7756 53340
rect 7692 53280 7756 53284
rect 7772 53340 7836 53344
rect 7772 53284 7776 53340
rect 7776 53284 7832 53340
rect 7832 53284 7836 53340
rect 7772 53280 7836 53284
rect 7852 53340 7916 53344
rect 7852 53284 7856 53340
rect 7856 53284 7912 53340
rect 7912 53284 7916 53340
rect 7852 53280 7916 53284
rect 12612 53340 12676 53344
rect 12612 53284 12616 53340
rect 12616 53284 12672 53340
rect 12672 53284 12676 53340
rect 12612 53280 12676 53284
rect 12692 53340 12756 53344
rect 12692 53284 12696 53340
rect 12696 53284 12752 53340
rect 12752 53284 12756 53340
rect 12692 53280 12756 53284
rect 12772 53340 12836 53344
rect 12772 53284 12776 53340
rect 12776 53284 12832 53340
rect 12832 53284 12836 53340
rect 12772 53280 12836 53284
rect 12852 53340 12916 53344
rect 12852 53284 12856 53340
rect 12856 53284 12912 53340
rect 12912 53284 12916 53340
rect 12852 53280 12916 53284
rect 17612 53340 17676 53344
rect 17612 53284 17616 53340
rect 17616 53284 17672 53340
rect 17672 53284 17676 53340
rect 17612 53280 17676 53284
rect 17692 53340 17756 53344
rect 17692 53284 17696 53340
rect 17696 53284 17752 53340
rect 17752 53284 17756 53340
rect 17692 53280 17756 53284
rect 17772 53340 17836 53344
rect 17772 53284 17776 53340
rect 17776 53284 17832 53340
rect 17832 53284 17836 53340
rect 17772 53280 17836 53284
rect 17852 53340 17916 53344
rect 17852 53284 17856 53340
rect 17856 53284 17912 53340
rect 17912 53284 17916 53340
rect 17852 53280 17916 53284
rect 1952 52796 2016 52800
rect 1952 52740 1956 52796
rect 1956 52740 2012 52796
rect 2012 52740 2016 52796
rect 1952 52736 2016 52740
rect 2032 52796 2096 52800
rect 2032 52740 2036 52796
rect 2036 52740 2092 52796
rect 2092 52740 2096 52796
rect 2032 52736 2096 52740
rect 2112 52796 2176 52800
rect 2112 52740 2116 52796
rect 2116 52740 2172 52796
rect 2172 52740 2176 52796
rect 2112 52736 2176 52740
rect 2192 52796 2256 52800
rect 2192 52740 2196 52796
rect 2196 52740 2252 52796
rect 2252 52740 2256 52796
rect 2192 52736 2256 52740
rect 6952 52796 7016 52800
rect 6952 52740 6956 52796
rect 6956 52740 7012 52796
rect 7012 52740 7016 52796
rect 6952 52736 7016 52740
rect 7032 52796 7096 52800
rect 7032 52740 7036 52796
rect 7036 52740 7092 52796
rect 7092 52740 7096 52796
rect 7032 52736 7096 52740
rect 7112 52796 7176 52800
rect 7112 52740 7116 52796
rect 7116 52740 7172 52796
rect 7172 52740 7176 52796
rect 7112 52736 7176 52740
rect 7192 52796 7256 52800
rect 7192 52740 7196 52796
rect 7196 52740 7252 52796
rect 7252 52740 7256 52796
rect 7192 52736 7256 52740
rect 11952 52796 12016 52800
rect 11952 52740 11956 52796
rect 11956 52740 12012 52796
rect 12012 52740 12016 52796
rect 11952 52736 12016 52740
rect 12032 52796 12096 52800
rect 12032 52740 12036 52796
rect 12036 52740 12092 52796
rect 12092 52740 12096 52796
rect 12032 52736 12096 52740
rect 12112 52796 12176 52800
rect 12112 52740 12116 52796
rect 12116 52740 12172 52796
rect 12172 52740 12176 52796
rect 12112 52736 12176 52740
rect 12192 52796 12256 52800
rect 12192 52740 12196 52796
rect 12196 52740 12252 52796
rect 12252 52740 12256 52796
rect 12192 52736 12256 52740
rect 16952 52796 17016 52800
rect 16952 52740 16956 52796
rect 16956 52740 17012 52796
rect 17012 52740 17016 52796
rect 16952 52736 17016 52740
rect 17032 52796 17096 52800
rect 17032 52740 17036 52796
rect 17036 52740 17092 52796
rect 17092 52740 17096 52796
rect 17032 52736 17096 52740
rect 17112 52796 17176 52800
rect 17112 52740 17116 52796
rect 17116 52740 17172 52796
rect 17172 52740 17176 52796
rect 17112 52736 17176 52740
rect 17192 52796 17256 52800
rect 17192 52740 17196 52796
rect 17196 52740 17252 52796
rect 17252 52740 17256 52796
rect 17192 52736 17256 52740
rect 8524 52532 8588 52596
rect 10916 52396 10980 52460
rect 2612 52252 2676 52256
rect 2612 52196 2616 52252
rect 2616 52196 2672 52252
rect 2672 52196 2676 52252
rect 2612 52192 2676 52196
rect 2692 52252 2756 52256
rect 2692 52196 2696 52252
rect 2696 52196 2752 52252
rect 2752 52196 2756 52252
rect 2692 52192 2756 52196
rect 2772 52252 2836 52256
rect 2772 52196 2776 52252
rect 2776 52196 2832 52252
rect 2832 52196 2836 52252
rect 2772 52192 2836 52196
rect 2852 52252 2916 52256
rect 2852 52196 2856 52252
rect 2856 52196 2912 52252
rect 2912 52196 2916 52252
rect 2852 52192 2916 52196
rect 7612 52252 7676 52256
rect 7612 52196 7616 52252
rect 7616 52196 7672 52252
rect 7672 52196 7676 52252
rect 7612 52192 7676 52196
rect 7692 52252 7756 52256
rect 7692 52196 7696 52252
rect 7696 52196 7752 52252
rect 7752 52196 7756 52252
rect 7692 52192 7756 52196
rect 7772 52252 7836 52256
rect 7772 52196 7776 52252
rect 7776 52196 7832 52252
rect 7832 52196 7836 52252
rect 7772 52192 7836 52196
rect 7852 52252 7916 52256
rect 7852 52196 7856 52252
rect 7856 52196 7912 52252
rect 7912 52196 7916 52252
rect 7852 52192 7916 52196
rect 12612 52252 12676 52256
rect 12612 52196 12616 52252
rect 12616 52196 12672 52252
rect 12672 52196 12676 52252
rect 12612 52192 12676 52196
rect 12692 52252 12756 52256
rect 12692 52196 12696 52252
rect 12696 52196 12752 52252
rect 12752 52196 12756 52252
rect 12692 52192 12756 52196
rect 12772 52252 12836 52256
rect 12772 52196 12776 52252
rect 12776 52196 12832 52252
rect 12832 52196 12836 52252
rect 12772 52192 12836 52196
rect 12852 52252 12916 52256
rect 12852 52196 12856 52252
rect 12856 52196 12912 52252
rect 12912 52196 12916 52252
rect 12852 52192 12916 52196
rect 17612 52252 17676 52256
rect 17612 52196 17616 52252
rect 17616 52196 17672 52252
rect 17672 52196 17676 52252
rect 17612 52192 17676 52196
rect 17692 52252 17756 52256
rect 17692 52196 17696 52252
rect 17696 52196 17752 52252
rect 17752 52196 17756 52252
rect 17692 52192 17756 52196
rect 17772 52252 17836 52256
rect 17772 52196 17776 52252
rect 17776 52196 17832 52252
rect 17832 52196 17836 52252
rect 17772 52192 17836 52196
rect 17852 52252 17916 52256
rect 17852 52196 17856 52252
rect 17856 52196 17912 52252
rect 17912 52196 17916 52252
rect 17852 52192 17916 52196
rect 8156 51852 8220 51916
rect 1952 51708 2016 51712
rect 1952 51652 1956 51708
rect 1956 51652 2012 51708
rect 2012 51652 2016 51708
rect 1952 51648 2016 51652
rect 2032 51708 2096 51712
rect 2032 51652 2036 51708
rect 2036 51652 2092 51708
rect 2092 51652 2096 51708
rect 2032 51648 2096 51652
rect 2112 51708 2176 51712
rect 2112 51652 2116 51708
rect 2116 51652 2172 51708
rect 2172 51652 2176 51708
rect 2112 51648 2176 51652
rect 2192 51708 2256 51712
rect 2192 51652 2196 51708
rect 2196 51652 2252 51708
rect 2252 51652 2256 51708
rect 2192 51648 2256 51652
rect 6952 51708 7016 51712
rect 6952 51652 6956 51708
rect 6956 51652 7012 51708
rect 7012 51652 7016 51708
rect 6952 51648 7016 51652
rect 7032 51708 7096 51712
rect 7032 51652 7036 51708
rect 7036 51652 7092 51708
rect 7092 51652 7096 51708
rect 7032 51648 7096 51652
rect 7112 51708 7176 51712
rect 7112 51652 7116 51708
rect 7116 51652 7172 51708
rect 7172 51652 7176 51708
rect 7112 51648 7176 51652
rect 7192 51708 7256 51712
rect 7192 51652 7196 51708
rect 7196 51652 7252 51708
rect 7252 51652 7256 51708
rect 7192 51648 7256 51652
rect 11952 51708 12016 51712
rect 11952 51652 11956 51708
rect 11956 51652 12012 51708
rect 12012 51652 12016 51708
rect 11952 51648 12016 51652
rect 12032 51708 12096 51712
rect 12032 51652 12036 51708
rect 12036 51652 12092 51708
rect 12092 51652 12096 51708
rect 12032 51648 12096 51652
rect 12112 51708 12176 51712
rect 12112 51652 12116 51708
rect 12116 51652 12172 51708
rect 12172 51652 12176 51708
rect 12112 51648 12176 51652
rect 12192 51708 12256 51712
rect 12192 51652 12196 51708
rect 12196 51652 12252 51708
rect 12252 51652 12256 51708
rect 12192 51648 12256 51652
rect 16952 51708 17016 51712
rect 16952 51652 16956 51708
rect 16956 51652 17012 51708
rect 17012 51652 17016 51708
rect 16952 51648 17016 51652
rect 17032 51708 17096 51712
rect 17032 51652 17036 51708
rect 17036 51652 17092 51708
rect 17092 51652 17096 51708
rect 17032 51648 17096 51652
rect 17112 51708 17176 51712
rect 17112 51652 17116 51708
rect 17116 51652 17172 51708
rect 17172 51652 17176 51708
rect 17112 51648 17176 51652
rect 17192 51708 17256 51712
rect 17192 51652 17196 51708
rect 17196 51652 17252 51708
rect 17252 51652 17256 51708
rect 17192 51648 17256 51652
rect 13124 51308 13188 51372
rect 2612 51164 2676 51168
rect 2612 51108 2616 51164
rect 2616 51108 2672 51164
rect 2672 51108 2676 51164
rect 2612 51104 2676 51108
rect 2692 51164 2756 51168
rect 2692 51108 2696 51164
rect 2696 51108 2752 51164
rect 2752 51108 2756 51164
rect 2692 51104 2756 51108
rect 2772 51164 2836 51168
rect 2772 51108 2776 51164
rect 2776 51108 2832 51164
rect 2832 51108 2836 51164
rect 2772 51104 2836 51108
rect 2852 51164 2916 51168
rect 2852 51108 2856 51164
rect 2856 51108 2912 51164
rect 2912 51108 2916 51164
rect 2852 51104 2916 51108
rect 7612 51164 7676 51168
rect 7612 51108 7616 51164
rect 7616 51108 7672 51164
rect 7672 51108 7676 51164
rect 7612 51104 7676 51108
rect 7692 51164 7756 51168
rect 7692 51108 7696 51164
rect 7696 51108 7752 51164
rect 7752 51108 7756 51164
rect 7692 51104 7756 51108
rect 7772 51164 7836 51168
rect 7772 51108 7776 51164
rect 7776 51108 7832 51164
rect 7832 51108 7836 51164
rect 7772 51104 7836 51108
rect 7852 51164 7916 51168
rect 7852 51108 7856 51164
rect 7856 51108 7912 51164
rect 7912 51108 7916 51164
rect 7852 51104 7916 51108
rect 12612 51164 12676 51168
rect 12612 51108 12616 51164
rect 12616 51108 12672 51164
rect 12672 51108 12676 51164
rect 12612 51104 12676 51108
rect 12692 51164 12756 51168
rect 12692 51108 12696 51164
rect 12696 51108 12752 51164
rect 12752 51108 12756 51164
rect 12692 51104 12756 51108
rect 12772 51164 12836 51168
rect 12772 51108 12776 51164
rect 12776 51108 12832 51164
rect 12832 51108 12836 51164
rect 12772 51104 12836 51108
rect 12852 51164 12916 51168
rect 12852 51108 12856 51164
rect 12856 51108 12912 51164
rect 12912 51108 12916 51164
rect 12852 51104 12916 51108
rect 17612 51164 17676 51168
rect 17612 51108 17616 51164
rect 17616 51108 17672 51164
rect 17672 51108 17676 51164
rect 17612 51104 17676 51108
rect 17692 51164 17756 51168
rect 17692 51108 17696 51164
rect 17696 51108 17752 51164
rect 17752 51108 17756 51164
rect 17692 51104 17756 51108
rect 17772 51164 17836 51168
rect 17772 51108 17776 51164
rect 17776 51108 17832 51164
rect 17832 51108 17836 51164
rect 17772 51104 17836 51108
rect 17852 51164 17916 51168
rect 17852 51108 17856 51164
rect 17856 51108 17912 51164
rect 17912 51108 17916 51164
rect 17852 51104 17916 51108
rect 7420 50764 7484 50828
rect 10732 50688 10796 50692
rect 10732 50632 10746 50688
rect 10746 50632 10796 50688
rect 10732 50628 10796 50632
rect 1952 50620 2016 50624
rect 1952 50564 1956 50620
rect 1956 50564 2012 50620
rect 2012 50564 2016 50620
rect 1952 50560 2016 50564
rect 2032 50620 2096 50624
rect 2032 50564 2036 50620
rect 2036 50564 2092 50620
rect 2092 50564 2096 50620
rect 2032 50560 2096 50564
rect 2112 50620 2176 50624
rect 2112 50564 2116 50620
rect 2116 50564 2172 50620
rect 2172 50564 2176 50620
rect 2112 50560 2176 50564
rect 2192 50620 2256 50624
rect 2192 50564 2196 50620
rect 2196 50564 2252 50620
rect 2252 50564 2256 50620
rect 2192 50560 2256 50564
rect 6952 50620 7016 50624
rect 6952 50564 6956 50620
rect 6956 50564 7012 50620
rect 7012 50564 7016 50620
rect 6952 50560 7016 50564
rect 7032 50620 7096 50624
rect 7032 50564 7036 50620
rect 7036 50564 7092 50620
rect 7092 50564 7096 50620
rect 7032 50560 7096 50564
rect 7112 50620 7176 50624
rect 7112 50564 7116 50620
rect 7116 50564 7172 50620
rect 7172 50564 7176 50620
rect 7112 50560 7176 50564
rect 7192 50620 7256 50624
rect 7192 50564 7196 50620
rect 7196 50564 7252 50620
rect 7252 50564 7256 50620
rect 7192 50560 7256 50564
rect 11952 50620 12016 50624
rect 11952 50564 11956 50620
rect 11956 50564 12012 50620
rect 12012 50564 12016 50620
rect 11952 50560 12016 50564
rect 12032 50620 12096 50624
rect 12032 50564 12036 50620
rect 12036 50564 12092 50620
rect 12092 50564 12096 50620
rect 12032 50560 12096 50564
rect 12112 50620 12176 50624
rect 12112 50564 12116 50620
rect 12116 50564 12172 50620
rect 12172 50564 12176 50620
rect 12112 50560 12176 50564
rect 12192 50620 12256 50624
rect 12192 50564 12196 50620
rect 12196 50564 12252 50620
rect 12252 50564 12256 50620
rect 12192 50560 12256 50564
rect 16952 50620 17016 50624
rect 16952 50564 16956 50620
rect 16956 50564 17012 50620
rect 17012 50564 17016 50620
rect 16952 50560 17016 50564
rect 17032 50620 17096 50624
rect 17032 50564 17036 50620
rect 17036 50564 17092 50620
rect 17092 50564 17096 50620
rect 17032 50560 17096 50564
rect 17112 50620 17176 50624
rect 17112 50564 17116 50620
rect 17116 50564 17172 50620
rect 17172 50564 17176 50620
rect 17112 50560 17176 50564
rect 17192 50620 17256 50624
rect 17192 50564 17196 50620
rect 17196 50564 17252 50620
rect 17252 50564 17256 50620
rect 17192 50560 17256 50564
rect 2612 50076 2676 50080
rect 2612 50020 2616 50076
rect 2616 50020 2672 50076
rect 2672 50020 2676 50076
rect 2612 50016 2676 50020
rect 2692 50076 2756 50080
rect 2692 50020 2696 50076
rect 2696 50020 2752 50076
rect 2752 50020 2756 50076
rect 2692 50016 2756 50020
rect 2772 50076 2836 50080
rect 2772 50020 2776 50076
rect 2776 50020 2832 50076
rect 2832 50020 2836 50076
rect 2772 50016 2836 50020
rect 2852 50076 2916 50080
rect 2852 50020 2856 50076
rect 2856 50020 2912 50076
rect 2912 50020 2916 50076
rect 2852 50016 2916 50020
rect 7612 50076 7676 50080
rect 7612 50020 7616 50076
rect 7616 50020 7672 50076
rect 7672 50020 7676 50076
rect 7612 50016 7676 50020
rect 7692 50076 7756 50080
rect 7692 50020 7696 50076
rect 7696 50020 7752 50076
rect 7752 50020 7756 50076
rect 7692 50016 7756 50020
rect 7772 50076 7836 50080
rect 7772 50020 7776 50076
rect 7776 50020 7832 50076
rect 7832 50020 7836 50076
rect 7772 50016 7836 50020
rect 7852 50076 7916 50080
rect 7852 50020 7856 50076
rect 7856 50020 7912 50076
rect 7912 50020 7916 50076
rect 7852 50016 7916 50020
rect 12612 50076 12676 50080
rect 12612 50020 12616 50076
rect 12616 50020 12672 50076
rect 12672 50020 12676 50076
rect 12612 50016 12676 50020
rect 12692 50076 12756 50080
rect 12692 50020 12696 50076
rect 12696 50020 12752 50076
rect 12752 50020 12756 50076
rect 12692 50016 12756 50020
rect 12772 50076 12836 50080
rect 12772 50020 12776 50076
rect 12776 50020 12832 50076
rect 12832 50020 12836 50076
rect 12772 50016 12836 50020
rect 12852 50076 12916 50080
rect 12852 50020 12856 50076
rect 12856 50020 12912 50076
rect 12912 50020 12916 50076
rect 12852 50016 12916 50020
rect 17612 50076 17676 50080
rect 17612 50020 17616 50076
rect 17616 50020 17672 50076
rect 17672 50020 17676 50076
rect 17612 50016 17676 50020
rect 17692 50076 17756 50080
rect 17692 50020 17696 50076
rect 17696 50020 17752 50076
rect 17752 50020 17756 50076
rect 17692 50016 17756 50020
rect 17772 50076 17836 50080
rect 17772 50020 17776 50076
rect 17776 50020 17832 50076
rect 17832 50020 17836 50076
rect 17772 50016 17836 50020
rect 17852 50076 17916 50080
rect 17852 50020 17856 50076
rect 17856 50020 17912 50076
rect 17912 50020 17916 50076
rect 17852 50016 17916 50020
rect 4476 49736 4540 49740
rect 4476 49680 4490 49736
rect 4490 49680 4540 49736
rect 4476 49676 4540 49680
rect 15884 49540 15948 49604
rect 1952 49532 2016 49536
rect 1952 49476 1956 49532
rect 1956 49476 2012 49532
rect 2012 49476 2016 49532
rect 1952 49472 2016 49476
rect 2032 49532 2096 49536
rect 2032 49476 2036 49532
rect 2036 49476 2092 49532
rect 2092 49476 2096 49532
rect 2032 49472 2096 49476
rect 2112 49532 2176 49536
rect 2112 49476 2116 49532
rect 2116 49476 2172 49532
rect 2172 49476 2176 49532
rect 2112 49472 2176 49476
rect 2192 49532 2256 49536
rect 2192 49476 2196 49532
rect 2196 49476 2252 49532
rect 2252 49476 2256 49532
rect 2192 49472 2256 49476
rect 6952 49532 7016 49536
rect 6952 49476 6956 49532
rect 6956 49476 7012 49532
rect 7012 49476 7016 49532
rect 6952 49472 7016 49476
rect 7032 49532 7096 49536
rect 7032 49476 7036 49532
rect 7036 49476 7092 49532
rect 7092 49476 7096 49532
rect 7032 49472 7096 49476
rect 7112 49532 7176 49536
rect 7112 49476 7116 49532
rect 7116 49476 7172 49532
rect 7172 49476 7176 49532
rect 7112 49472 7176 49476
rect 7192 49532 7256 49536
rect 7192 49476 7196 49532
rect 7196 49476 7252 49532
rect 7252 49476 7256 49532
rect 7192 49472 7256 49476
rect 11952 49532 12016 49536
rect 11952 49476 11956 49532
rect 11956 49476 12012 49532
rect 12012 49476 12016 49532
rect 11952 49472 12016 49476
rect 12032 49532 12096 49536
rect 12032 49476 12036 49532
rect 12036 49476 12092 49532
rect 12092 49476 12096 49532
rect 12032 49472 12096 49476
rect 12112 49532 12176 49536
rect 12112 49476 12116 49532
rect 12116 49476 12172 49532
rect 12172 49476 12176 49532
rect 12112 49472 12176 49476
rect 12192 49532 12256 49536
rect 12192 49476 12196 49532
rect 12196 49476 12252 49532
rect 12252 49476 12256 49532
rect 12192 49472 12256 49476
rect 16952 49532 17016 49536
rect 16952 49476 16956 49532
rect 16956 49476 17012 49532
rect 17012 49476 17016 49532
rect 16952 49472 17016 49476
rect 17032 49532 17096 49536
rect 17032 49476 17036 49532
rect 17036 49476 17092 49532
rect 17092 49476 17096 49532
rect 17032 49472 17096 49476
rect 17112 49532 17176 49536
rect 17112 49476 17116 49532
rect 17116 49476 17172 49532
rect 17172 49476 17176 49532
rect 17112 49472 17176 49476
rect 17192 49532 17256 49536
rect 17192 49476 17196 49532
rect 17196 49476 17252 49532
rect 17252 49476 17256 49532
rect 17192 49472 17256 49476
rect 2612 48988 2676 48992
rect 2612 48932 2616 48988
rect 2616 48932 2672 48988
rect 2672 48932 2676 48988
rect 2612 48928 2676 48932
rect 2692 48988 2756 48992
rect 2692 48932 2696 48988
rect 2696 48932 2752 48988
rect 2752 48932 2756 48988
rect 2692 48928 2756 48932
rect 2772 48988 2836 48992
rect 2772 48932 2776 48988
rect 2776 48932 2832 48988
rect 2832 48932 2836 48988
rect 2772 48928 2836 48932
rect 2852 48988 2916 48992
rect 2852 48932 2856 48988
rect 2856 48932 2912 48988
rect 2912 48932 2916 48988
rect 2852 48928 2916 48932
rect 7612 48988 7676 48992
rect 7612 48932 7616 48988
rect 7616 48932 7672 48988
rect 7672 48932 7676 48988
rect 7612 48928 7676 48932
rect 7692 48988 7756 48992
rect 7692 48932 7696 48988
rect 7696 48932 7752 48988
rect 7752 48932 7756 48988
rect 7692 48928 7756 48932
rect 7772 48988 7836 48992
rect 7772 48932 7776 48988
rect 7776 48932 7832 48988
rect 7832 48932 7836 48988
rect 7772 48928 7836 48932
rect 7852 48988 7916 48992
rect 7852 48932 7856 48988
rect 7856 48932 7912 48988
rect 7912 48932 7916 48988
rect 7852 48928 7916 48932
rect 12612 48988 12676 48992
rect 12612 48932 12616 48988
rect 12616 48932 12672 48988
rect 12672 48932 12676 48988
rect 12612 48928 12676 48932
rect 12692 48988 12756 48992
rect 12692 48932 12696 48988
rect 12696 48932 12752 48988
rect 12752 48932 12756 48988
rect 12692 48928 12756 48932
rect 12772 48988 12836 48992
rect 12772 48932 12776 48988
rect 12776 48932 12832 48988
rect 12832 48932 12836 48988
rect 12772 48928 12836 48932
rect 12852 48988 12916 48992
rect 12852 48932 12856 48988
rect 12856 48932 12912 48988
rect 12912 48932 12916 48988
rect 12852 48928 12916 48932
rect 17612 48988 17676 48992
rect 17612 48932 17616 48988
rect 17616 48932 17672 48988
rect 17672 48932 17676 48988
rect 17612 48928 17676 48932
rect 17692 48988 17756 48992
rect 17692 48932 17696 48988
rect 17696 48932 17752 48988
rect 17752 48932 17756 48988
rect 17692 48928 17756 48932
rect 17772 48988 17836 48992
rect 17772 48932 17776 48988
rect 17776 48932 17832 48988
rect 17832 48932 17836 48988
rect 17772 48928 17836 48932
rect 17852 48988 17916 48992
rect 17852 48932 17856 48988
rect 17856 48932 17912 48988
rect 17912 48932 17916 48988
rect 17852 48928 17916 48932
rect 1952 48444 2016 48448
rect 1952 48388 1956 48444
rect 1956 48388 2012 48444
rect 2012 48388 2016 48444
rect 1952 48384 2016 48388
rect 2032 48444 2096 48448
rect 2032 48388 2036 48444
rect 2036 48388 2092 48444
rect 2092 48388 2096 48444
rect 2032 48384 2096 48388
rect 2112 48444 2176 48448
rect 2112 48388 2116 48444
rect 2116 48388 2172 48444
rect 2172 48388 2176 48444
rect 2112 48384 2176 48388
rect 2192 48444 2256 48448
rect 2192 48388 2196 48444
rect 2196 48388 2252 48444
rect 2252 48388 2256 48444
rect 2192 48384 2256 48388
rect 6952 48444 7016 48448
rect 6952 48388 6956 48444
rect 6956 48388 7012 48444
rect 7012 48388 7016 48444
rect 6952 48384 7016 48388
rect 7032 48444 7096 48448
rect 7032 48388 7036 48444
rect 7036 48388 7092 48444
rect 7092 48388 7096 48444
rect 7032 48384 7096 48388
rect 7112 48444 7176 48448
rect 7112 48388 7116 48444
rect 7116 48388 7172 48444
rect 7172 48388 7176 48444
rect 7112 48384 7176 48388
rect 7192 48444 7256 48448
rect 7192 48388 7196 48444
rect 7196 48388 7252 48444
rect 7252 48388 7256 48444
rect 7192 48384 7256 48388
rect 11952 48444 12016 48448
rect 11952 48388 11956 48444
rect 11956 48388 12012 48444
rect 12012 48388 12016 48444
rect 11952 48384 12016 48388
rect 12032 48444 12096 48448
rect 12032 48388 12036 48444
rect 12036 48388 12092 48444
rect 12092 48388 12096 48444
rect 12032 48384 12096 48388
rect 12112 48444 12176 48448
rect 12112 48388 12116 48444
rect 12116 48388 12172 48444
rect 12172 48388 12176 48444
rect 12112 48384 12176 48388
rect 12192 48444 12256 48448
rect 12192 48388 12196 48444
rect 12196 48388 12252 48444
rect 12252 48388 12256 48444
rect 12192 48384 12256 48388
rect 16068 48376 16132 48380
rect 16068 48320 16082 48376
rect 16082 48320 16132 48376
rect 16068 48316 16132 48320
rect 16952 48444 17016 48448
rect 16952 48388 16956 48444
rect 16956 48388 17012 48444
rect 17012 48388 17016 48444
rect 16952 48384 17016 48388
rect 17032 48444 17096 48448
rect 17032 48388 17036 48444
rect 17036 48388 17092 48444
rect 17092 48388 17096 48444
rect 17032 48384 17096 48388
rect 17112 48444 17176 48448
rect 17112 48388 17116 48444
rect 17116 48388 17172 48444
rect 17172 48388 17176 48444
rect 17112 48384 17176 48388
rect 17192 48444 17256 48448
rect 17192 48388 17196 48444
rect 17196 48388 17252 48444
rect 17252 48388 17256 48444
rect 17192 48384 17256 48388
rect 4660 48180 4724 48244
rect 2612 47900 2676 47904
rect 2612 47844 2616 47900
rect 2616 47844 2672 47900
rect 2672 47844 2676 47900
rect 2612 47840 2676 47844
rect 2692 47900 2756 47904
rect 2692 47844 2696 47900
rect 2696 47844 2752 47900
rect 2752 47844 2756 47900
rect 2692 47840 2756 47844
rect 2772 47900 2836 47904
rect 2772 47844 2776 47900
rect 2776 47844 2832 47900
rect 2832 47844 2836 47900
rect 2772 47840 2836 47844
rect 2852 47900 2916 47904
rect 2852 47844 2856 47900
rect 2856 47844 2912 47900
rect 2912 47844 2916 47900
rect 2852 47840 2916 47844
rect 7612 47900 7676 47904
rect 7612 47844 7616 47900
rect 7616 47844 7672 47900
rect 7672 47844 7676 47900
rect 7612 47840 7676 47844
rect 7692 47900 7756 47904
rect 7692 47844 7696 47900
rect 7696 47844 7752 47900
rect 7752 47844 7756 47900
rect 7692 47840 7756 47844
rect 7772 47900 7836 47904
rect 7772 47844 7776 47900
rect 7776 47844 7832 47900
rect 7832 47844 7836 47900
rect 7772 47840 7836 47844
rect 7852 47900 7916 47904
rect 7852 47844 7856 47900
rect 7856 47844 7912 47900
rect 7912 47844 7916 47900
rect 7852 47840 7916 47844
rect 12612 47900 12676 47904
rect 12612 47844 12616 47900
rect 12616 47844 12672 47900
rect 12672 47844 12676 47900
rect 12612 47840 12676 47844
rect 12692 47900 12756 47904
rect 12692 47844 12696 47900
rect 12696 47844 12752 47900
rect 12752 47844 12756 47900
rect 12692 47840 12756 47844
rect 12772 47900 12836 47904
rect 12772 47844 12776 47900
rect 12776 47844 12832 47900
rect 12832 47844 12836 47900
rect 12772 47840 12836 47844
rect 12852 47900 12916 47904
rect 12852 47844 12856 47900
rect 12856 47844 12912 47900
rect 12912 47844 12916 47900
rect 12852 47840 12916 47844
rect 17612 47900 17676 47904
rect 17612 47844 17616 47900
rect 17616 47844 17672 47900
rect 17672 47844 17676 47900
rect 17612 47840 17676 47844
rect 17692 47900 17756 47904
rect 17692 47844 17696 47900
rect 17696 47844 17752 47900
rect 17752 47844 17756 47900
rect 17692 47840 17756 47844
rect 17772 47900 17836 47904
rect 17772 47844 17776 47900
rect 17776 47844 17832 47900
rect 17832 47844 17836 47900
rect 17772 47840 17836 47844
rect 17852 47900 17916 47904
rect 17852 47844 17856 47900
rect 17856 47844 17912 47900
rect 17912 47844 17916 47900
rect 17852 47840 17916 47844
rect 1952 47356 2016 47360
rect 1952 47300 1956 47356
rect 1956 47300 2012 47356
rect 2012 47300 2016 47356
rect 1952 47296 2016 47300
rect 2032 47356 2096 47360
rect 2032 47300 2036 47356
rect 2036 47300 2092 47356
rect 2092 47300 2096 47356
rect 2032 47296 2096 47300
rect 2112 47356 2176 47360
rect 2112 47300 2116 47356
rect 2116 47300 2172 47356
rect 2172 47300 2176 47356
rect 2112 47296 2176 47300
rect 2192 47356 2256 47360
rect 2192 47300 2196 47356
rect 2196 47300 2252 47356
rect 2252 47300 2256 47356
rect 2192 47296 2256 47300
rect 6952 47356 7016 47360
rect 6952 47300 6956 47356
rect 6956 47300 7012 47356
rect 7012 47300 7016 47356
rect 6952 47296 7016 47300
rect 7032 47356 7096 47360
rect 7032 47300 7036 47356
rect 7036 47300 7092 47356
rect 7092 47300 7096 47356
rect 7032 47296 7096 47300
rect 7112 47356 7176 47360
rect 7112 47300 7116 47356
rect 7116 47300 7172 47356
rect 7172 47300 7176 47356
rect 7112 47296 7176 47300
rect 7192 47356 7256 47360
rect 7192 47300 7196 47356
rect 7196 47300 7252 47356
rect 7252 47300 7256 47356
rect 7192 47296 7256 47300
rect 11952 47356 12016 47360
rect 11952 47300 11956 47356
rect 11956 47300 12012 47356
rect 12012 47300 12016 47356
rect 11952 47296 12016 47300
rect 12032 47356 12096 47360
rect 12032 47300 12036 47356
rect 12036 47300 12092 47356
rect 12092 47300 12096 47356
rect 12032 47296 12096 47300
rect 12112 47356 12176 47360
rect 12112 47300 12116 47356
rect 12116 47300 12172 47356
rect 12172 47300 12176 47356
rect 12112 47296 12176 47300
rect 12192 47356 12256 47360
rect 12192 47300 12196 47356
rect 12196 47300 12252 47356
rect 12252 47300 12256 47356
rect 12192 47296 12256 47300
rect 16952 47356 17016 47360
rect 16952 47300 16956 47356
rect 16956 47300 17012 47356
rect 17012 47300 17016 47356
rect 16952 47296 17016 47300
rect 17032 47356 17096 47360
rect 17032 47300 17036 47356
rect 17036 47300 17092 47356
rect 17092 47300 17096 47356
rect 17032 47296 17096 47300
rect 17112 47356 17176 47360
rect 17112 47300 17116 47356
rect 17116 47300 17172 47356
rect 17172 47300 17176 47356
rect 17112 47296 17176 47300
rect 17192 47356 17256 47360
rect 17192 47300 17196 47356
rect 17196 47300 17252 47356
rect 17252 47300 17256 47356
rect 17192 47296 17256 47300
rect 3188 47228 3252 47292
rect 2612 46812 2676 46816
rect 2612 46756 2616 46812
rect 2616 46756 2672 46812
rect 2672 46756 2676 46812
rect 2612 46752 2676 46756
rect 2692 46812 2756 46816
rect 2692 46756 2696 46812
rect 2696 46756 2752 46812
rect 2752 46756 2756 46812
rect 2692 46752 2756 46756
rect 2772 46812 2836 46816
rect 2772 46756 2776 46812
rect 2776 46756 2832 46812
rect 2832 46756 2836 46812
rect 2772 46752 2836 46756
rect 2852 46812 2916 46816
rect 2852 46756 2856 46812
rect 2856 46756 2912 46812
rect 2912 46756 2916 46812
rect 2852 46752 2916 46756
rect 7612 46812 7676 46816
rect 7612 46756 7616 46812
rect 7616 46756 7672 46812
rect 7672 46756 7676 46812
rect 7612 46752 7676 46756
rect 7692 46812 7756 46816
rect 7692 46756 7696 46812
rect 7696 46756 7752 46812
rect 7752 46756 7756 46812
rect 7692 46752 7756 46756
rect 7772 46812 7836 46816
rect 7772 46756 7776 46812
rect 7776 46756 7832 46812
rect 7832 46756 7836 46812
rect 7772 46752 7836 46756
rect 7852 46812 7916 46816
rect 7852 46756 7856 46812
rect 7856 46756 7912 46812
rect 7912 46756 7916 46812
rect 7852 46752 7916 46756
rect 12612 46812 12676 46816
rect 12612 46756 12616 46812
rect 12616 46756 12672 46812
rect 12672 46756 12676 46812
rect 12612 46752 12676 46756
rect 12692 46812 12756 46816
rect 12692 46756 12696 46812
rect 12696 46756 12752 46812
rect 12752 46756 12756 46812
rect 12692 46752 12756 46756
rect 12772 46812 12836 46816
rect 12772 46756 12776 46812
rect 12776 46756 12832 46812
rect 12832 46756 12836 46812
rect 12772 46752 12836 46756
rect 12852 46812 12916 46816
rect 12852 46756 12856 46812
rect 12856 46756 12912 46812
rect 12912 46756 12916 46812
rect 12852 46752 12916 46756
rect 17612 46812 17676 46816
rect 17612 46756 17616 46812
rect 17616 46756 17672 46812
rect 17672 46756 17676 46812
rect 17612 46752 17676 46756
rect 17692 46812 17756 46816
rect 17692 46756 17696 46812
rect 17696 46756 17752 46812
rect 17752 46756 17756 46812
rect 17692 46752 17756 46756
rect 17772 46812 17836 46816
rect 17772 46756 17776 46812
rect 17776 46756 17832 46812
rect 17832 46756 17836 46812
rect 17772 46752 17836 46756
rect 17852 46812 17916 46816
rect 17852 46756 17856 46812
rect 17856 46756 17912 46812
rect 17912 46756 17916 46812
rect 17852 46752 17916 46756
rect 1952 46268 2016 46272
rect 1952 46212 1956 46268
rect 1956 46212 2012 46268
rect 2012 46212 2016 46268
rect 1952 46208 2016 46212
rect 2032 46268 2096 46272
rect 2032 46212 2036 46268
rect 2036 46212 2092 46268
rect 2092 46212 2096 46268
rect 2032 46208 2096 46212
rect 2112 46268 2176 46272
rect 2112 46212 2116 46268
rect 2116 46212 2172 46268
rect 2172 46212 2176 46268
rect 2112 46208 2176 46212
rect 2192 46268 2256 46272
rect 2192 46212 2196 46268
rect 2196 46212 2252 46268
rect 2252 46212 2256 46268
rect 2192 46208 2256 46212
rect 6952 46268 7016 46272
rect 6952 46212 6956 46268
rect 6956 46212 7012 46268
rect 7012 46212 7016 46268
rect 6952 46208 7016 46212
rect 7032 46268 7096 46272
rect 7032 46212 7036 46268
rect 7036 46212 7092 46268
rect 7092 46212 7096 46268
rect 7032 46208 7096 46212
rect 7112 46268 7176 46272
rect 7112 46212 7116 46268
rect 7116 46212 7172 46268
rect 7172 46212 7176 46268
rect 7112 46208 7176 46212
rect 7192 46268 7256 46272
rect 7192 46212 7196 46268
rect 7196 46212 7252 46268
rect 7252 46212 7256 46268
rect 7192 46208 7256 46212
rect 11952 46268 12016 46272
rect 11952 46212 11956 46268
rect 11956 46212 12012 46268
rect 12012 46212 12016 46268
rect 11952 46208 12016 46212
rect 12032 46268 12096 46272
rect 12032 46212 12036 46268
rect 12036 46212 12092 46268
rect 12092 46212 12096 46268
rect 12032 46208 12096 46212
rect 12112 46268 12176 46272
rect 12112 46212 12116 46268
rect 12116 46212 12172 46268
rect 12172 46212 12176 46268
rect 12112 46208 12176 46212
rect 12192 46268 12256 46272
rect 12192 46212 12196 46268
rect 12196 46212 12252 46268
rect 12252 46212 12256 46268
rect 12192 46208 12256 46212
rect 16952 46268 17016 46272
rect 16952 46212 16956 46268
rect 16956 46212 17012 46268
rect 17012 46212 17016 46268
rect 16952 46208 17016 46212
rect 17032 46268 17096 46272
rect 17032 46212 17036 46268
rect 17036 46212 17092 46268
rect 17092 46212 17096 46268
rect 17032 46208 17096 46212
rect 17112 46268 17176 46272
rect 17112 46212 17116 46268
rect 17116 46212 17172 46268
rect 17172 46212 17176 46268
rect 17112 46208 17176 46212
rect 17192 46268 17256 46272
rect 17192 46212 17196 46268
rect 17196 46212 17252 46268
rect 17252 46212 17256 46268
rect 17192 46208 17256 46212
rect 2612 45724 2676 45728
rect 2612 45668 2616 45724
rect 2616 45668 2672 45724
rect 2672 45668 2676 45724
rect 2612 45664 2676 45668
rect 2692 45724 2756 45728
rect 2692 45668 2696 45724
rect 2696 45668 2752 45724
rect 2752 45668 2756 45724
rect 2692 45664 2756 45668
rect 2772 45724 2836 45728
rect 2772 45668 2776 45724
rect 2776 45668 2832 45724
rect 2832 45668 2836 45724
rect 2772 45664 2836 45668
rect 2852 45724 2916 45728
rect 2852 45668 2856 45724
rect 2856 45668 2912 45724
rect 2912 45668 2916 45724
rect 2852 45664 2916 45668
rect 7612 45724 7676 45728
rect 7612 45668 7616 45724
rect 7616 45668 7672 45724
rect 7672 45668 7676 45724
rect 7612 45664 7676 45668
rect 7692 45724 7756 45728
rect 7692 45668 7696 45724
rect 7696 45668 7752 45724
rect 7752 45668 7756 45724
rect 7692 45664 7756 45668
rect 7772 45724 7836 45728
rect 7772 45668 7776 45724
rect 7776 45668 7832 45724
rect 7832 45668 7836 45724
rect 7772 45664 7836 45668
rect 7852 45724 7916 45728
rect 7852 45668 7856 45724
rect 7856 45668 7912 45724
rect 7912 45668 7916 45724
rect 7852 45664 7916 45668
rect 12612 45724 12676 45728
rect 12612 45668 12616 45724
rect 12616 45668 12672 45724
rect 12672 45668 12676 45724
rect 12612 45664 12676 45668
rect 12692 45724 12756 45728
rect 12692 45668 12696 45724
rect 12696 45668 12752 45724
rect 12752 45668 12756 45724
rect 12692 45664 12756 45668
rect 12772 45724 12836 45728
rect 12772 45668 12776 45724
rect 12776 45668 12832 45724
rect 12832 45668 12836 45724
rect 12772 45664 12836 45668
rect 12852 45724 12916 45728
rect 12852 45668 12856 45724
rect 12856 45668 12912 45724
rect 12912 45668 12916 45724
rect 12852 45664 12916 45668
rect 17612 45724 17676 45728
rect 17612 45668 17616 45724
rect 17616 45668 17672 45724
rect 17672 45668 17676 45724
rect 17612 45664 17676 45668
rect 17692 45724 17756 45728
rect 17692 45668 17696 45724
rect 17696 45668 17752 45724
rect 17752 45668 17756 45724
rect 17692 45664 17756 45668
rect 17772 45724 17836 45728
rect 17772 45668 17776 45724
rect 17776 45668 17832 45724
rect 17832 45668 17836 45724
rect 17772 45664 17836 45668
rect 17852 45724 17916 45728
rect 17852 45668 17856 45724
rect 17856 45668 17912 45724
rect 17912 45668 17916 45724
rect 17852 45664 17916 45668
rect 1952 45180 2016 45184
rect 1952 45124 1956 45180
rect 1956 45124 2012 45180
rect 2012 45124 2016 45180
rect 1952 45120 2016 45124
rect 2032 45180 2096 45184
rect 2032 45124 2036 45180
rect 2036 45124 2092 45180
rect 2092 45124 2096 45180
rect 2032 45120 2096 45124
rect 2112 45180 2176 45184
rect 2112 45124 2116 45180
rect 2116 45124 2172 45180
rect 2172 45124 2176 45180
rect 2112 45120 2176 45124
rect 2192 45180 2256 45184
rect 2192 45124 2196 45180
rect 2196 45124 2252 45180
rect 2252 45124 2256 45180
rect 2192 45120 2256 45124
rect 6952 45180 7016 45184
rect 6952 45124 6956 45180
rect 6956 45124 7012 45180
rect 7012 45124 7016 45180
rect 6952 45120 7016 45124
rect 7032 45180 7096 45184
rect 7032 45124 7036 45180
rect 7036 45124 7092 45180
rect 7092 45124 7096 45180
rect 7032 45120 7096 45124
rect 7112 45180 7176 45184
rect 7112 45124 7116 45180
rect 7116 45124 7172 45180
rect 7172 45124 7176 45180
rect 7112 45120 7176 45124
rect 7192 45180 7256 45184
rect 7192 45124 7196 45180
rect 7196 45124 7252 45180
rect 7252 45124 7256 45180
rect 7192 45120 7256 45124
rect 11952 45180 12016 45184
rect 11952 45124 11956 45180
rect 11956 45124 12012 45180
rect 12012 45124 12016 45180
rect 11952 45120 12016 45124
rect 12032 45180 12096 45184
rect 12032 45124 12036 45180
rect 12036 45124 12092 45180
rect 12092 45124 12096 45180
rect 12032 45120 12096 45124
rect 12112 45180 12176 45184
rect 12112 45124 12116 45180
rect 12116 45124 12172 45180
rect 12172 45124 12176 45180
rect 12112 45120 12176 45124
rect 12192 45180 12256 45184
rect 12192 45124 12196 45180
rect 12196 45124 12252 45180
rect 12252 45124 12256 45180
rect 12192 45120 12256 45124
rect 16952 45180 17016 45184
rect 16952 45124 16956 45180
rect 16956 45124 17012 45180
rect 17012 45124 17016 45180
rect 16952 45120 17016 45124
rect 17032 45180 17096 45184
rect 17032 45124 17036 45180
rect 17036 45124 17092 45180
rect 17092 45124 17096 45180
rect 17032 45120 17096 45124
rect 17112 45180 17176 45184
rect 17112 45124 17116 45180
rect 17116 45124 17172 45180
rect 17172 45124 17176 45180
rect 17112 45120 17176 45124
rect 17192 45180 17256 45184
rect 17192 45124 17196 45180
rect 17196 45124 17252 45180
rect 17252 45124 17256 45180
rect 17192 45120 17256 45124
rect 2612 44636 2676 44640
rect 2612 44580 2616 44636
rect 2616 44580 2672 44636
rect 2672 44580 2676 44636
rect 2612 44576 2676 44580
rect 2692 44636 2756 44640
rect 2692 44580 2696 44636
rect 2696 44580 2752 44636
rect 2752 44580 2756 44636
rect 2692 44576 2756 44580
rect 2772 44636 2836 44640
rect 2772 44580 2776 44636
rect 2776 44580 2832 44636
rect 2832 44580 2836 44636
rect 2772 44576 2836 44580
rect 2852 44636 2916 44640
rect 2852 44580 2856 44636
rect 2856 44580 2912 44636
rect 2912 44580 2916 44636
rect 2852 44576 2916 44580
rect 7612 44636 7676 44640
rect 7612 44580 7616 44636
rect 7616 44580 7672 44636
rect 7672 44580 7676 44636
rect 7612 44576 7676 44580
rect 7692 44636 7756 44640
rect 7692 44580 7696 44636
rect 7696 44580 7752 44636
rect 7752 44580 7756 44636
rect 7692 44576 7756 44580
rect 7772 44636 7836 44640
rect 7772 44580 7776 44636
rect 7776 44580 7832 44636
rect 7832 44580 7836 44636
rect 7772 44576 7836 44580
rect 7852 44636 7916 44640
rect 7852 44580 7856 44636
rect 7856 44580 7912 44636
rect 7912 44580 7916 44636
rect 7852 44576 7916 44580
rect 12612 44636 12676 44640
rect 12612 44580 12616 44636
rect 12616 44580 12672 44636
rect 12672 44580 12676 44636
rect 12612 44576 12676 44580
rect 12692 44636 12756 44640
rect 12692 44580 12696 44636
rect 12696 44580 12752 44636
rect 12752 44580 12756 44636
rect 12692 44576 12756 44580
rect 12772 44636 12836 44640
rect 12772 44580 12776 44636
rect 12776 44580 12832 44636
rect 12832 44580 12836 44636
rect 12772 44576 12836 44580
rect 12852 44636 12916 44640
rect 12852 44580 12856 44636
rect 12856 44580 12912 44636
rect 12912 44580 12916 44636
rect 12852 44576 12916 44580
rect 17612 44636 17676 44640
rect 17612 44580 17616 44636
rect 17616 44580 17672 44636
rect 17672 44580 17676 44636
rect 17612 44576 17676 44580
rect 17692 44636 17756 44640
rect 17692 44580 17696 44636
rect 17696 44580 17752 44636
rect 17752 44580 17756 44636
rect 17692 44576 17756 44580
rect 17772 44636 17836 44640
rect 17772 44580 17776 44636
rect 17776 44580 17832 44636
rect 17832 44580 17836 44636
rect 17772 44576 17836 44580
rect 17852 44636 17916 44640
rect 17852 44580 17856 44636
rect 17856 44580 17912 44636
rect 17912 44580 17916 44636
rect 17852 44576 17916 44580
rect 1952 44092 2016 44096
rect 1952 44036 1956 44092
rect 1956 44036 2012 44092
rect 2012 44036 2016 44092
rect 1952 44032 2016 44036
rect 2032 44092 2096 44096
rect 2032 44036 2036 44092
rect 2036 44036 2092 44092
rect 2092 44036 2096 44092
rect 2032 44032 2096 44036
rect 2112 44092 2176 44096
rect 2112 44036 2116 44092
rect 2116 44036 2172 44092
rect 2172 44036 2176 44092
rect 2112 44032 2176 44036
rect 2192 44092 2256 44096
rect 2192 44036 2196 44092
rect 2196 44036 2252 44092
rect 2252 44036 2256 44092
rect 2192 44032 2256 44036
rect 6952 44092 7016 44096
rect 6952 44036 6956 44092
rect 6956 44036 7012 44092
rect 7012 44036 7016 44092
rect 6952 44032 7016 44036
rect 7032 44092 7096 44096
rect 7032 44036 7036 44092
rect 7036 44036 7092 44092
rect 7092 44036 7096 44092
rect 7032 44032 7096 44036
rect 7112 44092 7176 44096
rect 7112 44036 7116 44092
rect 7116 44036 7172 44092
rect 7172 44036 7176 44092
rect 7112 44032 7176 44036
rect 7192 44092 7256 44096
rect 7192 44036 7196 44092
rect 7196 44036 7252 44092
rect 7252 44036 7256 44092
rect 7192 44032 7256 44036
rect 11952 44092 12016 44096
rect 11952 44036 11956 44092
rect 11956 44036 12012 44092
rect 12012 44036 12016 44092
rect 11952 44032 12016 44036
rect 12032 44092 12096 44096
rect 12032 44036 12036 44092
rect 12036 44036 12092 44092
rect 12092 44036 12096 44092
rect 12032 44032 12096 44036
rect 12112 44092 12176 44096
rect 12112 44036 12116 44092
rect 12116 44036 12172 44092
rect 12172 44036 12176 44092
rect 12112 44032 12176 44036
rect 12192 44092 12256 44096
rect 12192 44036 12196 44092
rect 12196 44036 12252 44092
rect 12252 44036 12256 44092
rect 12192 44032 12256 44036
rect 16952 44092 17016 44096
rect 16952 44036 16956 44092
rect 16956 44036 17012 44092
rect 17012 44036 17016 44092
rect 16952 44032 17016 44036
rect 17032 44092 17096 44096
rect 17032 44036 17036 44092
rect 17036 44036 17092 44092
rect 17092 44036 17096 44092
rect 17032 44032 17096 44036
rect 17112 44092 17176 44096
rect 17112 44036 17116 44092
rect 17116 44036 17172 44092
rect 17172 44036 17176 44092
rect 17112 44032 17176 44036
rect 17192 44092 17256 44096
rect 17192 44036 17196 44092
rect 17196 44036 17252 44092
rect 17252 44036 17256 44092
rect 17192 44032 17256 44036
rect 2612 43548 2676 43552
rect 2612 43492 2616 43548
rect 2616 43492 2672 43548
rect 2672 43492 2676 43548
rect 2612 43488 2676 43492
rect 2692 43548 2756 43552
rect 2692 43492 2696 43548
rect 2696 43492 2752 43548
rect 2752 43492 2756 43548
rect 2692 43488 2756 43492
rect 2772 43548 2836 43552
rect 2772 43492 2776 43548
rect 2776 43492 2832 43548
rect 2832 43492 2836 43548
rect 2772 43488 2836 43492
rect 2852 43548 2916 43552
rect 2852 43492 2856 43548
rect 2856 43492 2912 43548
rect 2912 43492 2916 43548
rect 2852 43488 2916 43492
rect 7612 43548 7676 43552
rect 7612 43492 7616 43548
rect 7616 43492 7672 43548
rect 7672 43492 7676 43548
rect 7612 43488 7676 43492
rect 7692 43548 7756 43552
rect 7692 43492 7696 43548
rect 7696 43492 7752 43548
rect 7752 43492 7756 43548
rect 7692 43488 7756 43492
rect 7772 43548 7836 43552
rect 7772 43492 7776 43548
rect 7776 43492 7832 43548
rect 7832 43492 7836 43548
rect 7772 43488 7836 43492
rect 7852 43548 7916 43552
rect 7852 43492 7856 43548
rect 7856 43492 7912 43548
rect 7912 43492 7916 43548
rect 7852 43488 7916 43492
rect 12612 43548 12676 43552
rect 12612 43492 12616 43548
rect 12616 43492 12672 43548
rect 12672 43492 12676 43548
rect 12612 43488 12676 43492
rect 12692 43548 12756 43552
rect 12692 43492 12696 43548
rect 12696 43492 12752 43548
rect 12752 43492 12756 43548
rect 12692 43488 12756 43492
rect 12772 43548 12836 43552
rect 12772 43492 12776 43548
rect 12776 43492 12832 43548
rect 12832 43492 12836 43548
rect 12772 43488 12836 43492
rect 12852 43548 12916 43552
rect 12852 43492 12856 43548
rect 12856 43492 12912 43548
rect 12912 43492 12916 43548
rect 12852 43488 12916 43492
rect 17612 43548 17676 43552
rect 17612 43492 17616 43548
rect 17616 43492 17672 43548
rect 17672 43492 17676 43548
rect 17612 43488 17676 43492
rect 17692 43548 17756 43552
rect 17692 43492 17696 43548
rect 17696 43492 17752 43548
rect 17752 43492 17756 43548
rect 17692 43488 17756 43492
rect 17772 43548 17836 43552
rect 17772 43492 17776 43548
rect 17776 43492 17832 43548
rect 17832 43492 17836 43548
rect 17772 43488 17836 43492
rect 17852 43548 17916 43552
rect 17852 43492 17856 43548
rect 17856 43492 17912 43548
rect 17912 43492 17916 43548
rect 17852 43488 17916 43492
rect 7420 43284 7484 43348
rect 1952 43004 2016 43008
rect 1952 42948 1956 43004
rect 1956 42948 2012 43004
rect 2012 42948 2016 43004
rect 1952 42944 2016 42948
rect 2032 43004 2096 43008
rect 2032 42948 2036 43004
rect 2036 42948 2092 43004
rect 2092 42948 2096 43004
rect 2032 42944 2096 42948
rect 2112 43004 2176 43008
rect 2112 42948 2116 43004
rect 2116 42948 2172 43004
rect 2172 42948 2176 43004
rect 2112 42944 2176 42948
rect 2192 43004 2256 43008
rect 2192 42948 2196 43004
rect 2196 42948 2252 43004
rect 2252 42948 2256 43004
rect 2192 42944 2256 42948
rect 6952 43004 7016 43008
rect 6952 42948 6956 43004
rect 6956 42948 7012 43004
rect 7012 42948 7016 43004
rect 6952 42944 7016 42948
rect 7032 43004 7096 43008
rect 7032 42948 7036 43004
rect 7036 42948 7092 43004
rect 7092 42948 7096 43004
rect 7032 42944 7096 42948
rect 7112 43004 7176 43008
rect 7112 42948 7116 43004
rect 7116 42948 7172 43004
rect 7172 42948 7176 43004
rect 7112 42944 7176 42948
rect 7192 43004 7256 43008
rect 7192 42948 7196 43004
rect 7196 42948 7252 43004
rect 7252 42948 7256 43004
rect 7192 42944 7256 42948
rect 11952 43004 12016 43008
rect 11952 42948 11956 43004
rect 11956 42948 12012 43004
rect 12012 42948 12016 43004
rect 11952 42944 12016 42948
rect 12032 43004 12096 43008
rect 12032 42948 12036 43004
rect 12036 42948 12092 43004
rect 12092 42948 12096 43004
rect 12032 42944 12096 42948
rect 12112 43004 12176 43008
rect 12112 42948 12116 43004
rect 12116 42948 12172 43004
rect 12172 42948 12176 43004
rect 12112 42944 12176 42948
rect 12192 43004 12256 43008
rect 12192 42948 12196 43004
rect 12196 42948 12252 43004
rect 12252 42948 12256 43004
rect 12192 42944 12256 42948
rect 16952 43004 17016 43008
rect 16952 42948 16956 43004
rect 16956 42948 17012 43004
rect 17012 42948 17016 43004
rect 16952 42944 17016 42948
rect 17032 43004 17096 43008
rect 17032 42948 17036 43004
rect 17036 42948 17092 43004
rect 17092 42948 17096 43004
rect 17032 42944 17096 42948
rect 17112 43004 17176 43008
rect 17112 42948 17116 43004
rect 17116 42948 17172 43004
rect 17172 42948 17176 43004
rect 17112 42944 17176 42948
rect 17192 43004 17256 43008
rect 17192 42948 17196 43004
rect 17196 42948 17252 43004
rect 17252 42948 17256 43004
rect 17192 42944 17256 42948
rect 6500 42876 6564 42940
rect 11284 42740 11348 42804
rect 11468 42740 11532 42804
rect 2612 42460 2676 42464
rect 2612 42404 2616 42460
rect 2616 42404 2672 42460
rect 2672 42404 2676 42460
rect 2612 42400 2676 42404
rect 2692 42460 2756 42464
rect 2692 42404 2696 42460
rect 2696 42404 2752 42460
rect 2752 42404 2756 42460
rect 2692 42400 2756 42404
rect 2772 42460 2836 42464
rect 2772 42404 2776 42460
rect 2776 42404 2832 42460
rect 2832 42404 2836 42460
rect 2772 42400 2836 42404
rect 2852 42460 2916 42464
rect 2852 42404 2856 42460
rect 2856 42404 2912 42460
rect 2912 42404 2916 42460
rect 2852 42400 2916 42404
rect 7612 42460 7676 42464
rect 7612 42404 7616 42460
rect 7616 42404 7672 42460
rect 7672 42404 7676 42460
rect 7612 42400 7676 42404
rect 7692 42460 7756 42464
rect 7692 42404 7696 42460
rect 7696 42404 7752 42460
rect 7752 42404 7756 42460
rect 7692 42400 7756 42404
rect 7772 42460 7836 42464
rect 7772 42404 7776 42460
rect 7776 42404 7832 42460
rect 7832 42404 7836 42460
rect 7772 42400 7836 42404
rect 7852 42460 7916 42464
rect 7852 42404 7856 42460
rect 7856 42404 7912 42460
rect 7912 42404 7916 42460
rect 7852 42400 7916 42404
rect 12612 42460 12676 42464
rect 12612 42404 12616 42460
rect 12616 42404 12672 42460
rect 12672 42404 12676 42460
rect 12612 42400 12676 42404
rect 12692 42460 12756 42464
rect 12692 42404 12696 42460
rect 12696 42404 12752 42460
rect 12752 42404 12756 42460
rect 12692 42400 12756 42404
rect 12772 42460 12836 42464
rect 12772 42404 12776 42460
rect 12776 42404 12832 42460
rect 12832 42404 12836 42460
rect 12772 42400 12836 42404
rect 12852 42460 12916 42464
rect 12852 42404 12856 42460
rect 12856 42404 12912 42460
rect 12912 42404 12916 42460
rect 12852 42400 12916 42404
rect 17612 42460 17676 42464
rect 17612 42404 17616 42460
rect 17616 42404 17672 42460
rect 17672 42404 17676 42460
rect 17612 42400 17676 42404
rect 17692 42460 17756 42464
rect 17692 42404 17696 42460
rect 17696 42404 17752 42460
rect 17752 42404 17756 42460
rect 17692 42400 17756 42404
rect 17772 42460 17836 42464
rect 17772 42404 17776 42460
rect 17776 42404 17832 42460
rect 17832 42404 17836 42460
rect 17772 42400 17836 42404
rect 17852 42460 17916 42464
rect 17852 42404 17856 42460
rect 17856 42404 17912 42460
rect 17912 42404 17916 42460
rect 17852 42400 17916 42404
rect 1952 41916 2016 41920
rect 1952 41860 1956 41916
rect 1956 41860 2012 41916
rect 2012 41860 2016 41916
rect 1952 41856 2016 41860
rect 2032 41916 2096 41920
rect 2032 41860 2036 41916
rect 2036 41860 2092 41916
rect 2092 41860 2096 41916
rect 2032 41856 2096 41860
rect 2112 41916 2176 41920
rect 2112 41860 2116 41916
rect 2116 41860 2172 41916
rect 2172 41860 2176 41916
rect 2112 41856 2176 41860
rect 2192 41916 2256 41920
rect 2192 41860 2196 41916
rect 2196 41860 2252 41916
rect 2252 41860 2256 41916
rect 2192 41856 2256 41860
rect 6952 41916 7016 41920
rect 6952 41860 6956 41916
rect 6956 41860 7012 41916
rect 7012 41860 7016 41916
rect 6952 41856 7016 41860
rect 7032 41916 7096 41920
rect 7032 41860 7036 41916
rect 7036 41860 7092 41916
rect 7092 41860 7096 41916
rect 7032 41856 7096 41860
rect 7112 41916 7176 41920
rect 7112 41860 7116 41916
rect 7116 41860 7172 41916
rect 7172 41860 7176 41916
rect 7112 41856 7176 41860
rect 7192 41916 7256 41920
rect 7192 41860 7196 41916
rect 7196 41860 7252 41916
rect 7252 41860 7256 41916
rect 7192 41856 7256 41860
rect 11952 41916 12016 41920
rect 11952 41860 11956 41916
rect 11956 41860 12012 41916
rect 12012 41860 12016 41916
rect 11952 41856 12016 41860
rect 12032 41916 12096 41920
rect 12032 41860 12036 41916
rect 12036 41860 12092 41916
rect 12092 41860 12096 41916
rect 12032 41856 12096 41860
rect 12112 41916 12176 41920
rect 12112 41860 12116 41916
rect 12116 41860 12172 41916
rect 12172 41860 12176 41916
rect 12112 41856 12176 41860
rect 12192 41916 12256 41920
rect 12192 41860 12196 41916
rect 12196 41860 12252 41916
rect 12252 41860 12256 41916
rect 12192 41856 12256 41860
rect 16952 41916 17016 41920
rect 16952 41860 16956 41916
rect 16956 41860 17012 41916
rect 17012 41860 17016 41916
rect 16952 41856 17016 41860
rect 17032 41916 17096 41920
rect 17032 41860 17036 41916
rect 17036 41860 17092 41916
rect 17092 41860 17096 41916
rect 17032 41856 17096 41860
rect 17112 41916 17176 41920
rect 17112 41860 17116 41916
rect 17116 41860 17172 41916
rect 17172 41860 17176 41916
rect 17112 41856 17176 41860
rect 17192 41916 17256 41920
rect 17192 41860 17196 41916
rect 17196 41860 17252 41916
rect 17252 41860 17256 41916
rect 17192 41856 17256 41860
rect 2612 41372 2676 41376
rect 2612 41316 2616 41372
rect 2616 41316 2672 41372
rect 2672 41316 2676 41372
rect 2612 41312 2676 41316
rect 2692 41372 2756 41376
rect 2692 41316 2696 41372
rect 2696 41316 2752 41372
rect 2752 41316 2756 41372
rect 2692 41312 2756 41316
rect 2772 41372 2836 41376
rect 2772 41316 2776 41372
rect 2776 41316 2832 41372
rect 2832 41316 2836 41372
rect 2772 41312 2836 41316
rect 2852 41372 2916 41376
rect 2852 41316 2856 41372
rect 2856 41316 2912 41372
rect 2912 41316 2916 41372
rect 2852 41312 2916 41316
rect 7612 41372 7676 41376
rect 7612 41316 7616 41372
rect 7616 41316 7672 41372
rect 7672 41316 7676 41372
rect 7612 41312 7676 41316
rect 7692 41372 7756 41376
rect 7692 41316 7696 41372
rect 7696 41316 7752 41372
rect 7752 41316 7756 41372
rect 7692 41312 7756 41316
rect 7772 41372 7836 41376
rect 7772 41316 7776 41372
rect 7776 41316 7832 41372
rect 7832 41316 7836 41372
rect 7772 41312 7836 41316
rect 7852 41372 7916 41376
rect 7852 41316 7856 41372
rect 7856 41316 7912 41372
rect 7912 41316 7916 41372
rect 7852 41312 7916 41316
rect 12612 41372 12676 41376
rect 12612 41316 12616 41372
rect 12616 41316 12672 41372
rect 12672 41316 12676 41372
rect 12612 41312 12676 41316
rect 12692 41372 12756 41376
rect 12692 41316 12696 41372
rect 12696 41316 12752 41372
rect 12752 41316 12756 41372
rect 12692 41312 12756 41316
rect 12772 41372 12836 41376
rect 12772 41316 12776 41372
rect 12776 41316 12832 41372
rect 12832 41316 12836 41372
rect 12772 41312 12836 41316
rect 12852 41372 12916 41376
rect 12852 41316 12856 41372
rect 12856 41316 12912 41372
rect 12912 41316 12916 41372
rect 12852 41312 12916 41316
rect 17612 41372 17676 41376
rect 17612 41316 17616 41372
rect 17616 41316 17672 41372
rect 17672 41316 17676 41372
rect 17612 41312 17676 41316
rect 17692 41372 17756 41376
rect 17692 41316 17696 41372
rect 17696 41316 17752 41372
rect 17752 41316 17756 41372
rect 17692 41312 17756 41316
rect 17772 41372 17836 41376
rect 17772 41316 17776 41372
rect 17776 41316 17832 41372
rect 17832 41316 17836 41372
rect 17772 41312 17836 41316
rect 17852 41372 17916 41376
rect 17852 41316 17856 41372
rect 17856 41316 17912 41372
rect 17912 41316 17916 41372
rect 17852 41312 17916 41316
rect 1952 40828 2016 40832
rect 1952 40772 1956 40828
rect 1956 40772 2012 40828
rect 2012 40772 2016 40828
rect 1952 40768 2016 40772
rect 2032 40828 2096 40832
rect 2032 40772 2036 40828
rect 2036 40772 2092 40828
rect 2092 40772 2096 40828
rect 2032 40768 2096 40772
rect 2112 40828 2176 40832
rect 2112 40772 2116 40828
rect 2116 40772 2172 40828
rect 2172 40772 2176 40828
rect 2112 40768 2176 40772
rect 2192 40828 2256 40832
rect 2192 40772 2196 40828
rect 2196 40772 2252 40828
rect 2252 40772 2256 40828
rect 2192 40768 2256 40772
rect 6952 40828 7016 40832
rect 6952 40772 6956 40828
rect 6956 40772 7012 40828
rect 7012 40772 7016 40828
rect 6952 40768 7016 40772
rect 7032 40828 7096 40832
rect 7032 40772 7036 40828
rect 7036 40772 7092 40828
rect 7092 40772 7096 40828
rect 7032 40768 7096 40772
rect 7112 40828 7176 40832
rect 7112 40772 7116 40828
rect 7116 40772 7172 40828
rect 7172 40772 7176 40828
rect 7112 40768 7176 40772
rect 7192 40828 7256 40832
rect 7192 40772 7196 40828
rect 7196 40772 7252 40828
rect 7252 40772 7256 40828
rect 7192 40768 7256 40772
rect 11952 40828 12016 40832
rect 11952 40772 11956 40828
rect 11956 40772 12012 40828
rect 12012 40772 12016 40828
rect 11952 40768 12016 40772
rect 12032 40828 12096 40832
rect 12032 40772 12036 40828
rect 12036 40772 12092 40828
rect 12092 40772 12096 40828
rect 12032 40768 12096 40772
rect 12112 40828 12176 40832
rect 12112 40772 12116 40828
rect 12116 40772 12172 40828
rect 12172 40772 12176 40828
rect 12112 40768 12176 40772
rect 12192 40828 12256 40832
rect 12192 40772 12196 40828
rect 12196 40772 12252 40828
rect 12252 40772 12256 40828
rect 12192 40768 12256 40772
rect 16952 40828 17016 40832
rect 16952 40772 16956 40828
rect 16956 40772 17012 40828
rect 17012 40772 17016 40828
rect 16952 40768 17016 40772
rect 17032 40828 17096 40832
rect 17032 40772 17036 40828
rect 17036 40772 17092 40828
rect 17092 40772 17096 40828
rect 17032 40768 17096 40772
rect 17112 40828 17176 40832
rect 17112 40772 17116 40828
rect 17116 40772 17172 40828
rect 17172 40772 17176 40828
rect 17112 40768 17176 40772
rect 17192 40828 17256 40832
rect 17192 40772 17196 40828
rect 17196 40772 17252 40828
rect 17252 40772 17256 40828
rect 17192 40768 17256 40772
rect 9076 40564 9140 40628
rect 9260 40428 9324 40492
rect 2612 40284 2676 40288
rect 2612 40228 2616 40284
rect 2616 40228 2672 40284
rect 2672 40228 2676 40284
rect 2612 40224 2676 40228
rect 2692 40284 2756 40288
rect 2692 40228 2696 40284
rect 2696 40228 2752 40284
rect 2752 40228 2756 40284
rect 2692 40224 2756 40228
rect 2772 40284 2836 40288
rect 2772 40228 2776 40284
rect 2776 40228 2832 40284
rect 2832 40228 2836 40284
rect 2772 40224 2836 40228
rect 2852 40284 2916 40288
rect 2852 40228 2856 40284
rect 2856 40228 2912 40284
rect 2912 40228 2916 40284
rect 2852 40224 2916 40228
rect 7612 40284 7676 40288
rect 7612 40228 7616 40284
rect 7616 40228 7672 40284
rect 7672 40228 7676 40284
rect 7612 40224 7676 40228
rect 7692 40284 7756 40288
rect 7692 40228 7696 40284
rect 7696 40228 7752 40284
rect 7752 40228 7756 40284
rect 7692 40224 7756 40228
rect 7772 40284 7836 40288
rect 7772 40228 7776 40284
rect 7776 40228 7832 40284
rect 7832 40228 7836 40284
rect 7772 40224 7836 40228
rect 7852 40284 7916 40288
rect 7852 40228 7856 40284
rect 7856 40228 7912 40284
rect 7912 40228 7916 40284
rect 7852 40224 7916 40228
rect 12612 40284 12676 40288
rect 12612 40228 12616 40284
rect 12616 40228 12672 40284
rect 12672 40228 12676 40284
rect 12612 40224 12676 40228
rect 12692 40284 12756 40288
rect 12692 40228 12696 40284
rect 12696 40228 12752 40284
rect 12752 40228 12756 40284
rect 12692 40224 12756 40228
rect 12772 40284 12836 40288
rect 12772 40228 12776 40284
rect 12776 40228 12832 40284
rect 12832 40228 12836 40284
rect 12772 40224 12836 40228
rect 12852 40284 12916 40288
rect 12852 40228 12856 40284
rect 12856 40228 12912 40284
rect 12912 40228 12916 40284
rect 12852 40224 12916 40228
rect 17612 40284 17676 40288
rect 17612 40228 17616 40284
rect 17616 40228 17672 40284
rect 17672 40228 17676 40284
rect 17612 40224 17676 40228
rect 17692 40284 17756 40288
rect 17692 40228 17696 40284
rect 17696 40228 17752 40284
rect 17752 40228 17756 40284
rect 17692 40224 17756 40228
rect 17772 40284 17836 40288
rect 17772 40228 17776 40284
rect 17776 40228 17832 40284
rect 17832 40228 17836 40284
rect 17772 40224 17836 40228
rect 17852 40284 17916 40288
rect 17852 40228 17856 40284
rect 17856 40228 17912 40284
rect 17912 40228 17916 40284
rect 17852 40224 17916 40228
rect 1952 39740 2016 39744
rect 1952 39684 1956 39740
rect 1956 39684 2012 39740
rect 2012 39684 2016 39740
rect 1952 39680 2016 39684
rect 2032 39740 2096 39744
rect 2032 39684 2036 39740
rect 2036 39684 2092 39740
rect 2092 39684 2096 39740
rect 2032 39680 2096 39684
rect 2112 39740 2176 39744
rect 2112 39684 2116 39740
rect 2116 39684 2172 39740
rect 2172 39684 2176 39740
rect 2112 39680 2176 39684
rect 2192 39740 2256 39744
rect 2192 39684 2196 39740
rect 2196 39684 2252 39740
rect 2252 39684 2256 39740
rect 2192 39680 2256 39684
rect 6952 39740 7016 39744
rect 6952 39684 6956 39740
rect 6956 39684 7012 39740
rect 7012 39684 7016 39740
rect 6952 39680 7016 39684
rect 7032 39740 7096 39744
rect 7032 39684 7036 39740
rect 7036 39684 7092 39740
rect 7092 39684 7096 39740
rect 7032 39680 7096 39684
rect 7112 39740 7176 39744
rect 7112 39684 7116 39740
rect 7116 39684 7172 39740
rect 7172 39684 7176 39740
rect 7112 39680 7176 39684
rect 7192 39740 7256 39744
rect 7192 39684 7196 39740
rect 7196 39684 7252 39740
rect 7252 39684 7256 39740
rect 7192 39680 7256 39684
rect 11952 39740 12016 39744
rect 11952 39684 11956 39740
rect 11956 39684 12012 39740
rect 12012 39684 12016 39740
rect 11952 39680 12016 39684
rect 12032 39740 12096 39744
rect 12032 39684 12036 39740
rect 12036 39684 12092 39740
rect 12092 39684 12096 39740
rect 12032 39680 12096 39684
rect 12112 39740 12176 39744
rect 12112 39684 12116 39740
rect 12116 39684 12172 39740
rect 12172 39684 12176 39740
rect 12112 39680 12176 39684
rect 12192 39740 12256 39744
rect 12192 39684 12196 39740
rect 12196 39684 12252 39740
rect 12252 39684 12256 39740
rect 12192 39680 12256 39684
rect 16952 39740 17016 39744
rect 16952 39684 16956 39740
rect 16956 39684 17012 39740
rect 17012 39684 17016 39740
rect 16952 39680 17016 39684
rect 17032 39740 17096 39744
rect 17032 39684 17036 39740
rect 17036 39684 17092 39740
rect 17092 39684 17096 39740
rect 17032 39680 17096 39684
rect 17112 39740 17176 39744
rect 17112 39684 17116 39740
rect 17116 39684 17172 39740
rect 17172 39684 17176 39740
rect 17112 39680 17176 39684
rect 17192 39740 17256 39744
rect 17192 39684 17196 39740
rect 17196 39684 17252 39740
rect 17252 39684 17256 39740
rect 17192 39680 17256 39684
rect 2612 39196 2676 39200
rect 2612 39140 2616 39196
rect 2616 39140 2672 39196
rect 2672 39140 2676 39196
rect 2612 39136 2676 39140
rect 2692 39196 2756 39200
rect 2692 39140 2696 39196
rect 2696 39140 2752 39196
rect 2752 39140 2756 39196
rect 2692 39136 2756 39140
rect 2772 39196 2836 39200
rect 2772 39140 2776 39196
rect 2776 39140 2832 39196
rect 2832 39140 2836 39196
rect 2772 39136 2836 39140
rect 2852 39196 2916 39200
rect 2852 39140 2856 39196
rect 2856 39140 2912 39196
rect 2912 39140 2916 39196
rect 2852 39136 2916 39140
rect 7612 39196 7676 39200
rect 7612 39140 7616 39196
rect 7616 39140 7672 39196
rect 7672 39140 7676 39196
rect 7612 39136 7676 39140
rect 7692 39196 7756 39200
rect 7692 39140 7696 39196
rect 7696 39140 7752 39196
rect 7752 39140 7756 39196
rect 7692 39136 7756 39140
rect 7772 39196 7836 39200
rect 7772 39140 7776 39196
rect 7776 39140 7832 39196
rect 7832 39140 7836 39196
rect 7772 39136 7836 39140
rect 7852 39196 7916 39200
rect 7852 39140 7856 39196
rect 7856 39140 7912 39196
rect 7912 39140 7916 39196
rect 7852 39136 7916 39140
rect 12612 39196 12676 39200
rect 12612 39140 12616 39196
rect 12616 39140 12672 39196
rect 12672 39140 12676 39196
rect 12612 39136 12676 39140
rect 12692 39196 12756 39200
rect 12692 39140 12696 39196
rect 12696 39140 12752 39196
rect 12752 39140 12756 39196
rect 12692 39136 12756 39140
rect 12772 39196 12836 39200
rect 12772 39140 12776 39196
rect 12776 39140 12832 39196
rect 12832 39140 12836 39196
rect 12772 39136 12836 39140
rect 12852 39196 12916 39200
rect 12852 39140 12856 39196
rect 12856 39140 12912 39196
rect 12912 39140 12916 39196
rect 12852 39136 12916 39140
rect 17612 39196 17676 39200
rect 17612 39140 17616 39196
rect 17616 39140 17672 39196
rect 17672 39140 17676 39196
rect 17612 39136 17676 39140
rect 17692 39196 17756 39200
rect 17692 39140 17696 39196
rect 17696 39140 17752 39196
rect 17752 39140 17756 39196
rect 17692 39136 17756 39140
rect 17772 39196 17836 39200
rect 17772 39140 17776 39196
rect 17776 39140 17832 39196
rect 17832 39140 17836 39196
rect 17772 39136 17836 39140
rect 17852 39196 17916 39200
rect 17852 39140 17856 39196
rect 17856 39140 17912 39196
rect 17912 39140 17916 39196
rect 17852 39136 17916 39140
rect 1952 38652 2016 38656
rect 1952 38596 1956 38652
rect 1956 38596 2012 38652
rect 2012 38596 2016 38652
rect 1952 38592 2016 38596
rect 2032 38652 2096 38656
rect 2032 38596 2036 38652
rect 2036 38596 2092 38652
rect 2092 38596 2096 38652
rect 2032 38592 2096 38596
rect 2112 38652 2176 38656
rect 2112 38596 2116 38652
rect 2116 38596 2172 38652
rect 2172 38596 2176 38652
rect 2112 38592 2176 38596
rect 2192 38652 2256 38656
rect 2192 38596 2196 38652
rect 2196 38596 2252 38652
rect 2252 38596 2256 38652
rect 2192 38592 2256 38596
rect 6952 38652 7016 38656
rect 6952 38596 6956 38652
rect 6956 38596 7012 38652
rect 7012 38596 7016 38652
rect 6952 38592 7016 38596
rect 7032 38652 7096 38656
rect 7032 38596 7036 38652
rect 7036 38596 7092 38652
rect 7092 38596 7096 38652
rect 7032 38592 7096 38596
rect 7112 38652 7176 38656
rect 7112 38596 7116 38652
rect 7116 38596 7172 38652
rect 7172 38596 7176 38652
rect 7112 38592 7176 38596
rect 7192 38652 7256 38656
rect 7192 38596 7196 38652
rect 7196 38596 7252 38652
rect 7252 38596 7256 38652
rect 7192 38592 7256 38596
rect 11952 38652 12016 38656
rect 11952 38596 11956 38652
rect 11956 38596 12012 38652
rect 12012 38596 12016 38652
rect 11952 38592 12016 38596
rect 12032 38652 12096 38656
rect 12032 38596 12036 38652
rect 12036 38596 12092 38652
rect 12092 38596 12096 38652
rect 12032 38592 12096 38596
rect 12112 38652 12176 38656
rect 12112 38596 12116 38652
rect 12116 38596 12172 38652
rect 12172 38596 12176 38652
rect 12112 38592 12176 38596
rect 12192 38652 12256 38656
rect 12192 38596 12196 38652
rect 12196 38596 12252 38652
rect 12252 38596 12256 38652
rect 12192 38592 12256 38596
rect 16952 38652 17016 38656
rect 16952 38596 16956 38652
rect 16956 38596 17012 38652
rect 17012 38596 17016 38652
rect 16952 38592 17016 38596
rect 17032 38652 17096 38656
rect 17032 38596 17036 38652
rect 17036 38596 17092 38652
rect 17092 38596 17096 38652
rect 17032 38592 17096 38596
rect 17112 38652 17176 38656
rect 17112 38596 17116 38652
rect 17116 38596 17172 38652
rect 17172 38596 17176 38652
rect 17112 38592 17176 38596
rect 17192 38652 17256 38656
rect 17192 38596 17196 38652
rect 17196 38596 17252 38652
rect 17252 38596 17256 38652
rect 17192 38592 17256 38596
rect 2612 38108 2676 38112
rect 2612 38052 2616 38108
rect 2616 38052 2672 38108
rect 2672 38052 2676 38108
rect 2612 38048 2676 38052
rect 2692 38108 2756 38112
rect 2692 38052 2696 38108
rect 2696 38052 2752 38108
rect 2752 38052 2756 38108
rect 2692 38048 2756 38052
rect 2772 38108 2836 38112
rect 2772 38052 2776 38108
rect 2776 38052 2832 38108
rect 2832 38052 2836 38108
rect 2772 38048 2836 38052
rect 2852 38108 2916 38112
rect 2852 38052 2856 38108
rect 2856 38052 2912 38108
rect 2912 38052 2916 38108
rect 2852 38048 2916 38052
rect 7612 38108 7676 38112
rect 7612 38052 7616 38108
rect 7616 38052 7672 38108
rect 7672 38052 7676 38108
rect 7612 38048 7676 38052
rect 7692 38108 7756 38112
rect 7692 38052 7696 38108
rect 7696 38052 7752 38108
rect 7752 38052 7756 38108
rect 7692 38048 7756 38052
rect 7772 38108 7836 38112
rect 7772 38052 7776 38108
rect 7776 38052 7832 38108
rect 7832 38052 7836 38108
rect 7772 38048 7836 38052
rect 7852 38108 7916 38112
rect 7852 38052 7856 38108
rect 7856 38052 7912 38108
rect 7912 38052 7916 38108
rect 7852 38048 7916 38052
rect 12612 38108 12676 38112
rect 12612 38052 12616 38108
rect 12616 38052 12672 38108
rect 12672 38052 12676 38108
rect 12612 38048 12676 38052
rect 12692 38108 12756 38112
rect 12692 38052 12696 38108
rect 12696 38052 12752 38108
rect 12752 38052 12756 38108
rect 12692 38048 12756 38052
rect 12772 38108 12836 38112
rect 12772 38052 12776 38108
rect 12776 38052 12832 38108
rect 12832 38052 12836 38108
rect 12772 38048 12836 38052
rect 12852 38108 12916 38112
rect 12852 38052 12856 38108
rect 12856 38052 12912 38108
rect 12912 38052 12916 38108
rect 12852 38048 12916 38052
rect 17612 38108 17676 38112
rect 17612 38052 17616 38108
rect 17616 38052 17672 38108
rect 17672 38052 17676 38108
rect 17612 38048 17676 38052
rect 17692 38108 17756 38112
rect 17692 38052 17696 38108
rect 17696 38052 17752 38108
rect 17752 38052 17756 38108
rect 17692 38048 17756 38052
rect 17772 38108 17836 38112
rect 17772 38052 17776 38108
rect 17776 38052 17832 38108
rect 17832 38052 17836 38108
rect 17772 38048 17836 38052
rect 17852 38108 17916 38112
rect 17852 38052 17856 38108
rect 17856 38052 17912 38108
rect 17912 38052 17916 38108
rect 17852 38048 17916 38052
rect 1952 37564 2016 37568
rect 1952 37508 1956 37564
rect 1956 37508 2012 37564
rect 2012 37508 2016 37564
rect 1952 37504 2016 37508
rect 2032 37564 2096 37568
rect 2032 37508 2036 37564
rect 2036 37508 2092 37564
rect 2092 37508 2096 37564
rect 2032 37504 2096 37508
rect 2112 37564 2176 37568
rect 2112 37508 2116 37564
rect 2116 37508 2172 37564
rect 2172 37508 2176 37564
rect 2112 37504 2176 37508
rect 2192 37564 2256 37568
rect 2192 37508 2196 37564
rect 2196 37508 2252 37564
rect 2252 37508 2256 37564
rect 2192 37504 2256 37508
rect 6952 37564 7016 37568
rect 6952 37508 6956 37564
rect 6956 37508 7012 37564
rect 7012 37508 7016 37564
rect 6952 37504 7016 37508
rect 7032 37564 7096 37568
rect 7032 37508 7036 37564
rect 7036 37508 7092 37564
rect 7092 37508 7096 37564
rect 7032 37504 7096 37508
rect 7112 37564 7176 37568
rect 7112 37508 7116 37564
rect 7116 37508 7172 37564
rect 7172 37508 7176 37564
rect 7112 37504 7176 37508
rect 7192 37564 7256 37568
rect 7192 37508 7196 37564
rect 7196 37508 7252 37564
rect 7252 37508 7256 37564
rect 7192 37504 7256 37508
rect 11952 37564 12016 37568
rect 11952 37508 11956 37564
rect 11956 37508 12012 37564
rect 12012 37508 12016 37564
rect 11952 37504 12016 37508
rect 12032 37564 12096 37568
rect 12032 37508 12036 37564
rect 12036 37508 12092 37564
rect 12092 37508 12096 37564
rect 12032 37504 12096 37508
rect 12112 37564 12176 37568
rect 12112 37508 12116 37564
rect 12116 37508 12172 37564
rect 12172 37508 12176 37564
rect 12112 37504 12176 37508
rect 12192 37564 12256 37568
rect 12192 37508 12196 37564
rect 12196 37508 12252 37564
rect 12252 37508 12256 37564
rect 12192 37504 12256 37508
rect 16952 37564 17016 37568
rect 16952 37508 16956 37564
rect 16956 37508 17012 37564
rect 17012 37508 17016 37564
rect 16952 37504 17016 37508
rect 17032 37564 17096 37568
rect 17032 37508 17036 37564
rect 17036 37508 17092 37564
rect 17092 37508 17096 37564
rect 17032 37504 17096 37508
rect 17112 37564 17176 37568
rect 17112 37508 17116 37564
rect 17116 37508 17172 37564
rect 17172 37508 17176 37564
rect 17112 37504 17176 37508
rect 17192 37564 17256 37568
rect 17192 37508 17196 37564
rect 17196 37508 17252 37564
rect 17252 37508 17256 37564
rect 17192 37504 17256 37508
rect 15148 37300 15212 37364
rect 2612 37020 2676 37024
rect 2612 36964 2616 37020
rect 2616 36964 2672 37020
rect 2672 36964 2676 37020
rect 2612 36960 2676 36964
rect 2692 37020 2756 37024
rect 2692 36964 2696 37020
rect 2696 36964 2752 37020
rect 2752 36964 2756 37020
rect 2692 36960 2756 36964
rect 2772 37020 2836 37024
rect 2772 36964 2776 37020
rect 2776 36964 2832 37020
rect 2832 36964 2836 37020
rect 2772 36960 2836 36964
rect 2852 37020 2916 37024
rect 2852 36964 2856 37020
rect 2856 36964 2912 37020
rect 2912 36964 2916 37020
rect 2852 36960 2916 36964
rect 7612 37020 7676 37024
rect 7612 36964 7616 37020
rect 7616 36964 7672 37020
rect 7672 36964 7676 37020
rect 7612 36960 7676 36964
rect 7692 37020 7756 37024
rect 7692 36964 7696 37020
rect 7696 36964 7752 37020
rect 7752 36964 7756 37020
rect 7692 36960 7756 36964
rect 7772 37020 7836 37024
rect 7772 36964 7776 37020
rect 7776 36964 7832 37020
rect 7832 36964 7836 37020
rect 7772 36960 7836 36964
rect 7852 37020 7916 37024
rect 7852 36964 7856 37020
rect 7856 36964 7912 37020
rect 7912 36964 7916 37020
rect 7852 36960 7916 36964
rect 12612 37020 12676 37024
rect 12612 36964 12616 37020
rect 12616 36964 12672 37020
rect 12672 36964 12676 37020
rect 12612 36960 12676 36964
rect 12692 37020 12756 37024
rect 12692 36964 12696 37020
rect 12696 36964 12752 37020
rect 12752 36964 12756 37020
rect 12692 36960 12756 36964
rect 12772 37020 12836 37024
rect 12772 36964 12776 37020
rect 12776 36964 12832 37020
rect 12832 36964 12836 37020
rect 12772 36960 12836 36964
rect 12852 37020 12916 37024
rect 12852 36964 12856 37020
rect 12856 36964 12912 37020
rect 12912 36964 12916 37020
rect 12852 36960 12916 36964
rect 17612 37020 17676 37024
rect 17612 36964 17616 37020
rect 17616 36964 17672 37020
rect 17672 36964 17676 37020
rect 17612 36960 17676 36964
rect 17692 37020 17756 37024
rect 17692 36964 17696 37020
rect 17696 36964 17752 37020
rect 17752 36964 17756 37020
rect 17692 36960 17756 36964
rect 17772 37020 17836 37024
rect 17772 36964 17776 37020
rect 17776 36964 17832 37020
rect 17832 36964 17836 37020
rect 17772 36960 17836 36964
rect 17852 37020 17916 37024
rect 17852 36964 17856 37020
rect 17856 36964 17912 37020
rect 17912 36964 17916 37020
rect 17852 36960 17916 36964
rect 1952 36476 2016 36480
rect 1952 36420 1956 36476
rect 1956 36420 2012 36476
rect 2012 36420 2016 36476
rect 1952 36416 2016 36420
rect 2032 36476 2096 36480
rect 2032 36420 2036 36476
rect 2036 36420 2092 36476
rect 2092 36420 2096 36476
rect 2032 36416 2096 36420
rect 2112 36476 2176 36480
rect 2112 36420 2116 36476
rect 2116 36420 2172 36476
rect 2172 36420 2176 36476
rect 2112 36416 2176 36420
rect 2192 36476 2256 36480
rect 2192 36420 2196 36476
rect 2196 36420 2252 36476
rect 2252 36420 2256 36476
rect 2192 36416 2256 36420
rect 6952 36476 7016 36480
rect 6952 36420 6956 36476
rect 6956 36420 7012 36476
rect 7012 36420 7016 36476
rect 6952 36416 7016 36420
rect 7032 36476 7096 36480
rect 7032 36420 7036 36476
rect 7036 36420 7092 36476
rect 7092 36420 7096 36476
rect 7032 36416 7096 36420
rect 7112 36476 7176 36480
rect 7112 36420 7116 36476
rect 7116 36420 7172 36476
rect 7172 36420 7176 36476
rect 7112 36416 7176 36420
rect 7192 36476 7256 36480
rect 7192 36420 7196 36476
rect 7196 36420 7252 36476
rect 7252 36420 7256 36476
rect 7192 36416 7256 36420
rect 11952 36476 12016 36480
rect 11952 36420 11956 36476
rect 11956 36420 12012 36476
rect 12012 36420 12016 36476
rect 11952 36416 12016 36420
rect 12032 36476 12096 36480
rect 12032 36420 12036 36476
rect 12036 36420 12092 36476
rect 12092 36420 12096 36476
rect 12032 36416 12096 36420
rect 12112 36476 12176 36480
rect 12112 36420 12116 36476
rect 12116 36420 12172 36476
rect 12172 36420 12176 36476
rect 12112 36416 12176 36420
rect 12192 36476 12256 36480
rect 12192 36420 12196 36476
rect 12196 36420 12252 36476
rect 12252 36420 12256 36476
rect 12192 36416 12256 36420
rect 16952 36476 17016 36480
rect 16952 36420 16956 36476
rect 16956 36420 17012 36476
rect 17012 36420 17016 36476
rect 16952 36416 17016 36420
rect 17032 36476 17096 36480
rect 17032 36420 17036 36476
rect 17036 36420 17092 36476
rect 17092 36420 17096 36476
rect 17032 36416 17096 36420
rect 17112 36476 17176 36480
rect 17112 36420 17116 36476
rect 17116 36420 17172 36476
rect 17172 36420 17176 36476
rect 17112 36416 17176 36420
rect 17192 36476 17256 36480
rect 17192 36420 17196 36476
rect 17196 36420 17252 36476
rect 17252 36420 17256 36476
rect 17192 36416 17256 36420
rect 9812 36348 9876 36412
rect 2612 35932 2676 35936
rect 2612 35876 2616 35932
rect 2616 35876 2672 35932
rect 2672 35876 2676 35932
rect 2612 35872 2676 35876
rect 2692 35932 2756 35936
rect 2692 35876 2696 35932
rect 2696 35876 2752 35932
rect 2752 35876 2756 35932
rect 2692 35872 2756 35876
rect 2772 35932 2836 35936
rect 2772 35876 2776 35932
rect 2776 35876 2832 35932
rect 2832 35876 2836 35932
rect 2772 35872 2836 35876
rect 2852 35932 2916 35936
rect 2852 35876 2856 35932
rect 2856 35876 2912 35932
rect 2912 35876 2916 35932
rect 2852 35872 2916 35876
rect 7612 35932 7676 35936
rect 7612 35876 7616 35932
rect 7616 35876 7672 35932
rect 7672 35876 7676 35932
rect 7612 35872 7676 35876
rect 7692 35932 7756 35936
rect 7692 35876 7696 35932
rect 7696 35876 7752 35932
rect 7752 35876 7756 35932
rect 7692 35872 7756 35876
rect 7772 35932 7836 35936
rect 7772 35876 7776 35932
rect 7776 35876 7832 35932
rect 7832 35876 7836 35932
rect 7772 35872 7836 35876
rect 7852 35932 7916 35936
rect 7852 35876 7856 35932
rect 7856 35876 7912 35932
rect 7912 35876 7916 35932
rect 7852 35872 7916 35876
rect 12612 35932 12676 35936
rect 12612 35876 12616 35932
rect 12616 35876 12672 35932
rect 12672 35876 12676 35932
rect 12612 35872 12676 35876
rect 12692 35932 12756 35936
rect 12692 35876 12696 35932
rect 12696 35876 12752 35932
rect 12752 35876 12756 35932
rect 12692 35872 12756 35876
rect 12772 35932 12836 35936
rect 12772 35876 12776 35932
rect 12776 35876 12832 35932
rect 12832 35876 12836 35932
rect 12772 35872 12836 35876
rect 12852 35932 12916 35936
rect 12852 35876 12856 35932
rect 12856 35876 12912 35932
rect 12912 35876 12916 35932
rect 12852 35872 12916 35876
rect 17612 35932 17676 35936
rect 17612 35876 17616 35932
rect 17616 35876 17672 35932
rect 17672 35876 17676 35932
rect 17612 35872 17676 35876
rect 17692 35932 17756 35936
rect 17692 35876 17696 35932
rect 17696 35876 17752 35932
rect 17752 35876 17756 35932
rect 17692 35872 17756 35876
rect 17772 35932 17836 35936
rect 17772 35876 17776 35932
rect 17776 35876 17832 35932
rect 17832 35876 17836 35932
rect 17772 35872 17836 35876
rect 17852 35932 17916 35936
rect 17852 35876 17856 35932
rect 17856 35876 17912 35932
rect 17912 35876 17916 35932
rect 17852 35872 17916 35876
rect 10916 35668 10980 35732
rect 3372 35532 3436 35596
rect 1952 35388 2016 35392
rect 1952 35332 1956 35388
rect 1956 35332 2012 35388
rect 2012 35332 2016 35388
rect 1952 35328 2016 35332
rect 2032 35388 2096 35392
rect 2032 35332 2036 35388
rect 2036 35332 2092 35388
rect 2092 35332 2096 35388
rect 2032 35328 2096 35332
rect 2112 35388 2176 35392
rect 2112 35332 2116 35388
rect 2116 35332 2172 35388
rect 2172 35332 2176 35388
rect 2112 35328 2176 35332
rect 2192 35388 2256 35392
rect 2192 35332 2196 35388
rect 2196 35332 2252 35388
rect 2252 35332 2256 35388
rect 2192 35328 2256 35332
rect 6952 35388 7016 35392
rect 6952 35332 6956 35388
rect 6956 35332 7012 35388
rect 7012 35332 7016 35388
rect 6952 35328 7016 35332
rect 7032 35388 7096 35392
rect 7032 35332 7036 35388
rect 7036 35332 7092 35388
rect 7092 35332 7096 35388
rect 7032 35328 7096 35332
rect 7112 35388 7176 35392
rect 7112 35332 7116 35388
rect 7116 35332 7172 35388
rect 7172 35332 7176 35388
rect 7112 35328 7176 35332
rect 7192 35388 7256 35392
rect 7192 35332 7196 35388
rect 7196 35332 7252 35388
rect 7252 35332 7256 35388
rect 7192 35328 7256 35332
rect 11952 35388 12016 35392
rect 11952 35332 11956 35388
rect 11956 35332 12012 35388
rect 12012 35332 12016 35388
rect 11952 35328 12016 35332
rect 12032 35388 12096 35392
rect 12032 35332 12036 35388
rect 12036 35332 12092 35388
rect 12092 35332 12096 35388
rect 12032 35328 12096 35332
rect 12112 35388 12176 35392
rect 12112 35332 12116 35388
rect 12116 35332 12172 35388
rect 12172 35332 12176 35388
rect 12112 35328 12176 35332
rect 12192 35388 12256 35392
rect 12192 35332 12196 35388
rect 12196 35332 12252 35388
rect 12252 35332 12256 35388
rect 12192 35328 12256 35332
rect 16952 35388 17016 35392
rect 16952 35332 16956 35388
rect 16956 35332 17012 35388
rect 17012 35332 17016 35388
rect 16952 35328 17016 35332
rect 17032 35388 17096 35392
rect 17032 35332 17036 35388
rect 17036 35332 17092 35388
rect 17092 35332 17096 35388
rect 17032 35328 17096 35332
rect 17112 35388 17176 35392
rect 17112 35332 17116 35388
rect 17116 35332 17172 35388
rect 17172 35332 17176 35388
rect 17112 35328 17176 35332
rect 17192 35388 17256 35392
rect 17192 35332 17196 35388
rect 17196 35332 17252 35388
rect 17252 35332 17256 35388
rect 17192 35328 17256 35332
rect 2612 34844 2676 34848
rect 2612 34788 2616 34844
rect 2616 34788 2672 34844
rect 2672 34788 2676 34844
rect 2612 34784 2676 34788
rect 2692 34844 2756 34848
rect 2692 34788 2696 34844
rect 2696 34788 2752 34844
rect 2752 34788 2756 34844
rect 2692 34784 2756 34788
rect 2772 34844 2836 34848
rect 2772 34788 2776 34844
rect 2776 34788 2832 34844
rect 2832 34788 2836 34844
rect 2772 34784 2836 34788
rect 2852 34844 2916 34848
rect 2852 34788 2856 34844
rect 2856 34788 2912 34844
rect 2912 34788 2916 34844
rect 2852 34784 2916 34788
rect 7612 34844 7676 34848
rect 7612 34788 7616 34844
rect 7616 34788 7672 34844
rect 7672 34788 7676 34844
rect 7612 34784 7676 34788
rect 7692 34844 7756 34848
rect 7692 34788 7696 34844
rect 7696 34788 7752 34844
rect 7752 34788 7756 34844
rect 7692 34784 7756 34788
rect 7772 34844 7836 34848
rect 7772 34788 7776 34844
rect 7776 34788 7832 34844
rect 7832 34788 7836 34844
rect 7772 34784 7836 34788
rect 7852 34844 7916 34848
rect 7852 34788 7856 34844
rect 7856 34788 7912 34844
rect 7912 34788 7916 34844
rect 7852 34784 7916 34788
rect 12612 34844 12676 34848
rect 12612 34788 12616 34844
rect 12616 34788 12672 34844
rect 12672 34788 12676 34844
rect 12612 34784 12676 34788
rect 12692 34844 12756 34848
rect 12692 34788 12696 34844
rect 12696 34788 12752 34844
rect 12752 34788 12756 34844
rect 12692 34784 12756 34788
rect 12772 34844 12836 34848
rect 12772 34788 12776 34844
rect 12776 34788 12832 34844
rect 12832 34788 12836 34844
rect 12772 34784 12836 34788
rect 12852 34844 12916 34848
rect 12852 34788 12856 34844
rect 12856 34788 12912 34844
rect 12912 34788 12916 34844
rect 12852 34784 12916 34788
rect 17612 34844 17676 34848
rect 17612 34788 17616 34844
rect 17616 34788 17672 34844
rect 17672 34788 17676 34844
rect 17612 34784 17676 34788
rect 17692 34844 17756 34848
rect 17692 34788 17696 34844
rect 17696 34788 17752 34844
rect 17752 34788 17756 34844
rect 17692 34784 17756 34788
rect 17772 34844 17836 34848
rect 17772 34788 17776 34844
rect 17776 34788 17832 34844
rect 17832 34788 17836 34844
rect 17772 34784 17836 34788
rect 17852 34844 17916 34848
rect 17852 34788 17856 34844
rect 17856 34788 17912 34844
rect 17912 34788 17916 34844
rect 17852 34784 17916 34788
rect 1952 34300 2016 34304
rect 1952 34244 1956 34300
rect 1956 34244 2012 34300
rect 2012 34244 2016 34300
rect 1952 34240 2016 34244
rect 2032 34300 2096 34304
rect 2032 34244 2036 34300
rect 2036 34244 2092 34300
rect 2092 34244 2096 34300
rect 2032 34240 2096 34244
rect 2112 34300 2176 34304
rect 2112 34244 2116 34300
rect 2116 34244 2172 34300
rect 2172 34244 2176 34300
rect 2112 34240 2176 34244
rect 2192 34300 2256 34304
rect 2192 34244 2196 34300
rect 2196 34244 2252 34300
rect 2252 34244 2256 34300
rect 2192 34240 2256 34244
rect 6952 34300 7016 34304
rect 6952 34244 6956 34300
rect 6956 34244 7012 34300
rect 7012 34244 7016 34300
rect 6952 34240 7016 34244
rect 7032 34300 7096 34304
rect 7032 34244 7036 34300
rect 7036 34244 7092 34300
rect 7092 34244 7096 34300
rect 7032 34240 7096 34244
rect 7112 34300 7176 34304
rect 7112 34244 7116 34300
rect 7116 34244 7172 34300
rect 7172 34244 7176 34300
rect 7112 34240 7176 34244
rect 7192 34300 7256 34304
rect 7192 34244 7196 34300
rect 7196 34244 7252 34300
rect 7252 34244 7256 34300
rect 7192 34240 7256 34244
rect 11952 34300 12016 34304
rect 11952 34244 11956 34300
rect 11956 34244 12012 34300
rect 12012 34244 12016 34300
rect 11952 34240 12016 34244
rect 12032 34300 12096 34304
rect 12032 34244 12036 34300
rect 12036 34244 12092 34300
rect 12092 34244 12096 34300
rect 12032 34240 12096 34244
rect 12112 34300 12176 34304
rect 12112 34244 12116 34300
rect 12116 34244 12172 34300
rect 12172 34244 12176 34300
rect 12112 34240 12176 34244
rect 12192 34300 12256 34304
rect 12192 34244 12196 34300
rect 12196 34244 12252 34300
rect 12252 34244 12256 34300
rect 12192 34240 12256 34244
rect 16952 34300 17016 34304
rect 16952 34244 16956 34300
rect 16956 34244 17012 34300
rect 17012 34244 17016 34300
rect 16952 34240 17016 34244
rect 17032 34300 17096 34304
rect 17032 34244 17036 34300
rect 17036 34244 17092 34300
rect 17092 34244 17096 34300
rect 17032 34240 17096 34244
rect 17112 34300 17176 34304
rect 17112 34244 17116 34300
rect 17116 34244 17172 34300
rect 17172 34244 17176 34300
rect 17112 34240 17176 34244
rect 17192 34300 17256 34304
rect 17192 34244 17196 34300
rect 17196 34244 17252 34300
rect 17252 34244 17256 34300
rect 17192 34240 17256 34244
rect 2612 33756 2676 33760
rect 2612 33700 2616 33756
rect 2616 33700 2672 33756
rect 2672 33700 2676 33756
rect 2612 33696 2676 33700
rect 2692 33756 2756 33760
rect 2692 33700 2696 33756
rect 2696 33700 2752 33756
rect 2752 33700 2756 33756
rect 2692 33696 2756 33700
rect 2772 33756 2836 33760
rect 2772 33700 2776 33756
rect 2776 33700 2832 33756
rect 2832 33700 2836 33756
rect 2772 33696 2836 33700
rect 2852 33756 2916 33760
rect 2852 33700 2856 33756
rect 2856 33700 2912 33756
rect 2912 33700 2916 33756
rect 2852 33696 2916 33700
rect 7612 33756 7676 33760
rect 7612 33700 7616 33756
rect 7616 33700 7672 33756
rect 7672 33700 7676 33756
rect 7612 33696 7676 33700
rect 7692 33756 7756 33760
rect 7692 33700 7696 33756
rect 7696 33700 7752 33756
rect 7752 33700 7756 33756
rect 7692 33696 7756 33700
rect 7772 33756 7836 33760
rect 7772 33700 7776 33756
rect 7776 33700 7832 33756
rect 7832 33700 7836 33756
rect 7772 33696 7836 33700
rect 7852 33756 7916 33760
rect 7852 33700 7856 33756
rect 7856 33700 7912 33756
rect 7912 33700 7916 33756
rect 7852 33696 7916 33700
rect 12612 33756 12676 33760
rect 12612 33700 12616 33756
rect 12616 33700 12672 33756
rect 12672 33700 12676 33756
rect 12612 33696 12676 33700
rect 12692 33756 12756 33760
rect 12692 33700 12696 33756
rect 12696 33700 12752 33756
rect 12752 33700 12756 33756
rect 12692 33696 12756 33700
rect 12772 33756 12836 33760
rect 12772 33700 12776 33756
rect 12776 33700 12832 33756
rect 12832 33700 12836 33756
rect 12772 33696 12836 33700
rect 12852 33756 12916 33760
rect 12852 33700 12856 33756
rect 12856 33700 12912 33756
rect 12912 33700 12916 33756
rect 12852 33696 12916 33700
rect 17612 33756 17676 33760
rect 17612 33700 17616 33756
rect 17616 33700 17672 33756
rect 17672 33700 17676 33756
rect 17612 33696 17676 33700
rect 17692 33756 17756 33760
rect 17692 33700 17696 33756
rect 17696 33700 17752 33756
rect 17752 33700 17756 33756
rect 17692 33696 17756 33700
rect 17772 33756 17836 33760
rect 17772 33700 17776 33756
rect 17776 33700 17832 33756
rect 17832 33700 17836 33756
rect 17772 33696 17836 33700
rect 17852 33756 17916 33760
rect 17852 33700 17856 33756
rect 17856 33700 17912 33756
rect 17912 33700 17916 33756
rect 17852 33696 17916 33700
rect 1952 33212 2016 33216
rect 1952 33156 1956 33212
rect 1956 33156 2012 33212
rect 2012 33156 2016 33212
rect 1952 33152 2016 33156
rect 2032 33212 2096 33216
rect 2032 33156 2036 33212
rect 2036 33156 2092 33212
rect 2092 33156 2096 33212
rect 2032 33152 2096 33156
rect 2112 33212 2176 33216
rect 2112 33156 2116 33212
rect 2116 33156 2172 33212
rect 2172 33156 2176 33212
rect 2112 33152 2176 33156
rect 2192 33212 2256 33216
rect 2192 33156 2196 33212
rect 2196 33156 2252 33212
rect 2252 33156 2256 33212
rect 2192 33152 2256 33156
rect 6952 33212 7016 33216
rect 6952 33156 6956 33212
rect 6956 33156 7012 33212
rect 7012 33156 7016 33212
rect 6952 33152 7016 33156
rect 7032 33212 7096 33216
rect 7032 33156 7036 33212
rect 7036 33156 7092 33212
rect 7092 33156 7096 33212
rect 7032 33152 7096 33156
rect 7112 33212 7176 33216
rect 7112 33156 7116 33212
rect 7116 33156 7172 33212
rect 7172 33156 7176 33212
rect 7112 33152 7176 33156
rect 7192 33212 7256 33216
rect 7192 33156 7196 33212
rect 7196 33156 7252 33212
rect 7252 33156 7256 33212
rect 7192 33152 7256 33156
rect 11952 33212 12016 33216
rect 11952 33156 11956 33212
rect 11956 33156 12012 33212
rect 12012 33156 12016 33212
rect 11952 33152 12016 33156
rect 12032 33212 12096 33216
rect 12032 33156 12036 33212
rect 12036 33156 12092 33212
rect 12092 33156 12096 33212
rect 12032 33152 12096 33156
rect 12112 33212 12176 33216
rect 12112 33156 12116 33212
rect 12116 33156 12172 33212
rect 12172 33156 12176 33212
rect 12112 33152 12176 33156
rect 12192 33212 12256 33216
rect 12192 33156 12196 33212
rect 12196 33156 12252 33212
rect 12252 33156 12256 33212
rect 12192 33152 12256 33156
rect 16952 33212 17016 33216
rect 16952 33156 16956 33212
rect 16956 33156 17012 33212
rect 17012 33156 17016 33212
rect 16952 33152 17016 33156
rect 17032 33212 17096 33216
rect 17032 33156 17036 33212
rect 17036 33156 17092 33212
rect 17092 33156 17096 33212
rect 17032 33152 17096 33156
rect 17112 33212 17176 33216
rect 17112 33156 17116 33212
rect 17116 33156 17172 33212
rect 17172 33156 17176 33212
rect 17112 33152 17176 33156
rect 17192 33212 17256 33216
rect 17192 33156 17196 33212
rect 17196 33156 17252 33212
rect 17252 33156 17256 33212
rect 17192 33152 17256 33156
rect 8708 33084 8772 33148
rect 9076 32948 9140 33012
rect 2612 32668 2676 32672
rect 2612 32612 2616 32668
rect 2616 32612 2672 32668
rect 2672 32612 2676 32668
rect 2612 32608 2676 32612
rect 2692 32668 2756 32672
rect 2692 32612 2696 32668
rect 2696 32612 2752 32668
rect 2752 32612 2756 32668
rect 2692 32608 2756 32612
rect 2772 32668 2836 32672
rect 2772 32612 2776 32668
rect 2776 32612 2832 32668
rect 2832 32612 2836 32668
rect 2772 32608 2836 32612
rect 2852 32668 2916 32672
rect 2852 32612 2856 32668
rect 2856 32612 2912 32668
rect 2912 32612 2916 32668
rect 2852 32608 2916 32612
rect 7612 32668 7676 32672
rect 7612 32612 7616 32668
rect 7616 32612 7672 32668
rect 7672 32612 7676 32668
rect 7612 32608 7676 32612
rect 7692 32668 7756 32672
rect 7692 32612 7696 32668
rect 7696 32612 7752 32668
rect 7752 32612 7756 32668
rect 7692 32608 7756 32612
rect 7772 32668 7836 32672
rect 7772 32612 7776 32668
rect 7776 32612 7832 32668
rect 7832 32612 7836 32668
rect 7772 32608 7836 32612
rect 7852 32668 7916 32672
rect 7852 32612 7856 32668
rect 7856 32612 7912 32668
rect 7912 32612 7916 32668
rect 7852 32608 7916 32612
rect 12612 32668 12676 32672
rect 12612 32612 12616 32668
rect 12616 32612 12672 32668
rect 12672 32612 12676 32668
rect 12612 32608 12676 32612
rect 12692 32668 12756 32672
rect 12692 32612 12696 32668
rect 12696 32612 12752 32668
rect 12752 32612 12756 32668
rect 12692 32608 12756 32612
rect 12772 32668 12836 32672
rect 12772 32612 12776 32668
rect 12776 32612 12832 32668
rect 12832 32612 12836 32668
rect 12772 32608 12836 32612
rect 12852 32668 12916 32672
rect 12852 32612 12856 32668
rect 12856 32612 12912 32668
rect 12912 32612 12916 32668
rect 12852 32608 12916 32612
rect 17612 32668 17676 32672
rect 17612 32612 17616 32668
rect 17616 32612 17672 32668
rect 17672 32612 17676 32668
rect 17612 32608 17676 32612
rect 17692 32668 17756 32672
rect 17692 32612 17696 32668
rect 17696 32612 17752 32668
rect 17752 32612 17756 32668
rect 17692 32608 17756 32612
rect 17772 32668 17836 32672
rect 17772 32612 17776 32668
rect 17776 32612 17832 32668
rect 17832 32612 17836 32668
rect 17772 32608 17836 32612
rect 17852 32668 17916 32672
rect 17852 32612 17856 32668
rect 17856 32612 17912 32668
rect 17912 32612 17916 32668
rect 17852 32608 17916 32612
rect 1952 32124 2016 32128
rect 1952 32068 1956 32124
rect 1956 32068 2012 32124
rect 2012 32068 2016 32124
rect 1952 32064 2016 32068
rect 2032 32124 2096 32128
rect 2032 32068 2036 32124
rect 2036 32068 2092 32124
rect 2092 32068 2096 32124
rect 2032 32064 2096 32068
rect 2112 32124 2176 32128
rect 2112 32068 2116 32124
rect 2116 32068 2172 32124
rect 2172 32068 2176 32124
rect 2112 32064 2176 32068
rect 2192 32124 2256 32128
rect 2192 32068 2196 32124
rect 2196 32068 2252 32124
rect 2252 32068 2256 32124
rect 2192 32064 2256 32068
rect 6952 32124 7016 32128
rect 6952 32068 6956 32124
rect 6956 32068 7012 32124
rect 7012 32068 7016 32124
rect 6952 32064 7016 32068
rect 7032 32124 7096 32128
rect 7032 32068 7036 32124
rect 7036 32068 7092 32124
rect 7092 32068 7096 32124
rect 7032 32064 7096 32068
rect 7112 32124 7176 32128
rect 7112 32068 7116 32124
rect 7116 32068 7172 32124
rect 7172 32068 7176 32124
rect 7112 32064 7176 32068
rect 7192 32124 7256 32128
rect 7192 32068 7196 32124
rect 7196 32068 7252 32124
rect 7252 32068 7256 32124
rect 7192 32064 7256 32068
rect 11952 32124 12016 32128
rect 11952 32068 11956 32124
rect 11956 32068 12012 32124
rect 12012 32068 12016 32124
rect 11952 32064 12016 32068
rect 12032 32124 12096 32128
rect 12032 32068 12036 32124
rect 12036 32068 12092 32124
rect 12092 32068 12096 32124
rect 12032 32064 12096 32068
rect 12112 32124 12176 32128
rect 12112 32068 12116 32124
rect 12116 32068 12172 32124
rect 12172 32068 12176 32124
rect 12112 32064 12176 32068
rect 12192 32124 12256 32128
rect 12192 32068 12196 32124
rect 12196 32068 12252 32124
rect 12252 32068 12256 32124
rect 12192 32064 12256 32068
rect 16952 32124 17016 32128
rect 16952 32068 16956 32124
rect 16956 32068 17012 32124
rect 17012 32068 17016 32124
rect 16952 32064 17016 32068
rect 17032 32124 17096 32128
rect 17032 32068 17036 32124
rect 17036 32068 17092 32124
rect 17092 32068 17096 32124
rect 17032 32064 17096 32068
rect 17112 32124 17176 32128
rect 17112 32068 17116 32124
rect 17116 32068 17172 32124
rect 17172 32068 17176 32124
rect 17112 32064 17176 32068
rect 17192 32124 17256 32128
rect 17192 32068 17196 32124
rect 17196 32068 17252 32124
rect 17252 32068 17256 32124
rect 17192 32064 17256 32068
rect 4844 31724 4908 31788
rect 2612 31580 2676 31584
rect 2612 31524 2616 31580
rect 2616 31524 2672 31580
rect 2672 31524 2676 31580
rect 2612 31520 2676 31524
rect 2692 31580 2756 31584
rect 2692 31524 2696 31580
rect 2696 31524 2752 31580
rect 2752 31524 2756 31580
rect 2692 31520 2756 31524
rect 2772 31580 2836 31584
rect 2772 31524 2776 31580
rect 2776 31524 2832 31580
rect 2832 31524 2836 31580
rect 2772 31520 2836 31524
rect 2852 31580 2916 31584
rect 2852 31524 2856 31580
rect 2856 31524 2912 31580
rect 2912 31524 2916 31580
rect 2852 31520 2916 31524
rect 7612 31580 7676 31584
rect 7612 31524 7616 31580
rect 7616 31524 7672 31580
rect 7672 31524 7676 31580
rect 7612 31520 7676 31524
rect 7692 31580 7756 31584
rect 7692 31524 7696 31580
rect 7696 31524 7752 31580
rect 7752 31524 7756 31580
rect 7692 31520 7756 31524
rect 7772 31580 7836 31584
rect 7772 31524 7776 31580
rect 7776 31524 7832 31580
rect 7832 31524 7836 31580
rect 7772 31520 7836 31524
rect 7852 31580 7916 31584
rect 7852 31524 7856 31580
rect 7856 31524 7912 31580
rect 7912 31524 7916 31580
rect 7852 31520 7916 31524
rect 12612 31580 12676 31584
rect 12612 31524 12616 31580
rect 12616 31524 12672 31580
rect 12672 31524 12676 31580
rect 12612 31520 12676 31524
rect 12692 31580 12756 31584
rect 12692 31524 12696 31580
rect 12696 31524 12752 31580
rect 12752 31524 12756 31580
rect 12692 31520 12756 31524
rect 12772 31580 12836 31584
rect 12772 31524 12776 31580
rect 12776 31524 12832 31580
rect 12832 31524 12836 31580
rect 12772 31520 12836 31524
rect 12852 31580 12916 31584
rect 12852 31524 12856 31580
rect 12856 31524 12912 31580
rect 12912 31524 12916 31580
rect 12852 31520 12916 31524
rect 17612 31580 17676 31584
rect 17612 31524 17616 31580
rect 17616 31524 17672 31580
rect 17672 31524 17676 31580
rect 17612 31520 17676 31524
rect 17692 31580 17756 31584
rect 17692 31524 17696 31580
rect 17696 31524 17752 31580
rect 17752 31524 17756 31580
rect 17692 31520 17756 31524
rect 17772 31580 17836 31584
rect 17772 31524 17776 31580
rect 17776 31524 17832 31580
rect 17832 31524 17836 31580
rect 17772 31520 17836 31524
rect 17852 31580 17916 31584
rect 17852 31524 17856 31580
rect 17856 31524 17912 31580
rect 17912 31524 17916 31580
rect 17852 31520 17916 31524
rect 1952 31036 2016 31040
rect 1952 30980 1956 31036
rect 1956 30980 2012 31036
rect 2012 30980 2016 31036
rect 1952 30976 2016 30980
rect 2032 31036 2096 31040
rect 2032 30980 2036 31036
rect 2036 30980 2092 31036
rect 2092 30980 2096 31036
rect 2032 30976 2096 30980
rect 2112 31036 2176 31040
rect 2112 30980 2116 31036
rect 2116 30980 2172 31036
rect 2172 30980 2176 31036
rect 2112 30976 2176 30980
rect 2192 31036 2256 31040
rect 2192 30980 2196 31036
rect 2196 30980 2252 31036
rect 2252 30980 2256 31036
rect 2192 30976 2256 30980
rect 6952 31036 7016 31040
rect 6952 30980 6956 31036
rect 6956 30980 7012 31036
rect 7012 30980 7016 31036
rect 6952 30976 7016 30980
rect 7032 31036 7096 31040
rect 7032 30980 7036 31036
rect 7036 30980 7092 31036
rect 7092 30980 7096 31036
rect 7032 30976 7096 30980
rect 7112 31036 7176 31040
rect 7112 30980 7116 31036
rect 7116 30980 7172 31036
rect 7172 30980 7176 31036
rect 7112 30976 7176 30980
rect 7192 31036 7256 31040
rect 7192 30980 7196 31036
rect 7196 30980 7252 31036
rect 7252 30980 7256 31036
rect 7192 30976 7256 30980
rect 11952 31036 12016 31040
rect 11952 30980 11956 31036
rect 11956 30980 12012 31036
rect 12012 30980 12016 31036
rect 11952 30976 12016 30980
rect 12032 31036 12096 31040
rect 12032 30980 12036 31036
rect 12036 30980 12092 31036
rect 12092 30980 12096 31036
rect 12032 30976 12096 30980
rect 12112 31036 12176 31040
rect 12112 30980 12116 31036
rect 12116 30980 12172 31036
rect 12172 30980 12176 31036
rect 12112 30976 12176 30980
rect 12192 31036 12256 31040
rect 12192 30980 12196 31036
rect 12196 30980 12252 31036
rect 12252 30980 12256 31036
rect 12192 30976 12256 30980
rect 16952 31036 17016 31040
rect 16952 30980 16956 31036
rect 16956 30980 17012 31036
rect 17012 30980 17016 31036
rect 16952 30976 17016 30980
rect 17032 31036 17096 31040
rect 17032 30980 17036 31036
rect 17036 30980 17092 31036
rect 17092 30980 17096 31036
rect 17032 30976 17096 30980
rect 17112 31036 17176 31040
rect 17112 30980 17116 31036
rect 17116 30980 17172 31036
rect 17172 30980 17176 31036
rect 17112 30976 17176 30980
rect 17192 31036 17256 31040
rect 17192 30980 17196 31036
rect 17196 30980 17252 31036
rect 17252 30980 17256 31036
rect 17192 30976 17256 30980
rect 2612 30492 2676 30496
rect 2612 30436 2616 30492
rect 2616 30436 2672 30492
rect 2672 30436 2676 30492
rect 2612 30432 2676 30436
rect 2692 30492 2756 30496
rect 2692 30436 2696 30492
rect 2696 30436 2752 30492
rect 2752 30436 2756 30492
rect 2692 30432 2756 30436
rect 2772 30492 2836 30496
rect 2772 30436 2776 30492
rect 2776 30436 2832 30492
rect 2832 30436 2836 30492
rect 2772 30432 2836 30436
rect 2852 30492 2916 30496
rect 2852 30436 2856 30492
rect 2856 30436 2912 30492
rect 2912 30436 2916 30492
rect 2852 30432 2916 30436
rect 7612 30492 7676 30496
rect 7612 30436 7616 30492
rect 7616 30436 7672 30492
rect 7672 30436 7676 30492
rect 7612 30432 7676 30436
rect 7692 30492 7756 30496
rect 7692 30436 7696 30492
rect 7696 30436 7752 30492
rect 7752 30436 7756 30492
rect 7692 30432 7756 30436
rect 7772 30492 7836 30496
rect 7772 30436 7776 30492
rect 7776 30436 7832 30492
rect 7832 30436 7836 30492
rect 7772 30432 7836 30436
rect 7852 30492 7916 30496
rect 7852 30436 7856 30492
rect 7856 30436 7912 30492
rect 7912 30436 7916 30492
rect 7852 30432 7916 30436
rect 12612 30492 12676 30496
rect 12612 30436 12616 30492
rect 12616 30436 12672 30492
rect 12672 30436 12676 30492
rect 12612 30432 12676 30436
rect 12692 30492 12756 30496
rect 12692 30436 12696 30492
rect 12696 30436 12752 30492
rect 12752 30436 12756 30492
rect 12692 30432 12756 30436
rect 12772 30492 12836 30496
rect 12772 30436 12776 30492
rect 12776 30436 12832 30492
rect 12832 30436 12836 30492
rect 12772 30432 12836 30436
rect 12852 30492 12916 30496
rect 12852 30436 12856 30492
rect 12856 30436 12912 30492
rect 12912 30436 12916 30492
rect 12852 30432 12916 30436
rect 17612 30492 17676 30496
rect 17612 30436 17616 30492
rect 17616 30436 17672 30492
rect 17672 30436 17676 30492
rect 17612 30432 17676 30436
rect 17692 30492 17756 30496
rect 17692 30436 17696 30492
rect 17696 30436 17752 30492
rect 17752 30436 17756 30492
rect 17692 30432 17756 30436
rect 17772 30492 17836 30496
rect 17772 30436 17776 30492
rect 17776 30436 17832 30492
rect 17832 30436 17836 30492
rect 17772 30432 17836 30436
rect 17852 30492 17916 30496
rect 17852 30436 17856 30492
rect 17856 30436 17912 30492
rect 17912 30436 17916 30492
rect 17852 30432 17916 30436
rect 1952 29948 2016 29952
rect 1952 29892 1956 29948
rect 1956 29892 2012 29948
rect 2012 29892 2016 29948
rect 1952 29888 2016 29892
rect 2032 29948 2096 29952
rect 2032 29892 2036 29948
rect 2036 29892 2092 29948
rect 2092 29892 2096 29948
rect 2032 29888 2096 29892
rect 2112 29948 2176 29952
rect 2112 29892 2116 29948
rect 2116 29892 2172 29948
rect 2172 29892 2176 29948
rect 2112 29888 2176 29892
rect 2192 29948 2256 29952
rect 2192 29892 2196 29948
rect 2196 29892 2252 29948
rect 2252 29892 2256 29948
rect 2192 29888 2256 29892
rect 6952 29948 7016 29952
rect 6952 29892 6956 29948
rect 6956 29892 7012 29948
rect 7012 29892 7016 29948
rect 6952 29888 7016 29892
rect 7032 29948 7096 29952
rect 7032 29892 7036 29948
rect 7036 29892 7092 29948
rect 7092 29892 7096 29948
rect 7032 29888 7096 29892
rect 7112 29948 7176 29952
rect 7112 29892 7116 29948
rect 7116 29892 7172 29948
rect 7172 29892 7176 29948
rect 7112 29888 7176 29892
rect 7192 29948 7256 29952
rect 7192 29892 7196 29948
rect 7196 29892 7252 29948
rect 7252 29892 7256 29948
rect 7192 29888 7256 29892
rect 11952 29948 12016 29952
rect 11952 29892 11956 29948
rect 11956 29892 12012 29948
rect 12012 29892 12016 29948
rect 11952 29888 12016 29892
rect 12032 29948 12096 29952
rect 12032 29892 12036 29948
rect 12036 29892 12092 29948
rect 12092 29892 12096 29948
rect 12032 29888 12096 29892
rect 12112 29948 12176 29952
rect 12112 29892 12116 29948
rect 12116 29892 12172 29948
rect 12172 29892 12176 29948
rect 12112 29888 12176 29892
rect 12192 29948 12256 29952
rect 12192 29892 12196 29948
rect 12196 29892 12252 29948
rect 12252 29892 12256 29948
rect 12192 29888 12256 29892
rect 16952 29948 17016 29952
rect 16952 29892 16956 29948
rect 16956 29892 17012 29948
rect 17012 29892 17016 29948
rect 16952 29888 17016 29892
rect 17032 29948 17096 29952
rect 17032 29892 17036 29948
rect 17036 29892 17092 29948
rect 17092 29892 17096 29948
rect 17032 29888 17096 29892
rect 17112 29948 17176 29952
rect 17112 29892 17116 29948
rect 17116 29892 17172 29948
rect 17172 29892 17176 29948
rect 17112 29888 17176 29892
rect 17192 29948 17256 29952
rect 17192 29892 17196 29948
rect 17196 29892 17252 29948
rect 17252 29892 17256 29948
rect 17192 29888 17256 29892
rect 14964 29820 15028 29884
rect 2612 29404 2676 29408
rect 2612 29348 2616 29404
rect 2616 29348 2672 29404
rect 2672 29348 2676 29404
rect 2612 29344 2676 29348
rect 2692 29404 2756 29408
rect 2692 29348 2696 29404
rect 2696 29348 2752 29404
rect 2752 29348 2756 29404
rect 2692 29344 2756 29348
rect 2772 29404 2836 29408
rect 2772 29348 2776 29404
rect 2776 29348 2832 29404
rect 2832 29348 2836 29404
rect 2772 29344 2836 29348
rect 2852 29404 2916 29408
rect 2852 29348 2856 29404
rect 2856 29348 2912 29404
rect 2912 29348 2916 29404
rect 2852 29344 2916 29348
rect 7612 29404 7676 29408
rect 7612 29348 7616 29404
rect 7616 29348 7672 29404
rect 7672 29348 7676 29404
rect 7612 29344 7676 29348
rect 7692 29404 7756 29408
rect 7692 29348 7696 29404
rect 7696 29348 7752 29404
rect 7752 29348 7756 29404
rect 7692 29344 7756 29348
rect 7772 29404 7836 29408
rect 7772 29348 7776 29404
rect 7776 29348 7832 29404
rect 7832 29348 7836 29404
rect 7772 29344 7836 29348
rect 7852 29404 7916 29408
rect 7852 29348 7856 29404
rect 7856 29348 7912 29404
rect 7912 29348 7916 29404
rect 7852 29344 7916 29348
rect 12612 29404 12676 29408
rect 12612 29348 12616 29404
rect 12616 29348 12672 29404
rect 12672 29348 12676 29404
rect 12612 29344 12676 29348
rect 12692 29404 12756 29408
rect 12692 29348 12696 29404
rect 12696 29348 12752 29404
rect 12752 29348 12756 29404
rect 12692 29344 12756 29348
rect 12772 29404 12836 29408
rect 12772 29348 12776 29404
rect 12776 29348 12832 29404
rect 12832 29348 12836 29404
rect 12772 29344 12836 29348
rect 12852 29404 12916 29408
rect 12852 29348 12856 29404
rect 12856 29348 12912 29404
rect 12912 29348 12916 29404
rect 12852 29344 12916 29348
rect 17612 29404 17676 29408
rect 17612 29348 17616 29404
rect 17616 29348 17672 29404
rect 17672 29348 17676 29404
rect 17612 29344 17676 29348
rect 17692 29404 17756 29408
rect 17692 29348 17696 29404
rect 17696 29348 17752 29404
rect 17752 29348 17756 29404
rect 17692 29344 17756 29348
rect 17772 29404 17836 29408
rect 17772 29348 17776 29404
rect 17776 29348 17832 29404
rect 17832 29348 17836 29404
rect 17772 29344 17836 29348
rect 17852 29404 17916 29408
rect 17852 29348 17856 29404
rect 17856 29348 17912 29404
rect 17912 29348 17916 29404
rect 17852 29344 17916 29348
rect 1952 28860 2016 28864
rect 1952 28804 1956 28860
rect 1956 28804 2012 28860
rect 2012 28804 2016 28860
rect 1952 28800 2016 28804
rect 2032 28860 2096 28864
rect 2032 28804 2036 28860
rect 2036 28804 2092 28860
rect 2092 28804 2096 28860
rect 2032 28800 2096 28804
rect 2112 28860 2176 28864
rect 2112 28804 2116 28860
rect 2116 28804 2172 28860
rect 2172 28804 2176 28860
rect 2112 28800 2176 28804
rect 2192 28860 2256 28864
rect 2192 28804 2196 28860
rect 2196 28804 2252 28860
rect 2252 28804 2256 28860
rect 2192 28800 2256 28804
rect 6952 28860 7016 28864
rect 6952 28804 6956 28860
rect 6956 28804 7012 28860
rect 7012 28804 7016 28860
rect 6952 28800 7016 28804
rect 7032 28860 7096 28864
rect 7032 28804 7036 28860
rect 7036 28804 7092 28860
rect 7092 28804 7096 28860
rect 7032 28800 7096 28804
rect 7112 28860 7176 28864
rect 7112 28804 7116 28860
rect 7116 28804 7172 28860
rect 7172 28804 7176 28860
rect 7112 28800 7176 28804
rect 7192 28860 7256 28864
rect 7192 28804 7196 28860
rect 7196 28804 7252 28860
rect 7252 28804 7256 28860
rect 7192 28800 7256 28804
rect 11952 28860 12016 28864
rect 11952 28804 11956 28860
rect 11956 28804 12012 28860
rect 12012 28804 12016 28860
rect 11952 28800 12016 28804
rect 12032 28860 12096 28864
rect 12032 28804 12036 28860
rect 12036 28804 12092 28860
rect 12092 28804 12096 28860
rect 12032 28800 12096 28804
rect 12112 28860 12176 28864
rect 12112 28804 12116 28860
rect 12116 28804 12172 28860
rect 12172 28804 12176 28860
rect 12112 28800 12176 28804
rect 12192 28860 12256 28864
rect 12192 28804 12196 28860
rect 12196 28804 12252 28860
rect 12252 28804 12256 28860
rect 12192 28800 12256 28804
rect 16952 28860 17016 28864
rect 16952 28804 16956 28860
rect 16956 28804 17012 28860
rect 17012 28804 17016 28860
rect 16952 28800 17016 28804
rect 17032 28860 17096 28864
rect 17032 28804 17036 28860
rect 17036 28804 17092 28860
rect 17092 28804 17096 28860
rect 17032 28800 17096 28804
rect 17112 28860 17176 28864
rect 17112 28804 17116 28860
rect 17116 28804 17172 28860
rect 17172 28804 17176 28860
rect 17112 28800 17176 28804
rect 17192 28860 17256 28864
rect 17192 28804 17196 28860
rect 17196 28804 17252 28860
rect 17252 28804 17256 28860
rect 17192 28800 17256 28804
rect 8340 28460 8404 28524
rect 2612 28316 2676 28320
rect 2612 28260 2616 28316
rect 2616 28260 2672 28316
rect 2672 28260 2676 28316
rect 2612 28256 2676 28260
rect 2692 28316 2756 28320
rect 2692 28260 2696 28316
rect 2696 28260 2752 28316
rect 2752 28260 2756 28316
rect 2692 28256 2756 28260
rect 2772 28316 2836 28320
rect 2772 28260 2776 28316
rect 2776 28260 2832 28316
rect 2832 28260 2836 28316
rect 2772 28256 2836 28260
rect 2852 28316 2916 28320
rect 2852 28260 2856 28316
rect 2856 28260 2912 28316
rect 2912 28260 2916 28316
rect 2852 28256 2916 28260
rect 7612 28316 7676 28320
rect 7612 28260 7616 28316
rect 7616 28260 7672 28316
rect 7672 28260 7676 28316
rect 7612 28256 7676 28260
rect 7692 28316 7756 28320
rect 7692 28260 7696 28316
rect 7696 28260 7752 28316
rect 7752 28260 7756 28316
rect 7692 28256 7756 28260
rect 7772 28316 7836 28320
rect 7772 28260 7776 28316
rect 7776 28260 7832 28316
rect 7832 28260 7836 28316
rect 7772 28256 7836 28260
rect 7852 28316 7916 28320
rect 7852 28260 7856 28316
rect 7856 28260 7912 28316
rect 7912 28260 7916 28316
rect 7852 28256 7916 28260
rect 12612 28316 12676 28320
rect 12612 28260 12616 28316
rect 12616 28260 12672 28316
rect 12672 28260 12676 28316
rect 12612 28256 12676 28260
rect 12692 28316 12756 28320
rect 12692 28260 12696 28316
rect 12696 28260 12752 28316
rect 12752 28260 12756 28316
rect 12692 28256 12756 28260
rect 12772 28316 12836 28320
rect 12772 28260 12776 28316
rect 12776 28260 12832 28316
rect 12832 28260 12836 28316
rect 12772 28256 12836 28260
rect 12852 28316 12916 28320
rect 12852 28260 12856 28316
rect 12856 28260 12912 28316
rect 12912 28260 12916 28316
rect 12852 28256 12916 28260
rect 17612 28316 17676 28320
rect 17612 28260 17616 28316
rect 17616 28260 17672 28316
rect 17672 28260 17676 28316
rect 17612 28256 17676 28260
rect 17692 28316 17756 28320
rect 17692 28260 17696 28316
rect 17696 28260 17752 28316
rect 17752 28260 17756 28316
rect 17692 28256 17756 28260
rect 17772 28316 17836 28320
rect 17772 28260 17776 28316
rect 17776 28260 17832 28316
rect 17832 28260 17836 28316
rect 17772 28256 17836 28260
rect 17852 28316 17916 28320
rect 17852 28260 17856 28316
rect 17856 28260 17912 28316
rect 17912 28260 17916 28316
rect 17852 28256 17916 28260
rect 1952 27772 2016 27776
rect 1952 27716 1956 27772
rect 1956 27716 2012 27772
rect 2012 27716 2016 27772
rect 1952 27712 2016 27716
rect 2032 27772 2096 27776
rect 2032 27716 2036 27772
rect 2036 27716 2092 27772
rect 2092 27716 2096 27772
rect 2032 27712 2096 27716
rect 2112 27772 2176 27776
rect 2112 27716 2116 27772
rect 2116 27716 2172 27772
rect 2172 27716 2176 27772
rect 2112 27712 2176 27716
rect 2192 27772 2256 27776
rect 2192 27716 2196 27772
rect 2196 27716 2252 27772
rect 2252 27716 2256 27772
rect 2192 27712 2256 27716
rect 6952 27772 7016 27776
rect 6952 27716 6956 27772
rect 6956 27716 7012 27772
rect 7012 27716 7016 27772
rect 6952 27712 7016 27716
rect 7032 27772 7096 27776
rect 7032 27716 7036 27772
rect 7036 27716 7092 27772
rect 7092 27716 7096 27772
rect 7032 27712 7096 27716
rect 7112 27772 7176 27776
rect 7112 27716 7116 27772
rect 7116 27716 7172 27772
rect 7172 27716 7176 27772
rect 7112 27712 7176 27716
rect 7192 27772 7256 27776
rect 7192 27716 7196 27772
rect 7196 27716 7252 27772
rect 7252 27716 7256 27772
rect 7192 27712 7256 27716
rect 11952 27772 12016 27776
rect 11952 27716 11956 27772
rect 11956 27716 12012 27772
rect 12012 27716 12016 27772
rect 11952 27712 12016 27716
rect 12032 27772 12096 27776
rect 12032 27716 12036 27772
rect 12036 27716 12092 27772
rect 12092 27716 12096 27772
rect 12032 27712 12096 27716
rect 12112 27772 12176 27776
rect 12112 27716 12116 27772
rect 12116 27716 12172 27772
rect 12172 27716 12176 27772
rect 12112 27712 12176 27716
rect 12192 27772 12256 27776
rect 12192 27716 12196 27772
rect 12196 27716 12252 27772
rect 12252 27716 12256 27772
rect 12192 27712 12256 27716
rect 16952 27772 17016 27776
rect 16952 27716 16956 27772
rect 16956 27716 17012 27772
rect 17012 27716 17016 27772
rect 16952 27712 17016 27716
rect 17032 27772 17096 27776
rect 17032 27716 17036 27772
rect 17036 27716 17092 27772
rect 17092 27716 17096 27772
rect 17032 27712 17096 27716
rect 17112 27772 17176 27776
rect 17112 27716 17116 27772
rect 17116 27716 17172 27772
rect 17172 27716 17176 27772
rect 17112 27712 17176 27716
rect 17192 27772 17256 27776
rect 17192 27716 17196 27772
rect 17196 27716 17252 27772
rect 17252 27716 17256 27772
rect 17192 27712 17256 27716
rect 2612 27228 2676 27232
rect 2612 27172 2616 27228
rect 2616 27172 2672 27228
rect 2672 27172 2676 27228
rect 2612 27168 2676 27172
rect 2692 27228 2756 27232
rect 2692 27172 2696 27228
rect 2696 27172 2752 27228
rect 2752 27172 2756 27228
rect 2692 27168 2756 27172
rect 2772 27228 2836 27232
rect 2772 27172 2776 27228
rect 2776 27172 2832 27228
rect 2832 27172 2836 27228
rect 2772 27168 2836 27172
rect 2852 27228 2916 27232
rect 2852 27172 2856 27228
rect 2856 27172 2912 27228
rect 2912 27172 2916 27228
rect 2852 27168 2916 27172
rect 7612 27228 7676 27232
rect 7612 27172 7616 27228
rect 7616 27172 7672 27228
rect 7672 27172 7676 27228
rect 7612 27168 7676 27172
rect 7692 27228 7756 27232
rect 7692 27172 7696 27228
rect 7696 27172 7752 27228
rect 7752 27172 7756 27228
rect 7692 27168 7756 27172
rect 7772 27228 7836 27232
rect 7772 27172 7776 27228
rect 7776 27172 7832 27228
rect 7832 27172 7836 27228
rect 7772 27168 7836 27172
rect 7852 27228 7916 27232
rect 7852 27172 7856 27228
rect 7856 27172 7912 27228
rect 7912 27172 7916 27228
rect 7852 27168 7916 27172
rect 12612 27228 12676 27232
rect 12612 27172 12616 27228
rect 12616 27172 12672 27228
rect 12672 27172 12676 27228
rect 12612 27168 12676 27172
rect 12692 27228 12756 27232
rect 12692 27172 12696 27228
rect 12696 27172 12752 27228
rect 12752 27172 12756 27228
rect 12692 27168 12756 27172
rect 12772 27228 12836 27232
rect 12772 27172 12776 27228
rect 12776 27172 12832 27228
rect 12832 27172 12836 27228
rect 12772 27168 12836 27172
rect 12852 27228 12916 27232
rect 12852 27172 12856 27228
rect 12856 27172 12912 27228
rect 12912 27172 12916 27228
rect 12852 27168 12916 27172
rect 17612 27228 17676 27232
rect 17612 27172 17616 27228
rect 17616 27172 17672 27228
rect 17672 27172 17676 27228
rect 17612 27168 17676 27172
rect 17692 27228 17756 27232
rect 17692 27172 17696 27228
rect 17696 27172 17752 27228
rect 17752 27172 17756 27228
rect 17692 27168 17756 27172
rect 17772 27228 17836 27232
rect 17772 27172 17776 27228
rect 17776 27172 17832 27228
rect 17832 27172 17836 27228
rect 17772 27168 17836 27172
rect 17852 27228 17916 27232
rect 17852 27172 17856 27228
rect 17856 27172 17912 27228
rect 17912 27172 17916 27228
rect 17852 27168 17916 27172
rect 9444 26964 9508 27028
rect 9260 26828 9324 26892
rect 1952 26684 2016 26688
rect 1952 26628 1956 26684
rect 1956 26628 2012 26684
rect 2012 26628 2016 26684
rect 1952 26624 2016 26628
rect 2032 26684 2096 26688
rect 2032 26628 2036 26684
rect 2036 26628 2092 26684
rect 2092 26628 2096 26684
rect 2032 26624 2096 26628
rect 2112 26684 2176 26688
rect 2112 26628 2116 26684
rect 2116 26628 2172 26684
rect 2172 26628 2176 26684
rect 2112 26624 2176 26628
rect 2192 26684 2256 26688
rect 2192 26628 2196 26684
rect 2196 26628 2252 26684
rect 2252 26628 2256 26684
rect 2192 26624 2256 26628
rect 6952 26684 7016 26688
rect 6952 26628 6956 26684
rect 6956 26628 7012 26684
rect 7012 26628 7016 26684
rect 6952 26624 7016 26628
rect 7032 26684 7096 26688
rect 7032 26628 7036 26684
rect 7036 26628 7092 26684
rect 7092 26628 7096 26684
rect 7032 26624 7096 26628
rect 7112 26684 7176 26688
rect 7112 26628 7116 26684
rect 7116 26628 7172 26684
rect 7172 26628 7176 26684
rect 7112 26624 7176 26628
rect 7192 26684 7256 26688
rect 7192 26628 7196 26684
rect 7196 26628 7252 26684
rect 7252 26628 7256 26684
rect 7192 26624 7256 26628
rect 11952 26684 12016 26688
rect 11952 26628 11956 26684
rect 11956 26628 12012 26684
rect 12012 26628 12016 26684
rect 11952 26624 12016 26628
rect 12032 26684 12096 26688
rect 12032 26628 12036 26684
rect 12036 26628 12092 26684
rect 12092 26628 12096 26684
rect 12032 26624 12096 26628
rect 12112 26684 12176 26688
rect 12112 26628 12116 26684
rect 12116 26628 12172 26684
rect 12172 26628 12176 26684
rect 12112 26624 12176 26628
rect 12192 26684 12256 26688
rect 12192 26628 12196 26684
rect 12196 26628 12252 26684
rect 12252 26628 12256 26684
rect 12192 26624 12256 26628
rect 16952 26684 17016 26688
rect 16952 26628 16956 26684
rect 16956 26628 17012 26684
rect 17012 26628 17016 26684
rect 16952 26624 17016 26628
rect 17032 26684 17096 26688
rect 17032 26628 17036 26684
rect 17036 26628 17092 26684
rect 17092 26628 17096 26684
rect 17032 26624 17096 26628
rect 17112 26684 17176 26688
rect 17112 26628 17116 26684
rect 17116 26628 17172 26684
rect 17172 26628 17176 26684
rect 17112 26624 17176 26628
rect 17192 26684 17256 26688
rect 17192 26628 17196 26684
rect 17196 26628 17252 26684
rect 17252 26628 17256 26684
rect 17192 26624 17256 26628
rect 2612 26140 2676 26144
rect 2612 26084 2616 26140
rect 2616 26084 2672 26140
rect 2672 26084 2676 26140
rect 2612 26080 2676 26084
rect 2692 26140 2756 26144
rect 2692 26084 2696 26140
rect 2696 26084 2752 26140
rect 2752 26084 2756 26140
rect 2692 26080 2756 26084
rect 2772 26140 2836 26144
rect 2772 26084 2776 26140
rect 2776 26084 2832 26140
rect 2832 26084 2836 26140
rect 2772 26080 2836 26084
rect 2852 26140 2916 26144
rect 2852 26084 2856 26140
rect 2856 26084 2912 26140
rect 2912 26084 2916 26140
rect 2852 26080 2916 26084
rect 7612 26140 7676 26144
rect 7612 26084 7616 26140
rect 7616 26084 7672 26140
rect 7672 26084 7676 26140
rect 7612 26080 7676 26084
rect 7692 26140 7756 26144
rect 7692 26084 7696 26140
rect 7696 26084 7752 26140
rect 7752 26084 7756 26140
rect 7692 26080 7756 26084
rect 7772 26140 7836 26144
rect 7772 26084 7776 26140
rect 7776 26084 7832 26140
rect 7832 26084 7836 26140
rect 7772 26080 7836 26084
rect 7852 26140 7916 26144
rect 7852 26084 7856 26140
rect 7856 26084 7912 26140
rect 7912 26084 7916 26140
rect 7852 26080 7916 26084
rect 11284 26148 11348 26212
rect 12612 26140 12676 26144
rect 12612 26084 12616 26140
rect 12616 26084 12672 26140
rect 12672 26084 12676 26140
rect 12612 26080 12676 26084
rect 12692 26140 12756 26144
rect 12692 26084 12696 26140
rect 12696 26084 12752 26140
rect 12752 26084 12756 26140
rect 12692 26080 12756 26084
rect 12772 26140 12836 26144
rect 12772 26084 12776 26140
rect 12776 26084 12832 26140
rect 12832 26084 12836 26140
rect 12772 26080 12836 26084
rect 12852 26140 12916 26144
rect 12852 26084 12856 26140
rect 12856 26084 12912 26140
rect 12912 26084 12916 26140
rect 12852 26080 12916 26084
rect 17612 26140 17676 26144
rect 17612 26084 17616 26140
rect 17616 26084 17672 26140
rect 17672 26084 17676 26140
rect 17612 26080 17676 26084
rect 17692 26140 17756 26144
rect 17692 26084 17696 26140
rect 17696 26084 17752 26140
rect 17752 26084 17756 26140
rect 17692 26080 17756 26084
rect 17772 26140 17836 26144
rect 17772 26084 17776 26140
rect 17776 26084 17832 26140
rect 17832 26084 17836 26140
rect 17772 26080 17836 26084
rect 17852 26140 17916 26144
rect 17852 26084 17856 26140
rect 17856 26084 17912 26140
rect 17912 26084 17916 26140
rect 17852 26080 17916 26084
rect 8340 26072 8404 26076
rect 8340 26016 8354 26072
rect 8354 26016 8404 26072
rect 8340 26012 8404 26016
rect 10180 26072 10244 26076
rect 10180 26016 10194 26072
rect 10194 26016 10244 26072
rect 10180 26012 10244 26016
rect 11652 26012 11716 26076
rect 1952 25596 2016 25600
rect 1952 25540 1956 25596
rect 1956 25540 2012 25596
rect 2012 25540 2016 25596
rect 1952 25536 2016 25540
rect 2032 25596 2096 25600
rect 2032 25540 2036 25596
rect 2036 25540 2092 25596
rect 2092 25540 2096 25596
rect 2032 25536 2096 25540
rect 2112 25596 2176 25600
rect 2112 25540 2116 25596
rect 2116 25540 2172 25596
rect 2172 25540 2176 25596
rect 2112 25536 2176 25540
rect 2192 25596 2256 25600
rect 2192 25540 2196 25596
rect 2196 25540 2252 25596
rect 2252 25540 2256 25596
rect 2192 25536 2256 25540
rect 6952 25596 7016 25600
rect 6952 25540 6956 25596
rect 6956 25540 7012 25596
rect 7012 25540 7016 25596
rect 6952 25536 7016 25540
rect 7032 25596 7096 25600
rect 7032 25540 7036 25596
rect 7036 25540 7092 25596
rect 7092 25540 7096 25596
rect 7032 25536 7096 25540
rect 7112 25596 7176 25600
rect 7112 25540 7116 25596
rect 7116 25540 7172 25596
rect 7172 25540 7176 25596
rect 7112 25536 7176 25540
rect 7192 25596 7256 25600
rect 7192 25540 7196 25596
rect 7196 25540 7252 25596
rect 7252 25540 7256 25596
rect 7192 25536 7256 25540
rect 11952 25596 12016 25600
rect 11952 25540 11956 25596
rect 11956 25540 12012 25596
rect 12012 25540 12016 25596
rect 11952 25536 12016 25540
rect 12032 25596 12096 25600
rect 12032 25540 12036 25596
rect 12036 25540 12092 25596
rect 12092 25540 12096 25596
rect 12032 25536 12096 25540
rect 12112 25596 12176 25600
rect 12112 25540 12116 25596
rect 12116 25540 12172 25596
rect 12172 25540 12176 25596
rect 12112 25536 12176 25540
rect 12192 25596 12256 25600
rect 12192 25540 12196 25596
rect 12196 25540 12252 25596
rect 12252 25540 12256 25596
rect 12192 25536 12256 25540
rect 16952 25596 17016 25600
rect 16952 25540 16956 25596
rect 16956 25540 17012 25596
rect 17012 25540 17016 25596
rect 16952 25536 17016 25540
rect 17032 25596 17096 25600
rect 17032 25540 17036 25596
rect 17036 25540 17092 25596
rect 17092 25540 17096 25596
rect 17032 25536 17096 25540
rect 17112 25596 17176 25600
rect 17112 25540 17116 25596
rect 17116 25540 17172 25596
rect 17172 25540 17176 25596
rect 17112 25536 17176 25540
rect 17192 25596 17256 25600
rect 17192 25540 17196 25596
rect 17196 25540 17252 25596
rect 17252 25540 17256 25596
rect 17192 25536 17256 25540
rect 10364 25392 10428 25396
rect 10364 25336 10378 25392
rect 10378 25336 10428 25392
rect 10364 25332 10428 25336
rect 2612 25052 2676 25056
rect 2612 24996 2616 25052
rect 2616 24996 2672 25052
rect 2672 24996 2676 25052
rect 2612 24992 2676 24996
rect 2692 25052 2756 25056
rect 2692 24996 2696 25052
rect 2696 24996 2752 25052
rect 2752 24996 2756 25052
rect 2692 24992 2756 24996
rect 2772 25052 2836 25056
rect 2772 24996 2776 25052
rect 2776 24996 2832 25052
rect 2832 24996 2836 25052
rect 2772 24992 2836 24996
rect 2852 25052 2916 25056
rect 2852 24996 2856 25052
rect 2856 24996 2912 25052
rect 2912 24996 2916 25052
rect 2852 24992 2916 24996
rect 7612 25052 7676 25056
rect 7612 24996 7616 25052
rect 7616 24996 7672 25052
rect 7672 24996 7676 25052
rect 7612 24992 7676 24996
rect 7692 25052 7756 25056
rect 7692 24996 7696 25052
rect 7696 24996 7752 25052
rect 7752 24996 7756 25052
rect 7692 24992 7756 24996
rect 7772 25052 7836 25056
rect 7772 24996 7776 25052
rect 7776 24996 7832 25052
rect 7832 24996 7836 25052
rect 7772 24992 7836 24996
rect 7852 25052 7916 25056
rect 7852 24996 7856 25052
rect 7856 24996 7912 25052
rect 7912 24996 7916 25052
rect 7852 24992 7916 24996
rect 12612 25052 12676 25056
rect 12612 24996 12616 25052
rect 12616 24996 12672 25052
rect 12672 24996 12676 25052
rect 12612 24992 12676 24996
rect 12692 25052 12756 25056
rect 12692 24996 12696 25052
rect 12696 24996 12752 25052
rect 12752 24996 12756 25052
rect 12692 24992 12756 24996
rect 12772 25052 12836 25056
rect 12772 24996 12776 25052
rect 12776 24996 12832 25052
rect 12832 24996 12836 25052
rect 12772 24992 12836 24996
rect 12852 25052 12916 25056
rect 12852 24996 12856 25052
rect 12856 24996 12912 25052
rect 12912 24996 12916 25052
rect 12852 24992 12916 24996
rect 17612 25052 17676 25056
rect 17612 24996 17616 25052
rect 17616 24996 17672 25052
rect 17672 24996 17676 25052
rect 17612 24992 17676 24996
rect 17692 25052 17756 25056
rect 17692 24996 17696 25052
rect 17696 24996 17752 25052
rect 17752 24996 17756 25052
rect 17692 24992 17756 24996
rect 17772 25052 17836 25056
rect 17772 24996 17776 25052
rect 17776 24996 17832 25052
rect 17832 24996 17836 25052
rect 17772 24992 17836 24996
rect 17852 25052 17916 25056
rect 17852 24996 17856 25052
rect 17856 24996 17912 25052
rect 17912 24996 17916 25052
rect 17852 24992 17916 24996
rect 1716 24788 1780 24852
rect 13308 24788 13372 24852
rect 13124 24652 13188 24716
rect 1952 24508 2016 24512
rect 1952 24452 1956 24508
rect 1956 24452 2012 24508
rect 2012 24452 2016 24508
rect 1952 24448 2016 24452
rect 2032 24508 2096 24512
rect 2032 24452 2036 24508
rect 2036 24452 2092 24508
rect 2092 24452 2096 24508
rect 2032 24448 2096 24452
rect 2112 24508 2176 24512
rect 2112 24452 2116 24508
rect 2116 24452 2172 24508
rect 2172 24452 2176 24508
rect 2112 24448 2176 24452
rect 2192 24508 2256 24512
rect 2192 24452 2196 24508
rect 2196 24452 2252 24508
rect 2252 24452 2256 24508
rect 2192 24448 2256 24452
rect 6952 24508 7016 24512
rect 6952 24452 6956 24508
rect 6956 24452 7012 24508
rect 7012 24452 7016 24508
rect 6952 24448 7016 24452
rect 7032 24508 7096 24512
rect 7032 24452 7036 24508
rect 7036 24452 7092 24508
rect 7092 24452 7096 24508
rect 7032 24448 7096 24452
rect 7112 24508 7176 24512
rect 7112 24452 7116 24508
rect 7116 24452 7172 24508
rect 7172 24452 7176 24508
rect 7112 24448 7176 24452
rect 7192 24508 7256 24512
rect 7192 24452 7196 24508
rect 7196 24452 7252 24508
rect 7252 24452 7256 24508
rect 7192 24448 7256 24452
rect 11952 24508 12016 24512
rect 11952 24452 11956 24508
rect 11956 24452 12012 24508
rect 12012 24452 12016 24508
rect 11952 24448 12016 24452
rect 12032 24508 12096 24512
rect 12032 24452 12036 24508
rect 12036 24452 12092 24508
rect 12092 24452 12096 24508
rect 12032 24448 12096 24452
rect 12112 24508 12176 24512
rect 12112 24452 12116 24508
rect 12116 24452 12172 24508
rect 12172 24452 12176 24508
rect 12112 24448 12176 24452
rect 12192 24508 12256 24512
rect 12192 24452 12196 24508
rect 12196 24452 12252 24508
rect 12252 24452 12256 24508
rect 12192 24448 12256 24452
rect 16952 24508 17016 24512
rect 16952 24452 16956 24508
rect 16956 24452 17012 24508
rect 17012 24452 17016 24508
rect 16952 24448 17016 24452
rect 17032 24508 17096 24512
rect 17032 24452 17036 24508
rect 17036 24452 17092 24508
rect 17092 24452 17096 24508
rect 17032 24448 17096 24452
rect 17112 24508 17176 24512
rect 17112 24452 17116 24508
rect 17116 24452 17172 24508
rect 17172 24452 17176 24508
rect 17112 24448 17176 24452
rect 17192 24508 17256 24512
rect 17192 24452 17196 24508
rect 17196 24452 17252 24508
rect 17252 24452 17256 24508
rect 17192 24448 17256 24452
rect 2612 23964 2676 23968
rect 2612 23908 2616 23964
rect 2616 23908 2672 23964
rect 2672 23908 2676 23964
rect 2612 23904 2676 23908
rect 2692 23964 2756 23968
rect 2692 23908 2696 23964
rect 2696 23908 2752 23964
rect 2752 23908 2756 23964
rect 2692 23904 2756 23908
rect 2772 23964 2836 23968
rect 2772 23908 2776 23964
rect 2776 23908 2832 23964
rect 2832 23908 2836 23964
rect 2772 23904 2836 23908
rect 2852 23964 2916 23968
rect 2852 23908 2856 23964
rect 2856 23908 2912 23964
rect 2912 23908 2916 23964
rect 2852 23904 2916 23908
rect 7612 23964 7676 23968
rect 7612 23908 7616 23964
rect 7616 23908 7672 23964
rect 7672 23908 7676 23964
rect 7612 23904 7676 23908
rect 7692 23964 7756 23968
rect 7692 23908 7696 23964
rect 7696 23908 7752 23964
rect 7752 23908 7756 23964
rect 7692 23904 7756 23908
rect 7772 23964 7836 23968
rect 7772 23908 7776 23964
rect 7776 23908 7832 23964
rect 7832 23908 7836 23964
rect 7772 23904 7836 23908
rect 7852 23964 7916 23968
rect 7852 23908 7856 23964
rect 7856 23908 7912 23964
rect 7912 23908 7916 23964
rect 7852 23904 7916 23908
rect 12612 23964 12676 23968
rect 12612 23908 12616 23964
rect 12616 23908 12672 23964
rect 12672 23908 12676 23964
rect 12612 23904 12676 23908
rect 12692 23964 12756 23968
rect 12692 23908 12696 23964
rect 12696 23908 12752 23964
rect 12752 23908 12756 23964
rect 12692 23904 12756 23908
rect 12772 23964 12836 23968
rect 12772 23908 12776 23964
rect 12776 23908 12832 23964
rect 12832 23908 12836 23964
rect 12772 23904 12836 23908
rect 12852 23964 12916 23968
rect 12852 23908 12856 23964
rect 12856 23908 12912 23964
rect 12912 23908 12916 23964
rect 12852 23904 12916 23908
rect 17612 23964 17676 23968
rect 17612 23908 17616 23964
rect 17616 23908 17672 23964
rect 17672 23908 17676 23964
rect 17612 23904 17676 23908
rect 17692 23964 17756 23968
rect 17692 23908 17696 23964
rect 17696 23908 17752 23964
rect 17752 23908 17756 23964
rect 17692 23904 17756 23908
rect 17772 23964 17836 23968
rect 17772 23908 17776 23964
rect 17776 23908 17832 23964
rect 17832 23908 17836 23964
rect 17772 23904 17836 23908
rect 17852 23964 17916 23968
rect 17852 23908 17856 23964
rect 17856 23908 17912 23964
rect 17912 23908 17916 23964
rect 17852 23904 17916 23908
rect 4292 23564 4356 23628
rect 1952 23420 2016 23424
rect 1952 23364 1956 23420
rect 1956 23364 2012 23420
rect 2012 23364 2016 23420
rect 1952 23360 2016 23364
rect 2032 23420 2096 23424
rect 2032 23364 2036 23420
rect 2036 23364 2092 23420
rect 2092 23364 2096 23420
rect 2032 23360 2096 23364
rect 2112 23420 2176 23424
rect 2112 23364 2116 23420
rect 2116 23364 2172 23420
rect 2172 23364 2176 23420
rect 2112 23360 2176 23364
rect 2192 23420 2256 23424
rect 2192 23364 2196 23420
rect 2196 23364 2252 23420
rect 2252 23364 2256 23420
rect 2192 23360 2256 23364
rect 6952 23420 7016 23424
rect 6952 23364 6956 23420
rect 6956 23364 7012 23420
rect 7012 23364 7016 23420
rect 6952 23360 7016 23364
rect 7032 23420 7096 23424
rect 7032 23364 7036 23420
rect 7036 23364 7092 23420
rect 7092 23364 7096 23420
rect 7032 23360 7096 23364
rect 7112 23420 7176 23424
rect 7112 23364 7116 23420
rect 7116 23364 7172 23420
rect 7172 23364 7176 23420
rect 7112 23360 7176 23364
rect 7192 23420 7256 23424
rect 7192 23364 7196 23420
rect 7196 23364 7252 23420
rect 7252 23364 7256 23420
rect 7192 23360 7256 23364
rect 11952 23420 12016 23424
rect 11952 23364 11956 23420
rect 11956 23364 12012 23420
rect 12012 23364 12016 23420
rect 11952 23360 12016 23364
rect 12032 23420 12096 23424
rect 12032 23364 12036 23420
rect 12036 23364 12092 23420
rect 12092 23364 12096 23420
rect 12032 23360 12096 23364
rect 12112 23420 12176 23424
rect 12112 23364 12116 23420
rect 12116 23364 12172 23420
rect 12172 23364 12176 23420
rect 12112 23360 12176 23364
rect 12192 23420 12256 23424
rect 12192 23364 12196 23420
rect 12196 23364 12252 23420
rect 12252 23364 12256 23420
rect 12192 23360 12256 23364
rect 16952 23420 17016 23424
rect 16952 23364 16956 23420
rect 16956 23364 17012 23420
rect 17012 23364 17016 23420
rect 16952 23360 17016 23364
rect 17032 23420 17096 23424
rect 17032 23364 17036 23420
rect 17036 23364 17092 23420
rect 17092 23364 17096 23420
rect 17032 23360 17096 23364
rect 17112 23420 17176 23424
rect 17112 23364 17116 23420
rect 17116 23364 17172 23420
rect 17172 23364 17176 23420
rect 17112 23360 17176 23364
rect 17192 23420 17256 23424
rect 17192 23364 17196 23420
rect 17196 23364 17252 23420
rect 17252 23364 17256 23420
rect 17192 23360 17256 23364
rect 2612 22876 2676 22880
rect 2612 22820 2616 22876
rect 2616 22820 2672 22876
rect 2672 22820 2676 22876
rect 2612 22816 2676 22820
rect 2692 22876 2756 22880
rect 2692 22820 2696 22876
rect 2696 22820 2752 22876
rect 2752 22820 2756 22876
rect 2692 22816 2756 22820
rect 2772 22876 2836 22880
rect 2772 22820 2776 22876
rect 2776 22820 2832 22876
rect 2832 22820 2836 22876
rect 2772 22816 2836 22820
rect 2852 22876 2916 22880
rect 2852 22820 2856 22876
rect 2856 22820 2912 22876
rect 2912 22820 2916 22876
rect 2852 22816 2916 22820
rect 7612 22876 7676 22880
rect 7612 22820 7616 22876
rect 7616 22820 7672 22876
rect 7672 22820 7676 22876
rect 7612 22816 7676 22820
rect 7692 22876 7756 22880
rect 7692 22820 7696 22876
rect 7696 22820 7752 22876
rect 7752 22820 7756 22876
rect 7692 22816 7756 22820
rect 7772 22876 7836 22880
rect 7772 22820 7776 22876
rect 7776 22820 7832 22876
rect 7832 22820 7836 22876
rect 7772 22816 7836 22820
rect 7852 22876 7916 22880
rect 7852 22820 7856 22876
rect 7856 22820 7912 22876
rect 7912 22820 7916 22876
rect 7852 22816 7916 22820
rect 12612 22876 12676 22880
rect 12612 22820 12616 22876
rect 12616 22820 12672 22876
rect 12672 22820 12676 22876
rect 12612 22816 12676 22820
rect 12692 22876 12756 22880
rect 12692 22820 12696 22876
rect 12696 22820 12752 22876
rect 12752 22820 12756 22876
rect 12692 22816 12756 22820
rect 12772 22876 12836 22880
rect 12772 22820 12776 22876
rect 12776 22820 12832 22876
rect 12832 22820 12836 22876
rect 12772 22816 12836 22820
rect 12852 22876 12916 22880
rect 12852 22820 12856 22876
rect 12856 22820 12912 22876
rect 12912 22820 12916 22876
rect 12852 22816 12916 22820
rect 17612 22876 17676 22880
rect 17612 22820 17616 22876
rect 17616 22820 17672 22876
rect 17672 22820 17676 22876
rect 17612 22816 17676 22820
rect 17692 22876 17756 22880
rect 17692 22820 17696 22876
rect 17696 22820 17752 22876
rect 17752 22820 17756 22876
rect 17692 22816 17756 22820
rect 17772 22876 17836 22880
rect 17772 22820 17776 22876
rect 17776 22820 17832 22876
rect 17832 22820 17836 22876
rect 17772 22816 17836 22820
rect 17852 22876 17916 22880
rect 17852 22820 17856 22876
rect 17856 22820 17912 22876
rect 17912 22820 17916 22876
rect 17852 22816 17916 22820
rect 14412 22476 14476 22540
rect 1952 22332 2016 22336
rect 1952 22276 1956 22332
rect 1956 22276 2012 22332
rect 2012 22276 2016 22332
rect 1952 22272 2016 22276
rect 2032 22332 2096 22336
rect 2032 22276 2036 22332
rect 2036 22276 2092 22332
rect 2092 22276 2096 22332
rect 2032 22272 2096 22276
rect 2112 22332 2176 22336
rect 2112 22276 2116 22332
rect 2116 22276 2172 22332
rect 2172 22276 2176 22332
rect 2112 22272 2176 22276
rect 2192 22332 2256 22336
rect 2192 22276 2196 22332
rect 2196 22276 2252 22332
rect 2252 22276 2256 22332
rect 2192 22272 2256 22276
rect 6952 22332 7016 22336
rect 6952 22276 6956 22332
rect 6956 22276 7012 22332
rect 7012 22276 7016 22332
rect 6952 22272 7016 22276
rect 7032 22332 7096 22336
rect 7032 22276 7036 22332
rect 7036 22276 7092 22332
rect 7092 22276 7096 22332
rect 7032 22272 7096 22276
rect 7112 22332 7176 22336
rect 7112 22276 7116 22332
rect 7116 22276 7172 22332
rect 7172 22276 7176 22332
rect 7112 22272 7176 22276
rect 7192 22332 7256 22336
rect 7192 22276 7196 22332
rect 7196 22276 7252 22332
rect 7252 22276 7256 22332
rect 7192 22272 7256 22276
rect 11952 22332 12016 22336
rect 11952 22276 11956 22332
rect 11956 22276 12012 22332
rect 12012 22276 12016 22332
rect 11952 22272 12016 22276
rect 12032 22332 12096 22336
rect 12032 22276 12036 22332
rect 12036 22276 12092 22332
rect 12092 22276 12096 22332
rect 12032 22272 12096 22276
rect 12112 22332 12176 22336
rect 12112 22276 12116 22332
rect 12116 22276 12172 22332
rect 12172 22276 12176 22332
rect 12112 22272 12176 22276
rect 12192 22332 12256 22336
rect 12192 22276 12196 22332
rect 12196 22276 12252 22332
rect 12252 22276 12256 22332
rect 12192 22272 12256 22276
rect 16952 22332 17016 22336
rect 16952 22276 16956 22332
rect 16956 22276 17012 22332
rect 17012 22276 17016 22332
rect 16952 22272 17016 22276
rect 17032 22332 17096 22336
rect 17032 22276 17036 22332
rect 17036 22276 17092 22332
rect 17092 22276 17096 22332
rect 17032 22272 17096 22276
rect 17112 22332 17176 22336
rect 17112 22276 17116 22332
rect 17116 22276 17172 22332
rect 17172 22276 17176 22332
rect 17112 22272 17176 22276
rect 17192 22332 17256 22336
rect 17192 22276 17196 22332
rect 17196 22276 17252 22332
rect 17252 22276 17256 22332
rect 17192 22272 17256 22276
rect 4476 21932 4540 21996
rect 2612 21788 2676 21792
rect 2612 21732 2616 21788
rect 2616 21732 2672 21788
rect 2672 21732 2676 21788
rect 2612 21728 2676 21732
rect 2692 21788 2756 21792
rect 2692 21732 2696 21788
rect 2696 21732 2752 21788
rect 2752 21732 2756 21788
rect 2692 21728 2756 21732
rect 2772 21788 2836 21792
rect 2772 21732 2776 21788
rect 2776 21732 2832 21788
rect 2832 21732 2836 21788
rect 2772 21728 2836 21732
rect 2852 21788 2916 21792
rect 2852 21732 2856 21788
rect 2856 21732 2912 21788
rect 2912 21732 2916 21788
rect 2852 21728 2916 21732
rect 7612 21788 7676 21792
rect 7612 21732 7616 21788
rect 7616 21732 7672 21788
rect 7672 21732 7676 21788
rect 7612 21728 7676 21732
rect 7692 21788 7756 21792
rect 7692 21732 7696 21788
rect 7696 21732 7752 21788
rect 7752 21732 7756 21788
rect 7692 21728 7756 21732
rect 7772 21788 7836 21792
rect 7772 21732 7776 21788
rect 7776 21732 7832 21788
rect 7832 21732 7836 21788
rect 7772 21728 7836 21732
rect 7852 21788 7916 21792
rect 7852 21732 7856 21788
rect 7856 21732 7912 21788
rect 7912 21732 7916 21788
rect 7852 21728 7916 21732
rect 12612 21788 12676 21792
rect 12612 21732 12616 21788
rect 12616 21732 12672 21788
rect 12672 21732 12676 21788
rect 12612 21728 12676 21732
rect 12692 21788 12756 21792
rect 12692 21732 12696 21788
rect 12696 21732 12752 21788
rect 12752 21732 12756 21788
rect 12692 21728 12756 21732
rect 12772 21788 12836 21792
rect 12772 21732 12776 21788
rect 12776 21732 12832 21788
rect 12832 21732 12836 21788
rect 12772 21728 12836 21732
rect 12852 21788 12916 21792
rect 12852 21732 12856 21788
rect 12856 21732 12912 21788
rect 12912 21732 12916 21788
rect 12852 21728 12916 21732
rect 17612 21788 17676 21792
rect 17612 21732 17616 21788
rect 17616 21732 17672 21788
rect 17672 21732 17676 21788
rect 17612 21728 17676 21732
rect 17692 21788 17756 21792
rect 17692 21732 17696 21788
rect 17696 21732 17752 21788
rect 17752 21732 17756 21788
rect 17692 21728 17756 21732
rect 17772 21788 17836 21792
rect 17772 21732 17776 21788
rect 17776 21732 17832 21788
rect 17832 21732 17836 21788
rect 17772 21728 17836 21732
rect 17852 21788 17916 21792
rect 17852 21732 17856 21788
rect 17856 21732 17912 21788
rect 17912 21732 17916 21788
rect 17852 21728 17916 21732
rect 1952 21244 2016 21248
rect 1952 21188 1956 21244
rect 1956 21188 2012 21244
rect 2012 21188 2016 21244
rect 1952 21184 2016 21188
rect 2032 21244 2096 21248
rect 2032 21188 2036 21244
rect 2036 21188 2092 21244
rect 2092 21188 2096 21244
rect 2032 21184 2096 21188
rect 2112 21244 2176 21248
rect 2112 21188 2116 21244
rect 2116 21188 2172 21244
rect 2172 21188 2176 21244
rect 2112 21184 2176 21188
rect 2192 21244 2256 21248
rect 2192 21188 2196 21244
rect 2196 21188 2252 21244
rect 2252 21188 2256 21244
rect 2192 21184 2256 21188
rect 6952 21244 7016 21248
rect 6952 21188 6956 21244
rect 6956 21188 7012 21244
rect 7012 21188 7016 21244
rect 6952 21184 7016 21188
rect 7032 21244 7096 21248
rect 7032 21188 7036 21244
rect 7036 21188 7092 21244
rect 7092 21188 7096 21244
rect 7032 21184 7096 21188
rect 7112 21244 7176 21248
rect 7112 21188 7116 21244
rect 7116 21188 7172 21244
rect 7172 21188 7176 21244
rect 7112 21184 7176 21188
rect 7192 21244 7256 21248
rect 7192 21188 7196 21244
rect 7196 21188 7252 21244
rect 7252 21188 7256 21244
rect 7192 21184 7256 21188
rect 11952 21244 12016 21248
rect 11952 21188 11956 21244
rect 11956 21188 12012 21244
rect 12012 21188 12016 21244
rect 11952 21184 12016 21188
rect 12032 21244 12096 21248
rect 12032 21188 12036 21244
rect 12036 21188 12092 21244
rect 12092 21188 12096 21244
rect 12032 21184 12096 21188
rect 12112 21244 12176 21248
rect 12112 21188 12116 21244
rect 12116 21188 12172 21244
rect 12172 21188 12176 21244
rect 12112 21184 12176 21188
rect 12192 21244 12256 21248
rect 12192 21188 12196 21244
rect 12196 21188 12252 21244
rect 12252 21188 12256 21244
rect 12192 21184 12256 21188
rect 16952 21244 17016 21248
rect 16952 21188 16956 21244
rect 16956 21188 17012 21244
rect 17012 21188 17016 21244
rect 16952 21184 17016 21188
rect 17032 21244 17096 21248
rect 17032 21188 17036 21244
rect 17036 21188 17092 21244
rect 17092 21188 17096 21244
rect 17032 21184 17096 21188
rect 17112 21244 17176 21248
rect 17112 21188 17116 21244
rect 17116 21188 17172 21244
rect 17172 21188 17176 21244
rect 17112 21184 17176 21188
rect 17192 21244 17256 21248
rect 17192 21188 17196 21244
rect 17196 21188 17252 21244
rect 17252 21188 17256 21244
rect 17192 21184 17256 21188
rect 16436 20980 16500 21044
rect 4476 20708 4540 20772
rect 2612 20700 2676 20704
rect 2612 20644 2616 20700
rect 2616 20644 2672 20700
rect 2672 20644 2676 20700
rect 2612 20640 2676 20644
rect 2692 20700 2756 20704
rect 2692 20644 2696 20700
rect 2696 20644 2752 20700
rect 2752 20644 2756 20700
rect 2692 20640 2756 20644
rect 2772 20700 2836 20704
rect 2772 20644 2776 20700
rect 2776 20644 2832 20700
rect 2832 20644 2836 20700
rect 2772 20640 2836 20644
rect 2852 20700 2916 20704
rect 2852 20644 2856 20700
rect 2856 20644 2912 20700
rect 2912 20644 2916 20700
rect 2852 20640 2916 20644
rect 7612 20700 7676 20704
rect 7612 20644 7616 20700
rect 7616 20644 7672 20700
rect 7672 20644 7676 20700
rect 7612 20640 7676 20644
rect 7692 20700 7756 20704
rect 7692 20644 7696 20700
rect 7696 20644 7752 20700
rect 7752 20644 7756 20700
rect 7692 20640 7756 20644
rect 7772 20700 7836 20704
rect 7772 20644 7776 20700
rect 7776 20644 7832 20700
rect 7832 20644 7836 20700
rect 7772 20640 7836 20644
rect 7852 20700 7916 20704
rect 7852 20644 7856 20700
rect 7856 20644 7912 20700
rect 7912 20644 7916 20700
rect 7852 20640 7916 20644
rect 12612 20700 12676 20704
rect 12612 20644 12616 20700
rect 12616 20644 12672 20700
rect 12672 20644 12676 20700
rect 12612 20640 12676 20644
rect 12692 20700 12756 20704
rect 12692 20644 12696 20700
rect 12696 20644 12752 20700
rect 12752 20644 12756 20700
rect 12692 20640 12756 20644
rect 12772 20700 12836 20704
rect 12772 20644 12776 20700
rect 12776 20644 12832 20700
rect 12832 20644 12836 20700
rect 12772 20640 12836 20644
rect 12852 20700 12916 20704
rect 12852 20644 12856 20700
rect 12856 20644 12912 20700
rect 12912 20644 12916 20700
rect 12852 20640 12916 20644
rect 17612 20700 17676 20704
rect 17612 20644 17616 20700
rect 17616 20644 17672 20700
rect 17672 20644 17676 20700
rect 17612 20640 17676 20644
rect 17692 20700 17756 20704
rect 17692 20644 17696 20700
rect 17696 20644 17752 20700
rect 17752 20644 17756 20700
rect 17692 20640 17756 20644
rect 17772 20700 17836 20704
rect 17772 20644 17776 20700
rect 17776 20644 17832 20700
rect 17832 20644 17836 20700
rect 17772 20640 17836 20644
rect 17852 20700 17916 20704
rect 17852 20644 17856 20700
rect 17856 20644 17912 20700
rect 17912 20644 17916 20700
rect 17852 20640 17916 20644
rect 1952 20156 2016 20160
rect 1952 20100 1956 20156
rect 1956 20100 2012 20156
rect 2012 20100 2016 20156
rect 1952 20096 2016 20100
rect 2032 20156 2096 20160
rect 2032 20100 2036 20156
rect 2036 20100 2092 20156
rect 2092 20100 2096 20156
rect 2032 20096 2096 20100
rect 2112 20156 2176 20160
rect 2112 20100 2116 20156
rect 2116 20100 2172 20156
rect 2172 20100 2176 20156
rect 2112 20096 2176 20100
rect 2192 20156 2256 20160
rect 2192 20100 2196 20156
rect 2196 20100 2252 20156
rect 2252 20100 2256 20156
rect 2192 20096 2256 20100
rect 6952 20156 7016 20160
rect 6952 20100 6956 20156
rect 6956 20100 7012 20156
rect 7012 20100 7016 20156
rect 6952 20096 7016 20100
rect 7032 20156 7096 20160
rect 7032 20100 7036 20156
rect 7036 20100 7092 20156
rect 7092 20100 7096 20156
rect 7032 20096 7096 20100
rect 7112 20156 7176 20160
rect 7112 20100 7116 20156
rect 7116 20100 7172 20156
rect 7172 20100 7176 20156
rect 7112 20096 7176 20100
rect 7192 20156 7256 20160
rect 7192 20100 7196 20156
rect 7196 20100 7252 20156
rect 7252 20100 7256 20156
rect 7192 20096 7256 20100
rect 11952 20156 12016 20160
rect 11952 20100 11956 20156
rect 11956 20100 12012 20156
rect 12012 20100 12016 20156
rect 11952 20096 12016 20100
rect 12032 20156 12096 20160
rect 12032 20100 12036 20156
rect 12036 20100 12092 20156
rect 12092 20100 12096 20156
rect 12032 20096 12096 20100
rect 12112 20156 12176 20160
rect 12112 20100 12116 20156
rect 12116 20100 12172 20156
rect 12172 20100 12176 20156
rect 12112 20096 12176 20100
rect 12192 20156 12256 20160
rect 12192 20100 12196 20156
rect 12196 20100 12252 20156
rect 12252 20100 12256 20156
rect 12192 20096 12256 20100
rect 16952 20156 17016 20160
rect 16952 20100 16956 20156
rect 16956 20100 17012 20156
rect 17012 20100 17016 20156
rect 16952 20096 17016 20100
rect 17032 20156 17096 20160
rect 17032 20100 17036 20156
rect 17036 20100 17092 20156
rect 17092 20100 17096 20156
rect 17032 20096 17096 20100
rect 17112 20156 17176 20160
rect 17112 20100 17116 20156
rect 17116 20100 17172 20156
rect 17172 20100 17176 20156
rect 17112 20096 17176 20100
rect 17192 20156 17256 20160
rect 17192 20100 17196 20156
rect 17196 20100 17252 20156
rect 17252 20100 17256 20156
rect 17192 20096 17256 20100
rect 6500 19892 6564 19956
rect 2612 19612 2676 19616
rect 2612 19556 2616 19612
rect 2616 19556 2672 19612
rect 2672 19556 2676 19612
rect 2612 19552 2676 19556
rect 2692 19612 2756 19616
rect 2692 19556 2696 19612
rect 2696 19556 2752 19612
rect 2752 19556 2756 19612
rect 2692 19552 2756 19556
rect 2772 19612 2836 19616
rect 2772 19556 2776 19612
rect 2776 19556 2832 19612
rect 2832 19556 2836 19612
rect 2772 19552 2836 19556
rect 2852 19612 2916 19616
rect 2852 19556 2856 19612
rect 2856 19556 2912 19612
rect 2912 19556 2916 19612
rect 2852 19552 2916 19556
rect 7612 19612 7676 19616
rect 7612 19556 7616 19612
rect 7616 19556 7672 19612
rect 7672 19556 7676 19612
rect 7612 19552 7676 19556
rect 7692 19612 7756 19616
rect 7692 19556 7696 19612
rect 7696 19556 7752 19612
rect 7752 19556 7756 19612
rect 7692 19552 7756 19556
rect 7772 19612 7836 19616
rect 7772 19556 7776 19612
rect 7776 19556 7832 19612
rect 7832 19556 7836 19612
rect 7772 19552 7836 19556
rect 7852 19612 7916 19616
rect 7852 19556 7856 19612
rect 7856 19556 7912 19612
rect 7912 19556 7916 19612
rect 7852 19552 7916 19556
rect 12612 19612 12676 19616
rect 12612 19556 12616 19612
rect 12616 19556 12672 19612
rect 12672 19556 12676 19612
rect 12612 19552 12676 19556
rect 12692 19612 12756 19616
rect 12692 19556 12696 19612
rect 12696 19556 12752 19612
rect 12752 19556 12756 19612
rect 12692 19552 12756 19556
rect 12772 19612 12836 19616
rect 12772 19556 12776 19612
rect 12776 19556 12832 19612
rect 12832 19556 12836 19612
rect 12772 19552 12836 19556
rect 12852 19612 12916 19616
rect 12852 19556 12856 19612
rect 12856 19556 12912 19612
rect 12912 19556 12916 19612
rect 12852 19552 12916 19556
rect 17612 19612 17676 19616
rect 17612 19556 17616 19612
rect 17616 19556 17672 19612
rect 17672 19556 17676 19612
rect 17612 19552 17676 19556
rect 17692 19612 17756 19616
rect 17692 19556 17696 19612
rect 17696 19556 17752 19612
rect 17752 19556 17756 19612
rect 17692 19552 17756 19556
rect 17772 19612 17836 19616
rect 17772 19556 17776 19612
rect 17776 19556 17832 19612
rect 17832 19556 17836 19612
rect 17772 19552 17836 19556
rect 17852 19612 17916 19616
rect 17852 19556 17856 19612
rect 17856 19556 17912 19612
rect 17912 19556 17916 19612
rect 17852 19552 17916 19556
rect 1952 19068 2016 19072
rect 1952 19012 1956 19068
rect 1956 19012 2012 19068
rect 2012 19012 2016 19068
rect 1952 19008 2016 19012
rect 2032 19068 2096 19072
rect 2032 19012 2036 19068
rect 2036 19012 2092 19068
rect 2092 19012 2096 19068
rect 2032 19008 2096 19012
rect 2112 19068 2176 19072
rect 2112 19012 2116 19068
rect 2116 19012 2172 19068
rect 2172 19012 2176 19068
rect 2112 19008 2176 19012
rect 2192 19068 2256 19072
rect 2192 19012 2196 19068
rect 2196 19012 2252 19068
rect 2252 19012 2256 19068
rect 2192 19008 2256 19012
rect 6952 19068 7016 19072
rect 6952 19012 6956 19068
rect 6956 19012 7012 19068
rect 7012 19012 7016 19068
rect 6952 19008 7016 19012
rect 7032 19068 7096 19072
rect 7032 19012 7036 19068
rect 7036 19012 7092 19068
rect 7092 19012 7096 19068
rect 7032 19008 7096 19012
rect 7112 19068 7176 19072
rect 7112 19012 7116 19068
rect 7116 19012 7172 19068
rect 7172 19012 7176 19068
rect 7112 19008 7176 19012
rect 7192 19068 7256 19072
rect 7192 19012 7196 19068
rect 7196 19012 7252 19068
rect 7252 19012 7256 19068
rect 7192 19008 7256 19012
rect 11952 19068 12016 19072
rect 11952 19012 11956 19068
rect 11956 19012 12012 19068
rect 12012 19012 12016 19068
rect 11952 19008 12016 19012
rect 12032 19068 12096 19072
rect 12032 19012 12036 19068
rect 12036 19012 12092 19068
rect 12092 19012 12096 19068
rect 12032 19008 12096 19012
rect 12112 19068 12176 19072
rect 12112 19012 12116 19068
rect 12116 19012 12172 19068
rect 12172 19012 12176 19068
rect 12112 19008 12176 19012
rect 12192 19068 12256 19072
rect 12192 19012 12196 19068
rect 12196 19012 12252 19068
rect 12252 19012 12256 19068
rect 12192 19008 12256 19012
rect 16952 19068 17016 19072
rect 16952 19012 16956 19068
rect 16956 19012 17012 19068
rect 17012 19012 17016 19068
rect 16952 19008 17016 19012
rect 17032 19068 17096 19072
rect 17032 19012 17036 19068
rect 17036 19012 17092 19068
rect 17092 19012 17096 19068
rect 17032 19008 17096 19012
rect 17112 19068 17176 19072
rect 17112 19012 17116 19068
rect 17116 19012 17172 19068
rect 17172 19012 17176 19068
rect 17112 19008 17176 19012
rect 17192 19068 17256 19072
rect 17192 19012 17196 19068
rect 17196 19012 17252 19068
rect 17252 19012 17256 19068
rect 17192 19008 17256 19012
rect 2612 18524 2676 18528
rect 2612 18468 2616 18524
rect 2616 18468 2672 18524
rect 2672 18468 2676 18524
rect 2612 18464 2676 18468
rect 2692 18524 2756 18528
rect 2692 18468 2696 18524
rect 2696 18468 2752 18524
rect 2752 18468 2756 18524
rect 2692 18464 2756 18468
rect 2772 18524 2836 18528
rect 2772 18468 2776 18524
rect 2776 18468 2832 18524
rect 2832 18468 2836 18524
rect 2772 18464 2836 18468
rect 2852 18524 2916 18528
rect 2852 18468 2856 18524
rect 2856 18468 2912 18524
rect 2912 18468 2916 18524
rect 2852 18464 2916 18468
rect 7612 18524 7676 18528
rect 7612 18468 7616 18524
rect 7616 18468 7672 18524
rect 7672 18468 7676 18524
rect 7612 18464 7676 18468
rect 7692 18524 7756 18528
rect 7692 18468 7696 18524
rect 7696 18468 7752 18524
rect 7752 18468 7756 18524
rect 7692 18464 7756 18468
rect 7772 18524 7836 18528
rect 7772 18468 7776 18524
rect 7776 18468 7832 18524
rect 7832 18468 7836 18524
rect 7772 18464 7836 18468
rect 7852 18524 7916 18528
rect 7852 18468 7856 18524
rect 7856 18468 7912 18524
rect 7912 18468 7916 18524
rect 7852 18464 7916 18468
rect 12612 18524 12676 18528
rect 12612 18468 12616 18524
rect 12616 18468 12672 18524
rect 12672 18468 12676 18524
rect 12612 18464 12676 18468
rect 12692 18524 12756 18528
rect 12692 18468 12696 18524
rect 12696 18468 12752 18524
rect 12752 18468 12756 18524
rect 12692 18464 12756 18468
rect 12772 18524 12836 18528
rect 12772 18468 12776 18524
rect 12776 18468 12832 18524
rect 12832 18468 12836 18524
rect 12772 18464 12836 18468
rect 12852 18524 12916 18528
rect 12852 18468 12856 18524
rect 12856 18468 12912 18524
rect 12912 18468 12916 18524
rect 12852 18464 12916 18468
rect 17612 18524 17676 18528
rect 17612 18468 17616 18524
rect 17616 18468 17672 18524
rect 17672 18468 17676 18524
rect 17612 18464 17676 18468
rect 17692 18524 17756 18528
rect 17692 18468 17696 18524
rect 17696 18468 17752 18524
rect 17752 18468 17756 18524
rect 17692 18464 17756 18468
rect 17772 18524 17836 18528
rect 17772 18468 17776 18524
rect 17776 18468 17832 18524
rect 17832 18468 17836 18524
rect 17772 18464 17836 18468
rect 17852 18524 17916 18528
rect 17852 18468 17856 18524
rect 17856 18468 17912 18524
rect 17912 18468 17916 18524
rect 17852 18464 17916 18468
rect 1952 17980 2016 17984
rect 1952 17924 1956 17980
rect 1956 17924 2012 17980
rect 2012 17924 2016 17980
rect 1952 17920 2016 17924
rect 2032 17980 2096 17984
rect 2032 17924 2036 17980
rect 2036 17924 2092 17980
rect 2092 17924 2096 17980
rect 2032 17920 2096 17924
rect 2112 17980 2176 17984
rect 2112 17924 2116 17980
rect 2116 17924 2172 17980
rect 2172 17924 2176 17980
rect 2112 17920 2176 17924
rect 2192 17980 2256 17984
rect 2192 17924 2196 17980
rect 2196 17924 2252 17980
rect 2252 17924 2256 17980
rect 2192 17920 2256 17924
rect 6952 17980 7016 17984
rect 6952 17924 6956 17980
rect 6956 17924 7012 17980
rect 7012 17924 7016 17980
rect 6952 17920 7016 17924
rect 7032 17980 7096 17984
rect 7032 17924 7036 17980
rect 7036 17924 7092 17980
rect 7092 17924 7096 17980
rect 7032 17920 7096 17924
rect 7112 17980 7176 17984
rect 7112 17924 7116 17980
rect 7116 17924 7172 17980
rect 7172 17924 7176 17980
rect 7112 17920 7176 17924
rect 7192 17980 7256 17984
rect 7192 17924 7196 17980
rect 7196 17924 7252 17980
rect 7252 17924 7256 17980
rect 7192 17920 7256 17924
rect 11952 17980 12016 17984
rect 11952 17924 11956 17980
rect 11956 17924 12012 17980
rect 12012 17924 12016 17980
rect 11952 17920 12016 17924
rect 12032 17980 12096 17984
rect 12032 17924 12036 17980
rect 12036 17924 12092 17980
rect 12092 17924 12096 17980
rect 12032 17920 12096 17924
rect 12112 17980 12176 17984
rect 12112 17924 12116 17980
rect 12116 17924 12172 17980
rect 12172 17924 12176 17980
rect 12112 17920 12176 17924
rect 12192 17980 12256 17984
rect 12192 17924 12196 17980
rect 12196 17924 12252 17980
rect 12252 17924 12256 17980
rect 12192 17920 12256 17924
rect 16952 17980 17016 17984
rect 16952 17924 16956 17980
rect 16956 17924 17012 17980
rect 17012 17924 17016 17980
rect 16952 17920 17016 17924
rect 17032 17980 17096 17984
rect 17032 17924 17036 17980
rect 17036 17924 17092 17980
rect 17092 17924 17096 17980
rect 17032 17920 17096 17924
rect 17112 17980 17176 17984
rect 17112 17924 17116 17980
rect 17116 17924 17172 17980
rect 17172 17924 17176 17980
rect 17112 17920 17176 17924
rect 17192 17980 17256 17984
rect 17192 17924 17196 17980
rect 17196 17924 17252 17980
rect 17252 17924 17256 17980
rect 17192 17920 17256 17924
rect 2612 17436 2676 17440
rect 2612 17380 2616 17436
rect 2616 17380 2672 17436
rect 2672 17380 2676 17436
rect 2612 17376 2676 17380
rect 2692 17436 2756 17440
rect 2692 17380 2696 17436
rect 2696 17380 2752 17436
rect 2752 17380 2756 17436
rect 2692 17376 2756 17380
rect 2772 17436 2836 17440
rect 2772 17380 2776 17436
rect 2776 17380 2832 17436
rect 2832 17380 2836 17436
rect 2772 17376 2836 17380
rect 2852 17436 2916 17440
rect 2852 17380 2856 17436
rect 2856 17380 2912 17436
rect 2912 17380 2916 17436
rect 2852 17376 2916 17380
rect 7612 17436 7676 17440
rect 7612 17380 7616 17436
rect 7616 17380 7672 17436
rect 7672 17380 7676 17436
rect 7612 17376 7676 17380
rect 7692 17436 7756 17440
rect 7692 17380 7696 17436
rect 7696 17380 7752 17436
rect 7752 17380 7756 17436
rect 7692 17376 7756 17380
rect 7772 17436 7836 17440
rect 7772 17380 7776 17436
rect 7776 17380 7832 17436
rect 7832 17380 7836 17436
rect 7772 17376 7836 17380
rect 7852 17436 7916 17440
rect 7852 17380 7856 17436
rect 7856 17380 7912 17436
rect 7912 17380 7916 17436
rect 7852 17376 7916 17380
rect 12612 17436 12676 17440
rect 12612 17380 12616 17436
rect 12616 17380 12672 17436
rect 12672 17380 12676 17436
rect 12612 17376 12676 17380
rect 12692 17436 12756 17440
rect 12692 17380 12696 17436
rect 12696 17380 12752 17436
rect 12752 17380 12756 17436
rect 12692 17376 12756 17380
rect 12772 17436 12836 17440
rect 12772 17380 12776 17436
rect 12776 17380 12832 17436
rect 12832 17380 12836 17436
rect 12772 17376 12836 17380
rect 12852 17436 12916 17440
rect 12852 17380 12856 17436
rect 12856 17380 12912 17436
rect 12912 17380 12916 17436
rect 12852 17376 12916 17380
rect 17612 17436 17676 17440
rect 17612 17380 17616 17436
rect 17616 17380 17672 17436
rect 17672 17380 17676 17436
rect 17612 17376 17676 17380
rect 17692 17436 17756 17440
rect 17692 17380 17696 17436
rect 17696 17380 17752 17436
rect 17752 17380 17756 17436
rect 17692 17376 17756 17380
rect 17772 17436 17836 17440
rect 17772 17380 17776 17436
rect 17776 17380 17832 17436
rect 17832 17380 17836 17436
rect 17772 17376 17836 17380
rect 17852 17436 17916 17440
rect 17852 17380 17856 17436
rect 17856 17380 17912 17436
rect 17912 17380 17916 17436
rect 17852 17376 17916 17380
rect 1952 16892 2016 16896
rect 1952 16836 1956 16892
rect 1956 16836 2012 16892
rect 2012 16836 2016 16892
rect 1952 16832 2016 16836
rect 2032 16892 2096 16896
rect 2032 16836 2036 16892
rect 2036 16836 2092 16892
rect 2092 16836 2096 16892
rect 2032 16832 2096 16836
rect 2112 16892 2176 16896
rect 2112 16836 2116 16892
rect 2116 16836 2172 16892
rect 2172 16836 2176 16892
rect 2112 16832 2176 16836
rect 2192 16892 2256 16896
rect 2192 16836 2196 16892
rect 2196 16836 2252 16892
rect 2252 16836 2256 16892
rect 2192 16832 2256 16836
rect 6952 16892 7016 16896
rect 6952 16836 6956 16892
rect 6956 16836 7012 16892
rect 7012 16836 7016 16892
rect 6952 16832 7016 16836
rect 7032 16892 7096 16896
rect 7032 16836 7036 16892
rect 7036 16836 7092 16892
rect 7092 16836 7096 16892
rect 7032 16832 7096 16836
rect 7112 16892 7176 16896
rect 7112 16836 7116 16892
rect 7116 16836 7172 16892
rect 7172 16836 7176 16892
rect 7112 16832 7176 16836
rect 7192 16892 7256 16896
rect 7192 16836 7196 16892
rect 7196 16836 7252 16892
rect 7252 16836 7256 16892
rect 7192 16832 7256 16836
rect 11952 16892 12016 16896
rect 11952 16836 11956 16892
rect 11956 16836 12012 16892
rect 12012 16836 12016 16892
rect 11952 16832 12016 16836
rect 12032 16892 12096 16896
rect 12032 16836 12036 16892
rect 12036 16836 12092 16892
rect 12092 16836 12096 16892
rect 12032 16832 12096 16836
rect 12112 16892 12176 16896
rect 12112 16836 12116 16892
rect 12116 16836 12172 16892
rect 12172 16836 12176 16892
rect 12112 16832 12176 16836
rect 12192 16892 12256 16896
rect 12192 16836 12196 16892
rect 12196 16836 12252 16892
rect 12252 16836 12256 16892
rect 12192 16832 12256 16836
rect 16952 16892 17016 16896
rect 16952 16836 16956 16892
rect 16956 16836 17012 16892
rect 17012 16836 17016 16892
rect 16952 16832 17016 16836
rect 17032 16892 17096 16896
rect 17032 16836 17036 16892
rect 17036 16836 17092 16892
rect 17092 16836 17096 16892
rect 17032 16832 17096 16836
rect 17112 16892 17176 16896
rect 17112 16836 17116 16892
rect 17116 16836 17172 16892
rect 17172 16836 17176 16892
rect 17112 16832 17176 16836
rect 17192 16892 17256 16896
rect 17192 16836 17196 16892
rect 17196 16836 17252 16892
rect 17252 16836 17256 16892
rect 17192 16832 17256 16836
rect 6316 16628 6380 16692
rect 14596 16492 14660 16556
rect 2612 16348 2676 16352
rect 2612 16292 2616 16348
rect 2616 16292 2672 16348
rect 2672 16292 2676 16348
rect 2612 16288 2676 16292
rect 2692 16348 2756 16352
rect 2692 16292 2696 16348
rect 2696 16292 2752 16348
rect 2752 16292 2756 16348
rect 2692 16288 2756 16292
rect 2772 16348 2836 16352
rect 2772 16292 2776 16348
rect 2776 16292 2832 16348
rect 2832 16292 2836 16348
rect 2772 16288 2836 16292
rect 2852 16348 2916 16352
rect 2852 16292 2856 16348
rect 2856 16292 2912 16348
rect 2912 16292 2916 16348
rect 2852 16288 2916 16292
rect 7612 16348 7676 16352
rect 7612 16292 7616 16348
rect 7616 16292 7672 16348
rect 7672 16292 7676 16348
rect 7612 16288 7676 16292
rect 7692 16348 7756 16352
rect 7692 16292 7696 16348
rect 7696 16292 7752 16348
rect 7752 16292 7756 16348
rect 7692 16288 7756 16292
rect 7772 16348 7836 16352
rect 7772 16292 7776 16348
rect 7776 16292 7832 16348
rect 7832 16292 7836 16348
rect 7772 16288 7836 16292
rect 7852 16348 7916 16352
rect 7852 16292 7856 16348
rect 7856 16292 7912 16348
rect 7912 16292 7916 16348
rect 7852 16288 7916 16292
rect 12612 16348 12676 16352
rect 12612 16292 12616 16348
rect 12616 16292 12672 16348
rect 12672 16292 12676 16348
rect 12612 16288 12676 16292
rect 12692 16348 12756 16352
rect 12692 16292 12696 16348
rect 12696 16292 12752 16348
rect 12752 16292 12756 16348
rect 12692 16288 12756 16292
rect 12772 16348 12836 16352
rect 12772 16292 12776 16348
rect 12776 16292 12832 16348
rect 12832 16292 12836 16348
rect 12772 16288 12836 16292
rect 12852 16348 12916 16352
rect 12852 16292 12856 16348
rect 12856 16292 12912 16348
rect 12912 16292 12916 16348
rect 12852 16288 12916 16292
rect 17612 16348 17676 16352
rect 17612 16292 17616 16348
rect 17616 16292 17672 16348
rect 17672 16292 17676 16348
rect 17612 16288 17676 16292
rect 17692 16348 17756 16352
rect 17692 16292 17696 16348
rect 17696 16292 17752 16348
rect 17752 16292 17756 16348
rect 17692 16288 17756 16292
rect 17772 16348 17836 16352
rect 17772 16292 17776 16348
rect 17776 16292 17832 16348
rect 17832 16292 17836 16348
rect 17772 16288 17836 16292
rect 17852 16348 17916 16352
rect 17852 16292 17856 16348
rect 17856 16292 17912 16348
rect 17912 16292 17916 16348
rect 17852 16288 17916 16292
rect 1952 15804 2016 15808
rect 1952 15748 1956 15804
rect 1956 15748 2012 15804
rect 2012 15748 2016 15804
rect 1952 15744 2016 15748
rect 2032 15804 2096 15808
rect 2032 15748 2036 15804
rect 2036 15748 2092 15804
rect 2092 15748 2096 15804
rect 2032 15744 2096 15748
rect 2112 15804 2176 15808
rect 2112 15748 2116 15804
rect 2116 15748 2172 15804
rect 2172 15748 2176 15804
rect 2112 15744 2176 15748
rect 2192 15804 2256 15808
rect 2192 15748 2196 15804
rect 2196 15748 2252 15804
rect 2252 15748 2256 15804
rect 2192 15744 2256 15748
rect 6952 15804 7016 15808
rect 6952 15748 6956 15804
rect 6956 15748 7012 15804
rect 7012 15748 7016 15804
rect 6952 15744 7016 15748
rect 7032 15804 7096 15808
rect 7032 15748 7036 15804
rect 7036 15748 7092 15804
rect 7092 15748 7096 15804
rect 7032 15744 7096 15748
rect 7112 15804 7176 15808
rect 7112 15748 7116 15804
rect 7116 15748 7172 15804
rect 7172 15748 7176 15804
rect 7112 15744 7176 15748
rect 7192 15804 7256 15808
rect 7192 15748 7196 15804
rect 7196 15748 7252 15804
rect 7252 15748 7256 15804
rect 7192 15744 7256 15748
rect 11952 15804 12016 15808
rect 11952 15748 11956 15804
rect 11956 15748 12012 15804
rect 12012 15748 12016 15804
rect 11952 15744 12016 15748
rect 12032 15804 12096 15808
rect 12032 15748 12036 15804
rect 12036 15748 12092 15804
rect 12092 15748 12096 15804
rect 12032 15744 12096 15748
rect 12112 15804 12176 15808
rect 12112 15748 12116 15804
rect 12116 15748 12172 15804
rect 12172 15748 12176 15804
rect 12112 15744 12176 15748
rect 12192 15804 12256 15808
rect 12192 15748 12196 15804
rect 12196 15748 12252 15804
rect 12252 15748 12256 15804
rect 12192 15744 12256 15748
rect 16952 15804 17016 15808
rect 16952 15748 16956 15804
rect 16956 15748 17012 15804
rect 17012 15748 17016 15804
rect 16952 15744 17016 15748
rect 17032 15804 17096 15808
rect 17032 15748 17036 15804
rect 17036 15748 17092 15804
rect 17092 15748 17096 15804
rect 17032 15744 17096 15748
rect 17112 15804 17176 15808
rect 17112 15748 17116 15804
rect 17116 15748 17172 15804
rect 17172 15748 17176 15804
rect 17112 15744 17176 15748
rect 17192 15804 17256 15808
rect 17192 15748 17196 15804
rect 17196 15748 17252 15804
rect 17252 15748 17256 15804
rect 17192 15744 17256 15748
rect 11284 15540 11348 15604
rect 2612 15260 2676 15264
rect 2612 15204 2616 15260
rect 2616 15204 2672 15260
rect 2672 15204 2676 15260
rect 2612 15200 2676 15204
rect 2692 15260 2756 15264
rect 2692 15204 2696 15260
rect 2696 15204 2752 15260
rect 2752 15204 2756 15260
rect 2692 15200 2756 15204
rect 2772 15260 2836 15264
rect 2772 15204 2776 15260
rect 2776 15204 2832 15260
rect 2832 15204 2836 15260
rect 2772 15200 2836 15204
rect 2852 15260 2916 15264
rect 2852 15204 2856 15260
rect 2856 15204 2912 15260
rect 2912 15204 2916 15260
rect 2852 15200 2916 15204
rect 7612 15260 7676 15264
rect 7612 15204 7616 15260
rect 7616 15204 7672 15260
rect 7672 15204 7676 15260
rect 7612 15200 7676 15204
rect 7692 15260 7756 15264
rect 7692 15204 7696 15260
rect 7696 15204 7752 15260
rect 7752 15204 7756 15260
rect 7692 15200 7756 15204
rect 7772 15260 7836 15264
rect 7772 15204 7776 15260
rect 7776 15204 7832 15260
rect 7832 15204 7836 15260
rect 7772 15200 7836 15204
rect 7852 15260 7916 15264
rect 7852 15204 7856 15260
rect 7856 15204 7912 15260
rect 7912 15204 7916 15260
rect 7852 15200 7916 15204
rect 12612 15260 12676 15264
rect 12612 15204 12616 15260
rect 12616 15204 12672 15260
rect 12672 15204 12676 15260
rect 12612 15200 12676 15204
rect 12692 15260 12756 15264
rect 12692 15204 12696 15260
rect 12696 15204 12752 15260
rect 12752 15204 12756 15260
rect 12692 15200 12756 15204
rect 12772 15260 12836 15264
rect 12772 15204 12776 15260
rect 12776 15204 12832 15260
rect 12832 15204 12836 15260
rect 12772 15200 12836 15204
rect 12852 15260 12916 15264
rect 12852 15204 12856 15260
rect 12856 15204 12912 15260
rect 12912 15204 12916 15260
rect 12852 15200 12916 15204
rect 17612 15260 17676 15264
rect 17612 15204 17616 15260
rect 17616 15204 17672 15260
rect 17672 15204 17676 15260
rect 17612 15200 17676 15204
rect 17692 15260 17756 15264
rect 17692 15204 17696 15260
rect 17696 15204 17752 15260
rect 17752 15204 17756 15260
rect 17692 15200 17756 15204
rect 17772 15260 17836 15264
rect 17772 15204 17776 15260
rect 17776 15204 17832 15260
rect 17832 15204 17836 15260
rect 17772 15200 17836 15204
rect 17852 15260 17916 15264
rect 17852 15204 17856 15260
rect 17856 15204 17912 15260
rect 17912 15204 17916 15260
rect 17852 15200 17916 15204
rect 8524 15132 8588 15196
rect 3924 14996 3988 15060
rect 1532 14860 1596 14924
rect 1952 14716 2016 14720
rect 1952 14660 1956 14716
rect 1956 14660 2012 14716
rect 2012 14660 2016 14716
rect 1952 14656 2016 14660
rect 2032 14716 2096 14720
rect 2032 14660 2036 14716
rect 2036 14660 2092 14716
rect 2092 14660 2096 14716
rect 2032 14656 2096 14660
rect 2112 14716 2176 14720
rect 2112 14660 2116 14716
rect 2116 14660 2172 14716
rect 2172 14660 2176 14716
rect 2112 14656 2176 14660
rect 2192 14716 2256 14720
rect 2192 14660 2196 14716
rect 2196 14660 2252 14716
rect 2252 14660 2256 14716
rect 2192 14656 2256 14660
rect 6952 14716 7016 14720
rect 6952 14660 6956 14716
rect 6956 14660 7012 14716
rect 7012 14660 7016 14716
rect 6952 14656 7016 14660
rect 7032 14716 7096 14720
rect 7032 14660 7036 14716
rect 7036 14660 7092 14716
rect 7092 14660 7096 14716
rect 7032 14656 7096 14660
rect 7112 14716 7176 14720
rect 7112 14660 7116 14716
rect 7116 14660 7172 14716
rect 7172 14660 7176 14716
rect 7112 14656 7176 14660
rect 7192 14716 7256 14720
rect 7192 14660 7196 14716
rect 7196 14660 7252 14716
rect 7252 14660 7256 14716
rect 7192 14656 7256 14660
rect 11952 14716 12016 14720
rect 11952 14660 11956 14716
rect 11956 14660 12012 14716
rect 12012 14660 12016 14716
rect 11952 14656 12016 14660
rect 12032 14716 12096 14720
rect 12032 14660 12036 14716
rect 12036 14660 12092 14716
rect 12092 14660 12096 14716
rect 12032 14656 12096 14660
rect 12112 14716 12176 14720
rect 12112 14660 12116 14716
rect 12116 14660 12172 14716
rect 12172 14660 12176 14716
rect 12112 14656 12176 14660
rect 12192 14716 12256 14720
rect 12192 14660 12196 14716
rect 12196 14660 12252 14716
rect 12252 14660 12256 14716
rect 12192 14656 12256 14660
rect 16952 14716 17016 14720
rect 16952 14660 16956 14716
rect 16956 14660 17012 14716
rect 17012 14660 17016 14716
rect 16952 14656 17016 14660
rect 17032 14716 17096 14720
rect 17032 14660 17036 14716
rect 17036 14660 17092 14716
rect 17092 14660 17096 14716
rect 17032 14656 17096 14660
rect 17112 14716 17176 14720
rect 17112 14660 17116 14716
rect 17116 14660 17172 14716
rect 17172 14660 17176 14716
rect 17112 14656 17176 14660
rect 17192 14716 17256 14720
rect 17192 14660 17196 14716
rect 17196 14660 17252 14716
rect 17252 14660 17256 14716
rect 17192 14656 17256 14660
rect 2612 14172 2676 14176
rect 2612 14116 2616 14172
rect 2616 14116 2672 14172
rect 2672 14116 2676 14172
rect 2612 14112 2676 14116
rect 2692 14172 2756 14176
rect 2692 14116 2696 14172
rect 2696 14116 2752 14172
rect 2752 14116 2756 14172
rect 2692 14112 2756 14116
rect 2772 14172 2836 14176
rect 2772 14116 2776 14172
rect 2776 14116 2832 14172
rect 2832 14116 2836 14172
rect 2772 14112 2836 14116
rect 2852 14172 2916 14176
rect 2852 14116 2856 14172
rect 2856 14116 2912 14172
rect 2912 14116 2916 14172
rect 2852 14112 2916 14116
rect 7612 14172 7676 14176
rect 7612 14116 7616 14172
rect 7616 14116 7672 14172
rect 7672 14116 7676 14172
rect 7612 14112 7676 14116
rect 7692 14172 7756 14176
rect 7692 14116 7696 14172
rect 7696 14116 7752 14172
rect 7752 14116 7756 14172
rect 7692 14112 7756 14116
rect 7772 14172 7836 14176
rect 7772 14116 7776 14172
rect 7776 14116 7832 14172
rect 7832 14116 7836 14172
rect 7772 14112 7836 14116
rect 7852 14172 7916 14176
rect 7852 14116 7856 14172
rect 7856 14116 7912 14172
rect 7912 14116 7916 14172
rect 7852 14112 7916 14116
rect 12612 14172 12676 14176
rect 12612 14116 12616 14172
rect 12616 14116 12672 14172
rect 12672 14116 12676 14172
rect 12612 14112 12676 14116
rect 12692 14172 12756 14176
rect 12692 14116 12696 14172
rect 12696 14116 12752 14172
rect 12752 14116 12756 14172
rect 12692 14112 12756 14116
rect 12772 14172 12836 14176
rect 12772 14116 12776 14172
rect 12776 14116 12832 14172
rect 12832 14116 12836 14172
rect 12772 14112 12836 14116
rect 12852 14172 12916 14176
rect 12852 14116 12856 14172
rect 12856 14116 12912 14172
rect 12912 14116 12916 14172
rect 12852 14112 12916 14116
rect 17612 14172 17676 14176
rect 17612 14116 17616 14172
rect 17616 14116 17672 14172
rect 17672 14116 17676 14172
rect 17612 14112 17676 14116
rect 17692 14172 17756 14176
rect 17692 14116 17696 14172
rect 17696 14116 17752 14172
rect 17752 14116 17756 14172
rect 17692 14112 17756 14116
rect 17772 14172 17836 14176
rect 17772 14116 17776 14172
rect 17776 14116 17832 14172
rect 17832 14116 17836 14172
rect 17772 14112 17836 14116
rect 17852 14172 17916 14176
rect 17852 14116 17856 14172
rect 17856 14116 17912 14172
rect 17912 14116 17916 14172
rect 17852 14112 17916 14116
rect 1952 13628 2016 13632
rect 1952 13572 1956 13628
rect 1956 13572 2012 13628
rect 2012 13572 2016 13628
rect 1952 13568 2016 13572
rect 2032 13628 2096 13632
rect 2032 13572 2036 13628
rect 2036 13572 2092 13628
rect 2092 13572 2096 13628
rect 2032 13568 2096 13572
rect 2112 13628 2176 13632
rect 2112 13572 2116 13628
rect 2116 13572 2172 13628
rect 2172 13572 2176 13628
rect 2112 13568 2176 13572
rect 2192 13628 2256 13632
rect 2192 13572 2196 13628
rect 2196 13572 2252 13628
rect 2252 13572 2256 13628
rect 2192 13568 2256 13572
rect 6952 13628 7016 13632
rect 6952 13572 6956 13628
rect 6956 13572 7012 13628
rect 7012 13572 7016 13628
rect 6952 13568 7016 13572
rect 7032 13628 7096 13632
rect 7032 13572 7036 13628
rect 7036 13572 7092 13628
rect 7092 13572 7096 13628
rect 7032 13568 7096 13572
rect 7112 13628 7176 13632
rect 7112 13572 7116 13628
rect 7116 13572 7172 13628
rect 7172 13572 7176 13628
rect 7112 13568 7176 13572
rect 7192 13628 7256 13632
rect 7192 13572 7196 13628
rect 7196 13572 7252 13628
rect 7252 13572 7256 13628
rect 7192 13568 7256 13572
rect 11952 13628 12016 13632
rect 11952 13572 11956 13628
rect 11956 13572 12012 13628
rect 12012 13572 12016 13628
rect 11952 13568 12016 13572
rect 12032 13628 12096 13632
rect 12032 13572 12036 13628
rect 12036 13572 12092 13628
rect 12092 13572 12096 13628
rect 12032 13568 12096 13572
rect 12112 13628 12176 13632
rect 12112 13572 12116 13628
rect 12116 13572 12172 13628
rect 12172 13572 12176 13628
rect 12112 13568 12176 13572
rect 12192 13628 12256 13632
rect 12192 13572 12196 13628
rect 12196 13572 12252 13628
rect 12252 13572 12256 13628
rect 12192 13568 12256 13572
rect 16952 13628 17016 13632
rect 16952 13572 16956 13628
rect 16956 13572 17012 13628
rect 17012 13572 17016 13628
rect 16952 13568 17016 13572
rect 17032 13628 17096 13632
rect 17032 13572 17036 13628
rect 17036 13572 17092 13628
rect 17092 13572 17096 13628
rect 17032 13568 17096 13572
rect 17112 13628 17176 13632
rect 17112 13572 17116 13628
rect 17116 13572 17172 13628
rect 17172 13572 17176 13628
rect 17112 13568 17176 13572
rect 17192 13628 17256 13632
rect 17192 13572 17196 13628
rect 17196 13572 17252 13628
rect 17252 13572 17256 13628
rect 17192 13568 17256 13572
rect 11468 13228 11532 13292
rect 2612 13084 2676 13088
rect 2612 13028 2616 13084
rect 2616 13028 2672 13084
rect 2672 13028 2676 13084
rect 2612 13024 2676 13028
rect 2692 13084 2756 13088
rect 2692 13028 2696 13084
rect 2696 13028 2752 13084
rect 2752 13028 2756 13084
rect 2692 13024 2756 13028
rect 2772 13084 2836 13088
rect 2772 13028 2776 13084
rect 2776 13028 2832 13084
rect 2832 13028 2836 13084
rect 2772 13024 2836 13028
rect 2852 13084 2916 13088
rect 2852 13028 2856 13084
rect 2856 13028 2912 13084
rect 2912 13028 2916 13084
rect 2852 13024 2916 13028
rect 7612 13084 7676 13088
rect 7612 13028 7616 13084
rect 7616 13028 7672 13084
rect 7672 13028 7676 13084
rect 7612 13024 7676 13028
rect 7692 13084 7756 13088
rect 7692 13028 7696 13084
rect 7696 13028 7752 13084
rect 7752 13028 7756 13084
rect 7692 13024 7756 13028
rect 7772 13084 7836 13088
rect 7772 13028 7776 13084
rect 7776 13028 7832 13084
rect 7832 13028 7836 13084
rect 7772 13024 7836 13028
rect 7852 13084 7916 13088
rect 7852 13028 7856 13084
rect 7856 13028 7912 13084
rect 7912 13028 7916 13084
rect 7852 13024 7916 13028
rect 12612 13084 12676 13088
rect 12612 13028 12616 13084
rect 12616 13028 12672 13084
rect 12672 13028 12676 13084
rect 12612 13024 12676 13028
rect 12692 13084 12756 13088
rect 12692 13028 12696 13084
rect 12696 13028 12752 13084
rect 12752 13028 12756 13084
rect 12692 13024 12756 13028
rect 12772 13084 12836 13088
rect 12772 13028 12776 13084
rect 12776 13028 12832 13084
rect 12832 13028 12836 13084
rect 12772 13024 12836 13028
rect 12852 13084 12916 13088
rect 12852 13028 12856 13084
rect 12856 13028 12912 13084
rect 12912 13028 12916 13084
rect 12852 13024 12916 13028
rect 17612 13084 17676 13088
rect 17612 13028 17616 13084
rect 17616 13028 17672 13084
rect 17672 13028 17676 13084
rect 17612 13024 17676 13028
rect 17692 13084 17756 13088
rect 17692 13028 17696 13084
rect 17696 13028 17752 13084
rect 17752 13028 17756 13084
rect 17692 13024 17756 13028
rect 17772 13084 17836 13088
rect 17772 13028 17776 13084
rect 17776 13028 17832 13084
rect 17832 13028 17836 13084
rect 17772 13024 17836 13028
rect 17852 13084 17916 13088
rect 17852 13028 17856 13084
rect 17856 13028 17912 13084
rect 17912 13028 17916 13084
rect 17852 13024 17916 13028
rect 1952 12540 2016 12544
rect 1952 12484 1956 12540
rect 1956 12484 2012 12540
rect 2012 12484 2016 12540
rect 1952 12480 2016 12484
rect 2032 12540 2096 12544
rect 2032 12484 2036 12540
rect 2036 12484 2092 12540
rect 2092 12484 2096 12540
rect 2032 12480 2096 12484
rect 2112 12540 2176 12544
rect 2112 12484 2116 12540
rect 2116 12484 2172 12540
rect 2172 12484 2176 12540
rect 2112 12480 2176 12484
rect 2192 12540 2256 12544
rect 2192 12484 2196 12540
rect 2196 12484 2252 12540
rect 2252 12484 2256 12540
rect 2192 12480 2256 12484
rect 6952 12540 7016 12544
rect 6952 12484 6956 12540
rect 6956 12484 7012 12540
rect 7012 12484 7016 12540
rect 6952 12480 7016 12484
rect 7032 12540 7096 12544
rect 7032 12484 7036 12540
rect 7036 12484 7092 12540
rect 7092 12484 7096 12540
rect 7032 12480 7096 12484
rect 7112 12540 7176 12544
rect 7112 12484 7116 12540
rect 7116 12484 7172 12540
rect 7172 12484 7176 12540
rect 7112 12480 7176 12484
rect 7192 12540 7256 12544
rect 7192 12484 7196 12540
rect 7196 12484 7252 12540
rect 7252 12484 7256 12540
rect 7192 12480 7256 12484
rect 11952 12540 12016 12544
rect 11952 12484 11956 12540
rect 11956 12484 12012 12540
rect 12012 12484 12016 12540
rect 11952 12480 12016 12484
rect 12032 12540 12096 12544
rect 12032 12484 12036 12540
rect 12036 12484 12092 12540
rect 12092 12484 12096 12540
rect 12032 12480 12096 12484
rect 12112 12540 12176 12544
rect 12112 12484 12116 12540
rect 12116 12484 12172 12540
rect 12172 12484 12176 12540
rect 12112 12480 12176 12484
rect 12192 12540 12256 12544
rect 12192 12484 12196 12540
rect 12196 12484 12252 12540
rect 12252 12484 12256 12540
rect 12192 12480 12256 12484
rect 16952 12540 17016 12544
rect 16952 12484 16956 12540
rect 16956 12484 17012 12540
rect 17012 12484 17016 12540
rect 16952 12480 17016 12484
rect 17032 12540 17096 12544
rect 17032 12484 17036 12540
rect 17036 12484 17092 12540
rect 17092 12484 17096 12540
rect 17032 12480 17096 12484
rect 17112 12540 17176 12544
rect 17112 12484 17116 12540
rect 17116 12484 17172 12540
rect 17172 12484 17176 12540
rect 17112 12480 17176 12484
rect 17192 12540 17256 12544
rect 17192 12484 17196 12540
rect 17196 12484 17252 12540
rect 17252 12484 17256 12540
rect 17192 12480 17256 12484
rect 9076 12276 9140 12340
rect 13676 12140 13740 12204
rect 2612 11996 2676 12000
rect 2612 11940 2616 11996
rect 2616 11940 2672 11996
rect 2672 11940 2676 11996
rect 2612 11936 2676 11940
rect 2692 11996 2756 12000
rect 2692 11940 2696 11996
rect 2696 11940 2752 11996
rect 2752 11940 2756 11996
rect 2692 11936 2756 11940
rect 2772 11996 2836 12000
rect 2772 11940 2776 11996
rect 2776 11940 2832 11996
rect 2832 11940 2836 11996
rect 2772 11936 2836 11940
rect 2852 11996 2916 12000
rect 2852 11940 2856 11996
rect 2856 11940 2912 11996
rect 2912 11940 2916 11996
rect 2852 11936 2916 11940
rect 7612 11996 7676 12000
rect 7612 11940 7616 11996
rect 7616 11940 7672 11996
rect 7672 11940 7676 11996
rect 7612 11936 7676 11940
rect 7692 11996 7756 12000
rect 7692 11940 7696 11996
rect 7696 11940 7752 11996
rect 7752 11940 7756 11996
rect 7692 11936 7756 11940
rect 7772 11996 7836 12000
rect 7772 11940 7776 11996
rect 7776 11940 7832 11996
rect 7832 11940 7836 11996
rect 7772 11936 7836 11940
rect 7852 11996 7916 12000
rect 7852 11940 7856 11996
rect 7856 11940 7912 11996
rect 7912 11940 7916 11996
rect 7852 11936 7916 11940
rect 12612 11996 12676 12000
rect 12612 11940 12616 11996
rect 12616 11940 12672 11996
rect 12672 11940 12676 11996
rect 12612 11936 12676 11940
rect 12692 11996 12756 12000
rect 12692 11940 12696 11996
rect 12696 11940 12752 11996
rect 12752 11940 12756 11996
rect 12692 11936 12756 11940
rect 12772 11996 12836 12000
rect 12772 11940 12776 11996
rect 12776 11940 12832 11996
rect 12832 11940 12836 11996
rect 12772 11936 12836 11940
rect 12852 11996 12916 12000
rect 12852 11940 12856 11996
rect 12856 11940 12912 11996
rect 12912 11940 12916 11996
rect 12852 11936 12916 11940
rect 17612 11996 17676 12000
rect 17612 11940 17616 11996
rect 17616 11940 17672 11996
rect 17672 11940 17676 11996
rect 17612 11936 17676 11940
rect 17692 11996 17756 12000
rect 17692 11940 17696 11996
rect 17696 11940 17752 11996
rect 17752 11940 17756 11996
rect 17692 11936 17756 11940
rect 17772 11996 17836 12000
rect 17772 11940 17776 11996
rect 17776 11940 17832 11996
rect 17832 11940 17836 11996
rect 17772 11936 17836 11940
rect 17852 11996 17916 12000
rect 17852 11940 17856 11996
rect 17856 11940 17912 11996
rect 17912 11940 17916 11996
rect 17852 11936 17916 11940
rect 1952 11452 2016 11456
rect 1952 11396 1956 11452
rect 1956 11396 2012 11452
rect 2012 11396 2016 11452
rect 1952 11392 2016 11396
rect 2032 11452 2096 11456
rect 2032 11396 2036 11452
rect 2036 11396 2092 11452
rect 2092 11396 2096 11452
rect 2032 11392 2096 11396
rect 2112 11452 2176 11456
rect 2112 11396 2116 11452
rect 2116 11396 2172 11452
rect 2172 11396 2176 11452
rect 2112 11392 2176 11396
rect 2192 11452 2256 11456
rect 2192 11396 2196 11452
rect 2196 11396 2252 11452
rect 2252 11396 2256 11452
rect 2192 11392 2256 11396
rect 6952 11452 7016 11456
rect 6952 11396 6956 11452
rect 6956 11396 7012 11452
rect 7012 11396 7016 11452
rect 6952 11392 7016 11396
rect 7032 11452 7096 11456
rect 7032 11396 7036 11452
rect 7036 11396 7092 11452
rect 7092 11396 7096 11452
rect 7032 11392 7096 11396
rect 7112 11452 7176 11456
rect 7112 11396 7116 11452
rect 7116 11396 7172 11452
rect 7172 11396 7176 11452
rect 7112 11392 7176 11396
rect 7192 11452 7256 11456
rect 7192 11396 7196 11452
rect 7196 11396 7252 11452
rect 7252 11396 7256 11452
rect 7192 11392 7256 11396
rect 11952 11452 12016 11456
rect 11952 11396 11956 11452
rect 11956 11396 12012 11452
rect 12012 11396 12016 11452
rect 11952 11392 12016 11396
rect 12032 11452 12096 11456
rect 12032 11396 12036 11452
rect 12036 11396 12092 11452
rect 12092 11396 12096 11452
rect 12032 11392 12096 11396
rect 12112 11452 12176 11456
rect 12112 11396 12116 11452
rect 12116 11396 12172 11452
rect 12172 11396 12176 11452
rect 12112 11392 12176 11396
rect 12192 11452 12256 11456
rect 12192 11396 12196 11452
rect 12196 11396 12252 11452
rect 12252 11396 12256 11452
rect 12192 11392 12256 11396
rect 16952 11452 17016 11456
rect 16952 11396 16956 11452
rect 16956 11396 17012 11452
rect 17012 11396 17016 11452
rect 16952 11392 17016 11396
rect 17032 11452 17096 11456
rect 17032 11396 17036 11452
rect 17036 11396 17092 11452
rect 17092 11396 17096 11452
rect 17032 11392 17096 11396
rect 17112 11452 17176 11456
rect 17112 11396 17116 11452
rect 17116 11396 17172 11452
rect 17172 11396 17176 11452
rect 17112 11392 17176 11396
rect 17192 11452 17256 11456
rect 17192 11396 17196 11452
rect 17196 11396 17252 11452
rect 17252 11396 17256 11452
rect 17192 11392 17256 11396
rect 8892 11188 8956 11252
rect 15700 11052 15764 11116
rect 2612 10908 2676 10912
rect 2612 10852 2616 10908
rect 2616 10852 2672 10908
rect 2672 10852 2676 10908
rect 2612 10848 2676 10852
rect 2692 10908 2756 10912
rect 2692 10852 2696 10908
rect 2696 10852 2752 10908
rect 2752 10852 2756 10908
rect 2692 10848 2756 10852
rect 2772 10908 2836 10912
rect 2772 10852 2776 10908
rect 2776 10852 2832 10908
rect 2832 10852 2836 10908
rect 2772 10848 2836 10852
rect 2852 10908 2916 10912
rect 2852 10852 2856 10908
rect 2856 10852 2912 10908
rect 2912 10852 2916 10908
rect 2852 10848 2916 10852
rect 7612 10908 7676 10912
rect 7612 10852 7616 10908
rect 7616 10852 7672 10908
rect 7672 10852 7676 10908
rect 7612 10848 7676 10852
rect 7692 10908 7756 10912
rect 7692 10852 7696 10908
rect 7696 10852 7752 10908
rect 7752 10852 7756 10908
rect 7692 10848 7756 10852
rect 7772 10908 7836 10912
rect 7772 10852 7776 10908
rect 7776 10852 7832 10908
rect 7832 10852 7836 10908
rect 7772 10848 7836 10852
rect 7852 10908 7916 10912
rect 7852 10852 7856 10908
rect 7856 10852 7912 10908
rect 7912 10852 7916 10908
rect 7852 10848 7916 10852
rect 12612 10908 12676 10912
rect 12612 10852 12616 10908
rect 12616 10852 12672 10908
rect 12672 10852 12676 10908
rect 12612 10848 12676 10852
rect 12692 10908 12756 10912
rect 12692 10852 12696 10908
rect 12696 10852 12752 10908
rect 12752 10852 12756 10908
rect 12692 10848 12756 10852
rect 12772 10908 12836 10912
rect 12772 10852 12776 10908
rect 12776 10852 12832 10908
rect 12832 10852 12836 10908
rect 12772 10848 12836 10852
rect 12852 10908 12916 10912
rect 12852 10852 12856 10908
rect 12856 10852 12912 10908
rect 12912 10852 12916 10908
rect 12852 10848 12916 10852
rect 17612 10908 17676 10912
rect 17612 10852 17616 10908
rect 17616 10852 17672 10908
rect 17672 10852 17676 10908
rect 17612 10848 17676 10852
rect 17692 10908 17756 10912
rect 17692 10852 17696 10908
rect 17696 10852 17752 10908
rect 17752 10852 17756 10908
rect 17692 10848 17756 10852
rect 17772 10908 17836 10912
rect 17772 10852 17776 10908
rect 17776 10852 17832 10908
rect 17832 10852 17836 10908
rect 17772 10848 17836 10852
rect 17852 10908 17916 10912
rect 17852 10852 17856 10908
rect 17856 10852 17912 10908
rect 17912 10852 17916 10908
rect 17852 10848 17916 10852
rect 6132 10644 6196 10708
rect 15148 10508 15212 10572
rect 1952 10364 2016 10368
rect 1952 10308 1956 10364
rect 1956 10308 2012 10364
rect 2012 10308 2016 10364
rect 1952 10304 2016 10308
rect 2032 10364 2096 10368
rect 2032 10308 2036 10364
rect 2036 10308 2092 10364
rect 2092 10308 2096 10364
rect 2032 10304 2096 10308
rect 2112 10364 2176 10368
rect 2112 10308 2116 10364
rect 2116 10308 2172 10364
rect 2172 10308 2176 10364
rect 2112 10304 2176 10308
rect 2192 10364 2256 10368
rect 2192 10308 2196 10364
rect 2196 10308 2252 10364
rect 2252 10308 2256 10364
rect 2192 10304 2256 10308
rect 6952 10364 7016 10368
rect 6952 10308 6956 10364
rect 6956 10308 7012 10364
rect 7012 10308 7016 10364
rect 6952 10304 7016 10308
rect 7032 10364 7096 10368
rect 7032 10308 7036 10364
rect 7036 10308 7092 10364
rect 7092 10308 7096 10364
rect 7032 10304 7096 10308
rect 7112 10364 7176 10368
rect 7112 10308 7116 10364
rect 7116 10308 7172 10364
rect 7172 10308 7176 10364
rect 7112 10304 7176 10308
rect 7192 10364 7256 10368
rect 7192 10308 7196 10364
rect 7196 10308 7252 10364
rect 7252 10308 7256 10364
rect 7192 10304 7256 10308
rect 11952 10364 12016 10368
rect 11952 10308 11956 10364
rect 11956 10308 12012 10364
rect 12012 10308 12016 10364
rect 11952 10304 12016 10308
rect 12032 10364 12096 10368
rect 12032 10308 12036 10364
rect 12036 10308 12092 10364
rect 12092 10308 12096 10364
rect 12032 10304 12096 10308
rect 12112 10364 12176 10368
rect 12112 10308 12116 10364
rect 12116 10308 12172 10364
rect 12172 10308 12176 10364
rect 12112 10304 12176 10308
rect 12192 10364 12256 10368
rect 12192 10308 12196 10364
rect 12196 10308 12252 10364
rect 12252 10308 12256 10364
rect 12192 10304 12256 10308
rect 16952 10364 17016 10368
rect 16952 10308 16956 10364
rect 16956 10308 17012 10364
rect 17012 10308 17016 10364
rect 16952 10304 17016 10308
rect 17032 10364 17096 10368
rect 17032 10308 17036 10364
rect 17036 10308 17092 10364
rect 17092 10308 17096 10364
rect 17032 10304 17096 10308
rect 17112 10364 17176 10368
rect 17112 10308 17116 10364
rect 17116 10308 17172 10364
rect 17172 10308 17176 10364
rect 17112 10304 17176 10308
rect 17192 10364 17256 10368
rect 17192 10308 17196 10364
rect 17196 10308 17252 10364
rect 17252 10308 17256 10364
rect 17192 10304 17256 10308
rect 3188 9964 3252 10028
rect 2612 9820 2676 9824
rect 2612 9764 2616 9820
rect 2616 9764 2672 9820
rect 2672 9764 2676 9820
rect 2612 9760 2676 9764
rect 2692 9820 2756 9824
rect 2692 9764 2696 9820
rect 2696 9764 2752 9820
rect 2752 9764 2756 9820
rect 2692 9760 2756 9764
rect 2772 9820 2836 9824
rect 2772 9764 2776 9820
rect 2776 9764 2832 9820
rect 2832 9764 2836 9820
rect 2772 9760 2836 9764
rect 2852 9820 2916 9824
rect 2852 9764 2856 9820
rect 2856 9764 2912 9820
rect 2912 9764 2916 9820
rect 2852 9760 2916 9764
rect 7612 9820 7676 9824
rect 7612 9764 7616 9820
rect 7616 9764 7672 9820
rect 7672 9764 7676 9820
rect 7612 9760 7676 9764
rect 7692 9820 7756 9824
rect 7692 9764 7696 9820
rect 7696 9764 7752 9820
rect 7752 9764 7756 9820
rect 7692 9760 7756 9764
rect 7772 9820 7836 9824
rect 7772 9764 7776 9820
rect 7776 9764 7832 9820
rect 7832 9764 7836 9820
rect 7772 9760 7836 9764
rect 7852 9820 7916 9824
rect 7852 9764 7856 9820
rect 7856 9764 7912 9820
rect 7912 9764 7916 9820
rect 7852 9760 7916 9764
rect 12612 9820 12676 9824
rect 12612 9764 12616 9820
rect 12616 9764 12672 9820
rect 12672 9764 12676 9820
rect 12612 9760 12676 9764
rect 12692 9820 12756 9824
rect 12692 9764 12696 9820
rect 12696 9764 12752 9820
rect 12752 9764 12756 9820
rect 12692 9760 12756 9764
rect 12772 9820 12836 9824
rect 12772 9764 12776 9820
rect 12776 9764 12832 9820
rect 12832 9764 12836 9820
rect 12772 9760 12836 9764
rect 12852 9820 12916 9824
rect 12852 9764 12856 9820
rect 12856 9764 12912 9820
rect 12912 9764 12916 9820
rect 12852 9760 12916 9764
rect 17612 9820 17676 9824
rect 17612 9764 17616 9820
rect 17616 9764 17672 9820
rect 17672 9764 17676 9820
rect 17612 9760 17676 9764
rect 17692 9820 17756 9824
rect 17692 9764 17696 9820
rect 17696 9764 17752 9820
rect 17752 9764 17756 9820
rect 17692 9760 17756 9764
rect 17772 9820 17836 9824
rect 17772 9764 17776 9820
rect 17776 9764 17832 9820
rect 17832 9764 17836 9820
rect 17772 9760 17836 9764
rect 17852 9820 17916 9824
rect 17852 9764 17856 9820
rect 17856 9764 17912 9820
rect 17912 9764 17916 9820
rect 17852 9760 17916 9764
rect 6684 9616 6748 9620
rect 6684 9560 6698 9616
rect 6698 9560 6748 9616
rect 6684 9556 6748 9560
rect 1952 9276 2016 9280
rect 1952 9220 1956 9276
rect 1956 9220 2012 9276
rect 2012 9220 2016 9276
rect 1952 9216 2016 9220
rect 2032 9276 2096 9280
rect 2032 9220 2036 9276
rect 2036 9220 2092 9276
rect 2092 9220 2096 9276
rect 2032 9216 2096 9220
rect 2112 9276 2176 9280
rect 2112 9220 2116 9276
rect 2116 9220 2172 9276
rect 2172 9220 2176 9276
rect 2112 9216 2176 9220
rect 2192 9276 2256 9280
rect 2192 9220 2196 9276
rect 2196 9220 2252 9276
rect 2252 9220 2256 9276
rect 2192 9216 2256 9220
rect 6952 9276 7016 9280
rect 6952 9220 6956 9276
rect 6956 9220 7012 9276
rect 7012 9220 7016 9276
rect 6952 9216 7016 9220
rect 7032 9276 7096 9280
rect 7032 9220 7036 9276
rect 7036 9220 7092 9276
rect 7092 9220 7096 9276
rect 7032 9216 7096 9220
rect 7112 9276 7176 9280
rect 7112 9220 7116 9276
rect 7116 9220 7172 9276
rect 7172 9220 7176 9276
rect 7112 9216 7176 9220
rect 7192 9276 7256 9280
rect 7192 9220 7196 9276
rect 7196 9220 7252 9276
rect 7252 9220 7256 9276
rect 7192 9216 7256 9220
rect 11952 9276 12016 9280
rect 11952 9220 11956 9276
rect 11956 9220 12012 9276
rect 12012 9220 12016 9276
rect 11952 9216 12016 9220
rect 12032 9276 12096 9280
rect 12032 9220 12036 9276
rect 12036 9220 12092 9276
rect 12092 9220 12096 9276
rect 12032 9216 12096 9220
rect 12112 9276 12176 9280
rect 12112 9220 12116 9276
rect 12116 9220 12172 9276
rect 12172 9220 12176 9276
rect 12112 9216 12176 9220
rect 12192 9276 12256 9280
rect 12192 9220 12196 9276
rect 12196 9220 12252 9276
rect 12252 9220 12256 9276
rect 12192 9216 12256 9220
rect 16952 9276 17016 9280
rect 16952 9220 16956 9276
rect 16956 9220 17012 9276
rect 17012 9220 17016 9276
rect 16952 9216 17016 9220
rect 17032 9276 17096 9280
rect 17032 9220 17036 9276
rect 17036 9220 17092 9276
rect 17092 9220 17096 9276
rect 17032 9216 17096 9220
rect 17112 9276 17176 9280
rect 17112 9220 17116 9276
rect 17116 9220 17172 9276
rect 17172 9220 17176 9276
rect 17112 9216 17176 9220
rect 17192 9276 17256 9280
rect 17192 9220 17196 9276
rect 17196 9220 17252 9276
rect 17252 9220 17256 9276
rect 17192 9216 17256 9220
rect 2612 8732 2676 8736
rect 2612 8676 2616 8732
rect 2616 8676 2672 8732
rect 2672 8676 2676 8732
rect 2612 8672 2676 8676
rect 2692 8732 2756 8736
rect 2692 8676 2696 8732
rect 2696 8676 2752 8732
rect 2752 8676 2756 8732
rect 2692 8672 2756 8676
rect 2772 8732 2836 8736
rect 2772 8676 2776 8732
rect 2776 8676 2832 8732
rect 2832 8676 2836 8732
rect 2772 8672 2836 8676
rect 2852 8732 2916 8736
rect 2852 8676 2856 8732
rect 2856 8676 2912 8732
rect 2912 8676 2916 8732
rect 2852 8672 2916 8676
rect 7612 8732 7676 8736
rect 7612 8676 7616 8732
rect 7616 8676 7672 8732
rect 7672 8676 7676 8732
rect 7612 8672 7676 8676
rect 7692 8732 7756 8736
rect 7692 8676 7696 8732
rect 7696 8676 7752 8732
rect 7752 8676 7756 8732
rect 7692 8672 7756 8676
rect 7772 8732 7836 8736
rect 7772 8676 7776 8732
rect 7776 8676 7832 8732
rect 7832 8676 7836 8732
rect 7772 8672 7836 8676
rect 7852 8732 7916 8736
rect 7852 8676 7856 8732
rect 7856 8676 7912 8732
rect 7912 8676 7916 8732
rect 7852 8672 7916 8676
rect 12612 8732 12676 8736
rect 12612 8676 12616 8732
rect 12616 8676 12672 8732
rect 12672 8676 12676 8732
rect 12612 8672 12676 8676
rect 12692 8732 12756 8736
rect 12692 8676 12696 8732
rect 12696 8676 12752 8732
rect 12752 8676 12756 8732
rect 12692 8672 12756 8676
rect 12772 8732 12836 8736
rect 12772 8676 12776 8732
rect 12776 8676 12832 8732
rect 12832 8676 12836 8732
rect 12772 8672 12836 8676
rect 12852 8732 12916 8736
rect 12852 8676 12856 8732
rect 12856 8676 12912 8732
rect 12912 8676 12916 8732
rect 12852 8672 12916 8676
rect 17612 8732 17676 8736
rect 17612 8676 17616 8732
rect 17616 8676 17672 8732
rect 17672 8676 17676 8732
rect 17612 8672 17676 8676
rect 17692 8732 17756 8736
rect 17692 8676 17696 8732
rect 17696 8676 17752 8732
rect 17752 8676 17756 8732
rect 17692 8672 17756 8676
rect 17772 8732 17836 8736
rect 17772 8676 17776 8732
rect 17776 8676 17832 8732
rect 17832 8676 17836 8732
rect 17772 8672 17836 8676
rect 17852 8732 17916 8736
rect 17852 8676 17856 8732
rect 17856 8676 17912 8732
rect 17912 8676 17916 8732
rect 17852 8672 17916 8676
rect 14228 8256 14292 8260
rect 14228 8200 14242 8256
rect 14242 8200 14292 8256
rect 14228 8196 14292 8200
rect 1952 8188 2016 8192
rect 1952 8132 1956 8188
rect 1956 8132 2012 8188
rect 2012 8132 2016 8188
rect 1952 8128 2016 8132
rect 2032 8188 2096 8192
rect 2032 8132 2036 8188
rect 2036 8132 2092 8188
rect 2092 8132 2096 8188
rect 2032 8128 2096 8132
rect 2112 8188 2176 8192
rect 2112 8132 2116 8188
rect 2116 8132 2172 8188
rect 2172 8132 2176 8188
rect 2112 8128 2176 8132
rect 2192 8188 2256 8192
rect 2192 8132 2196 8188
rect 2196 8132 2252 8188
rect 2252 8132 2256 8188
rect 2192 8128 2256 8132
rect 6952 8188 7016 8192
rect 6952 8132 6956 8188
rect 6956 8132 7012 8188
rect 7012 8132 7016 8188
rect 6952 8128 7016 8132
rect 7032 8188 7096 8192
rect 7032 8132 7036 8188
rect 7036 8132 7092 8188
rect 7092 8132 7096 8188
rect 7032 8128 7096 8132
rect 7112 8188 7176 8192
rect 7112 8132 7116 8188
rect 7116 8132 7172 8188
rect 7172 8132 7176 8188
rect 7112 8128 7176 8132
rect 7192 8188 7256 8192
rect 7192 8132 7196 8188
rect 7196 8132 7252 8188
rect 7252 8132 7256 8188
rect 7192 8128 7256 8132
rect 11952 8188 12016 8192
rect 11952 8132 11956 8188
rect 11956 8132 12012 8188
rect 12012 8132 12016 8188
rect 11952 8128 12016 8132
rect 12032 8188 12096 8192
rect 12032 8132 12036 8188
rect 12036 8132 12092 8188
rect 12092 8132 12096 8188
rect 12032 8128 12096 8132
rect 12112 8188 12176 8192
rect 12112 8132 12116 8188
rect 12116 8132 12172 8188
rect 12172 8132 12176 8188
rect 12112 8128 12176 8132
rect 12192 8188 12256 8192
rect 12192 8132 12196 8188
rect 12196 8132 12252 8188
rect 12252 8132 12256 8188
rect 12192 8128 12256 8132
rect 16952 8188 17016 8192
rect 16952 8132 16956 8188
rect 16956 8132 17012 8188
rect 17012 8132 17016 8188
rect 16952 8128 17016 8132
rect 17032 8188 17096 8192
rect 17032 8132 17036 8188
rect 17036 8132 17092 8188
rect 17092 8132 17096 8188
rect 17032 8128 17096 8132
rect 17112 8188 17176 8192
rect 17112 8132 17116 8188
rect 17116 8132 17172 8188
rect 17172 8132 17176 8188
rect 17112 8128 17176 8132
rect 17192 8188 17256 8192
rect 17192 8132 17196 8188
rect 17196 8132 17252 8188
rect 17252 8132 17256 8188
rect 17192 8128 17256 8132
rect 9444 8060 9508 8124
rect 16620 7924 16684 7988
rect 2612 7644 2676 7648
rect 2612 7588 2616 7644
rect 2616 7588 2672 7644
rect 2672 7588 2676 7644
rect 2612 7584 2676 7588
rect 2692 7644 2756 7648
rect 2692 7588 2696 7644
rect 2696 7588 2752 7644
rect 2752 7588 2756 7644
rect 2692 7584 2756 7588
rect 2772 7644 2836 7648
rect 2772 7588 2776 7644
rect 2776 7588 2832 7644
rect 2832 7588 2836 7644
rect 2772 7584 2836 7588
rect 2852 7644 2916 7648
rect 2852 7588 2856 7644
rect 2856 7588 2912 7644
rect 2912 7588 2916 7644
rect 2852 7584 2916 7588
rect 7612 7644 7676 7648
rect 7612 7588 7616 7644
rect 7616 7588 7672 7644
rect 7672 7588 7676 7644
rect 7612 7584 7676 7588
rect 7692 7644 7756 7648
rect 7692 7588 7696 7644
rect 7696 7588 7752 7644
rect 7752 7588 7756 7644
rect 7692 7584 7756 7588
rect 7772 7644 7836 7648
rect 7772 7588 7776 7644
rect 7776 7588 7832 7644
rect 7832 7588 7836 7644
rect 7772 7584 7836 7588
rect 7852 7644 7916 7648
rect 7852 7588 7856 7644
rect 7856 7588 7912 7644
rect 7912 7588 7916 7644
rect 7852 7584 7916 7588
rect 12612 7644 12676 7648
rect 12612 7588 12616 7644
rect 12616 7588 12672 7644
rect 12672 7588 12676 7644
rect 12612 7584 12676 7588
rect 12692 7644 12756 7648
rect 12692 7588 12696 7644
rect 12696 7588 12752 7644
rect 12752 7588 12756 7644
rect 12692 7584 12756 7588
rect 12772 7644 12836 7648
rect 12772 7588 12776 7644
rect 12776 7588 12832 7644
rect 12832 7588 12836 7644
rect 12772 7584 12836 7588
rect 12852 7644 12916 7648
rect 12852 7588 12856 7644
rect 12856 7588 12912 7644
rect 12912 7588 12916 7644
rect 12852 7584 12916 7588
rect 17612 7644 17676 7648
rect 17612 7588 17616 7644
rect 17616 7588 17672 7644
rect 17672 7588 17676 7644
rect 17612 7584 17676 7588
rect 17692 7644 17756 7648
rect 17692 7588 17696 7644
rect 17696 7588 17752 7644
rect 17752 7588 17756 7644
rect 17692 7584 17756 7588
rect 17772 7644 17836 7648
rect 17772 7588 17776 7644
rect 17776 7588 17832 7644
rect 17832 7588 17836 7644
rect 17772 7584 17836 7588
rect 17852 7644 17916 7648
rect 17852 7588 17856 7644
rect 17856 7588 17912 7644
rect 17912 7588 17916 7644
rect 17852 7584 17916 7588
rect 4660 7244 4724 7308
rect 1952 7100 2016 7104
rect 1952 7044 1956 7100
rect 1956 7044 2012 7100
rect 2012 7044 2016 7100
rect 1952 7040 2016 7044
rect 2032 7100 2096 7104
rect 2032 7044 2036 7100
rect 2036 7044 2092 7100
rect 2092 7044 2096 7100
rect 2032 7040 2096 7044
rect 2112 7100 2176 7104
rect 2112 7044 2116 7100
rect 2116 7044 2172 7100
rect 2172 7044 2176 7100
rect 2112 7040 2176 7044
rect 2192 7100 2256 7104
rect 2192 7044 2196 7100
rect 2196 7044 2252 7100
rect 2252 7044 2256 7100
rect 2192 7040 2256 7044
rect 6952 7100 7016 7104
rect 6952 7044 6956 7100
rect 6956 7044 7012 7100
rect 7012 7044 7016 7100
rect 6952 7040 7016 7044
rect 7032 7100 7096 7104
rect 7032 7044 7036 7100
rect 7036 7044 7092 7100
rect 7092 7044 7096 7100
rect 7032 7040 7096 7044
rect 7112 7100 7176 7104
rect 7112 7044 7116 7100
rect 7116 7044 7172 7100
rect 7172 7044 7176 7100
rect 7112 7040 7176 7044
rect 7192 7100 7256 7104
rect 7192 7044 7196 7100
rect 7196 7044 7252 7100
rect 7252 7044 7256 7100
rect 7192 7040 7256 7044
rect 11952 7100 12016 7104
rect 11952 7044 11956 7100
rect 11956 7044 12012 7100
rect 12012 7044 12016 7100
rect 11952 7040 12016 7044
rect 12032 7100 12096 7104
rect 12032 7044 12036 7100
rect 12036 7044 12092 7100
rect 12092 7044 12096 7100
rect 12032 7040 12096 7044
rect 12112 7100 12176 7104
rect 12112 7044 12116 7100
rect 12116 7044 12172 7100
rect 12172 7044 12176 7100
rect 12112 7040 12176 7044
rect 12192 7100 12256 7104
rect 12192 7044 12196 7100
rect 12196 7044 12252 7100
rect 12252 7044 12256 7100
rect 12192 7040 12256 7044
rect 16952 7100 17016 7104
rect 16952 7044 16956 7100
rect 16956 7044 17012 7100
rect 17012 7044 17016 7100
rect 16952 7040 17016 7044
rect 17032 7100 17096 7104
rect 17032 7044 17036 7100
rect 17036 7044 17092 7100
rect 17092 7044 17096 7100
rect 17032 7040 17096 7044
rect 17112 7100 17176 7104
rect 17112 7044 17116 7100
rect 17116 7044 17172 7100
rect 17172 7044 17176 7100
rect 17112 7040 17176 7044
rect 17192 7100 17256 7104
rect 17192 7044 17196 7100
rect 17196 7044 17252 7100
rect 17252 7044 17256 7100
rect 17192 7040 17256 7044
rect 8156 6836 8220 6900
rect 9812 6700 9876 6764
rect 13308 6896 13372 6900
rect 13308 6840 13358 6896
rect 13358 6840 13372 6896
rect 13308 6836 13372 6840
rect 16068 6700 16132 6764
rect 2612 6556 2676 6560
rect 2612 6500 2616 6556
rect 2616 6500 2672 6556
rect 2672 6500 2676 6556
rect 2612 6496 2676 6500
rect 2692 6556 2756 6560
rect 2692 6500 2696 6556
rect 2696 6500 2752 6556
rect 2752 6500 2756 6556
rect 2692 6496 2756 6500
rect 2772 6556 2836 6560
rect 2772 6500 2776 6556
rect 2776 6500 2832 6556
rect 2832 6500 2836 6556
rect 2772 6496 2836 6500
rect 2852 6556 2916 6560
rect 2852 6500 2856 6556
rect 2856 6500 2912 6556
rect 2912 6500 2916 6556
rect 2852 6496 2916 6500
rect 7612 6556 7676 6560
rect 7612 6500 7616 6556
rect 7616 6500 7672 6556
rect 7672 6500 7676 6556
rect 7612 6496 7676 6500
rect 7692 6556 7756 6560
rect 7692 6500 7696 6556
rect 7696 6500 7752 6556
rect 7752 6500 7756 6556
rect 7692 6496 7756 6500
rect 7772 6556 7836 6560
rect 7772 6500 7776 6556
rect 7776 6500 7832 6556
rect 7832 6500 7836 6556
rect 7772 6496 7836 6500
rect 7852 6556 7916 6560
rect 7852 6500 7856 6556
rect 7856 6500 7912 6556
rect 7912 6500 7916 6556
rect 7852 6496 7916 6500
rect 12612 6556 12676 6560
rect 12612 6500 12616 6556
rect 12616 6500 12672 6556
rect 12672 6500 12676 6556
rect 12612 6496 12676 6500
rect 12692 6556 12756 6560
rect 12692 6500 12696 6556
rect 12696 6500 12752 6556
rect 12752 6500 12756 6556
rect 12692 6496 12756 6500
rect 12772 6556 12836 6560
rect 12772 6500 12776 6556
rect 12776 6500 12832 6556
rect 12832 6500 12836 6556
rect 12772 6496 12836 6500
rect 12852 6556 12916 6560
rect 12852 6500 12856 6556
rect 12856 6500 12912 6556
rect 12912 6500 12916 6556
rect 12852 6496 12916 6500
rect 17612 6556 17676 6560
rect 17612 6500 17616 6556
rect 17616 6500 17672 6556
rect 17672 6500 17676 6556
rect 17612 6496 17676 6500
rect 17692 6556 17756 6560
rect 17692 6500 17696 6556
rect 17696 6500 17752 6556
rect 17752 6500 17756 6556
rect 17692 6496 17756 6500
rect 17772 6556 17836 6560
rect 17772 6500 17776 6556
rect 17776 6500 17832 6556
rect 17832 6500 17836 6556
rect 17772 6496 17836 6500
rect 17852 6556 17916 6560
rect 17852 6500 17856 6556
rect 17856 6500 17912 6556
rect 17912 6500 17916 6556
rect 17852 6496 17916 6500
rect 1952 6012 2016 6016
rect 1952 5956 1956 6012
rect 1956 5956 2012 6012
rect 2012 5956 2016 6012
rect 1952 5952 2016 5956
rect 2032 6012 2096 6016
rect 2032 5956 2036 6012
rect 2036 5956 2092 6012
rect 2092 5956 2096 6012
rect 2032 5952 2096 5956
rect 2112 6012 2176 6016
rect 2112 5956 2116 6012
rect 2116 5956 2172 6012
rect 2172 5956 2176 6012
rect 2112 5952 2176 5956
rect 2192 6012 2256 6016
rect 2192 5956 2196 6012
rect 2196 5956 2252 6012
rect 2252 5956 2256 6012
rect 2192 5952 2256 5956
rect 6952 6012 7016 6016
rect 6952 5956 6956 6012
rect 6956 5956 7012 6012
rect 7012 5956 7016 6012
rect 6952 5952 7016 5956
rect 7032 6012 7096 6016
rect 7032 5956 7036 6012
rect 7036 5956 7092 6012
rect 7092 5956 7096 6012
rect 7032 5952 7096 5956
rect 7112 6012 7176 6016
rect 7112 5956 7116 6012
rect 7116 5956 7172 6012
rect 7172 5956 7176 6012
rect 7112 5952 7176 5956
rect 7192 6012 7256 6016
rect 7192 5956 7196 6012
rect 7196 5956 7252 6012
rect 7252 5956 7256 6012
rect 7192 5952 7256 5956
rect 11952 6012 12016 6016
rect 11952 5956 11956 6012
rect 11956 5956 12012 6012
rect 12012 5956 12016 6012
rect 11952 5952 12016 5956
rect 12032 6012 12096 6016
rect 12032 5956 12036 6012
rect 12036 5956 12092 6012
rect 12092 5956 12096 6012
rect 12032 5952 12096 5956
rect 12112 6012 12176 6016
rect 12112 5956 12116 6012
rect 12116 5956 12172 6012
rect 12172 5956 12176 6012
rect 12112 5952 12176 5956
rect 12192 6012 12256 6016
rect 12192 5956 12196 6012
rect 12196 5956 12252 6012
rect 12252 5956 12256 6012
rect 12192 5952 12256 5956
rect 16952 6012 17016 6016
rect 16952 5956 16956 6012
rect 16956 5956 17012 6012
rect 17012 5956 17016 6012
rect 16952 5952 17016 5956
rect 17032 6012 17096 6016
rect 17032 5956 17036 6012
rect 17036 5956 17092 6012
rect 17092 5956 17096 6012
rect 17032 5952 17096 5956
rect 17112 6012 17176 6016
rect 17112 5956 17116 6012
rect 17116 5956 17172 6012
rect 17172 5956 17176 6012
rect 17112 5952 17176 5956
rect 17192 6012 17256 6016
rect 17192 5956 17196 6012
rect 17196 5956 17252 6012
rect 17252 5956 17256 6012
rect 17192 5952 17256 5956
rect 2612 5468 2676 5472
rect 2612 5412 2616 5468
rect 2616 5412 2672 5468
rect 2672 5412 2676 5468
rect 2612 5408 2676 5412
rect 2692 5468 2756 5472
rect 2692 5412 2696 5468
rect 2696 5412 2752 5468
rect 2752 5412 2756 5468
rect 2692 5408 2756 5412
rect 2772 5468 2836 5472
rect 2772 5412 2776 5468
rect 2776 5412 2832 5468
rect 2832 5412 2836 5468
rect 2772 5408 2836 5412
rect 2852 5468 2916 5472
rect 2852 5412 2856 5468
rect 2856 5412 2912 5468
rect 2912 5412 2916 5468
rect 2852 5408 2916 5412
rect 7612 5468 7676 5472
rect 7612 5412 7616 5468
rect 7616 5412 7672 5468
rect 7672 5412 7676 5468
rect 7612 5408 7676 5412
rect 7692 5468 7756 5472
rect 7692 5412 7696 5468
rect 7696 5412 7752 5468
rect 7752 5412 7756 5468
rect 7692 5408 7756 5412
rect 7772 5468 7836 5472
rect 7772 5412 7776 5468
rect 7776 5412 7832 5468
rect 7832 5412 7836 5468
rect 7772 5408 7836 5412
rect 7852 5468 7916 5472
rect 7852 5412 7856 5468
rect 7856 5412 7912 5468
rect 7912 5412 7916 5468
rect 7852 5408 7916 5412
rect 12612 5468 12676 5472
rect 12612 5412 12616 5468
rect 12616 5412 12672 5468
rect 12672 5412 12676 5468
rect 12612 5408 12676 5412
rect 12692 5468 12756 5472
rect 12692 5412 12696 5468
rect 12696 5412 12752 5468
rect 12752 5412 12756 5468
rect 12692 5408 12756 5412
rect 12772 5468 12836 5472
rect 12772 5412 12776 5468
rect 12776 5412 12832 5468
rect 12832 5412 12836 5468
rect 12772 5408 12836 5412
rect 12852 5468 12916 5472
rect 12852 5412 12856 5468
rect 12856 5412 12912 5468
rect 12912 5412 12916 5468
rect 12852 5408 12916 5412
rect 17612 5468 17676 5472
rect 17612 5412 17616 5468
rect 17616 5412 17672 5468
rect 17672 5412 17676 5468
rect 17612 5408 17676 5412
rect 17692 5468 17756 5472
rect 17692 5412 17696 5468
rect 17696 5412 17752 5468
rect 17752 5412 17756 5468
rect 17692 5408 17756 5412
rect 17772 5468 17836 5472
rect 17772 5412 17776 5468
rect 17776 5412 17832 5468
rect 17832 5412 17836 5468
rect 17772 5408 17836 5412
rect 17852 5468 17916 5472
rect 17852 5412 17856 5468
rect 17856 5412 17912 5468
rect 17912 5412 17916 5468
rect 17852 5408 17916 5412
rect 10916 5204 10980 5268
rect 1952 4924 2016 4928
rect 1952 4868 1956 4924
rect 1956 4868 2012 4924
rect 2012 4868 2016 4924
rect 1952 4864 2016 4868
rect 2032 4924 2096 4928
rect 2032 4868 2036 4924
rect 2036 4868 2092 4924
rect 2092 4868 2096 4924
rect 2032 4864 2096 4868
rect 2112 4924 2176 4928
rect 2112 4868 2116 4924
rect 2116 4868 2172 4924
rect 2172 4868 2176 4924
rect 2112 4864 2176 4868
rect 2192 4924 2256 4928
rect 2192 4868 2196 4924
rect 2196 4868 2252 4924
rect 2252 4868 2256 4924
rect 2192 4864 2256 4868
rect 6952 4924 7016 4928
rect 6952 4868 6956 4924
rect 6956 4868 7012 4924
rect 7012 4868 7016 4924
rect 6952 4864 7016 4868
rect 7032 4924 7096 4928
rect 7032 4868 7036 4924
rect 7036 4868 7092 4924
rect 7092 4868 7096 4924
rect 7032 4864 7096 4868
rect 7112 4924 7176 4928
rect 7112 4868 7116 4924
rect 7116 4868 7172 4924
rect 7172 4868 7176 4924
rect 7112 4864 7176 4868
rect 7192 4924 7256 4928
rect 7192 4868 7196 4924
rect 7196 4868 7252 4924
rect 7252 4868 7256 4924
rect 7192 4864 7256 4868
rect 11952 4924 12016 4928
rect 11952 4868 11956 4924
rect 11956 4868 12012 4924
rect 12012 4868 12016 4924
rect 11952 4864 12016 4868
rect 12032 4924 12096 4928
rect 12032 4868 12036 4924
rect 12036 4868 12092 4924
rect 12092 4868 12096 4924
rect 12032 4864 12096 4868
rect 12112 4924 12176 4928
rect 12112 4868 12116 4924
rect 12116 4868 12172 4924
rect 12172 4868 12176 4924
rect 12112 4864 12176 4868
rect 12192 4924 12256 4928
rect 12192 4868 12196 4924
rect 12196 4868 12252 4924
rect 12252 4868 12256 4924
rect 12192 4864 12256 4868
rect 16952 4924 17016 4928
rect 16952 4868 16956 4924
rect 16956 4868 17012 4924
rect 17012 4868 17016 4924
rect 16952 4864 17016 4868
rect 17032 4924 17096 4928
rect 17032 4868 17036 4924
rect 17036 4868 17092 4924
rect 17092 4868 17096 4924
rect 17032 4864 17096 4868
rect 17112 4924 17176 4928
rect 17112 4868 17116 4924
rect 17116 4868 17172 4924
rect 17172 4868 17176 4924
rect 17112 4864 17176 4868
rect 17192 4924 17256 4928
rect 17192 4868 17196 4924
rect 17196 4868 17252 4924
rect 17252 4868 17256 4924
rect 17192 4864 17256 4868
rect 2612 4380 2676 4384
rect 2612 4324 2616 4380
rect 2616 4324 2672 4380
rect 2672 4324 2676 4380
rect 2612 4320 2676 4324
rect 2692 4380 2756 4384
rect 2692 4324 2696 4380
rect 2696 4324 2752 4380
rect 2752 4324 2756 4380
rect 2692 4320 2756 4324
rect 2772 4380 2836 4384
rect 2772 4324 2776 4380
rect 2776 4324 2832 4380
rect 2832 4324 2836 4380
rect 2772 4320 2836 4324
rect 2852 4380 2916 4384
rect 2852 4324 2856 4380
rect 2856 4324 2912 4380
rect 2912 4324 2916 4380
rect 2852 4320 2916 4324
rect 7612 4380 7676 4384
rect 7612 4324 7616 4380
rect 7616 4324 7672 4380
rect 7672 4324 7676 4380
rect 7612 4320 7676 4324
rect 7692 4380 7756 4384
rect 7692 4324 7696 4380
rect 7696 4324 7752 4380
rect 7752 4324 7756 4380
rect 7692 4320 7756 4324
rect 7772 4380 7836 4384
rect 7772 4324 7776 4380
rect 7776 4324 7832 4380
rect 7832 4324 7836 4380
rect 7772 4320 7836 4324
rect 7852 4380 7916 4384
rect 7852 4324 7856 4380
rect 7856 4324 7912 4380
rect 7912 4324 7916 4380
rect 7852 4320 7916 4324
rect 12612 4380 12676 4384
rect 12612 4324 12616 4380
rect 12616 4324 12672 4380
rect 12672 4324 12676 4380
rect 12612 4320 12676 4324
rect 12692 4380 12756 4384
rect 12692 4324 12696 4380
rect 12696 4324 12752 4380
rect 12752 4324 12756 4380
rect 12692 4320 12756 4324
rect 12772 4380 12836 4384
rect 12772 4324 12776 4380
rect 12776 4324 12832 4380
rect 12832 4324 12836 4380
rect 12772 4320 12836 4324
rect 12852 4380 12916 4384
rect 12852 4324 12856 4380
rect 12856 4324 12912 4380
rect 12912 4324 12916 4380
rect 12852 4320 12916 4324
rect 17612 4380 17676 4384
rect 17612 4324 17616 4380
rect 17616 4324 17672 4380
rect 17672 4324 17676 4380
rect 17612 4320 17676 4324
rect 17692 4380 17756 4384
rect 17692 4324 17696 4380
rect 17696 4324 17752 4380
rect 17752 4324 17756 4380
rect 17692 4320 17756 4324
rect 17772 4380 17836 4384
rect 17772 4324 17776 4380
rect 17776 4324 17832 4380
rect 17832 4324 17836 4380
rect 17772 4320 17836 4324
rect 17852 4380 17916 4384
rect 17852 4324 17856 4380
rect 17856 4324 17912 4380
rect 17912 4324 17916 4380
rect 17852 4320 17916 4324
rect 1952 3836 2016 3840
rect 1952 3780 1956 3836
rect 1956 3780 2012 3836
rect 2012 3780 2016 3836
rect 1952 3776 2016 3780
rect 2032 3836 2096 3840
rect 2032 3780 2036 3836
rect 2036 3780 2092 3836
rect 2092 3780 2096 3836
rect 2032 3776 2096 3780
rect 2112 3836 2176 3840
rect 2112 3780 2116 3836
rect 2116 3780 2172 3836
rect 2172 3780 2176 3836
rect 2112 3776 2176 3780
rect 2192 3836 2256 3840
rect 2192 3780 2196 3836
rect 2196 3780 2252 3836
rect 2252 3780 2256 3836
rect 2192 3776 2256 3780
rect 6952 3836 7016 3840
rect 6952 3780 6956 3836
rect 6956 3780 7012 3836
rect 7012 3780 7016 3836
rect 6952 3776 7016 3780
rect 7032 3836 7096 3840
rect 7032 3780 7036 3836
rect 7036 3780 7092 3836
rect 7092 3780 7096 3836
rect 7032 3776 7096 3780
rect 7112 3836 7176 3840
rect 7112 3780 7116 3836
rect 7116 3780 7172 3836
rect 7172 3780 7176 3836
rect 7112 3776 7176 3780
rect 7192 3836 7256 3840
rect 7192 3780 7196 3836
rect 7196 3780 7252 3836
rect 7252 3780 7256 3836
rect 7192 3776 7256 3780
rect 11952 3836 12016 3840
rect 11952 3780 11956 3836
rect 11956 3780 12012 3836
rect 12012 3780 12016 3836
rect 11952 3776 12016 3780
rect 12032 3836 12096 3840
rect 12032 3780 12036 3836
rect 12036 3780 12092 3836
rect 12092 3780 12096 3836
rect 12032 3776 12096 3780
rect 12112 3836 12176 3840
rect 12112 3780 12116 3836
rect 12116 3780 12172 3836
rect 12172 3780 12176 3836
rect 12112 3776 12176 3780
rect 12192 3836 12256 3840
rect 12192 3780 12196 3836
rect 12196 3780 12252 3836
rect 12252 3780 12256 3836
rect 12192 3776 12256 3780
rect 16952 3836 17016 3840
rect 16952 3780 16956 3836
rect 16956 3780 17012 3836
rect 17012 3780 17016 3836
rect 16952 3776 17016 3780
rect 17032 3836 17096 3840
rect 17032 3780 17036 3836
rect 17036 3780 17092 3836
rect 17092 3780 17096 3836
rect 17032 3776 17096 3780
rect 17112 3836 17176 3840
rect 17112 3780 17116 3836
rect 17116 3780 17172 3836
rect 17172 3780 17176 3836
rect 17112 3776 17176 3780
rect 17192 3836 17256 3840
rect 17192 3780 17196 3836
rect 17196 3780 17252 3836
rect 17252 3780 17256 3836
rect 17192 3776 17256 3780
rect 2612 3292 2676 3296
rect 2612 3236 2616 3292
rect 2616 3236 2672 3292
rect 2672 3236 2676 3292
rect 2612 3232 2676 3236
rect 2692 3292 2756 3296
rect 2692 3236 2696 3292
rect 2696 3236 2752 3292
rect 2752 3236 2756 3292
rect 2692 3232 2756 3236
rect 2772 3292 2836 3296
rect 2772 3236 2776 3292
rect 2776 3236 2832 3292
rect 2832 3236 2836 3292
rect 2772 3232 2836 3236
rect 2852 3292 2916 3296
rect 2852 3236 2856 3292
rect 2856 3236 2912 3292
rect 2912 3236 2916 3292
rect 2852 3232 2916 3236
rect 7612 3292 7676 3296
rect 7612 3236 7616 3292
rect 7616 3236 7672 3292
rect 7672 3236 7676 3292
rect 7612 3232 7676 3236
rect 7692 3292 7756 3296
rect 7692 3236 7696 3292
rect 7696 3236 7752 3292
rect 7752 3236 7756 3292
rect 7692 3232 7756 3236
rect 7772 3292 7836 3296
rect 7772 3236 7776 3292
rect 7776 3236 7832 3292
rect 7832 3236 7836 3292
rect 7772 3232 7836 3236
rect 7852 3292 7916 3296
rect 7852 3236 7856 3292
rect 7856 3236 7912 3292
rect 7912 3236 7916 3292
rect 7852 3232 7916 3236
rect 12612 3292 12676 3296
rect 12612 3236 12616 3292
rect 12616 3236 12672 3292
rect 12672 3236 12676 3292
rect 12612 3232 12676 3236
rect 12692 3292 12756 3296
rect 12692 3236 12696 3292
rect 12696 3236 12752 3292
rect 12752 3236 12756 3292
rect 12692 3232 12756 3236
rect 12772 3292 12836 3296
rect 12772 3236 12776 3292
rect 12776 3236 12832 3292
rect 12832 3236 12836 3292
rect 12772 3232 12836 3236
rect 12852 3292 12916 3296
rect 12852 3236 12856 3292
rect 12856 3236 12912 3292
rect 12912 3236 12916 3292
rect 12852 3232 12916 3236
rect 17612 3292 17676 3296
rect 17612 3236 17616 3292
rect 17616 3236 17672 3292
rect 17672 3236 17676 3292
rect 17612 3232 17676 3236
rect 17692 3292 17756 3296
rect 17692 3236 17696 3292
rect 17696 3236 17752 3292
rect 17752 3236 17756 3292
rect 17692 3232 17756 3236
rect 17772 3292 17836 3296
rect 17772 3236 17776 3292
rect 17776 3236 17832 3292
rect 17832 3236 17836 3292
rect 17772 3232 17836 3236
rect 17852 3292 17916 3296
rect 17852 3236 17856 3292
rect 17856 3236 17912 3292
rect 17912 3236 17916 3292
rect 17852 3232 17916 3236
rect 1952 2748 2016 2752
rect 1952 2692 1956 2748
rect 1956 2692 2012 2748
rect 2012 2692 2016 2748
rect 1952 2688 2016 2692
rect 2032 2748 2096 2752
rect 2032 2692 2036 2748
rect 2036 2692 2092 2748
rect 2092 2692 2096 2748
rect 2032 2688 2096 2692
rect 2112 2748 2176 2752
rect 2112 2692 2116 2748
rect 2116 2692 2172 2748
rect 2172 2692 2176 2748
rect 2112 2688 2176 2692
rect 2192 2748 2256 2752
rect 2192 2692 2196 2748
rect 2196 2692 2252 2748
rect 2252 2692 2256 2748
rect 2192 2688 2256 2692
rect 6952 2748 7016 2752
rect 6952 2692 6956 2748
rect 6956 2692 7012 2748
rect 7012 2692 7016 2748
rect 6952 2688 7016 2692
rect 7032 2748 7096 2752
rect 7032 2692 7036 2748
rect 7036 2692 7092 2748
rect 7092 2692 7096 2748
rect 7032 2688 7096 2692
rect 7112 2748 7176 2752
rect 7112 2692 7116 2748
rect 7116 2692 7172 2748
rect 7172 2692 7176 2748
rect 7112 2688 7176 2692
rect 7192 2748 7256 2752
rect 7192 2692 7196 2748
rect 7196 2692 7252 2748
rect 7252 2692 7256 2748
rect 7192 2688 7256 2692
rect 11952 2748 12016 2752
rect 11952 2692 11956 2748
rect 11956 2692 12012 2748
rect 12012 2692 12016 2748
rect 11952 2688 12016 2692
rect 12032 2748 12096 2752
rect 12032 2692 12036 2748
rect 12036 2692 12092 2748
rect 12092 2692 12096 2748
rect 12032 2688 12096 2692
rect 12112 2748 12176 2752
rect 12112 2692 12116 2748
rect 12116 2692 12172 2748
rect 12172 2692 12176 2748
rect 12112 2688 12176 2692
rect 12192 2748 12256 2752
rect 12192 2692 12196 2748
rect 12196 2692 12252 2748
rect 12252 2692 12256 2748
rect 12192 2688 12256 2692
rect 16952 2748 17016 2752
rect 16952 2692 16956 2748
rect 16956 2692 17012 2748
rect 17012 2692 17016 2748
rect 16952 2688 17016 2692
rect 17032 2748 17096 2752
rect 17032 2692 17036 2748
rect 17036 2692 17092 2748
rect 17092 2692 17096 2748
rect 17032 2688 17096 2692
rect 17112 2748 17176 2752
rect 17112 2692 17116 2748
rect 17116 2692 17172 2748
rect 17172 2692 17176 2748
rect 17112 2688 17176 2692
rect 17192 2748 17256 2752
rect 17192 2692 17196 2748
rect 17196 2692 17252 2748
rect 17252 2692 17256 2748
rect 17192 2688 17256 2692
rect 2612 2204 2676 2208
rect 2612 2148 2616 2204
rect 2616 2148 2672 2204
rect 2672 2148 2676 2204
rect 2612 2144 2676 2148
rect 2692 2204 2756 2208
rect 2692 2148 2696 2204
rect 2696 2148 2752 2204
rect 2752 2148 2756 2204
rect 2692 2144 2756 2148
rect 2772 2204 2836 2208
rect 2772 2148 2776 2204
rect 2776 2148 2832 2204
rect 2832 2148 2836 2204
rect 2772 2144 2836 2148
rect 2852 2204 2916 2208
rect 2852 2148 2856 2204
rect 2856 2148 2912 2204
rect 2912 2148 2916 2204
rect 2852 2144 2916 2148
rect 7612 2204 7676 2208
rect 7612 2148 7616 2204
rect 7616 2148 7672 2204
rect 7672 2148 7676 2204
rect 7612 2144 7676 2148
rect 7692 2204 7756 2208
rect 7692 2148 7696 2204
rect 7696 2148 7752 2204
rect 7752 2148 7756 2204
rect 7692 2144 7756 2148
rect 7772 2204 7836 2208
rect 7772 2148 7776 2204
rect 7776 2148 7832 2204
rect 7832 2148 7836 2204
rect 7772 2144 7836 2148
rect 7852 2204 7916 2208
rect 7852 2148 7856 2204
rect 7856 2148 7912 2204
rect 7912 2148 7916 2204
rect 7852 2144 7916 2148
rect 12612 2204 12676 2208
rect 12612 2148 12616 2204
rect 12616 2148 12672 2204
rect 12672 2148 12676 2204
rect 12612 2144 12676 2148
rect 12692 2204 12756 2208
rect 12692 2148 12696 2204
rect 12696 2148 12752 2204
rect 12752 2148 12756 2204
rect 12692 2144 12756 2148
rect 12772 2204 12836 2208
rect 12772 2148 12776 2204
rect 12776 2148 12832 2204
rect 12832 2148 12836 2204
rect 12772 2144 12836 2148
rect 12852 2204 12916 2208
rect 12852 2148 12856 2204
rect 12856 2148 12912 2204
rect 12912 2148 12916 2204
rect 12852 2144 12916 2148
rect 17612 2204 17676 2208
rect 17612 2148 17616 2204
rect 17616 2148 17672 2204
rect 17672 2148 17676 2204
rect 17612 2144 17676 2148
rect 17692 2204 17756 2208
rect 17692 2148 17696 2204
rect 17696 2148 17752 2204
rect 17752 2148 17756 2204
rect 17692 2144 17756 2148
rect 17772 2204 17836 2208
rect 17772 2148 17776 2204
rect 17776 2148 17832 2204
rect 17832 2148 17836 2204
rect 17772 2144 17836 2148
rect 17852 2204 17916 2208
rect 17852 2148 17856 2204
rect 17856 2148 17912 2204
rect 17912 2148 17916 2204
rect 17852 2144 17916 2148
<< metal4 >>
rect 1944 77824 2264 77840
rect 1944 77760 1952 77824
rect 2016 77760 2032 77824
rect 2096 77760 2112 77824
rect 2176 77760 2192 77824
rect 2256 77760 2264 77824
rect 1944 76736 2264 77760
rect 1944 76672 1952 76736
rect 2016 76672 2032 76736
rect 2096 76672 2112 76736
rect 2176 76672 2192 76736
rect 2256 76672 2264 76736
rect 1944 75648 2264 76672
rect 1944 75584 1952 75648
rect 2016 75584 2032 75648
rect 2096 75584 2112 75648
rect 2176 75584 2192 75648
rect 2256 75584 2264 75648
rect 1944 74560 2264 75584
rect 1944 74496 1952 74560
rect 2016 74496 2032 74560
rect 2096 74496 2112 74560
rect 2176 74496 2192 74560
rect 2256 74496 2264 74560
rect 1944 73472 2264 74496
rect 1944 73408 1952 73472
rect 2016 73408 2032 73472
rect 2096 73408 2112 73472
rect 2176 73408 2192 73472
rect 2256 73408 2264 73472
rect 1944 73294 2264 73408
rect 1944 73058 1986 73294
rect 2222 73058 2264 73294
rect 1944 72384 2264 73058
rect 1944 72320 1952 72384
rect 2016 72320 2032 72384
rect 2096 72320 2112 72384
rect 2176 72320 2192 72384
rect 2256 72320 2264 72384
rect 1944 71296 2264 72320
rect 1944 71232 1952 71296
rect 2016 71232 2032 71296
rect 2096 71232 2112 71296
rect 2176 71232 2192 71296
rect 2256 71232 2264 71296
rect 1944 70208 2264 71232
rect 1944 70144 1952 70208
rect 2016 70144 2032 70208
rect 2096 70144 2112 70208
rect 2176 70144 2192 70208
rect 2256 70144 2264 70208
rect 1715 69324 1781 69325
rect 1715 69260 1716 69324
rect 1780 69260 1781 69324
rect 1715 69259 1781 69260
rect 1531 55724 1597 55725
rect 1531 55660 1532 55724
rect 1596 55660 1597 55724
rect 1531 55659 1597 55660
rect 1534 14925 1594 55659
rect 1718 24853 1778 69259
rect 1944 69120 2264 70144
rect 1944 69056 1952 69120
rect 2016 69056 2032 69120
rect 2096 69056 2112 69120
rect 2176 69056 2192 69120
rect 2256 69056 2264 69120
rect 1944 68294 2264 69056
rect 1944 68058 1986 68294
rect 2222 68058 2264 68294
rect 1944 68032 2264 68058
rect 1944 67968 1952 68032
rect 2016 67968 2032 68032
rect 2096 67968 2112 68032
rect 2176 67968 2192 68032
rect 2256 67968 2264 68032
rect 1944 66944 2264 67968
rect 1944 66880 1952 66944
rect 2016 66880 2032 66944
rect 2096 66880 2112 66944
rect 2176 66880 2192 66944
rect 2256 66880 2264 66944
rect 1944 65856 2264 66880
rect 1944 65792 1952 65856
rect 2016 65792 2032 65856
rect 2096 65792 2112 65856
rect 2176 65792 2192 65856
rect 2256 65792 2264 65856
rect 1944 64768 2264 65792
rect 1944 64704 1952 64768
rect 2016 64704 2032 64768
rect 2096 64704 2112 64768
rect 2176 64704 2192 64768
rect 2256 64704 2264 64768
rect 1944 63680 2264 64704
rect 1944 63616 1952 63680
rect 2016 63616 2032 63680
rect 2096 63616 2112 63680
rect 2176 63616 2192 63680
rect 2256 63616 2264 63680
rect 1944 63294 2264 63616
rect 1944 63058 1986 63294
rect 2222 63058 2264 63294
rect 1944 62592 2264 63058
rect 1944 62528 1952 62592
rect 2016 62528 2032 62592
rect 2096 62528 2112 62592
rect 2176 62528 2192 62592
rect 2256 62528 2264 62592
rect 1944 61504 2264 62528
rect 1944 61440 1952 61504
rect 2016 61440 2032 61504
rect 2096 61440 2112 61504
rect 2176 61440 2192 61504
rect 2256 61440 2264 61504
rect 1944 60416 2264 61440
rect 1944 60352 1952 60416
rect 2016 60352 2032 60416
rect 2096 60352 2112 60416
rect 2176 60352 2192 60416
rect 2256 60352 2264 60416
rect 1944 59328 2264 60352
rect 1944 59264 1952 59328
rect 2016 59264 2032 59328
rect 2096 59264 2112 59328
rect 2176 59264 2192 59328
rect 2256 59264 2264 59328
rect 1944 58294 2264 59264
rect 1944 58240 1986 58294
rect 2222 58240 2264 58294
rect 1944 58176 1952 58240
rect 2256 58176 2264 58240
rect 1944 58058 1986 58176
rect 2222 58058 2264 58176
rect 1944 57152 2264 58058
rect 1944 57088 1952 57152
rect 2016 57088 2032 57152
rect 2096 57088 2112 57152
rect 2176 57088 2192 57152
rect 2256 57088 2264 57152
rect 1944 56064 2264 57088
rect 1944 56000 1952 56064
rect 2016 56000 2032 56064
rect 2096 56000 2112 56064
rect 2176 56000 2192 56064
rect 2256 56000 2264 56064
rect 1944 54976 2264 56000
rect 1944 54912 1952 54976
rect 2016 54912 2032 54976
rect 2096 54912 2112 54976
rect 2176 54912 2192 54976
rect 2256 54912 2264 54976
rect 1944 53888 2264 54912
rect 1944 53824 1952 53888
rect 2016 53824 2032 53888
rect 2096 53824 2112 53888
rect 2176 53824 2192 53888
rect 2256 53824 2264 53888
rect 1944 53294 2264 53824
rect 1944 53058 1986 53294
rect 2222 53058 2264 53294
rect 1944 52800 2264 53058
rect 1944 52736 1952 52800
rect 2016 52736 2032 52800
rect 2096 52736 2112 52800
rect 2176 52736 2192 52800
rect 2256 52736 2264 52800
rect 1944 51712 2264 52736
rect 1944 51648 1952 51712
rect 2016 51648 2032 51712
rect 2096 51648 2112 51712
rect 2176 51648 2192 51712
rect 2256 51648 2264 51712
rect 1944 50624 2264 51648
rect 1944 50560 1952 50624
rect 2016 50560 2032 50624
rect 2096 50560 2112 50624
rect 2176 50560 2192 50624
rect 2256 50560 2264 50624
rect 1944 49536 2264 50560
rect 1944 49472 1952 49536
rect 2016 49472 2032 49536
rect 2096 49472 2112 49536
rect 2176 49472 2192 49536
rect 2256 49472 2264 49536
rect 1944 48448 2264 49472
rect 1944 48384 1952 48448
rect 2016 48384 2032 48448
rect 2096 48384 2112 48448
rect 2176 48384 2192 48448
rect 2256 48384 2264 48448
rect 1944 48294 2264 48384
rect 1944 48058 1986 48294
rect 2222 48058 2264 48294
rect 1944 47360 2264 48058
rect 1944 47296 1952 47360
rect 2016 47296 2032 47360
rect 2096 47296 2112 47360
rect 2176 47296 2192 47360
rect 2256 47296 2264 47360
rect 1944 46272 2264 47296
rect 1944 46208 1952 46272
rect 2016 46208 2032 46272
rect 2096 46208 2112 46272
rect 2176 46208 2192 46272
rect 2256 46208 2264 46272
rect 1944 45184 2264 46208
rect 1944 45120 1952 45184
rect 2016 45120 2032 45184
rect 2096 45120 2112 45184
rect 2176 45120 2192 45184
rect 2256 45120 2264 45184
rect 1944 44096 2264 45120
rect 1944 44032 1952 44096
rect 2016 44032 2032 44096
rect 2096 44032 2112 44096
rect 2176 44032 2192 44096
rect 2256 44032 2264 44096
rect 1944 43294 2264 44032
rect 1944 43058 1986 43294
rect 2222 43058 2264 43294
rect 1944 43008 2264 43058
rect 1944 42944 1952 43008
rect 2016 42944 2032 43008
rect 2096 42944 2112 43008
rect 2176 42944 2192 43008
rect 2256 42944 2264 43008
rect 1944 41920 2264 42944
rect 1944 41856 1952 41920
rect 2016 41856 2032 41920
rect 2096 41856 2112 41920
rect 2176 41856 2192 41920
rect 2256 41856 2264 41920
rect 1944 40832 2264 41856
rect 1944 40768 1952 40832
rect 2016 40768 2032 40832
rect 2096 40768 2112 40832
rect 2176 40768 2192 40832
rect 2256 40768 2264 40832
rect 1944 39744 2264 40768
rect 1944 39680 1952 39744
rect 2016 39680 2032 39744
rect 2096 39680 2112 39744
rect 2176 39680 2192 39744
rect 2256 39680 2264 39744
rect 1944 38656 2264 39680
rect 1944 38592 1952 38656
rect 2016 38592 2032 38656
rect 2096 38592 2112 38656
rect 2176 38592 2192 38656
rect 2256 38592 2264 38656
rect 1944 38294 2264 38592
rect 1944 38058 1986 38294
rect 2222 38058 2264 38294
rect 1944 37568 2264 38058
rect 1944 37504 1952 37568
rect 2016 37504 2032 37568
rect 2096 37504 2112 37568
rect 2176 37504 2192 37568
rect 2256 37504 2264 37568
rect 1944 36480 2264 37504
rect 1944 36416 1952 36480
rect 2016 36416 2032 36480
rect 2096 36416 2112 36480
rect 2176 36416 2192 36480
rect 2256 36416 2264 36480
rect 1944 35392 2264 36416
rect 1944 35328 1952 35392
rect 2016 35328 2032 35392
rect 2096 35328 2112 35392
rect 2176 35328 2192 35392
rect 2256 35328 2264 35392
rect 1944 34304 2264 35328
rect 1944 34240 1952 34304
rect 2016 34240 2032 34304
rect 2096 34240 2112 34304
rect 2176 34240 2192 34304
rect 2256 34240 2264 34304
rect 1944 33294 2264 34240
rect 1944 33216 1986 33294
rect 2222 33216 2264 33294
rect 1944 33152 1952 33216
rect 2256 33152 2264 33216
rect 1944 33058 1986 33152
rect 2222 33058 2264 33152
rect 1944 32128 2264 33058
rect 1944 32064 1952 32128
rect 2016 32064 2032 32128
rect 2096 32064 2112 32128
rect 2176 32064 2192 32128
rect 2256 32064 2264 32128
rect 1944 31040 2264 32064
rect 1944 30976 1952 31040
rect 2016 30976 2032 31040
rect 2096 30976 2112 31040
rect 2176 30976 2192 31040
rect 2256 30976 2264 31040
rect 1944 29952 2264 30976
rect 1944 29888 1952 29952
rect 2016 29888 2032 29952
rect 2096 29888 2112 29952
rect 2176 29888 2192 29952
rect 2256 29888 2264 29952
rect 1944 28864 2264 29888
rect 1944 28800 1952 28864
rect 2016 28800 2032 28864
rect 2096 28800 2112 28864
rect 2176 28800 2192 28864
rect 2256 28800 2264 28864
rect 1944 28294 2264 28800
rect 1944 28058 1986 28294
rect 2222 28058 2264 28294
rect 1944 27776 2264 28058
rect 1944 27712 1952 27776
rect 2016 27712 2032 27776
rect 2096 27712 2112 27776
rect 2176 27712 2192 27776
rect 2256 27712 2264 27776
rect 1944 26688 2264 27712
rect 1944 26624 1952 26688
rect 2016 26624 2032 26688
rect 2096 26624 2112 26688
rect 2176 26624 2192 26688
rect 2256 26624 2264 26688
rect 1944 25600 2264 26624
rect 1944 25536 1952 25600
rect 2016 25536 2032 25600
rect 2096 25536 2112 25600
rect 2176 25536 2192 25600
rect 2256 25536 2264 25600
rect 1715 24852 1781 24853
rect 1715 24788 1716 24852
rect 1780 24788 1781 24852
rect 1715 24787 1781 24788
rect 1944 24512 2264 25536
rect 1944 24448 1952 24512
rect 2016 24448 2032 24512
rect 2096 24448 2112 24512
rect 2176 24448 2192 24512
rect 2256 24448 2264 24512
rect 1944 23424 2264 24448
rect 1944 23360 1952 23424
rect 2016 23360 2032 23424
rect 2096 23360 2112 23424
rect 2176 23360 2192 23424
rect 2256 23360 2264 23424
rect 1944 23294 2264 23360
rect 1944 23058 1986 23294
rect 2222 23058 2264 23294
rect 1944 22336 2264 23058
rect 1944 22272 1952 22336
rect 2016 22272 2032 22336
rect 2096 22272 2112 22336
rect 2176 22272 2192 22336
rect 2256 22272 2264 22336
rect 1944 21248 2264 22272
rect 1944 21184 1952 21248
rect 2016 21184 2032 21248
rect 2096 21184 2112 21248
rect 2176 21184 2192 21248
rect 2256 21184 2264 21248
rect 1944 20160 2264 21184
rect 1944 20096 1952 20160
rect 2016 20096 2032 20160
rect 2096 20096 2112 20160
rect 2176 20096 2192 20160
rect 2256 20096 2264 20160
rect 1944 19072 2264 20096
rect 1944 19008 1952 19072
rect 2016 19008 2032 19072
rect 2096 19008 2112 19072
rect 2176 19008 2192 19072
rect 2256 19008 2264 19072
rect 1944 18294 2264 19008
rect 1944 18058 1986 18294
rect 2222 18058 2264 18294
rect 1944 17984 2264 18058
rect 1944 17920 1952 17984
rect 2016 17920 2032 17984
rect 2096 17920 2112 17984
rect 2176 17920 2192 17984
rect 2256 17920 2264 17984
rect 1944 16896 2264 17920
rect 1944 16832 1952 16896
rect 2016 16832 2032 16896
rect 2096 16832 2112 16896
rect 2176 16832 2192 16896
rect 2256 16832 2264 16896
rect 1944 15808 2264 16832
rect 1944 15744 1952 15808
rect 2016 15744 2032 15808
rect 2096 15744 2112 15808
rect 2176 15744 2192 15808
rect 2256 15744 2264 15808
rect 1531 14924 1597 14925
rect 1531 14860 1532 14924
rect 1596 14860 1597 14924
rect 1531 14859 1597 14860
rect 1944 14720 2264 15744
rect 1944 14656 1952 14720
rect 2016 14656 2032 14720
rect 2096 14656 2112 14720
rect 2176 14656 2192 14720
rect 2256 14656 2264 14720
rect 1944 13632 2264 14656
rect 1944 13568 1952 13632
rect 2016 13568 2032 13632
rect 2096 13568 2112 13632
rect 2176 13568 2192 13632
rect 2256 13568 2264 13632
rect 1944 13294 2264 13568
rect 1944 13058 1986 13294
rect 2222 13058 2264 13294
rect 1944 12544 2264 13058
rect 1944 12480 1952 12544
rect 2016 12480 2032 12544
rect 2096 12480 2112 12544
rect 2176 12480 2192 12544
rect 2256 12480 2264 12544
rect 1944 11456 2264 12480
rect 1944 11392 1952 11456
rect 2016 11392 2032 11456
rect 2096 11392 2112 11456
rect 2176 11392 2192 11456
rect 2256 11392 2264 11456
rect 1944 10368 2264 11392
rect 1944 10304 1952 10368
rect 2016 10304 2032 10368
rect 2096 10304 2112 10368
rect 2176 10304 2192 10368
rect 2256 10304 2264 10368
rect 1944 9280 2264 10304
rect 1944 9216 1952 9280
rect 2016 9216 2032 9280
rect 2096 9216 2112 9280
rect 2176 9216 2192 9280
rect 2256 9216 2264 9280
rect 1944 8294 2264 9216
rect 1944 8192 1986 8294
rect 2222 8192 2264 8294
rect 1944 8128 1952 8192
rect 2256 8128 2264 8192
rect 1944 8058 1986 8128
rect 2222 8058 2264 8128
rect 1944 7104 2264 8058
rect 1944 7040 1952 7104
rect 2016 7040 2032 7104
rect 2096 7040 2112 7104
rect 2176 7040 2192 7104
rect 2256 7040 2264 7104
rect 1944 6016 2264 7040
rect 1944 5952 1952 6016
rect 2016 5952 2032 6016
rect 2096 5952 2112 6016
rect 2176 5952 2192 6016
rect 2256 5952 2264 6016
rect 1944 4928 2264 5952
rect 1944 4864 1952 4928
rect 2016 4864 2032 4928
rect 2096 4864 2112 4928
rect 2176 4864 2192 4928
rect 2256 4864 2264 4928
rect 1944 3840 2264 4864
rect 1944 3776 1952 3840
rect 2016 3776 2032 3840
rect 2096 3776 2112 3840
rect 2176 3776 2192 3840
rect 2256 3776 2264 3840
rect 1944 3294 2264 3776
rect 1944 3058 1986 3294
rect 2222 3058 2264 3294
rect 1944 2752 2264 3058
rect 1944 2688 1952 2752
rect 2016 2688 2032 2752
rect 2096 2688 2112 2752
rect 2176 2688 2192 2752
rect 2256 2688 2264 2752
rect 1944 2128 2264 2688
rect 2604 77280 2924 77840
rect 2604 77216 2612 77280
rect 2676 77216 2692 77280
rect 2756 77216 2772 77280
rect 2836 77216 2852 77280
rect 2916 77216 2924 77280
rect 2604 76192 2924 77216
rect 6944 77824 7264 77840
rect 6944 77760 6952 77824
rect 7016 77760 7032 77824
rect 7096 77760 7112 77824
rect 7176 77760 7192 77824
rect 7256 77760 7264 77824
rect 6944 76736 7264 77760
rect 6944 76672 6952 76736
rect 7016 76672 7032 76736
rect 7096 76672 7112 76736
rect 7176 76672 7192 76736
rect 7256 76672 7264 76736
rect 6131 76396 6197 76397
rect 6131 76332 6132 76396
rect 6196 76332 6197 76396
rect 6131 76331 6197 76332
rect 2604 76128 2612 76192
rect 2676 76128 2692 76192
rect 2756 76128 2772 76192
rect 2836 76128 2852 76192
rect 2916 76128 2924 76192
rect 2604 75104 2924 76128
rect 2604 75040 2612 75104
rect 2676 75040 2692 75104
rect 2756 75040 2772 75104
rect 2836 75040 2852 75104
rect 2916 75040 2924 75104
rect 2604 74016 2924 75040
rect 2604 73952 2612 74016
rect 2676 73954 2692 74016
rect 2756 73954 2772 74016
rect 2836 73954 2852 74016
rect 2916 73952 2924 74016
rect 2604 73718 2646 73952
rect 2882 73718 2924 73952
rect 2604 72928 2924 73718
rect 2604 72864 2612 72928
rect 2676 72864 2692 72928
rect 2756 72864 2772 72928
rect 2836 72864 2852 72928
rect 2916 72864 2924 72928
rect 2604 71840 2924 72864
rect 2604 71776 2612 71840
rect 2676 71776 2692 71840
rect 2756 71776 2772 71840
rect 2836 71776 2852 71840
rect 2916 71776 2924 71840
rect 2604 70752 2924 71776
rect 3371 70956 3437 70957
rect 3371 70892 3372 70956
rect 3436 70892 3437 70956
rect 3371 70891 3437 70892
rect 2604 70688 2612 70752
rect 2676 70688 2692 70752
rect 2756 70688 2772 70752
rect 2836 70688 2852 70752
rect 2916 70688 2924 70752
rect 2604 69664 2924 70688
rect 2604 69600 2612 69664
rect 2676 69600 2692 69664
rect 2756 69600 2772 69664
rect 2836 69600 2852 69664
rect 2916 69600 2924 69664
rect 2604 68954 2924 69600
rect 2604 68718 2646 68954
rect 2882 68718 2924 68954
rect 2604 68576 2924 68718
rect 2604 68512 2612 68576
rect 2676 68512 2692 68576
rect 2756 68512 2772 68576
rect 2836 68512 2852 68576
rect 2916 68512 2924 68576
rect 2604 67488 2924 68512
rect 2604 67424 2612 67488
rect 2676 67424 2692 67488
rect 2756 67424 2772 67488
rect 2836 67424 2852 67488
rect 2916 67424 2924 67488
rect 2604 66400 2924 67424
rect 2604 66336 2612 66400
rect 2676 66336 2692 66400
rect 2756 66336 2772 66400
rect 2836 66336 2852 66400
rect 2916 66336 2924 66400
rect 2604 65312 2924 66336
rect 2604 65248 2612 65312
rect 2676 65248 2692 65312
rect 2756 65248 2772 65312
rect 2836 65248 2852 65312
rect 2916 65248 2924 65312
rect 2604 64224 2924 65248
rect 2604 64160 2612 64224
rect 2676 64160 2692 64224
rect 2756 64160 2772 64224
rect 2836 64160 2852 64224
rect 2916 64160 2924 64224
rect 2604 63954 2924 64160
rect 2604 63718 2646 63954
rect 2882 63718 2924 63954
rect 2604 63136 2924 63718
rect 2604 63072 2612 63136
rect 2676 63072 2692 63136
rect 2756 63072 2772 63136
rect 2836 63072 2852 63136
rect 2916 63072 2924 63136
rect 2604 62048 2924 63072
rect 2604 61984 2612 62048
rect 2676 61984 2692 62048
rect 2756 61984 2772 62048
rect 2836 61984 2852 62048
rect 2916 61984 2924 62048
rect 2604 60960 2924 61984
rect 2604 60896 2612 60960
rect 2676 60896 2692 60960
rect 2756 60896 2772 60960
rect 2836 60896 2852 60960
rect 2916 60896 2924 60960
rect 2604 59872 2924 60896
rect 2604 59808 2612 59872
rect 2676 59808 2692 59872
rect 2756 59808 2772 59872
rect 2836 59808 2852 59872
rect 2916 59808 2924 59872
rect 2604 58954 2924 59808
rect 2604 58784 2646 58954
rect 2882 58784 2924 58954
rect 2604 58720 2612 58784
rect 2916 58720 2924 58784
rect 2604 58718 2646 58720
rect 2882 58718 2924 58720
rect 2604 57696 2924 58718
rect 2604 57632 2612 57696
rect 2676 57632 2692 57696
rect 2756 57632 2772 57696
rect 2836 57632 2852 57696
rect 2916 57632 2924 57696
rect 2604 56608 2924 57632
rect 2604 56544 2612 56608
rect 2676 56544 2692 56608
rect 2756 56544 2772 56608
rect 2836 56544 2852 56608
rect 2916 56544 2924 56608
rect 2604 55520 2924 56544
rect 2604 55456 2612 55520
rect 2676 55456 2692 55520
rect 2756 55456 2772 55520
rect 2836 55456 2852 55520
rect 2916 55456 2924 55520
rect 2604 54432 2924 55456
rect 2604 54368 2612 54432
rect 2676 54368 2692 54432
rect 2756 54368 2772 54432
rect 2836 54368 2852 54432
rect 2916 54368 2924 54432
rect 2604 53954 2924 54368
rect 2604 53718 2646 53954
rect 2882 53718 2924 53954
rect 2604 53344 2924 53718
rect 2604 53280 2612 53344
rect 2676 53280 2692 53344
rect 2756 53280 2772 53344
rect 2836 53280 2852 53344
rect 2916 53280 2924 53344
rect 2604 52256 2924 53280
rect 2604 52192 2612 52256
rect 2676 52192 2692 52256
rect 2756 52192 2772 52256
rect 2836 52192 2852 52256
rect 2916 52192 2924 52256
rect 2604 51168 2924 52192
rect 2604 51104 2612 51168
rect 2676 51104 2692 51168
rect 2756 51104 2772 51168
rect 2836 51104 2852 51168
rect 2916 51104 2924 51168
rect 2604 50080 2924 51104
rect 2604 50016 2612 50080
rect 2676 50016 2692 50080
rect 2756 50016 2772 50080
rect 2836 50016 2852 50080
rect 2916 50016 2924 50080
rect 2604 48992 2924 50016
rect 2604 48928 2612 48992
rect 2676 48954 2692 48992
rect 2756 48954 2772 48992
rect 2836 48954 2852 48992
rect 2916 48928 2924 48992
rect 2604 48718 2646 48928
rect 2882 48718 2924 48928
rect 2604 47904 2924 48718
rect 2604 47840 2612 47904
rect 2676 47840 2692 47904
rect 2756 47840 2772 47904
rect 2836 47840 2852 47904
rect 2916 47840 2924 47904
rect 2604 46816 2924 47840
rect 3187 47292 3253 47293
rect 3187 47228 3188 47292
rect 3252 47228 3253 47292
rect 3187 47227 3253 47228
rect 2604 46752 2612 46816
rect 2676 46752 2692 46816
rect 2756 46752 2772 46816
rect 2836 46752 2852 46816
rect 2916 46752 2924 46816
rect 2604 45728 2924 46752
rect 2604 45664 2612 45728
rect 2676 45664 2692 45728
rect 2756 45664 2772 45728
rect 2836 45664 2852 45728
rect 2916 45664 2924 45728
rect 2604 44640 2924 45664
rect 2604 44576 2612 44640
rect 2676 44576 2692 44640
rect 2756 44576 2772 44640
rect 2836 44576 2852 44640
rect 2916 44576 2924 44640
rect 2604 43954 2924 44576
rect 2604 43718 2646 43954
rect 2882 43718 2924 43954
rect 2604 43552 2924 43718
rect 2604 43488 2612 43552
rect 2676 43488 2692 43552
rect 2756 43488 2772 43552
rect 2836 43488 2852 43552
rect 2916 43488 2924 43552
rect 2604 42464 2924 43488
rect 2604 42400 2612 42464
rect 2676 42400 2692 42464
rect 2756 42400 2772 42464
rect 2836 42400 2852 42464
rect 2916 42400 2924 42464
rect 2604 41376 2924 42400
rect 2604 41312 2612 41376
rect 2676 41312 2692 41376
rect 2756 41312 2772 41376
rect 2836 41312 2852 41376
rect 2916 41312 2924 41376
rect 2604 40288 2924 41312
rect 2604 40224 2612 40288
rect 2676 40224 2692 40288
rect 2756 40224 2772 40288
rect 2836 40224 2852 40288
rect 2916 40224 2924 40288
rect 2604 39200 2924 40224
rect 2604 39136 2612 39200
rect 2676 39136 2692 39200
rect 2756 39136 2772 39200
rect 2836 39136 2852 39200
rect 2916 39136 2924 39200
rect 2604 38954 2924 39136
rect 2604 38718 2646 38954
rect 2882 38718 2924 38954
rect 2604 38112 2924 38718
rect 2604 38048 2612 38112
rect 2676 38048 2692 38112
rect 2756 38048 2772 38112
rect 2836 38048 2852 38112
rect 2916 38048 2924 38112
rect 2604 37024 2924 38048
rect 2604 36960 2612 37024
rect 2676 36960 2692 37024
rect 2756 36960 2772 37024
rect 2836 36960 2852 37024
rect 2916 36960 2924 37024
rect 2604 35936 2924 36960
rect 2604 35872 2612 35936
rect 2676 35872 2692 35936
rect 2756 35872 2772 35936
rect 2836 35872 2852 35936
rect 2916 35872 2924 35936
rect 2604 34848 2924 35872
rect 2604 34784 2612 34848
rect 2676 34784 2692 34848
rect 2756 34784 2772 34848
rect 2836 34784 2852 34848
rect 2916 34784 2924 34848
rect 2604 33954 2924 34784
rect 2604 33760 2646 33954
rect 2882 33760 2924 33954
rect 2604 33696 2612 33760
rect 2676 33696 2692 33718
rect 2756 33696 2772 33718
rect 2836 33696 2852 33718
rect 2916 33696 2924 33760
rect 2604 32672 2924 33696
rect 2604 32608 2612 32672
rect 2676 32608 2692 32672
rect 2756 32608 2772 32672
rect 2836 32608 2852 32672
rect 2916 32608 2924 32672
rect 2604 31584 2924 32608
rect 2604 31520 2612 31584
rect 2676 31520 2692 31584
rect 2756 31520 2772 31584
rect 2836 31520 2852 31584
rect 2916 31520 2924 31584
rect 2604 30496 2924 31520
rect 2604 30432 2612 30496
rect 2676 30432 2692 30496
rect 2756 30432 2772 30496
rect 2836 30432 2852 30496
rect 2916 30432 2924 30496
rect 2604 29408 2924 30432
rect 2604 29344 2612 29408
rect 2676 29344 2692 29408
rect 2756 29344 2772 29408
rect 2836 29344 2852 29408
rect 2916 29344 2924 29408
rect 2604 28954 2924 29344
rect 2604 28718 2646 28954
rect 2882 28718 2924 28954
rect 2604 28320 2924 28718
rect 2604 28256 2612 28320
rect 2676 28256 2692 28320
rect 2756 28256 2772 28320
rect 2836 28256 2852 28320
rect 2916 28256 2924 28320
rect 2604 27232 2924 28256
rect 2604 27168 2612 27232
rect 2676 27168 2692 27232
rect 2756 27168 2772 27232
rect 2836 27168 2852 27232
rect 2916 27168 2924 27232
rect 2604 26144 2924 27168
rect 2604 26080 2612 26144
rect 2676 26080 2692 26144
rect 2756 26080 2772 26144
rect 2836 26080 2852 26144
rect 2916 26080 2924 26144
rect 2604 25056 2924 26080
rect 2604 24992 2612 25056
rect 2676 24992 2692 25056
rect 2756 24992 2772 25056
rect 2836 24992 2852 25056
rect 2916 24992 2924 25056
rect 2604 23968 2924 24992
rect 2604 23904 2612 23968
rect 2676 23954 2692 23968
rect 2756 23954 2772 23968
rect 2836 23954 2852 23968
rect 2916 23904 2924 23968
rect 2604 23718 2646 23904
rect 2882 23718 2924 23904
rect 2604 22880 2924 23718
rect 2604 22816 2612 22880
rect 2676 22816 2692 22880
rect 2756 22816 2772 22880
rect 2836 22816 2852 22880
rect 2916 22816 2924 22880
rect 2604 21792 2924 22816
rect 2604 21728 2612 21792
rect 2676 21728 2692 21792
rect 2756 21728 2772 21792
rect 2836 21728 2852 21792
rect 2916 21728 2924 21792
rect 2604 20704 2924 21728
rect 2604 20640 2612 20704
rect 2676 20640 2692 20704
rect 2756 20640 2772 20704
rect 2836 20640 2852 20704
rect 2916 20640 2924 20704
rect 2604 19616 2924 20640
rect 2604 19552 2612 19616
rect 2676 19552 2692 19616
rect 2756 19552 2772 19616
rect 2836 19552 2852 19616
rect 2916 19552 2924 19616
rect 2604 18954 2924 19552
rect 2604 18718 2646 18954
rect 2882 18718 2924 18954
rect 2604 18528 2924 18718
rect 2604 18464 2612 18528
rect 2676 18464 2692 18528
rect 2756 18464 2772 18528
rect 2836 18464 2852 18528
rect 2916 18464 2924 18528
rect 2604 17440 2924 18464
rect 2604 17376 2612 17440
rect 2676 17376 2692 17440
rect 2756 17376 2772 17440
rect 2836 17376 2852 17440
rect 2916 17376 2924 17440
rect 2604 16352 2924 17376
rect 2604 16288 2612 16352
rect 2676 16288 2692 16352
rect 2756 16288 2772 16352
rect 2836 16288 2852 16352
rect 2916 16288 2924 16352
rect 2604 15264 2924 16288
rect 2604 15200 2612 15264
rect 2676 15200 2692 15264
rect 2756 15200 2772 15264
rect 2836 15200 2852 15264
rect 2916 15200 2924 15264
rect 2604 14176 2924 15200
rect 2604 14112 2612 14176
rect 2676 14112 2692 14176
rect 2756 14112 2772 14176
rect 2836 14112 2852 14176
rect 2916 14112 2924 14176
rect 2604 13954 2924 14112
rect 2604 13718 2646 13954
rect 2882 13718 2924 13954
rect 2604 13088 2924 13718
rect 2604 13024 2612 13088
rect 2676 13024 2692 13088
rect 2756 13024 2772 13088
rect 2836 13024 2852 13088
rect 2916 13024 2924 13088
rect 2604 12000 2924 13024
rect 2604 11936 2612 12000
rect 2676 11936 2692 12000
rect 2756 11936 2772 12000
rect 2836 11936 2852 12000
rect 2916 11936 2924 12000
rect 2604 10912 2924 11936
rect 2604 10848 2612 10912
rect 2676 10848 2692 10912
rect 2756 10848 2772 10912
rect 2836 10848 2852 10912
rect 2916 10848 2924 10912
rect 2604 9824 2924 10848
rect 3190 10029 3250 47227
rect 3374 35597 3434 70891
rect 3923 65244 3989 65245
rect 3923 65180 3924 65244
rect 3988 65180 3989 65244
rect 3923 65179 3989 65180
rect 3371 35596 3437 35597
rect 3371 35532 3372 35596
rect 3436 35532 3437 35596
rect 3371 35531 3437 35532
rect 3926 15061 3986 65179
rect 4843 63340 4909 63341
rect 4843 63276 4844 63340
rect 4908 63276 4909 63340
rect 4843 63275 4909 63276
rect 4291 62252 4357 62253
rect 4291 62188 4292 62252
rect 4356 62188 4357 62252
rect 4291 62187 4357 62188
rect 4294 23629 4354 62187
rect 4475 49740 4541 49741
rect 4475 49676 4476 49740
rect 4540 49676 4541 49740
rect 4475 49675 4541 49676
rect 4291 23628 4357 23629
rect 4291 23564 4292 23628
rect 4356 23564 4357 23628
rect 4291 23563 4357 23564
rect 4478 21997 4538 49675
rect 4659 48244 4725 48245
rect 4659 48180 4660 48244
rect 4724 48180 4725 48244
rect 4659 48179 4725 48180
rect 4475 21996 4541 21997
rect 4475 21932 4476 21996
rect 4540 21932 4541 21996
rect 4475 21931 4541 21932
rect 4478 20773 4538 21931
rect 4475 20772 4541 20773
rect 4475 20708 4476 20772
rect 4540 20708 4541 20772
rect 4475 20707 4541 20708
rect 3923 15060 3989 15061
rect 3923 14996 3924 15060
rect 3988 14996 3989 15060
rect 3923 14995 3989 14996
rect 3187 10028 3253 10029
rect 3187 9964 3188 10028
rect 3252 9964 3253 10028
rect 3187 9963 3253 9964
rect 2604 9760 2612 9824
rect 2676 9760 2692 9824
rect 2756 9760 2772 9824
rect 2836 9760 2852 9824
rect 2916 9760 2924 9824
rect 2604 8954 2924 9760
rect 2604 8736 2646 8954
rect 2882 8736 2924 8954
rect 2604 8672 2612 8736
rect 2676 8672 2692 8718
rect 2756 8672 2772 8718
rect 2836 8672 2852 8718
rect 2916 8672 2924 8736
rect 2604 7648 2924 8672
rect 2604 7584 2612 7648
rect 2676 7584 2692 7648
rect 2756 7584 2772 7648
rect 2836 7584 2852 7648
rect 2916 7584 2924 7648
rect 2604 6560 2924 7584
rect 4662 7309 4722 48179
rect 4846 31789 4906 63275
rect 4843 31788 4909 31789
rect 4843 31724 4844 31788
rect 4908 31724 4909 31788
rect 4843 31723 4909 31724
rect 6134 10709 6194 76331
rect 6944 75648 7264 76672
rect 6944 75584 6952 75648
rect 7016 75584 7032 75648
rect 7096 75584 7112 75648
rect 7176 75584 7192 75648
rect 7256 75584 7264 75648
rect 6683 75172 6749 75173
rect 6683 75108 6684 75172
rect 6748 75108 6749 75172
rect 6683 75107 6749 75108
rect 6315 56676 6381 56677
rect 6315 56612 6316 56676
rect 6380 56612 6381 56676
rect 6315 56611 6381 56612
rect 6318 16693 6378 56611
rect 6499 42940 6565 42941
rect 6499 42876 6500 42940
rect 6564 42876 6565 42940
rect 6499 42875 6565 42876
rect 6502 19957 6562 42875
rect 6499 19956 6565 19957
rect 6499 19892 6500 19956
rect 6564 19892 6565 19956
rect 6499 19891 6565 19892
rect 6315 16692 6381 16693
rect 6315 16628 6316 16692
rect 6380 16628 6381 16692
rect 6315 16627 6381 16628
rect 6131 10708 6197 10709
rect 6131 10644 6132 10708
rect 6196 10644 6197 10708
rect 6131 10643 6197 10644
rect 6686 9621 6746 75107
rect 6944 74560 7264 75584
rect 6944 74496 6952 74560
rect 7016 74496 7032 74560
rect 7096 74496 7112 74560
rect 7176 74496 7192 74560
rect 7256 74496 7264 74560
rect 6944 73472 7264 74496
rect 6944 73408 6952 73472
rect 7016 73408 7032 73472
rect 7096 73408 7112 73472
rect 7176 73408 7192 73472
rect 7256 73408 7264 73472
rect 6944 73294 7264 73408
rect 6944 73058 6986 73294
rect 7222 73058 7264 73294
rect 6944 72384 7264 73058
rect 6944 72320 6952 72384
rect 7016 72320 7032 72384
rect 7096 72320 7112 72384
rect 7176 72320 7192 72384
rect 7256 72320 7264 72384
rect 6944 71296 7264 72320
rect 6944 71232 6952 71296
rect 7016 71232 7032 71296
rect 7096 71232 7112 71296
rect 7176 71232 7192 71296
rect 7256 71232 7264 71296
rect 6944 70208 7264 71232
rect 6944 70144 6952 70208
rect 7016 70144 7032 70208
rect 7096 70144 7112 70208
rect 7176 70144 7192 70208
rect 7256 70144 7264 70208
rect 6944 69120 7264 70144
rect 6944 69056 6952 69120
rect 7016 69056 7032 69120
rect 7096 69056 7112 69120
rect 7176 69056 7192 69120
rect 7256 69056 7264 69120
rect 6944 68294 7264 69056
rect 6944 68058 6986 68294
rect 7222 68058 7264 68294
rect 6944 68032 7264 68058
rect 6944 67968 6952 68032
rect 7016 67968 7032 68032
rect 7096 67968 7112 68032
rect 7176 67968 7192 68032
rect 7256 67968 7264 68032
rect 6944 66944 7264 67968
rect 6944 66880 6952 66944
rect 7016 66880 7032 66944
rect 7096 66880 7112 66944
rect 7176 66880 7192 66944
rect 7256 66880 7264 66944
rect 6944 65856 7264 66880
rect 6944 65792 6952 65856
rect 7016 65792 7032 65856
rect 7096 65792 7112 65856
rect 7176 65792 7192 65856
rect 7256 65792 7264 65856
rect 6944 64768 7264 65792
rect 6944 64704 6952 64768
rect 7016 64704 7032 64768
rect 7096 64704 7112 64768
rect 7176 64704 7192 64768
rect 7256 64704 7264 64768
rect 6944 63680 7264 64704
rect 6944 63616 6952 63680
rect 7016 63616 7032 63680
rect 7096 63616 7112 63680
rect 7176 63616 7192 63680
rect 7256 63616 7264 63680
rect 6944 63294 7264 63616
rect 6944 63058 6986 63294
rect 7222 63058 7264 63294
rect 6944 62592 7264 63058
rect 6944 62528 6952 62592
rect 7016 62528 7032 62592
rect 7096 62528 7112 62592
rect 7176 62528 7192 62592
rect 7256 62528 7264 62592
rect 6944 61504 7264 62528
rect 6944 61440 6952 61504
rect 7016 61440 7032 61504
rect 7096 61440 7112 61504
rect 7176 61440 7192 61504
rect 7256 61440 7264 61504
rect 6944 60416 7264 61440
rect 6944 60352 6952 60416
rect 7016 60352 7032 60416
rect 7096 60352 7112 60416
rect 7176 60352 7192 60416
rect 7256 60352 7264 60416
rect 6944 59328 7264 60352
rect 6944 59264 6952 59328
rect 7016 59264 7032 59328
rect 7096 59264 7112 59328
rect 7176 59264 7192 59328
rect 7256 59264 7264 59328
rect 6944 58294 7264 59264
rect 6944 58240 6986 58294
rect 7222 58240 7264 58294
rect 6944 58176 6952 58240
rect 7256 58176 7264 58240
rect 6944 58058 6986 58176
rect 7222 58058 7264 58176
rect 6944 57152 7264 58058
rect 6944 57088 6952 57152
rect 7016 57088 7032 57152
rect 7096 57088 7112 57152
rect 7176 57088 7192 57152
rect 7256 57088 7264 57152
rect 6944 56064 7264 57088
rect 6944 56000 6952 56064
rect 7016 56000 7032 56064
rect 7096 56000 7112 56064
rect 7176 56000 7192 56064
rect 7256 56000 7264 56064
rect 6944 54976 7264 56000
rect 6944 54912 6952 54976
rect 7016 54912 7032 54976
rect 7096 54912 7112 54976
rect 7176 54912 7192 54976
rect 7256 54912 7264 54976
rect 6944 53888 7264 54912
rect 6944 53824 6952 53888
rect 7016 53824 7032 53888
rect 7096 53824 7112 53888
rect 7176 53824 7192 53888
rect 7256 53824 7264 53888
rect 6944 53294 7264 53824
rect 6944 53058 6986 53294
rect 7222 53058 7264 53294
rect 6944 52800 7264 53058
rect 6944 52736 6952 52800
rect 7016 52736 7032 52800
rect 7096 52736 7112 52800
rect 7176 52736 7192 52800
rect 7256 52736 7264 52800
rect 6944 51712 7264 52736
rect 6944 51648 6952 51712
rect 7016 51648 7032 51712
rect 7096 51648 7112 51712
rect 7176 51648 7192 51712
rect 7256 51648 7264 51712
rect 6944 50624 7264 51648
rect 7604 77280 7924 77840
rect 7604 77216 7612 77280
rect 7676 77216 7692 77280
rect 7756 77216 7772 77280
rect 7836 77216 7852 77280
rect 7916 77216 7924 77280
rect 7604 76192 7924 77216
rect 11944 77824 12264 77840
rect 11944 77760 11952 77824
rect 12016 77760 12032 77824
rect 12096 77760 12112 77824
rect 12176 77760 12192 77824
rect 12256 77760 12264 77824
rect 11944 76736 12264 77760
rect 11944 76672 11952 76736
rect 12016 76672 12032 76736
rect 12096 76672 12112 76736
rect 12176 76672 12192 76736
rect 12256 76672 12264 76736
rect 11283 76260 11349 76261
rect 11283 76196 11284 76260
rect 11348 76196 11349 76260
rect 11283 76195 11349 76196
rect 7604 76128 7612 76192
rect 7676 76128 7692 76192
rect 7756 76128 7772 76192
rect 7836 76128 7852 76192
rect 7916 76128 7924 76192
rect 7604 75104 7924 76128
rect 8891 76124 8957 76125
rect 8891 76060 8892 76124
rect 8956 76060 8957 76124
rect 8891 76059 8957 76060
rect 7604 75040 7612 75104
rect 7676 75040 7692 75104
rect 7756 75040 7772 75104
rect 7836 75040 7852 75104
rect 7916 75040 7924 75104
rect 7604 74016 7924 75040
rect 7604 73952 7612 74016
rect 7676 73954 7692 74016
rect 7756 73954 7772 74016
rect 7836 73954 7852 74016
rect 7916 73952 7924 74016
rect 7604 73718 7646 73952
rect 7882 73718 7924 73952
rect 7604 72928 7924 73718
rect 7604 72864 7612 72928
rect 7676 72864 7692 72928
rect 7756 72864 7772 72928
rect 7836 72864 7852 72928
rect 7916 72864 7924 72928
rect 7604 71840 7924 72864
rect 7604 71776 7612 71840
rect 7676 71776 7692 71840
rect 7756 71776 7772 71840
rect 7836 71776 7852 71840
rect 7916 71776 7924 71840
rect 7604 70752 7924 71776
rect 7604 70688 7612 70752
rect 7676 70688 7692 70752
rect 7756 70688 7772 70752
rect 7836 70688 7852 70752
rect 7916 70688 7924 70752
rect 7604 69664 7924 70688
rect 7604 69600 7612 69664
rect 7676 69600 7692 69664
rect 7756 69600 7772 69664
rect 7836 69600 7852 69664
rect 7916 69600 7924 69664
rect 7604 68954 7924 69600
rect 7604 68718 7646 68954
rect 7882 68718 7924 68954
rect 7604 68576 7924 68718
rect 7604 68512 7612 68576
rect 7676 68512 7692 68576
rect 7756 68512 7772 68576
rect 7836 68512 7852 68576
rect 7916 68512 7924 68576
rect 7604 67488 7924 68512
rect 7604 67424 7612 67488
rect 7676 67424 7692 67488
rect 7756 67424 7772 67488
rect 7836 67424 7852 67488
rect 7916 67424 7924 67488
rect 7604 66400 7924 67424
rect 7604 66336 7612 66400
rect 7676 66336 7692 66400
rect 7756 66336 7772 66400
rect 7836 66336 7852 66400
rect 7916 66336 7924 66400
rect 7604 65312 7924 66336
rect 7604 65248 7612 65312
rect 7676 65248 7692 65312
rect 7756 65248 7772 65312
rect 7836 65248 7852 65312
rect 7916 65248 7924 65312
rect 7604 64224 7924 65248
rect 7604 64160 7612 64224
rect 7676 64160 7692 64224
rect 7756 64160 7772 64224
rect 7836 64160 7852 64224
rect 7916 64160 7924 64224
rect 7604 63954 7924 64160
rect 7604 63718 7646 63954
rect 7882 63718 7924 63954
rect 7604 63136 7924 63718
rect 7604 63072 7612 63136
rect 7676 63072 7692 63136
rect 7756 63072 7772 63136
rect 7836 63072 7852 63136
rect 7916 63072 7924 63136
rect 7604 62048 7924 63072
rect 8707 62660 8773 62661
rect 8707 62596 8708 62660
rect 8772 62596 8773 62660
rect 8707 62595 8773 62596
rect 7604 61984 7612 62048
rect 7676 61984 7692 62048
rect 7756 61984 7772 62048
rect 7836 61984 7852 62048
rect 7916 61984 7924 62048
rect 7604 60960 7924 61984
rect 7604 60896 7612 60960
rect 7676 60896 7692 60960
rect 7756 60896 7772 60960
rect 7836 60896 7852 60960
rect 7916 60896 7924 60960
rect 7604 59872 7924 60896
rect 7604 59808 7612 59872
rect 7676 59808 7692 59872
rect 7756 59808 7772 59872
rect 7836 59808 7852 59872
rect 7916 59808 7924 59872
rect 7604 58954 7924 59808
rect 7604 58784 7646 58954
rect 7882 58784 7924 58954
rect 7604 58720 7612 58784
rect 7916 58720 7924 58784
rect 7604 58718 7646 58720
rect 7882 58718 7924 58720
rect 7604 57696 7924 58718
rect 7604 57632 7612 57696
rect 7676 57632 7692 57696
rect 7756 57632 7772 57696
rect 7836 57632 7852 57696
rect 7916 57632 7924 57696
rect 7604 56608 7924 57632
rect 7604 56544 7612 56608
rect 7676 56544 7692 56608
rect 7756 56544 7772 56608
rect 7836 56544 7852 56608
rect 7916 56544 7924 56608
rect 7604 55520 7924 56544
rect 7604 55456 7612 55520
rect 7676 55456 7692 55520
rect 7756 55456 7772 55520
rect 7836 55456 7852 55520
rect 7916 55456 7924 55520
rect 7604 54432 7924 55456
rect 7604 54368 7612 54432
rect 7676 54368 7692 54432
rect 7756 54368 7772 54432
rect 7836 54368 7852 54432
rect 7916 54368 7924 54432
rect 7604 53954 7924 54368
rect 7604 53718 7646 53954
rect 7882 53718 7924 53954
rect 7604 53344 7924 53718
rect 7604 53280 7612 53344
rect 7676 53280 7692 53344
rect 7756 53280 7772 53344
rect 7836 53280 7852 53344
rect 7916 53280 7924 53344
rect 7604 52256 7924 53280
rect 8523 52596 8589 52597
rect 8523 52532 8524 52596
rect 8588 52532 8589 52596
rect 8523 52531 8589 52532
rect 7604 52192 7612 52256
rect 7676 52192 7692 52256
rect 7756 52192 7772 52256
rect 7836 52192 7852 52256
rect 7916 52192 7924 52256
rect 7604 51168 7924 52192
rect 8155 51916 8221 51917
rect 8155 51852 8156 51916
rect 8220 51852 8221 51916
rect 8155 51851 8221 51852
rect 7604 51104 7612 51168
rect 7676 51104 7692 51168
rect 7756 51104 7772 51168
rect 7836 51104 7852 51168
rect 7916 51104 7924 51168
rect 7419 50828 7485 50829
rect 7419 50764 7420 50828
rect 7484 50764 7485 50828
rect 7419 50763 7485 50764
rect 6944 50560 6952 50624
rect 7016 50560 7032 50624
rect 7096 50560 7112 50624
rect 7176 50560 7192 50624
rect 7256 50560 7264 50624
rect 6944 49536 7264 50560
rect 6944 49472 6952 49536
rect 7016 49472 7032 49536
rect 7096 49472 7112 49536
rect 7176 49472 7192 49536
rect 7256 49472 7264 49536
rect 6944 48448 7264 49472
rect 6944 48384 6952 48448
rect 7016 48384 7032 48448
rect 7096 48384 7112 48448
rect 7176 48384 7192 48448
rect 7256 48384 7264 48448
rect 6944 48294 7264 48384
rect 6944 48058 6986 48294
rect 7222 48058 7264 48294
rect 6944 47360 7264 48058
rect 6944 47296 6952 47360
rect 7016 47296 7032 47360
rect 7096 47296 7112 47360
rect 7176 47296 7192 47360
rect 7256 47296 7264 47360
rect 6944 46272 7264 47296
rect 6944 46208 6952 46272
rect 7016 46208 7032 46272
rect 7096 46208 7112 46272
rect 7176 46208 7192 46272
rect 7256 46208 7264 46272
rect 6944 45184 7264 46208
rect 6944 45120 6952 45184
rect 7016 45120 7032 45184
rect 7096 45120 7112 45184
rect 7176 45120 7192 45184
rect 7256 45120 7264 45184
rect 6944 44096 7264 45120
rect 6944 44032 6952 44096
rect 7016 44032 7032 44096
rect 7096 44032 7112 44096
rect 7176 44032 7192 44096
rect 7256 44032 7264 44096
rect 6944 43294 7264 44032
rect 7422 43349 7482 50763
rect 7604 50080 7924 51104
rect 7604 50016 7612 50080
rect 7676 50016 7692 50080
rect 7756 50016 7772 50080
rect 7836 50016 7852 50080
rect 7916 50016 7924 50080
rect 7604 48992 7924 50016
rect 7604 48928 7612 48992
rect 7676 48954 7692 48992
rect 7756 48954 7772 48992
rect 7836 48954 7852 48992
rect 7916 48928 7924 48992
rect 7604 48718 7646 48928
rect 7882 48718 7924 48928
rect 7604 47904 7924 48718
rect 7604 47840 7612 47904
rect 7676 47840 7692 47904
rect 7756 47840 7772 47904
rect 7836 47840 7852 47904
rect 7916 47840 7924 47904
rect 7604 46816 7924 47840
rect 7604 46752 7612 46816
rect 7676 46752 7692 46816
rect 7756 46752 7772 46816
rect 7836 46752 7852 46816
rect 7916 46752 7924 46816
rect 7604 45728 7924 46752
rect 7604 45664 7612 45728
rect 7676 45664 7692 45728
rect 7756 45664 7772 45728
rect 7836 45664 7852 45728
rect 7916 45664 7924 45728
rect 7604 44640 7924 45664
rect 7604 44576 7612 44640
rect 7676 44576 7692 44640
rect 7756 44576 7772 44640
rect 7836 44576 7852 44640
rect 7916 44576 7924 44640
rect 7604 43954 7924 44576
rect 7604 43718 7646 43954
rect 7882 43718 7924 43954
rect 7604 43552 7924 43718
rect 7604 43488 7612 43552
rect 7676 43488 7692 43552
rect 7756 43488 7772 43552
rect 7836 43488 7852 43552
rect 7916 43488 7924 43552
rect 6944 43058 6986 43294
rect 7222 43058 7264 43294
rect 7419 43348 7485 43349
rect 7419 43284 7420 43348
rect 7484 43284 7485 43348
rect 7419 43283 7485 43284
rect 6944 43008 7264 43058
rect 6944 42944 6952 43008
rect 7016 42944 7032 43008
rect 7096 42944 7112 43008
rect 7176 42944 7192 43008
rect 7256 42944 7264 43008
rect 6944 41920 7264 42944
rect 6944 41856 6952 41920
rect 7016 41856 7032 41920
rect 7096 41856 7112 41920
rect 7176 41856 7192 41920
rect 7256 41856 7264 41920
rect 6944 40832 7264 41856
rect 6944 40768 6952 40832
rect 7016 40768 7032 40832
rect 7096 40768 7112 40832
rect 7176 40768 7192 40832
rect 7256 40768 7264 40832
rect 6944 39744 7264 40768
rect 6944 39680 6952 39744
rect 7016 39680 7032 39744
rect 7096 39680 7112 39744
rect 7176 39680 7192 39744
rect 7256 39680 7264 39744
rect 6944 38656 7264 39680
rect 6944 38592 6952 38656
rect 7016 38592 7032 38656
rect 7096 38592 7112 38656
rect 7176 38592 7192 38656
rect 7256 38592 7264 38656
rect 6944 38294 7264 38592
rect 6944 38058 6986 38294
rect 7222 38058 7264 38294
rect 6944 37568 7264 38058
rect 6944 37504 6952 37568
rect 7016 37504 7032 37568
rect 7096 37504 7112 37568
rect 7176 37504 7192 37568
rect 7256 37504 7264 37568
rect 6944 36480 7264 37504
rect 6944 36416 6952 36480
rect 7016 36416 7032 36480
rect 7096 36416 7112 36480
rect 7176 36416 7192 36480
rect 7256 36416 7264 36480
rect 6944 35392 7264 36416
rect 6944 35328 6952 35392
rect 7016 35328 7032 35392
rect 7096 35328 7112 35392
rect 7176 35328 7192 35392
rect 7256 35328 7264 35392
rect 6944 34304 7264 35328
rect 6944 34240 6952 34304
rect 7016 34240 7032 34304
rect 7096 34240 7112 34304
rect 7176 34240 7192 34304
rect 7256 34240 7264 34304
rect 6944 33294 7264 34240
rect 6944 33216 6986 33294
rect 7222 33216 7264 33294
rect 6944 33152 6952 33216
rect 7256 33152 7264 33216
rect 6944 33058 6986 33152
rect 7222 33058 7264 33152
rect 6944 32128 7264 33058
rect 6944 32064 6952 32128
rect 7016 32064 7032 32128
rect 7096 32064 7112 32128
rect 7176 32064 7192 32128
rect 7256 32064 7264 32128
rect 6944 31040 7264 32064
rect 6944 30976 6952 31040
rect 7016 30976 7032 31040
rect 7096 30976 7112 31040
rect 7176 30976 7192 31040
rect 7256 30976 7264 31040
rect 6944 29952 7264 30976
rect 6944 29888 6952 29952
rect 7016 29888 7032 29952
rect 7096 29888 7112 29952
rect 7176 29888 7192 29952
rect 7256 29888 7264 29952
rect 6944 28864 7264 29888
rect 6944 28800 6952 28864
rect 7016 28800 7032 28864
rect 7096 28800 7112 28864
rect 7176 28800 7192 28864
rect 7256 28800 7264 28864
rect 6944 28294 7264 28800
rect 6944 28058 6986 28294
rect 7222 28058 7264 28294
rect 6944 27776 7264 28058
rect 6944 27712 6952 27776
rect 7016 27712 7032 27776
rect 7096 27712 7112 27776
rect 7176 27712 7192 27776
rect 7256 27712 7264 27776
rect 6944 26688 7264 27712
rect 6944 26624 6952 26688
rect 7016 26624 7032 26688
rect 7096 26624 7112 26688
rect 7176 26624 7192 26688
rect 7256 26624 7264 26688
rect 6944 25600 7264 26624
rect 6944 25536 6952 25600
rect 7016 25536 7032 25600
rect 7096 25536 7112 25600
rect 7176 25536 7192 25600
rect 7256 25536 7264 25600
rect 6944 24512 7264 25536
rect 6944 24448 6952 24512
rect 7016 24448 7032 24512
rect 7096 24448 7112 24512
rect 7176 24448 7192 24512
rect 7256 24448 7264 24512
rect 6944 23424 7264 24448
rect 6944 23360 6952 23424
rect 7016 23360 7032 23424
rect 7096 23360 7112 23424
rect 7176 23360 7192 23424
rect 7256 23360 7264 23424
rect 6944 23294 7264 23360
rect 6944 23058 6986 23294
rect 7222 23058 7264 23294
rect 6944 22336 7264 23058
rect 6944 22272 6952 22336
rect 7016 22272 7032 22336
rect 7096 22272 7112 22336
rect 7176 22272 7192 22336
rect 7256 22272 7264 22336
rect 6944 21248 7264 22272
rect 6944 21184 6952 21248
rect 7016 21184 7032 21248
rect 7096 21184 7112 21248
rect 7176 21184 7192 21248
rect 7256 21184 7264 21248
rect 6944 20160 7264 21184
rect 6944 20096 6952 20160
rect 7016 20096 7032 20160
rect 7096 20096 7112 20160
rect 7176 20096 7192 20160
rect 7256 20096 7264 20160
rect 6944 19072 7264 20096
rect 6944 19008 6952 19072
rect 7016 19008 7032 19072
rect 7096 19008 7112 19072
rect 7176 19008 7192 19072
rect 7256 19008 7264 19072
rect 6944 18294 7264 19008
rect 6944 18058 6986 18294
rect 7222 18058 7264 18294
rect 6944 17984 7264 18058
rect 6944 17920 6952 17984
rect 7016 17920 7032 17984
rect 7096 17920 7112 17984
rect 7176 17920 7192 17984
rect 7256 17920 7264 17984
rect 6944 16896 7264 17920
rect 6944 16832 6952 16896
rect 7016 16832 7032 16896
rect 7096 16832 7112 16896
rect 7176 16832 7192 16896
rect 7256 16832 7264 16896
rect 6944 15808 7264 16832
rect 6944 15744 6952 15808
rect 7016 15744 7032 15808
rect 7096 15744 7112 15808
rect 7176 15744 7192 15808
rect 7256 15744 7264 15808
rect 6944 14720 7264 15744
rect 6944 14656 6952 14720
rect 7016 14656 7032 14720
rect 7096 14656 7112 14720
rect 7176 14656 7192 14720
rect 7256 14656 7264 14720
rect 6944 13632 7264 14656
rect 6944 13568 6952 13632
rect 7016 13568 7032 13632
rect 7096 13568 7112 13632
rect 7176 13568 7192 13632
rect 7256 13568 7264 13632
rect 6944 13294 7264 13568
rect 6944 13058 6986 13294
rect 7222 13058 7264 13294
rect 6944 12544 7264 13058
rect 6944 12480 6952 12544
rect 7016 12480 7032 12544
rect 7096 12480 7112 12544
rect 7176 12480 7192 12544
rect 7256 12480 7264 12544
rect 6944 11456 7264 12480
rect 6944 11392 6952 11456
rect 7016 11392 7032 11456
rect 7096 11392 7112 11456
rect 7176 11392 7192 11456
rect 7256 11392 7264 11456
rect 6944 10368 7264 11392
rect 6944 10304 6952 10368
rect 7016 10304 7032 10368
rect 7096 10304 7112 10368
rect 7176 10304 7192 10368
rect 7256 10304 7264 10368
rect 6683 9620 6749 9621
rect 6683 9556 6684 9620
rect 6748 9556 6749 9620
rect 6683 9555 6749 9556
rect 6944 9280 7264 10304
rect 6944 9216 6952 9280
rect 7016 9216 7032 9280
rect 7096 9216 7112 9280
rect 7176 9216 7192 9280
rect 7256 9216 7264 9280
rect 6944 8294 7264 9216
rect 6944 8192 6986 8294
rect 7222 8192 7264 8294
rect 6944 8128 6952 8192
rect 7256 8128 7264 8192
rect 6944 8058 6986 8128
rect 7222 8058 7264 8128
rect 4659 7308 4725 7309
rect 4659 7244 4660 7308
rect 4724 7244 4725 7308
rect 4659 7243 4725 7244
rect 2604 6496 2612 6560
rect 2676 6496 2692 6560
rect 2756 6496 2772 6560
rect 2836 6496 2852 6560
rect 2916 6496 2924 6560
rect 2604 5472 2924 6496
rect 2604 5408 2612 5472
rect 2676 5408 2692 5472
rect 2756 5408 2772 5472
rect 2836 5408 2852 5472
rect 2916 5408 2924 5472
rect 2604 4384 2924 5408
rect 2604 4320 2612 4384
rect 2676 4320 2692 4384
rect 2756 4320 2772 4384
rect 2836 4320 2852 4384
rect 2916 4320 2924 4384
rect 2604 3954 2924 4320
rect 2604 3718 2646 3954
rect 2882 3718 2924 3954
rect 2604 3296 2924 3718
rect 2604 3232 2612 3296
rect 2676 3232 2692 3296
rect 2756 3232 2772 3296
rect 2836 3232 2852 3296
rect 2916 3232 2924 3296
rect 2604 2208 2924 3232
rect 2604 2144 2612 2208
rect 2676 2144 2692 2208
rect 2756 2144 2772 2208
rect 2836 2144 2852 2208
rect 2916 2144 2924 2208
rect 2604 2128 2924 2144
rect 6944 7104 7264 8058
rect 6944 7040 6952 7104
rect 7016 7040 7032 7104
rect 7096 7040 7112 7104
rect 7176 7040 7192 7104
rect 7256 7040 7264 7104
rect 6944 6016 7264 7040
rect 6944 5952 6952 6016
rect 7016 5952 7032 6016
rect 7096 5952 7112 6016
rect 7176 5952 7192 6016
rect 7256 5952 7264 6016
rect 6944 4928 7264 5952
rect 6944 4864 6952 4928
rect 7016 4864 7032 4928
rect 7096 4864 7112 4928
rect 7176 4864 7192 4928
rect 7256 4864 7264 4928
rect 6944 3840 7264 4864
rect 6944 3776 6952 3840
rect 7016 3776 7032 3840
rect 7096 3776 7112 3840
rect 7176 3776 7192 3840
rect 7256 3776 7264 3840
rect 6944 3294 7264 3776
rect 6944 3058 6986 3294
rect 7222 3058 7264 3294
rect 6944 2752 7264 3058
rect 6944 2688 6952 2752
rect 7016 2688 7032 2752
rect 7096 2688 7112 2752
rect 7176 2688 7192 2752
rect 7256 2688 7264 2752
rect 6944 2128 7264 2688
rect 7604 42464 7924 43488
rect 7604 42400 7612 42464
rect 7676 42400 7692 42464
rect 7756 42400 7772 42464
rect 7836 42400 7852 42464
rect 7916 42400 7924 42464
rect 7604 41376 7924 42400
rect 7604 41312 7612 41376
rect 7676 41312 7692 41376
rect 7756 41312 7772 41376
rect 7836 41312 7852 41376
rect 7916 41312 7924 41376
rect 7604 40288 7924 41312
rect 7604 40224 7612 40288
rect 7676 40224 7692 40288
rect 7756 40224 7772 40288
rect 7836 40224 7852 40288
rect 7916 40224 7924 40288
rect 7604 39200 7924 40224
rect 7604 39136 7612 39200
rect 7676 39136 7692 39200
rect 7756 39136 7772 39200
rect 7836 39136 7852 39200
rect 7916 39136 7924 39200
rect 7604 38954 7924 39136
rect 7604 38718 7646 38954
rect 7882 38718 7924 38954
rect 7604 38112 7924 38718
rect 7604 38048 7612 38112
rect 7676 38048 7692 38112
rect 7756 38048 7772 38112
rect 7836 38048 7852 38112
rect 7916 38048 7924 38112
rect 7604 37024 7924 38048
rect 7604 36960 7612 37024
rect 7676 36960 7692 37024
rect 7756 36960 7772 37024
rect 7836 36960 7852 37024
rect 7916 36960 7924 37024
rect 7604 35936 7924 36960
rect 7604 35872 7612 35936
rect 7676 35872 7692 35936
rect 7756 35872 7772 35936
rect 7836 35872 7852 35936
rect 7916 35872 7924 35936
rect 7604 34848 7924 35872
rect 7604 34784 7612 34848
rect 7676 34784 7692 34848
rect 7756 34784 7772 34848
rect 7836 34784 7852 34848
rect 7916 34784 7924 34848
rect 7604 33954 7924 34784
rect 7604 33760 7646 33954
rect 7882 33760 7924 33954
rect 7604 33696 7612 33760
rect 7676 33696 7692 33718
rect 7756 33696 7772 33718
rect 7836 33696 7852 33718
rect 7916 33696 7924 33760
rect 7604 32672 7924 33696
rect 7604 32608 7612 32672
rect 7676 32608 7692 32672
rect 7756 32608 7772 32672
rect 7836 32608 7852 32672
rect 7916 32608 7924 32672
rect 7604 31584 7924 32608
rect 7604 31520 7612 31584
rect 7676 31520 7692 31584
rect 7756 31520 7772 31584
rect 7836 31520 7852 31584
rect 7916 31520 7924 31584
rect 7604 30496 7924 31520
rect 7604 30432 7612 30496
rect 7676 30432 7692 30496
rect 7756 30432 7772 30496
rect 7836 30432 7852 30496
rect 7916 30432 7924 30496
rect 7604 29408 7924 30432
rect 7604 29344 7612 29408
rect 7676 29344 7692 29408
rect 7756 29344 7772 29408
rect 7836 29344 7852 29408
rect 7916 29344 7924 29408
rect 7604 28954 7924 29344
rect 7604 28718 7646 28954
rect 7882 28718 7924 28954
rect 7604 28320 7924 28718
rect 7604 28256 7612 28320
rect 7676 28256 7692 28320
rect 7756 28256 7772 28320
rect 7836 28256 7852 28320
rect 7916 28256 7924 28320
rect 7604 27232 7924 28256
rect 7604 27168 7612 27232
rect 7676 27168 7692 27232
rect 7756 27168 7772 27232
rect 7836 27168 7852 27232
rect 7916 27168 7924 27232
rect 7604 26144 7924 27168
rect 7604 26080 7612 26144
rect 7676 26080 7692 26144
rect 7756 26080 7772 26144
rect 7836 26080 7852 26144
rect 7916 26080 7924 26144
rect 7604 25056 7924 26080
rect 7604 24992 7612 25056
rect 7676 24992 7692 25056
rect 7756 24992 7772 25056
rect 7836 24992 7852 25056
rect 7916 24992 7924 25056
rect 7604 23968 7924 24992
rect 7604 23904 7612 23968
rect 7676 23954 7692 23968
rect 7756 23954 7772 23968
rect 7836 23954 7852 23968
rect 7916 23904 7924 23968
rect 7604 23718 7646 23904
rect 7882 23718 7924 23904
rect 7604 22880 7924 23718
rect 7604 22816 7612 22880
rect 7676 22816 7692 22880
rect 7756 22816 7772 22880
rect 7836 22816 7852 22880
rect 7916 22816 7924 22880
rect 7604 21792 7924 22816
rect 7604 21728 7612 21792
rect 7676 21728 7692 21792
rect 7756 21728 7772 21792
rect 7836 21728 7852 21792
rect 7916 21728 7924 21792
rect 7604 20704 7924 21728
rect 7604 20640 7612 20704
rect 7676 20640 7692 20704
rect 7756 20640 7772 20704
rect 7836 20640 7852 20704
rect 7916 20640 7924 20704
rect 7604 19616 7924 20640
rect 7604 19552 7612 19616
rect 7676 19552 7692 19616
rect 7756 19552 7772 19616
rect 7836 19552 7852 19616
rect 7916 19552 7924 19616
rect 7604 18954 7924 19552
rect 7604 18718 7646 18954
rect 7882 18718 7924 18954
rect 7604 18528 7924 18718
rect 7604 18464 7612 18528
rect 7676 18464 7692 18528
rect 7756 18464 7772 18528
rect 7836 18464 7852 18528
rect 7916 18464 7924 18528
rect 7604 17440 7924 18464
rect 7604 17376 7612 17440
rect 7676 17376 7692 17440
rect 7756 17376 7772 17440
rect 7836 17376 7852 17440
rect 7916 17376 7924 17440
rect 7604 16352 7924 17376
rect 7604 16288 7612 16352
rect 7676 16288 7692 16352
rect 7756 16288 7772 16352
rect 7836 16288 7852 16352
rect 7916 16288 7924 16352
rect 7604 15264 7924 16288
rect 7604 15200 7612 15264
rect 7676 15200 7692 15264
rect 7756 15200 7772 15264
rect 7836 15200 7852 15264
rect 7916 15200 7924 15264
rect 7604 14176 7924 15200
rect 7604 14112 7612 14176
rect 7676 14112 7692 14176
rect 7756 14112 7772 14176
rect 7836 14112 7852 14176
rect 7916 14112 7924 14176
rect 7604 13954 7924 14112
rect 7604 13718 7646 13954
rect 7882 13718 7924 13954
rect 7604 13088 7924 13718
rect 7604 13024 7612 13088
rect 7676 13024 7692 13088
rect 7756 13024 7772 13088
rect 7836 13024 7852 13088
rect 7916 13024 7924 13088
rect 7604 12000 7924 13024
rect 7604 11936 7612 12000
rect 7676 11936 7692 12000
rect 7756 11936 7772 12000
rect 7836 11936 7852 12000
rect 7916 11936 7924 12000
rect 7604 10912 7924 11936
rect 7604 10848 7612 10912
rect 7676 10848 7692 10912
rect 7756 10848 7772 10912
rect 7836 10848 7852 10912
rect 7916 10848 7924 10912
rect 7604 9824 7924 10848
rect 7604 9760 7612 9824
rect 7676 9760 7692 9824
rect 7756 9760 7772 9824
rect 7836 9760 7852 9824
rect 7916 9760 7924 9824
rect 7604 8954 7924 9760
rect 7604 8736 7646 8954
rect 7882 8736 7924 8954
rect 7604 8672 7612 8736
rect 7676 8672 7692 8718
rect 7756 8672 7772 8718
rect 7836 8672 7852 8718
rect 7916 8672 7924 8736
rect 7604 7648 7924 8672
rect 7604 7584 7612 7648
rect 7676 7584 7692 7648
rect 7756 7584 7772 7648
rect 7836 7584 7852 7648
rect 7916 7584 7924 7648
rect 7604 6560 7924 7584
rect 8158 6901 8218 51851
rect 8339 28524 8405 28525
rect 8339 28460 8340 28524
rect 8404 28460 8405 28524
rect 8339 28459 8405 28460
rect 8342 26077 8402 28459
rect 8339 26076 8405 26077
rect 8339 26012 8340 26076
rect 8404 26012 8405 26076
rect 8339 26011 8405 26012
rect 8526 15197 8586 52531
rect 8710 33149 8770 62595
rect 8707 33148 8773 33149
rect 8707 33084 8708 33148
rect 8772 33084 8773 33148
rect 8707 33083 8773 33084
rect 8523 15196 8589 15197
rect 8523 15132 8524 15196
rect 8588 15132 8589 15196
rect 8523 15131 8589 15132
rect 8894 11253 8954 76059
rect 10363 67692 10429 67693
rect 10363 67628 10364 67692
rect 10428 67628 10429 67692
rect 10363 67627 10429 67628
rect 9075 59940 9141 59941
rect 9075 59876 9076 59940
rect 9140 59876 9141 59940
rect 9075 59875 9141 59876
rect 9078 40629 9138 59875
rect 10179 54092 10245 54093
rect 10179 54028 10180 54092
rect 10244 54028 10245 54092
rect 10179 54027 10245 54028
rect 9075 40628 9141 40629
rect 9075 40564 9076 40628
rect 9140 40564 9141 40628
rect 9075 40563 9141 40564
rect 9259 40492 9325 40493
rect 9259 40428 9260 40492
rect 9324 40428 9325 40492
rect 9259 40427 9325 40428
rect 9075 33012 9141 33013
rect 9075 32948 9076 33012
rect 9140 32948 9141 33012
rect 9075 32947 9141 32948
rect 9078 12341 9138 32947
rect 9262 26893 9322 40427
rect 9811 36412 9877 36413
rect 9811 36348 9812 36412
rect 9876 36348 9877 36412
rect 9811 36347 9877 36348
rect 9443 27028 9509 27029
rect 9443 26964 9444 27028
rect 9508 26964 9509 27028
rect 9443 26963 9509 26964
rect 9259 26892 9325 26893
rect 9259 26828 9260 26892
rect 9324 26828 9325 26892
rect 9259 26827 9325 26828
rect 9075 12340 9141 12341
rect 9075 12276 9076 12340
rect 9140 12276 9141 12340
rect 9075 12275 9141 12276
rect 8891 11252 8957 11253
rect 8891 11188 8892 11252
rect 8956 11188 8957 11252
rect 8891 11187 8957 11188
rect 9446 8125 9506 26963
rect 9443 8124 9509 8125
rect 9443 8060 9444 8124
rect 9508 8060 9509 8124
rect 9443 8059 9509 8060
rect 8155 6900 8221 6901
rect 8155 6836 8156 6900
rect 8220 6836 8221 6900
rect 8155 6835 8221 6836
rect 9814 6765 9874 36347
rect 10182 26077 10242 54027
rect 10179 26076 10245 26077
rect 10179 26012 10180 26076
rect 10244 26012 10245 26076
rect 10179 26011 10245 26012
rect 10366 25397 10426 67627
rect 10915 52460 10981 52461
rect 10915 52396 10916 52460
rect 10980 52396 10981 52460
rect 10915 52395 10981 52396
rect 10731 50692 10797 50693
rect 10731 50628 10732 50692
rect 10796 50628 10797 50692
rect 10731 50627 10797 50628
rect 10734 31770 10794 50627
rect 10918 35733 10978 52395
rect 11286 42805 11346 76195
rect 11944 75648 12264 76672
rect 11944 75584 11952 75648
rect 12016 75584 12032 75648
rect 12096 75584 12112 75648
rect 12176 75584 12192 75648
rect 12256 75584 12264 75648
rect 11944 74560 12264 75584
rect 11944 74496 11952 74560
rect 12016 74496 12032 74560
rect 12096 74496 12112 74560
rect 12176 74496 12192 74560
rect 12256 74496 12264 74560
rect 11944 73472 12264 74496
rect 11944 73408 11952 73472
rect 12016 73408 12032 73472
rect 12096 73408 12112 73472
rect 12176 73408 12192 73472
rect 12256 73408 12264 73472
rect 11944 73294 12264 73408
rect 11944 73058 11986 73294
rect 12222 73058 12264 73294
rect 11944 72384 12264 73058
rect 11944 72320 11952 72384
rect 12016 72320 12032 72384
rect 12096 72320 12112 72384
rect 12176 72320 12192 72384
rect 12256 72320 12264 72384
rect 11944 71296 12264 72320
rect 11944 71232 11952 71296
rect 12016 71232 12032 71296
rect 12096 71232 12112 71296
rect 12176 71232 12192 71296
rect 12256 71232 12264 71296
rect 11944 70208 12264 71232
rect 11944 70144 11952 70208
rect 12016 70144 12032 70208
rect 12096 70144 12112 70208
rect 12176 70144 12192 70208
rect 12256 70144 12264 70208
rect 11944 69120 12264 70144
rect 11944 69056 11952 69120
rect 12016 69056 12032 69120
rect 12096 69056 12112 69120
rect 12176 69056 12192 69120
rect 12256 69056 12264 69120
rect 11944 68294 12264 69056
rect 11944 68058 11986 68294
rect 12222 68058 12264 68294
rect 11944 68032 12264 68058
rect 11944 67968 11952 68032
rect 12016 67968 12032 68032
rect 12096 67968 12112 68032
rect 12176 67968 12192 68032
rect 12256 67968 12264 68032
rect 11651 67692 11717 67693
rect 11651 67628 11652 67692
rect 11716 67628 11717 67692
rect 11651 67627 11717 67628
rect 11283 42804 11349 42805
rect 11283 42740 11284 42804
rect 11348 42740 11349 42804
rect 11283 42739 11349 42740
rect 11467 42804 11533 42805
rect 11467 42740 11468 42804
rect 11532 42740 11533 42804
rect 11467 42739 11533 42740
rect 10915 35732 10981 35733
rect 10915 35668 10916 35732
rect 10980 35668 10981 35732
rect 10915 35667 10981 35668
rect 10734 31710 10978 31770
rect 10363 25396 10429 25397
rect 10363 25332 10364 25396
rect 10428 25332 10429 25396
rect 10363 25331 10429 25332
rect 9811 6764 9877 6765
rect 9811 6700 9812 6764
rect 9876 6700 9877 6764
rect 9811 6699 9877 6700
rect 7604 6496 7612 6560
rect 7676 6496 7692 6560
rect 7756 6496 7772 6560
rect 7836 6496 7852 6560
rect 7916 6496 7924 6560
rect 7604 5472 7924 6496
rect 7604 5408 7612 5472
rect 7676 5408 7692 5472
rect 7756 5408 7772 5472
rect 7836 5408 7852 5472
rect 7916 5408 7924 5472
rect 7604 4384 7924 5408
rect 10918 5269 10978 31710
rect 11283 26212 11349 26213
rect 11283 26148 11284 26212
rect 11348 26148 11349 26212
rect 11283 26147 11349 26148
rect 11286 15605 11346 26147
rect 11283 15604 11349 15605
rect 11283 15540 11284 15604
rect 11348 15540 11349 15604
rect 11283 15539 11349 15540
rect 11470 13293 11530 42739
rect 11654 26077 11714 67627
rect 11944 66944 12264 67968
rect 11944 66880 11952 66944
rect 12016 66880 12032 66944
rect 12096 66880 12112 66944
rect 12176 66880 12192 66944
rect 12256 66880 12264 66944
rect 11944 65856 12264 66880
rect 11944 65792 11952 65856
rect 12016 65792 12032 65856
rect 12096 65792 12112 65856
rect 12176 65792 12192 65856
rect 12256 65792 12264 65856
rect 11944 64768 12264 65792
rect 11944 64704 11952 64768
rect 12016 64704 12032 64768
rect 12096 64704 12112 64768
rect 12176 64704 12192 64768
rect 12256 64704 12264 64768
rect 11944 63680 12264 64704
rect 11944 63616 11952 63680
rect 12016 63616 12032 63680
rect 12096 63616 12112 63680
rect 12176 63616 12192 63680
rect 12256 63616 12264 63680
rect 11944 63294 12264 63616
rect 11944 63058 11986 63294
rect 12222 63058 12264 63294
rect 11944 62592 12264 63058
rect 11944 62528 11952 62592
rect 12016 62528 12032 62592
rect 12096 62528 12112 62592
rect 12176 62528 12192 62592
rect 12256 62528 12264 62592
rect 11944 61504 12264 62528
rect 11944 61440 11952 61504
rect 12016 61440 12032 61504
rect 12096 61440 12112 61504
rect 12176 61440 12192 61504
rect 12256 61440 12264 61504
rect 11944 60416 12264 61440
rect 11944 60352 11952 60416
rect 12016 60352 12032 60416
rect 12096 60352 12112 60416
rect 12176 60352 12192 60416
rect 12256 60352 12264 60416
rect 11944 59328 12264 60352
rect 11944 59264 11952 59328
rect 12016 59264 12032 59328
rect 12096 59264 12112 59328
rect 12176 59264 12192 59328
rect 12256 59264 12264 59328
rect 11944 58294 12264 59264
rect 11944 58240 11986 58294
rect 12222 58240 12264 58294
rect 11944 58176 11952 58240
rect 12256 58176 12264 58240
rect 11944 58058 11986 58176
rect 12222 58058 12264 58176
rect 11944 57152 12264 58058
rect 11944 57088 11952 57152
rect 12016 57088 12032 57152
rect 12096 57088 12112 57152
rect 12176 57088 12192 57152
rect 12256 57088 12264 57152
rect 11944 56064 12264 57088
rect 11944 56000 11952 56064
rect 12016 56000 12032 56064
rect 12096 56000 12112 56064
rect 12176 56000 12192 56064
rect 12256 56000 12264 56064
rect 11944 54976 12264 56000
rect 11944 54912 11952 54976
rect 12016 54912 12032 54976
rect 12096 54912 12112 54976
rect 12176 54912 12192 54976
rect 12256 54912 12264 54976
rect 11944 53888 12264 54912
rect 11944 53824 11952 53888
rect 12016 53824 12032 53888
rect 12096 53824 12112 53888
rect 12176 53824 12192 53888
rect 12256 53824 12264 53888
rect 11944 53294 12264 53824
rect 11944 53058 11986 53294
rect 12222 53058 12264 53294
rect 11944 52800 12264 53058
rect 11944 52736 11952 52800
rect 12016 52736 12032 52800
rect 12096 52736 12112 52800
rect 12176 52736 12192 52800
rect 12256 52736 12264 52800
rect 11944 51712 12264 52736
rect 11944 51648 11952 51712
rect 12016 51648 12032 51712
rect 12096 51648 12112 51712
rect 12176 51648 12192 51712
rect 12256 51648 12264 51712
rect 11944 50624 12264 51648
rect 11944 50560 11952 50624
rect 12016 50560 12032 50624
rect 12096 50560 12112 50624
rect 12176 50560 12192 50624
rect 12256 50560 12264 50624
rect 11944 49536 12264 50560
rect 11944 49472 11952 49536
rect 12016 49472 12032 49536
rect 12096 49472 12112 49536
rect 12176 49472 12192 49536
rect 12256 49472 12264 49536
rect 11944 48448 12264 49472
rect 11944 48384 11952 48448
rect 12016 48384 12032 48448
rect 12096 48384 12112 48448
rect 12176 48384 12192 48448
rect 12256 48384 12264 48448
rect 11944 48294 12264 48384
rect 11944 48058 11986 48294
rect 12222 48058 12264 48294
rect 11944 47360 12264 48058
rect 11944 47296 11952 47360
rect 12016 47296 12032 47360
rect 12096 47296 12112 47360
rect 12176 47296 12192 47360
rect 12256 47296 12264 47360
rect 11944 46272 12264 47296
rect 11944 46208 11952 46272
rect 12016 46208 12032 46272
rect 12096 46208 12112 46272
rect 12176 46208 12192 46272
rect 12256 46208 12264 46272
rect 11944 45184 12264 46208
rect 11944 45120 11952 45184
rect 12016 45120 12032 45184
rect 12096 45120 12112 45184
rect 12176 45120 12192 45184
rect 12256 45120 12264 45184
rect 11944 44096 12264 45120
rect 11944 44032 11952 44096
rect 12016 44032 12032 44096
rect 12096 44032 12112 44096
rect 12176 44032 12192 44096
rect 12256 44032 12264 44096
rect 11944 43294 12264 44032
rect 11944 43058 11986 43294
rect 12222 43058 12264 43294
rect 11944 43008 12264 43058
rect 11944 42944 11952 43008
rect 12016 42944 12032 43008
rect 12096 42944 12112 43008
rect 12176 42944 12192 43008
rect 12256 42944 12264 43008
rect 11944 41920 12264 42944
rect 11944 41856 11952 41920
rect 12016 41856 12032 41920
rect 12096 41856 12112 41920
rect 12176 41856 12192 41920
rect 12256 41856 12264 41920
rect 11944 40832 12264 41856
rect 11944 40768 11952 40832
rect 12016 40768 12032 40832
rect 12096 40768 12112 40832
rect 12176 40768 12192 40832
rect 12256 40768 12264 40832
rect 11944 39744 12264 40768
rect 11944 39680 11952 39744
rect 12016 39680 12032 39744
rect 12096 39680 12112 39744
rect 12176 39680 12192 39744
rect 12256 39680 12264 39744
rect 11944 38656 12264 39680
rect 11944 38592 11952 38656
rect 12016 38592 12032 38656
rect 12096 38592 12112 38656
rect 12176 38592 12192 38656
rect 12256 38592 12264 38656
rect 11944 38294 12264 38592
rect 11944 38058 11986 38294
rect 12222 38058 12264 38294
rect 11944 37568 12264 38058
rect 11944 37504 11952 37568
rect 12016 37504 12032 37568
rect 12096 37504 12112 37568
rect 12176 37504 12192 37568
rect 12256 37504 12264 37568
rect 11944 36480 12264 37504
rect 11944 36416 11952 36480
rect 12016 36416 12032 36480
rect 12096 36416 12112 36480
rect 12176 36416 12192 36480
rect 12256 36416 12264 36480
rect 11944 35392 12264 36416
rect 11944 35328 11952 35392
rect 12016 35328 12032 35392
rect 12096 35328 12112 35392
rect 12176 35328 12192 35392
rect 12256 35328 12264 35392
rect 11944 34304 12264 35328
rect 11944 34240 11952 34304
rect 12016 34240 12032 34304
rect 12096 34240 12112 34304
rect 12176 34240 12192 34304
rect 12256 34240 12264 34304
rect 11944 33294 12264 34240
rect 11944 33216 11986 33294
rect 12222 33216 12264 33294
rect 11944 33152 11952 33216
rect 12256 33152 12264 33216
rect 11944 33058 11986 33152
rect 12222 33058 12264 33152
rect 11944 32128 12264 33058
rect 11944 32064 11952 32128
rect 12016 32064 12032 32128
rect 12096 32064 12112 32128
rect 12176 32064 12192 32128
rect 12256 32064 12264 32128
rect 11944 31040 12264 32064
rect 11944 30976 11952 31040
rect 12016 30976 12032 31040
rect 12096 30976 12112 31040
rect 12176 30976 12192 31040
rect 12256 30976 12264 31040
rect 11944 29952 12264 30976
rect 11944 29888 11952 29952
rect 12016 29888 12032 29952
rect 12096 29888 12112 29952
rect 12176 29888 12192 29952
rect 12256 29888 12264 29952
rect 11944 28864 12264 29888
rect 11944 28800 11952 28864
rect 12016 28800 12032 28864
rect 12096 28800 12112 28864
rect 12176 28800 12192 28864
rect 12256 28800 12264 28864
rect 11944 28294 12264 28800
rect 11944 28058 11986 28294
rect 12222 28058 12264 28294
rect 11944 27776 12264 28058
rect 11944 27712 11952 27776
rect 12016 27712 12032 27776
rect 12096 27712 12112 27776
rect 12176 27712 12192 27776
rect 12256 27712 12264 27776
rect 11944 26688 12264 27712
rect 11944 26624 11952 26688
rect 12016 26624 12032 26688
rect 12096 26624 12112 26688
rect 12176 26624 12192 26688
rect 12256 26624 12264 26688
rect 11651 26076 11717 26077
rect 11651 26012 11652 26076
rect 11716 26012 11717 26076
rect 11651 26011 11717 26012
rect 11944 25600 12264 26624
rect 11944 25536 11952 25600
rect 12016 25536 12032 25600
rect 12096 25536 12112 25600
rect 12176 25536 12192 25600
rect 12256 25536 12264 25600
rect 11944 24512 12264 25536
rect 11944 24448 11952 24512
rect 12016 24448 12032 24512
rect 12096 24448 12112 24512
rect 12176 24448 12192 24512
rect 12256 24448 12264 24512
rect 11944 23424 12264 24448
rect 11944 23360 11952 23424
rect 12016 23360 12032 23424
rect 12096 23360 12112 23424
rect 12176 23360 12192 23424
rect 12256 23360 12264 23424
rect 11944 23294 12264 23360
rect 11944 23058 11986 23294
rect 12222 23058 12264 23294
rect 11944 22336 12264 23058
rect 11944 22272 11952 22336
rect 12016 22272 12032 22336
rect 12096 22272 12112 22336
rect 12176 22272 12192 22336
rect 12256 22272 12264 22336
rect 11944 21248 12264 22272
rect 11944 21184 11952 21248
rect 12016 21184 12032 21248
rect 12096 21184 12112 21248
rect 12176 21184 12192 21248
rect 12256 21184 12264 21248
rect 11944 20160 12264 21184
rect 11944 20096 11952 20160
rect 12016 20096 12032 20160
rect 12096 20096 12112 20160
rect 12176 20096 12192 20160
rect 12256 20096 12264 20160
rect 11944 19072 12264 20096
rect 11944 19008 11952 19072
rect 12016 19008 12032 19072
rect 12096 19008 12112 19072
rect 12176 19008 12192 19072
rect 12256 19008 12264 19072
rect 11944 18294 12264 19008
rect 11944 18058 11986 18294
rect 12222 18058 12264 18294
rect 11944 17984 12264 18058
rect 11944 17920 11952 17984
rect 12016 17920 12032 17984
rect 12096 17920 12112 17984
rect 12176 17920 12192 17984
rect 12256 17920 12264 17984
rect 11944 16896 12264 17920
rect 11944 16832 11952 16896
rect 12016 16832 12032 16896
rect 12096 16832 12112 16896
rect 12176 16832 12192 16896
rect 12256 16832 12264 16896
rect 11944 15808 12264 16832
rect 11944 15744 11952 15808
rect 12016 15744 12032 15808
rect 12096 15744 12112 15808
rect 12176 15744 12192 15808
rect 12256 15744 12264 15808
rect 11944 14720 12264 15744
rect 11944 14656 11952 14720
rect 12016 14656 12032 14720
rect 12096 14656 12112 14720
rect 12176 14656 12192 14720
rect 12256 14656 12264 14720
rect 11944 13632 12264 14656
rect 11944 13568 11952 13632
rect 12016 13568 12032 13632
rect 12096 13568 12112 13632
rect 12176 13568 12192 13632
rect 12256 13568 12264 13632
rect 11944 13294 12264 13568
rect 11467 13292 11533 13293
rect 11467 13228 11468 13292
rect 11532 13228 11533 13292
rect 11467 13227 11533 13228
rect 11944 13058 11986 13294
rect 12222 13058 12264 13294
rect 11944 12544 12264 13058
rect 11944 12480 11952 12544
rect 12016 12480 12032 12544
rect 12096 12480 12112 12544
rect 12176 12480 12192 12544
rect 12256 12480 12264 12544
rect 11944 11456 12264 12480
rect 11944 11392 11952 11456
rect 12016 11392 12032 11456
rect 12096 11392 12112 11456
rect 12176 11392 12192 11456
rect 12256 11392 12264 11456
rect 11944 10368 12264 11392
rect 11944 10304 11952 10368
rect 12016 10304 12032 10368
rect 12096 10304 12112 10368
rect 12176 10304 12192 10368
rect 12256 10304 12264 10368
rect 11944 9280 12264 10304
rect 11944 9216 11952 9280
rect 12016 9216 12032 9280
rect 12096 9216 12112 9280
rect 12176 9216 12192 9280
rect 12256 9216 12264 9280
rect 11944 8294 12264 9216
rect 11944 8192 11986 8294
rect 12222 8192 12264 8294
rect 11944 8128 11952 8192
rect 12256 8128 12264 8192
rect 11944 8058 11986 8128
rect 12222 8058 12264 8128
rect 11944 7104 12264 8058
rect 11944 7040 11952 7104
rect 12016 7040 12032 7104
rect 12096 7040 12112 7104
rect 12176 7040 12192 7104
rect 12256 7040 12264 7104
rect 11944 6016 12264 7040
rect 11944 5952 11952 6016
rect 12016 5952 12032 6016
rect 12096 5952 12112 6016
rect 12176 5952 12192 6016
rect 12256 5952 12264 6016
rect 10915 5268 10981 5269
rect 10915 5204 10916 5268
rect 10980 5204 10981 5268
rect 10915 5203 10981 5204
rect 7604 4320 7612 4384
rect 7676 4320 7692 4384
rect 7756 4320 7772 4384
rect 7836 4320 7852 4384
rect 7916 4320 7924 4384
rect 7604 3954 7924 4320
rect 7604 3718 7646 3954
rect 7882 3718 7924 3954
rect 7604 3296 7924 3718
rect 7604 3232 7612 3296
rect 7676 3232 7692 3296
rect 7756 3232 7772 3296
rect 7836 3232 7852 3296
rect 7916 3232 7924 3296
rect 7604 2208 7924 3232
rect 7604 2144 7612 2208
rect 7676 2144 7692 2208
rect 7756 2144 7772 2208
rect 7836 2144 7852 2208
rect 7916 2144 7924 2208
rect 7604 2128 7924 2144
rect 11944 4928 12264 5952
rect 11944 4864 11952 4928
rect 12016 4864 12032 4928
rect 12096 4864 12112 4928
rect 12176 4864 12192 4928
rect 12256 4864 12264 4928
rect 11944 3840 12264 4864
rect 11944 3776 11952 3840
rect 12016 3776 12032 3840
rect 12096 3776 12112 3840
rect 12176 3776 12192 3840
rect 12256 3776 12264 3840
rect 11944 3294 12264 3776
rect 11944 3058 11986 3294
rect 12222 3058 12264 3294
rect 11944 2752 12264 3058
rect 11944 2688 11952 2752
rect 12016 2688 12032 2752
rect 12096 2688 12112 2752
rect 12176 2688 12192 2752
rect 12256 2688 12264 2752
rect 11944 2128 12264 2688
rect 12604 77280 12924 77840
rect 12604 77216 12612 77280
rect 12676 77216 12692 77280
rect 12756 77216 12772 77280
rect 12836 77216 12852 77280
rect 12916 77216 12924 77280
rect 12604 76192 12924 77216
rect 16944 77824 17264 77840
rect 16944 77760 16952 77824
rect 17016 77760 17032 77824
rect 17096 77760 17112 77824
rect 17176 77760 17192 77824
rect 17256 77760 17264 77824
rect 14595 76804 14661 76805
rect 14595 76740 14596 76804
rect 14660 76740 14661 76804
rect 14595 76739 14661 76740
rect 15883 76804 15949 76805
rect 15883 76740 15884 76804
rect 15948 76740 15949 76804
rect 15883 76739 15949 76740
rect 12604 76128 12612 76192
rect 12676 76128 12692 76192
rect 12756 76128 12772 76192
rect 12836 76128 12852 76192
rect 12916 76128 12924 76192
rect 12604 75104 12924 76128
rect 14227 75988 14293 75989
rect 14227 75924 14228 75988
rect 14292 75924 14293 75988
rect 14227 75923 14293 75924
rect 12604 75040 12612 75104
rect 12676 75040 12692 75104
rect 12756 75040 12772 75104
rect 12836 75040 12852 75104
rect 12916 75040 12924 75104
rect 12604 74016 12924 75040
rect 12604 73952 12612 74016
rect 12676 73954 12692 74016
rect 12756 73954 12772 74016
rect 12836 73954 12852 74016
rect 12916 73952 12924 74016
rect 12604 73718 12646 73952
rect 12882 73718 12924 73952
rect 12604 72928 12924 73718
rect 12604 72864 12612 72928
rect 12676 72864 12692 72928
rect 12756 72864 12772 72928
rect 12836 72864 12852 72928
rect 12916 72864 12924 72928
rect 12604 71840 12924 72864
rect 12604 71776 12612 71840
rect 12676 71776 12692 71840
rect 12756 71776 12772 71840
rect 12836 71776 12852 71840
rect 12916 71776 12924 71840
rect 12604 70752 12924 71776
rect 12604 70688 12612 70752
rect 12676 70688 12692 70752
rect 12756 70688 12772 70752
rect 12836 70688 12852 70752
rect 12916 70688 12924 70752
rect 12604 69664 12924 70688
rect 12604 69600 12612 69664
rect 12676 69600 12692 69664
rect 12756 69600 12772 69664
rect 12836 69600 12852 69664
rect 12916 69600 12924 69664
rect 12604 68954 12924 69600
rect 12604 68718 12646 68954
rect 12882 68718 12924 68954
rect 12604 68576 12924 68718
rect 12604 68512 12612 68576
rect 12676 68512 12692 68576
rect 12756 68512 12772 68576
rect 12836 68512 12852 68576
rect 12916 68512 12924 68576
rect 12604 67488 12924 68512
rect 12604 67424 12612 67488
rect 12676 67424 12692 67488
rect 12756 67424 12772 67488
rect 12836 67424 12852 67488
rect 12916 67424 12924 67488
rect 12604 66400 12924 67424
rect 12604 66336 12612 66400
rect 12676 66336 12692 66400
rect 12756 66336 12772 66400
rect 12836 66336 12852 66400
rect 12916 66336 12924 66400
rect 12604 65312 12924 66336
rect 12604 65248 12612 65312
rect 12676 65248 12692 65312
rect 12756 65248 12772 65312
rect 12836 65248 12852 65312
rect 12916 65248 12924 65312
rect 12604 64224 12924 65248
rect 12604 64160 12612 64224
rect 12676 64160 12692 64224
rect 12756 64160 12772 64224
rect 12836 64160 12852 64224
rect 12916 64160 12924 64224
rect 12604 63954 12924 64160
rect 12604 63718 12646 63954
rect 12882 63718 12924 63954
rect 12604 63136 12924 63718
rect 12604 63072 12612 63136
rect 12676 63072 12692 63136
rect 12756 63072 12772 63136
rect 12836 63072 12852 63136
rect 12916 63072 12924 63136
rect 12604 62048 12924 63072
rect 12604 61984 12612 62048
rect 12676 61984 12692 62048
rect 12756 61984 12772 62048
rect 12836 61984 12852 62048
rect 12916 61984 12924 62048
rect 12604 60960 12924 61984
rect 12604 60896 12612 60960
rect 12676 60896 12692 60960
rect 12756 60896 12772 60960
rect 12836 60896 12852 60960
rect 12916 60896 12924 60960
rect 12604 59872 12924 60896
rect 12604 59808 12612 59872
rect 12676 59808 12692 59872
rect 12756 59808 12772 59872
rect 12836 59808 12852 59872
rect 12916 59808 12924 59872
rect 12604 58954 12924 59808
rect 12604 58784 12646 58954
rect 12882 58784 12924 58954
rect 13675 58852 13741 58853
rect 13675 58788 13676 58852
rect 13740 58788 13741 58852
rect 13675 58787 13741 58788
rect 12604 58720 12612 58784
rect 12916 58720 12924 58784
rect 12604 58718 12646 58720
rect 12882 58718 12924 58720
rect 12604 57696 12924 58718
rect 12604 57632 12612 57696
rect 12676 57632 12692 57696
rect 12756 57632 12772 57696
rect 12836 57632 12852 57696
rect 12916 57632 12924 57696
rect 12604 56608 12924 57632
rect 12604 56544 12612 56608
rect 12676 56544 12692 56608
rect 12756 56544 12772 56608
rect 12836 56544 12852 56608
rect 12916 56544 12924 56608
rect 12604 55520 12924 56544
rect 12604 55456 12612 55520
rect 12676 55456 12692 55520
rect 12756 55456 12772 55520
rect 12836 55456 12852 55520
rect 12916 55456 12924 55520
rect 12604 54432 12924 55456
rect 12604 54368 12612 54432
rect 12676 54368 12692 54432
rect 12756 54368 12772 54432
rect 12836 54368 12852 54432
rect 12916 54368 12924 54432
rect 12604 53954 12924 54368
rect 12604 53718 12646 53954
rect 12882 53718 12924 53954
rect 12604 53344 12924 53718
rect 12604 53280 12612 53344
rect 12676 53280 12692 53344
rect 12756 53280 12772 53344
rect 12836 53280 12852 53344
rect 12916 53280 12924 53344
rect 12604 52256 12924 53280
rect 12604 52192 12612 52256
rect 12676 52192 12692 52256
rect 12756 52192 12772 52256
rect 12836 52192 12852 52256
rect 12916 52192 12924 52256
rect 12604 51168 12924 52192
rect 13123 51372 13189 51373
rect 13123 51308 13124 51372
rect 13188 51308 13189 51372
rect 13123 51307 13189 51308
rect 12604 51104 12612 51168
rect 12676 51104 12692 51168
rect 12756 51104 12772 51168
rect 12836 51104 12852 51168
rect 12916 51104 12924 51168
rect 12604 50080 12924 51104
rect 12604 50016 12612 50080
rect 12676 50016 12692 50080
rect 12756 50016 12772 50080
rect 12836 50016 12852 50080
rect 12916 50016 12924 50080
rect 12604 48992 12924 50016
rect 12604 48928 12612 48992
rect 12676 48954 12692 48992
rect 12756 48954 12772 48992
rect 12836 48954 12852 48992
rect 12916 48928 12924 48992
rect 12604 48718 12646 48928
rect 12882 48718 12924 48928
rect 12604 47904 12924 48718
rect 12604 47840 12612 47904
rect 12676 47840 12692 47904
rect 12756 47840 12772 47904
rect 12836 47840 12852 47904
rect 12916 47840 12924 47904
rect 12604 46816 12924 47840
rect 12604 46752 12612 46816
rect 12676 46752 12692 46816
rect 12756 46752 12772 46816
rect 12836 46752 12852 46816
rect 12916 46752 12924 46816
rect 12604 45728 12924 46752
rect 12604 45664 12612 45728
rect 12676 45664 12692 45728
rect 12756 45664 12772 45728
rect 12836 45664 12852 45728
rect 12916 45664 12924 45728
rect 12604 44640 12924 45664
rect 12604 44576 12612 44640
rect 12676 44576 12692 44640
rect 12756 44576 12772 44640
rect 12836 44576 12852 44640
rect 12916 44576 12924 44640
rect 12604 43954 12924 44576
rect 12604 43718 12646 43954
rect 12882 43718 12924 43954
rect 12604 43552 12924 43718
rect 12604 43488 12612 43552
rect 12676 43488 12692 43552
rect 12756 43488 12772 43552
rect 12836 43488 12852 43552
rect 12916 43488 12924 43552
rect 12604 42464 12924 43488
rect 12604 42400 12612 42464
rect 12676 42400 12692 42464
rect 12756 42400 12772 42464
rect 12836 42400 12852 42464
rect 12916 42400 12924 42464
rect 12604 41376 12924 42400
rect 12604 41312 12612 41376
rect 12676 41312 12692 41376
rect 12756 41312 12772 41376
rect 12836 41312 12852 41376
rect 12916 41312 12924 41376
rect 12604 40288 12924 41312
rect 12604 40224 12612 40288
rect 12676 40224 12692 40288
rect 12756 40224 12772 40288
rect 12836 40224 12852 40288
rect 12916 40224 12924 40288
rect 12604 39200 12924 40224
rect 12604 39136 12612 39200
rect 12676 39136 12692 39200
rect 12756 39136 12772 39200
rect 12836 39136 12852 39200
rect 12916 39136 12924 39200
rect 12604 38954 12924 39136
rect 12604 38718 12646 38954
rect 12882 38718 12924 38954
rect 12604 38112 12924 38718
rect 12604 38048 12612 38112
rect 12676 38048 12692 38112
rect 12756 38048 12772 38112
rect 12836 38048 12852 38112
rect 12916 38048 12924 38112
rect 12604 37024 12924 38048
rect 12604 36960 12612 37024
rect 12676 36960 12692 37024
rect 12756 36960 12772 37024
rect 12836 36960 12852 37024
rect 12916 36960 12924 37024
rect 12604 35936 12924 36960
rect 12604 35872 12612 35936
rect 12676 35872 12692 35936
rect 12756 35872 12772 35936
rect 12836 35872 12852 35936
rect 12916 35872 12924 35936
rect 12604 34848 12924 35872
rect 12604 34784 12612 34848
rect 12676 34784 12692 34848
rect 12756 34784 12772 34848
rect 12836 34784 12852 34848
rect 12916 34784 12924 34848
rect 12604 33954 12924 34784
rect 12604 33760 12646 33954
rect 12882 33760 12924 33954
rect 12604 33696 12612 33760
rect 12676 33696 12692 33718
rect 12756 33696 12772 33718
rect 12836 33696 12852 33718
rect 12916 33696 12924 33760
rect 12604 32672 12924 33696
rect 12604 32608 12612 32672
rect 12676 32608 12692 32672
rect 12756 32608 12772 32672
rect 12836 32608 12852 32672
rect 12916 32608 12924 32672
rect 12604 31584 12924 32608
rect 12604 31520 12612 31584
rect 12676 31520 12692 31584
rect 12756 31520 12772 31584
rect 12836 31520 12852 31584
rect 12916 31520 12924 31584
rect 12604 30496 12924 31520
rect 12604 30432 12612 30496
rect 12676 30432 12692 30496
rect 12756 30432 12772 30496
rect 12836 30432 12852 30496
rect 12916 30432 12924 30496
rect 12604 29408 12924 30432
rect 12604 29344 12612 29408
rect 12676 29344 12692 29408
rect 12756 29344 12772 29408
rect 12836 29344 12852 29408
rect 12916 29344 12924 29408
rect 12604 28954 12924 29344
rect 12604 28718 12646 28954
rect 12882 28718 12924 28954
rect 12604 28320 12924 28718
rect 12604 28256 12612 28320
rect 12676 28256 12692 28320
rect 12756 28256 12772 28320
rect 12836 28256 12852 28320
rect 12916 28256 12924 28320
rect 12604 27232 12924 28256
rect 12604 27168 12612 27232
rect 12676 27168 12692 27232
rect 12756 27168 12772 27232
rect 12836 27168 12852 27232
rect 12916 27168 12924 27232
rect 12604 26144 12924 27168
rect 12604 26080 12612 26144
rect 12676 26080 12692 26144
rect 12756 26080 12772 26144
rect 12836 26080 12852 26144
rect 12916 26080 12924 26144
rect 12604 25056 12924 26080
rect 12604 24992 12612 25056
rect 12676 24992 12692 25056
rect 12756 24992 12772 25056
rect 12836 24992 12852 25056
rect 12916 24992 12924 25056
rect 12604 23968 12924 24992
rect 13126 24717 13186 51307
rect 13307 24852 13373 24853
rect 13307 24788 13308 24852
rect 13372 24788 13373 24852
rect 13307 24787 13373 24788
rect 13123 24716 13189 24717
rect 13123 24652 13124 24716
rect 13188 24652 13189 24716
rect 13123 24651 13189 24652
rect 12604 23904 12612 23968
rect 12676 23954 12692 23968
rect 12756 23954 12772 23968
rect 12836 23954 12852 23968
rect 12916 23904 12924 23968
rect 12604 23718 12646 23904
rect 12882 23718 12924 23904
rect 12604 22880 12924 23718
rect 12604 22816 12612 22880
rect 12676 22816 12692 22880
rect 12756 22816 12772 22880
rect 12836 22816 12852 22880
rect 12916 22816 12924 22880
rect 12604 21792 12924 22816
rect 12604 21728 12612 21792
rect 12676 21728 12692 21792
rect 12756 21728 12772 21792
rect 12836 21728 12852 21792
rect 12916 21728 12924 21792
rect 12604 20704 12924 21728
rect 12604 20640 12612 20704
rect 12676 20640 12692 20704
rect 12756 20640 12772 20704
rect 12836 20640 12852 20704
rect 12916 20640 12924 20704
rect 12604 19616 12924 20640
rect 12604 19552 12612 19616
rect 12676 19552 12692 19616
rect 12756 19552 12772 19616
rect 12836 19552 12852 19616
rect 12916 19552 12924 19616
rect 12604 18954 12924 19552
rect 12604 18718 12646 18954
rect 12882 18718 12924 18954
rect 12604 18528 12924 18718
rect 12604 18464 12612 18528
rect 12676 18464 12692 18528
rect 12756 18464 12772 18528
rect 12836 18464 12852 18528
rect 12916 18464 12924 18528
rect 12604 17440 12924 18464
rect 12604 17376 12612 17440
rect 12676 17376 12692 17440
rect 12756 17376 12772 17440
rect 12836 17376 12852 17440
rect 12916 17376 12924 17440
rect 12604 16352 12924 17376
rect 12604 16288 12612 16352
rect 12676 16288 12692 16352
rect 12756 16288 12772 16352
rect 12836 16288 12852 16352
rect 12916 16288 12924 16352
rect 12604 15264 12924 16288
rect 12604 15200 12612 15264
rect 12676 15200 12692 15264
rect 12756 15200 12772 15264
rect 12836 15200 12852 15264
rect 12916 15200 12924 15264
rect 12604 14176 12924 15200
rect 12604 14112 12612 14176
rect 12676 14112 12692 14176
rect 12756 14112 12772 14176
rect 12836 14112 12852 14176
rect 12916 14112 12924 14176
rect 12604 13954 12924 14112
rect 12604 13718 12646 13954
rect 12882 13718 12924 13954
rect 12604 13088 12924 13718
rect 12604 13024 12612 13088
rect 12676 13024 12692 13088
rect 12756 13024 12772 13088
rect 12836 13024 12852 13088
rect 12916 13024 12924 13088
rect 12604 12000 12924 13024
rect 12604 11936 12612 12000
rect 12676 11936 12692 12000
rect 12756 11936 12772 12000
rect 12836 11936 12852 12000
rect 12916 11936 12924 12000
rect 12604 10912 12924 11936
rect 12604 10848 12612 10912
rect 12676 10848 12692 10912
rect 12756 10848 12772 10912
rect 12836 10848 12852 10912
rect 12916 10848 12924 10912
rect 12604 9824 12924 10848
rect 12604 9760 12612 9824
rect 12676 9760 12692 9824
rect 12756 9760 12772 9824
rect 12836 9760 12852 9824
rect 12916 9760 12924 9824
rect 12604 8954 12924 9760
rect 12604 8736 12646 8954
rect 12882 8736 12924 8954
rect 12604 8672 12612 8736
rect 12676 8672 12692 8718
rect 12756 8672 12772 8718
rect 12836 8672 12852 8718
rect 12916 8672 12924 8736
rect 12604 7648 12924 8672
rect 12604 7584 12612 7648
rect 12676 7584 12692 7648
rect 12756 7584 12772 7648
rect 12836 7584 12852 7648
rect 12916 7584 12924 7648
rect 12604 6560 12924 7584
rect 13310 6901 13370 24787
rect 13678 12205 13738 58787
rect 13675 12204 13741 12205
rect 13675 12140 13676 12204
rect 13740 12140 13741 12204
rect 13675 12139 13741 12140
rect 14230 8261 14290 75923
rect 14411 55724 14477 55725
rect 14411 55660 14412 55724
rect 14476 55660 14477 55724
rect 14411 55659 14477 55660
rect 14414 22541 14474 55659
rect 14411 22540 14477 22541
rect 14411 22476 14412 22540
rect 14476 22476 14477 22540
rect 14411 22475 14477 22476
rect 14598 16557 14658 76739
rect 14963 69052 15029 69053
rect 14963 68988 14964 69052
rect 15028 68988 15029 69052
rect 14963 68987 15029 68988
rect 14966 29885 15026 68987
rect 15699 65108 15765 65109
rect 15699 65044 15700 65108
rect 15764 65044 15765 65108
rect 15699 65043 15765 65044
rect 15147 37364 15213 37365
rect 15147 37300 15148 37364
rect 15212 37300 15213 37364
rect 15147 37299 15213 37300
rect 14963 29884 15029 29885
rect 14963 29820 14964 29884
rect 15028 29820 15029 29884
rect 14963 29819 15029 29820
rect 14595 16556 14661 16557
rect 14595 16492 14596 16556
rect 14660 16492 14661 16556
rect 14595 16491 14661 16492
rect 15150 10573 15210 37299
rect 15702 11117 15762 65043
rect 15886 49605 15946 76739
rect 16944 76736 17264 77760
rect 16944 76672 16952 76736
rect 17016 76672 17032 76736
rect 17096 76672 17112 76736
rect 17176 76672 17192 76736
rect 17256 76672 17264 76736
rect 16944 75648 17264 76672
rect 16944 75584 16952 75648
rect 17016 75584 17032 75648
rect 17096 75584 17112 75648
rect 17176 75584 17192 75648
rect 17256 75584 17264 75648
rect 16944 74560 17264 75584
rect 16944 74496 16952 74560
rect 17016 74496 17032 74560
rect 17096 74496 17112 74560
rect 17176 74496 17192 74560
rect 17256 74496 17264 74560
rect 16944 73472 17264 74496
rect 16944 73408 16952 73472
rect 17016 73408 17032 73472
rect 17096 73408 17112 73472
rect 17176 73408 17192 73472
rect 17256 73408 17264 73472
rect 16944 73294 17264 73408
rect 16944 73058 16986 73294
rect 17222 73058 17264 73294
rect 16944 72384 17264 73058
rect 16944 72320 16952 72384
rect 17016 72320 17032 72384
rect 17096 72320 17112 72384
rect 17176 72320 17192 72384
rect 17256 72320 17264 72384
rect 16944 71296 17264 72320
rect 16944 71232 16952 71296
rect 17016 71232 17032 71296
rect 17096 71232 17112 71296
rect 17176 71232 17192 71296
rect 17256 71232 17264 71296
rect 16944 70208 17264 71232
rect 16944 70144 16952 70208
rect 17016 70144 17032 70208
rect 17096 70144 17112 70208
rect 17176 70144 17192 70208
rect 17256 70144 17264 70208
rect 16944 69120 17264 70144
rect 16944 69056 16952 69120
rect 17016 69056 17032 69120
rect 17096 69056 17112 69120
rect 17176 69056 17192 69120
rect 17256 69056 17264 69120
rect 16944 68294 17264 69056
rect 16944 68058 16986 68294
rect 17222 68058 17264 68294
rect 16944 68032 17264 68058
rect 16944 67968 16952 68032
rect 17016 67968 17032 68032
rect 17096 67968 17112 68032
rect 17176 67968 17192 68032
rect 17256 67968 17264 68032
rect 16944 66944 17264 67968
rect 16944 66880 16952 66944
rect 17016 66880 17032 66944
rect 17096 66880 17112 66944
rect 17176 66880 17192 66944
rect 17256 66880 17264 66944
rect 16944 65856 17264 66880
rect 16944 65792 16952 65856
rect 17016 65792 17032 65856
rect 17096 65792 17112 65856
rect 17176 65792 17192 65856
rect 17256 65792 17264 65856
rect 16944 64768 17264 65792
rect 16944 64704 16952 64768
rect 17016 64704 17032 64768
rect 17096 64704 17112 64768
rect 17176 64704 17192 64768
rect 17256 64704 17264 64768
rect 16944 63680 17264 64704
rect 16944 63616 16952 63680
rect 17016 63616 17032 63680
rect 17096 63616 17112 63680
rect 17176 63616 17192 63680
rect 17256 63616 17264 63680
rect 16944 63294 17264 63616
rect 16944 63058 16986 63294
rect 17222 63058 17264 63294
rect 16944 62592 17264 63058
rect 16944 62528 16952 62592
rect 17016 62528 17032 62592
rect 17096 62528 17112 62592
rect 17176 62528 17192 62592
rect 17256 62528 17264 62592
rect 16944 61504 17264 62528
rect 16944 61440 16952 61504
rect 17016 61440 17032 61504
rect 17096 61440 17112 61504
rect 17176 61440 17192 61504
rect 17256 61440 17264 61504
rect 16944 60416 17264 61440
rect 16944 60352 16952 60416
rect 17016 60352 17032 60416
rect 17096 60352 17112 60416
rect 17176 60352 17192 60416
rect 17256 60352 17264 60416
rect 16435 60076 16501 60077
rect 16435 60012 16436 60076
rect 16500 60012 16501 60076
rect 16435 60011 16501 60012
rect 15883 49604 15949 49605
rect 15883 49540 15884 49604
rect 15948 49540 15949 49604
rect 15883 49539 15949 49540
rect 16067 48380 16133 48381
rect 16067 48316 16068 48380
rect 16132 48316 16133 48380
rect 16067 48315 16133 48316
rect 15699 11116 15765 11117
rect 15699 11052 15700 11116
rect 15764 11052 15765 11116
rect 15699 11051 15765 11052
rect 15147 10572 15213 10573
rect 15147 10508 15148 10572
rect 15212 10508 15213 10572
rect 15147 10507 15213 10508
rect 14227 8260 14293 8261
rect 14227 8196 14228 8260
rect 14292 8196 14293 8260
rect 14227 8195 14293 8196
rect 13307 6900 13373 6901
rect 13307 6836 13308 6900
rect 13372 6836 13373 6900
rect 13307 6835 13373 6836
rect 16070 6765 16130 48315
rect 16438 21045 16498 60011
rect 16944 59328 17264 60352
rect 16944 59264 16952 59328
rect 17016 59264 17032 59328
rect 17096 59264 17112 59328
rect 17176 59264 17192 59328
rect 17256 59264 17264 59328
rect 16944 58294 17264 59264
rect 16944 58240 16986 58294
rect 17222 58240 17264 58294
rect 16944 58176 16952 58240
rect 17256 58176 17264 58240
rect 16944 58058 16986 58176
rect 17222 58058 17264 58176
rect 16944 57152 17264 58058
rect 16944 57088 16952 57152
rect 17016 57088 17032 57152
rect 17096 57088 17112 57152
rect 17176 57088 17192 57152
rect 17256 57088 17264 57152
rect 16944 56064 17264 57088
rect 16944 56000 16952 56064
rect 17016 56000 17032 56064
rect 17096 56000 17112 56064
rect 17176 56000 17192 56064
rect 17256 56000 17264 56064
rect 16619 55724 16685 55725
rect 16619 55660 16620 55724
rect 16684 55660 16685 55724
rect 16619 55659 16685 55660
rect 16435 21044 16501 21045
rect 16435 20980 16436 21044
rect 16500 20980 16501 21044
rect 16435 20979 16501 20980
rect 16622 7989 16682 55659
rect 16944 54976 17264 56000
rect 16944 54912 16952 54976
rect 17016 54912 17032 54976
rect 17096 54912 17112 54976
rect 17176 54912 17192 54976
rect 17256 54912 17264 54976
rect 16944 53888 17264 54912
rect 16944 53824 16952 53888
rect 17016 53824 17032 53888
rect 17096 53824 17112 53888
rect 17176 53824 17192 53888
rect 17256 53824 17264 53888
rect 16944 53294 17264 53824
rect 16944 53058 16986 53294
rect 17222 53058 17264 53294
rect 16944 52800 17264 53058
rect 16944 52736 16952 52800
rect 17016 52736 17032 52800
rect 17096 52736 17112 52800
rect 17176 52736 17192 52800
rect 17256 52736 17264 52800
rect 16944 51712 17264 52736
rect 16944 51648 16952 51712
rect 17016 51648 17032 51712
rect 17096 51648 17112 51712
rect 17176 51648 17192 51712
rect 17256 51648 17264 51712
rect 16944 50624 17264 51648
rect 16944 50560 16952 50624
rect 17016 50560 17032 50624
rect 17096 50560 17112 50624
rect 17176 50560 17192 50624
rect 17256 50560 17264 50624
rect 16944 49536 17264 50560
rect 16944 49472 16952 49536
rect 17016 49472 17032 49536
rect 17096 49472 17112 49536
rect 17176 49472 17192 49536
rect 17256 49472 17264 49536
rect 16944 48448 17264 49472
rect 16944 48384 16952 48448
rect 17016 48384 17032 48448
rect 17096 48384 17112 48448
rect 17176 48384 17192 48448
rect 17256 48384 17264 48448
rect 16944 48294 17264 48384
rect 16944 48058 16986 48294
rect 17222 48058 17264 48294
rect 16944 47360 17264 48058
rect 16944 47296 16952 47360
rect 17016 47296 17032 47360
rect 17096 47296 17112 47360
rect 17176 47296 17192 47360
rect 17256 47296 17264 47360
rect 16944 46272 17264 47296
rect 16944 46208 16952 46272
rect 17016 46208 17032 46272
rect 17096 46208 17112 46272
rect 17176 46208 17192 46272
rect 17256 46208 17264 46272
rect 16944 45184 17264 46208
rect 16944 45120 16952 45184
rect 17016 45120 17032 45184
rect 17096 45120 17112 45184
rect 17176 45120 17192 45184
rect 17256 45120 17264 45184
rect 16944 44096 17264 45120
rect 16944 44032 16952 44096
rect 17016 44032 17032 44096
rect 17096 44032 17112 44096
rect 17176 44032 17192 44096
rect 17256 44032 17264 44096
rect 16944 43294 17264 44032
rect 16944 43058 16986 43294
rect 17222 43058 17264 43294
rect 16944 43008 17264 43058
rect 16944 42944 16952 43008
rect 17016 42944 17032 43008
rect 17096 42944 17112 43008
rect 17176 42944 17192 43008
rect 17256 42944 17264 43008
rect 16944 41920 17264 42944
rect 16944 41856 16952 41920
rect 17016 41856 17032 41920
rect 17096 41856 17112 41920
rect 17176 41856 17192 41920
rect 17256 41856 17264 41920
rect 16944 40832 17264 41856
rect 16944 40768 16952 40832
rect 17016 40768 17032 40832
rect 17096 40768 17112 40832
rect 17176 40768 17192 40832
rect 17256 40768 17264 40832
rect 16944 39744 17264 40768
rect 16944 39680 16952 39744
rect 17016 39680 17032 39744
rect 17096 39680 17112 39744
rect 17176 39680 17192 39744
rect 17256 39680 17264 39744
rect 16944 38656 17264 39680
rect 16944 38592 16952 38656
rect 17016 38592 17032 38656
rect 17096 38592 17112 38656
rect 17176 38592 17192 38656
rect 17256 38592 17264 38656
rect 16944 38294 17264 38592
rect 16944 38058 16986 38294
rect 17222 38058 17264 38294
rect 16944 37568 17264 38058
rect 16944 37504 16952 37568
rect 17016 37504 17032 37568
rect 17096 37504 17112 37568
rect 17176 37504 17192 37568
rect 17256 37504 17264 37568
rect 16944 36480 17264 37504
rect 16944 36416 16952 36480
rect 17016 36416 17032 36480
rect 17096 36416 17112 36480
rect 17176 36416 17192 36480
rect 17256 36416 17264 36480
rect 16944 35392 17264 36416
rect 16944 35328 16952 35392
rect 17016 35328 17032 35392
rect 17096 35328 17112 35392
rect 17176 35328 17192 35392
rect 17256 35328 17264 35392
rect 16944 34304 17264 35328
rect 16944 34240 16952 34304
rect 17016 34240 17032 34304
rect 17096 34240 17112 34304
rect 17176 34240 17192 34304
rect 17256 34240 17264 34304
rect 16944 33294 17264 34240
rect 16944 33216 16986 33294
rect 17222 33216 17264 33294
rect 16944 33152 16952 33216
rect 17256 33152 17264 33216
rect 16944 33058 16986 33152
rect 17222 33058 17264 33152
rect 16944 32128 17264 33058
rect 16944 32064 16952 32128
rect 17016 32064 17032 32128
rect 17096 32064 17112 32128
rect 17176 32064 17192 32128
rect 17256 32064 17264 32128
rect 16944 31040 17264 32064
rect 16944 30976 16952 31040
rect 17016 30976 17032 31040
rect 17096 30976 17112 31040
rect 17176 30976 17192 31040
rect 17256 30976 17264 31040
rect 16944 29952 17264 30976
rect 16944 29888 16952 29952
rect 17016 29888 17032 29952
rect 17096 29888 17112 29952
rect 17176 29888 17192 29952
rect 17256 29888 17264 29952
rect 16944 28864 17264 29888
rect 16944 28800 16952 28864
rect 17016 28800 17032 28864
rect 17096 28800 17112 28864
rect 17176 28800 17192 28864
rect 17256 28800 17264 28864
rect 16944 28294 17264 28800
rect 16944 28058 16986 28294
rect 17222 28058 17264 28294
rect 16944 27776 17264 28058
rect 16944 27712 16952 27776
rect 17016 27712 17032 27776
rect 17096 27712 17112 27776
rect 17176 27712 17192 27776
rect 17256 27712 17264 27776
rect 16944 26688 17264 27712
rect 16944 26624 16952 26688
rect 17016 26624 17032 26688
rect 17096 26624 17112 26688
rect 17176 26624 17192 26688
rect 17256 26624 17264 26688
rect 16944 25600 17264 26624
rect 16944 25536 16952 25600
rect 17016 25536 17032 25600
rect 17096 25536 17112 25600
rect 17176 25536 17192 25600
rect 17256 25536 17264 25600
rect 16944 24512 17264 25536
rect 16944 24448 16952 24512
rect 17016 24448 17032 24512
rect 17096 24448 17112 24512
rect 17176 24448 17192 24512
rect 17256 24448 17264 24512
rect 16944 23424 17264 24448
rect 16944 23360 16952 23424
rect 17016 23360 17032 23424
rect 17096 23360 17112 23424
rect 17176 23360 17192 23424
rect 17256 23360 17264 23424
rect 16944 23294 17264 23360
rect 16944 23058 16986 23294
rect 17222 23058 17264 23294
rect 16944 22336 17264 23058
rect 16944 22272 16952 22336
rect 17016 22272 17032 22336
rect 17096 22272 17112 22336
rect 17176 22272 17192 22336
rect 17256 22272 17264 22336
rect 16944 21248 17264 22272
rect 16944 21184 16952 21248
rect 17016 21184 17032 21248
rect 17096 21184 17112 21248
rect 17176 21184 17192 21248
rect 17256 21184 17264 21248
rect 16944 20160 17264 21184
rect 16944 20096 16952 20160
rect 17016 20096 17032 20160
rect 17096 20096 17112 20160
rect 17176 20096 17192 20160
rect 17256 20096 17264 20160
rect 16944 19072 17264 20096
rect 16944 19008 16952 19072
rect 17016 19008 17032 19072
rect 17096 19008 17112 19072
rect 17176 19008 17192 19072
rect 17256 19008 17264 19072
rect 16944 18294 17264 19008
rect 16944 18058 16986 18294
rect 17222 18058 17264 18294
rect 16944 17984 17264 18058
rect 16944 17920 16952 17984
rect 17016 17920 17032 17984
rect 17096 17920 17112 17984
rect 17176 17920 17192 17984
rect 17256 17920 17264 17984
rect 16944 16896 17264 17920
rect 16944 16832 16952 16896
rect 17016 16832 17032 16896
rect 17096 16832 17112 16896
rect 17176 16832 17192 16896
rect 17256 16832 17264 16896
rect 16944 15808 17264 16832
rect 16944 15744 16952 15808
rect 17016 15744 17032 15808
rect 17096 15744 17112 15808
rect 17176 15744 17192 15808
rect 17256 15744 17264 15808
rect 16944 14720 17264 15744
rect 16944 14656 16952 14720
rect 17016 14656 17032 14720
rect 17096 14656 17112 14720
rect 17176 14656 17192 14720
rect 17256 14656 17264 14720
rect 16944 13632 17264 14656
rect 16944 13568 16952 13632
rect 17016 13568 17032 13632
rect 17096 13568 17112 13632
rect 17176 13568 17192 13632
rect 17256 13568 17264 13632
rect 16944 13294 17264 13568
rect 16944 13058 16986 13294
rect 17222 13058 17264 13294
rect 16944 12544 17264 13058
rect 16944 12480 16952 12544
rect 17016 12480 17032 12544
rect 17096 12480 17112 12544
rect 17176 12480 17192 12544
rect 17256 12480 17264 12544
rect 16944 11456 17264 12480
rect 16944 11392 16952 11456
rect 17016 11392 17032 11456
rect 17096 11392 17112 11456
rect 17176 11392 17192 11456
rect 17256 11392 17264 11456
rect 16944 10368 17264 11392
rect 16944 10304 16952 10368
rect 17016 10304 17032 10368
rect 17096 10304 17112 10368
rect 17176 10304 17192 10368
rect 17256 10304 17264 10368
rect 16944 9280 17264 10304
rect 16944 9216 16952 9280
rect 17016 9216 17032 9280
rect 17096 9216 17112 9280
rect 17176 9216 17192 9280
rect 17256 9216 17264 9280
rect 16944 8294 17264 9216
rect 16944 8192 16986 8294
rect 17222 8192 17264 8294
rect 16944 8128 16952 8192
rect 17256 8128 17264 8192
rect 16944 8058 16986 8128
rect 17222 8058 17264 8128
rect 16619 7988 16685 7989
rect 16619 7924 16620 7988
rect 16684 7924 16685 7988
rect 16619 7923 16685 7924
rect 16944 7104 17264 8058
rect 16944 7040 16952 7104
rect 17016 7040 17032 7104
rect 17096 7040 17112 7104
rect 17176 7040 17192 7104
rect 17256 7040 17264 7104
rect 16067 6764 16133 6765
rect 16067 6700 16068 6764
rect 16132 6700 16133 6764
rect 16067 6699 16133 6700
rect 12604 6496 12612 6560
rect 12676 6496 12692 6560
rect 12756 6496 12772 6560
rect 12836 6496 12852 6560
rect 12916 6496 12924 6560
rect 12604 5472 12924 6496
rect 12604 5408 12612 5472
rect 12676 5408 12692 5472
rect 12756 5408 12772 5472
rect 12836 5408 12852 5472
rect 12916 5408 12924 5472
rect 12604 4384 12924 5408
rect 12604 4320 12612 4384
rect 12676 4320 12692 4384
rect 12756 4320 12772 4384
rect 12836 4320 12852 4384
rect 12916 4320 12924 4384
rect 12604 3954 12924 4320
rect 12604 3718 12646 3954
rect 12882 3718 12924 3954
rect 12604 3296 12924 3718
rect 12604 3232 12612 3296
rect 12676 3232 12692 3296
rect 12756 3232 12772 3296
rect 12836 3232 12852 3296
rect 12916 3232 12924 3296
rect 12604 2208 12924 3232
rect 12604 2144 12612 2208
rect 12676 2144 12692 2208
rect 12756 2144 12772 2208
rect 12836 2144 12852 2208
rect 12916 2144 12924 2208
rect 12604 2128 12924 2144
rect 16944 6016 17264 7040
rect 16944 5952 16952 6016
rect 17016 5952 17032 6016
rect 17096 5952 17112 6016
rect 17176 5952 17192 6016
rect 17256 5952 17264 6016
rect 16944 4928 17264 5952
rect 16944 4864 16952 4928
rect 17016 4864 17032 4928
rect 17096 4864 17112 4928
rect 17176 4864 17192 4928
rect 17256 4864 17264 4928
rect 16944 3840 17264 4864
rect 16944 3776 16952 3840
rect 17016 3776 17032 3840
rect 17096 3776 17112 3840
rect 17176 3776 17192 3840
rect 17256 3776 17264 3840
rect 16944 3294 17264 3776
rect 16944 3058 16986 3294
rect 17222 3058 17264 3294
rect 16944 2752 17264 3058
rect 16944 2688 16952 2752
rect 17016 2688 17032 2752
rect 17096 2688 17112 2752
rect 17176 2688 17192 2752
rect 17256 2688 17264 2752
rect 16944 2128 17264 2688
rect 17604 77280 17924 77840
rect 17604 77216 17612 77280
rect 17676 77216 17692 77280
rect 17756 77216 17772 77280
rect 17836 77216 17852 77280
rect 17916 77216 17924 77280
rect 17604 76192 17924 77216
rect 17604 76128 17612 76192
rect 17676 76128 17692 76192
rect 17756 76128 17772 76192
rect 17836 76128 17852 76192
rect 17916 76128 17924 76192
rect 17604 75104 17924 76128
rect 17604 75040 17612 75104
rect 17676 75040 17692 75104
rect 17756 75040 17772 75104
rect 17836 75040 17852 75104
rect 17916 75040 17924 75104
rect 17604 74016 17924 75040
rect 17604 73952 17612 74016
rect 17676 73954 17692 74016
rect 17756 73954 17772 74016
rect 17836 73954 17852 74016
rect 17916 73952 17924 74016
rect 17604 73718 17646 73952
rect 17882 73718 17924 73952
rect 17604 72928 17924 73718
rect 17604 72864 17612 72928
rect 17676 72864 17692 72928
rect 17756 72864 17772 72928
rect 17836 72864 17852 72928
rect 17916 72864 17924 72928
rect 17604 71840 17924 72864
rect 17604 71776 17612 71840
rect 17676 71776 17692 71840
rect 17756 71776 17772 71840
rect 17836 71776 17852 71840
rect 17916 71776 17924 71840
rect 17604 70752 17924 71776
rect 17604 70688 17612 70752
rect 17676 70688 17692 70752
rect 17756 70688 17772 70752
rect 17836 70688 17852 70752
rect 17916 70688 17924 70752
rect 17604 69664 17924 70688
rect 17604 69600 17612 69664
rect 17676 69600 17692 69664
rect 17756 69600 17772 69664
rect 17836 69600 17852 69664
rect 17916 69600 17924 69664
rect 17604 68954 17924 69600
rect 17604 68718 17646 68954
rect 17882 68718 17924 68954
rect 17604 68576 17924 68718
rect 17604 68512 17612 68576
rect 17676 68512 17692 68576
rect 17756 68512 17772 68576
rect 17836 68512 17852 68576
rect 17916 68512 17924 68576
rect 17604 67488 17924 68512
rect 17604 67424 17612 67488
rect 17676 67424 17692 67488
rect 17756 67424 17772 67488
rect 17836 67424 17852 67488
rect 17916 67424 17924 67488
rect 17604 66400 17924 67424
rect 17604 66336 17612 66400
rect 17676 66336 17692 66400
rect 17756 66336 17772 66400
rect 17836 66336 17852 66400
rect 17916 66336 17924 66400
rect 17604 65312 17924 66336
rect 17604 65248 17612 65312
rect 17676 65248 17692 65312
rect 17756 65248 17772 65312
rect 17836 65248 17852 65312
rect 17916 65248 17924 65312
rect 17604 64224 17924 65248
rect 17604 64160 17612 64224
rect 17676 64160 17692 64224
rect 17756 64160 17772 64224
rect 17836 64160 17852 64224
rect 17916 64160 17924 64224
rect 17604 63954 17924 64160
rect 17604 63718 17646 63954
rect 17882 63718 17924 63954
rect 17604 63136 17924 63718
rect 17604 63072 17612 63136
rect 17676 63072 17692 63136
rect 17756 63072 17772 63136
rect 17836 63072 17852 63136
rect 17916 63072 17924 63136
rect 17604 62048 17924 63072
rect 17604 61984 17612 62048
rect 17676 61984 17692 62048
rect 17756 61984 17772 62048
rect 17836 61984 17852 62048
rect 17916 61984 17924 62048
rect 17604 60960 17924 61984
rect 17604 60896 17612 60960
rect 17676 60896 17692 60960
rect 17756 60896 17772 60960
rect 17836 60896 17852 60960
rect 17916 60896 17924 60960
rect 17604 59872 17924 60896
rect 17604 59808 17612 59872
rect 17676 59808 17692 59872
rect 17756 59808 17772 59872
rect 17836 59808 17852 59872
rect 17916 59808 17924 59872
rect 17604 58954 17924 59808
rect 17604 58784 17646 58954
rect 17882 58784 17924 58954
rect 17604 58720 17612 58784
rect 17916 58720 17924 58784
rect 17604 58718 17646 58720
rect 17882 58718 17924 58720
rect 17604 57696 17924 58718
rect 17604 57632 17612 57696
rect 17676 57632 17692 57696
rect 17756 57632 17772 57696
rect 17836 57632 17852 57696
rect 17916 57632 17924 57696
rect 17604 56608 17924 57632
rect 17604 56544 17612 56608
rect 17676 56544 17692 56608
rect 17756 56544 17772 56608
rect 17836 56544 17852 56608
rect 17916 56544 17924 56608
rect 17604 55520 17924 56544
rect 17604 55456 17612 55520
rect 17676 55456 17692 55520
rect 17756 55456 17772 55520
rect 17836 55456 17852 55520
rect 17916 55456 17924 55520
rect 17604 54432 17924 55456
rect 17604 54368 17612 54432
rect 17676 54368 17692 54432
rect 17756 54368 17772 54432
rect 17836 54368 17852 54432
rect 17916 54368 17924 54432
rect 17604 53954 17924 54368
rect 17604 53718 17646 53954
rect 17882 53718 17924 53954
rect 17604 53344 17924 53718
rect 17604 53280 17612 53344
rect 17676 53280 17692 53344
rect 17756 53280 17772 53344
rect 17836 53280 17852 53344
rect 17916 53280 17924 53344
rect 17604 52256 17924 53280
rect 17604 52192 17612 52256
rect 17676 52192 17692 52256
rect 17756 52192 17772 52256
rect 17836 52192 17852 52256
rect 17916 52192 17924 52256
rect 17604 51168 17924 52192
rect 17604 51104 17612 51168
rect 17676 51104 17692 51168
rect 17756 51104 17772 51168
rect 17836 51104 17852 51168
rect 17916 51104 17924 51168
rect 17604 50080 17924 51104
rect 17604 50016 17612 50080
rect 17676 50016 17692 50080
rect 17756 50016 17772 50080
rect 17836 50016 17852 50080
rect 17916 50016 17924 50080
rect 17604 48992 17924 50016
rect 17604 48928 17612 48992
rect 17676 48954 17692 48992
rect 17756 48954 17772 48992
rect 17836 48954 17852 48992
rect 17916 48928 17924 48992
rect 17604 48718 17646 48928
rect 17882 48718 17924 48928
rect 17604 47904 17924 48718
rect 17604 47840 17612 47904
rect 17676 47840 17692 47904
rect 17756 47840 17772 47904
rect 17836 47840 17852 47904
rect 17916 47840 17924 47904
rect 17604 46816 17924 47840
rect 17604 46752 17612 46816
rect 17676 46752 17692 46816
rect 17756 46752 17772 46816
rect 17836 46752 17852 46816
rect 17916 46752 17924 46816
rect 17604 45728 17924 46752
rect 17604 45664 17612 45728
rect 17676 45664 17692 45728
rect 17756 45664 17772 45728
rect 17836 45664 17852 45728
rect 17916 45664 17924 45728
rect 17604 44640 17924 45664
rect 17604 44576 17612 44640
rect 17676 44576 17692 44640
rect 17756 44576 17772 44640
rect 17836 44576 17852 44640
rect 17916 44576 17924 44640
rect 17604 43954 17924 44576
rect 17604 43718 17646 43954
rect 17882 43718 17924 43954
rect 17604 43552 17924 43718
rect 17604 43488 17612 43552
rect 17676 43488 17692 43552
rect 17756 43488 17772 43552
rect 17836 43488 17852 43552
rect 17916 43488 17924 43552
rect 17604 42464 17924 43488
rect 17604 42400 17612 42464
rect 17676 42400 17692 42464
rect 17756 42400 17772 42464
rect 17836 42400 17852 42464
rect 17916 42400 17924 42464
rect 17604 41376 17924 42400
rect 17604 41312 17612 41376
rect 17676 41312 17692 41376
rect 17756 41312 17772 41376
rect 17836 41312 17852 41376
rect 17916 41312 17924 41376
rect 17604 40288 17924 41312
rect 17604 40224 17612 40288
rect 17676 40224 17692 40288
rect 17756 40224 17772 40288
rect 17836 40224 17852 40288
rect 17916 40224 17924 40288
rect 17604 39200 17924 40224
rect 17604 39136 17612 39200
rect 17676 39136 17692 39200
rect 17756 39136 17772 39200
rect 17836 39136 17852 39200
rect 17916 39136 17924 39200
rect 17604 38954 17924 39136
rect 17604 38718 17646 38954
rect 17882 38718 17924 38954
rect 17604 38112 17924 38718
rect 17604 38048 17612 38112
rect 17676 38048 17692 38112
rect 17756 38048 17772 38112
rect 17836 38048 17852 38112
rect 17916 38048 17924 38112
rect 17604 37024 17924 38048
rect 17604 36960 17612 37024
rect 17676 36960 17692 37024
rect 17756 36960 17772 37024
rect 17836 36960 17852 37024
rect 17916 36960 17924 37024
rect 17604 35936 17924 36960
rect 17604 35872 17612 35936
rect 17676 35872 17692 35936
rect 17756 35872 17772 35936
rect 17836 35872 17852 35936
rect 17916 35872 17924 35936
rect 17604 34848 17924 35872
rect 17604 34784 17612 34848
rect 17676 34784 17692 34848
rect 17756 34784 17772 34848
rect 17836 34784 17852 34848
rect 17916 34784 17924 34848
rect 17604 33954 17924 34784
rect 17604 33760 17646 33954
rect 17882 33760 17924 33954
rect 17604 33696 17612 33760
rect 17676 33696 17692 33718
rect 17756 33696 17772 33718
rect 17836 33696 17852 33718
rect 17916 33696 17924 33760
rect 17604 32672 17924 33696
rect 17604 32608 17612 32672
rect 17676 32608 17692 32672
rect 17756 32608 17772 32672
rect 17836 32608 17852 32672
rect 17916 32608 17924 32672
rect 17604 31584 17924 32608
rect 17604 31520 17612 31584
rect 17676 31520 17692 31584
rect 17756 31520 17772 31584
rect 17836 31520 17852 31584
rect 17916 31520 17924 31584
rect 17604 30496 17924 31520
rect 17604 30432 17612 30496
rect 17676 30432 17692 30496
rect 17756 30432 17772 30496
rect 17836 30432 17852 30496
rect 17916 30432 17924 30496
rect 17604 29408 17924 30432
rect 17604 29344 17612 29408
rect 17676 29344 17692 29408
rect 17756 29344 17772 29408
rect 17836 29344 17852 29408
rect 17916 29344 17924 29408
rect 17604 28954 17924 29344
rect 17604 28718 17646 28954
rect 17882 28718 17924 28954
rect 17604 28320 17924 28718
rect 17604 28256 17612 28320
rect 17676 28256 17692 28320
rect 17756 28256 17772 28320
rect 17836 28256 17852 28320
rect 17916 28256 17924 28320
rect 17604 27232 17924 28256
rect 17604 27168 17612 27232
rect 17676 27168 17692 27232
rect 17756 27168 17772 27232
rect 17836 27168 17852 27232
rect 17916 27168 17924 27232
rect 17604 26144 17924 27168
rect 17604 26080 17612 26144
rect 17676 26080 17692 26144
rect 17756 26080 17772 26144
rect 17836 26080 17852 26144
rect 17916 26080 17924 26144
rect 17604 25056 17924 26080
rect 17604 24992 17612 25056
rect 17676 24992 17692 25056
rect 17756 24992 17772 25056
rect 17836 24992 17852 25056
rect 17916 24992 17924 25056
rect 17604 23968 17924 24992
rect 17604 23904 17612 23968
rect 17676 23954 17692 23968
rect 17756 23954 17772 23968
rect 17836 23954 17852 23968
rect 17916 23904 17924 23968
rect 17604 23718 17646 23904
rect 17882 23718 17924 23904
rect 17604 22880 17924 23718
rect 17604 22816 17612 22880
rect 17676 22816 17692 22880
rect 17756 22816 17772 22880
rect 17836 22816 17852 22880
rect 17916 22816 17924 22880
rect 17604 21792 17924 22816
rect 17604 21728 17612 21792
rect 17676 21728 17692 21792
rect 17756 21728 17772 21792
rect 17836 21728 17852 21792
rect 17916 21728 17924 21792
rect 17604 20704 17924 21728
rect 17604 20640 17612 20704
rect 17676 20640 17692 20704
rect 17756 20640 17772 20704
rect 17836 20640 17852 20704
rect 17916 20640 17924 20704
rect 17604 19616 17924 20640
rect 17604 19552 17612 19616
rect 17676 19552 17692 19616
rect 17756 19552 17772 19616
rect 17836 19552 17852 19616
rect 17916 19552 17924 19616
rect 17604 18954 17924 19552
rect 17604 18718 17646 18954
rect 17882 18718 17924 18954
rect 17604 18528 17924 18718
rect 17604 18464 17612 18528
rect 17676 18464 17692 18528
rect 17756 18464 17772 18528
rect 17836 18464 17852 18528
rect 17916 18464 17924 18528
rect 17604 17440 17924 18464
rect 17604 17376 17612 17440
rect 17676 17376 17692 17440
rect 17756 17376 17772 17440
rect 17836 17376 17852 17440
rect 17916 17376 17924 17440
rect 17604 16352 17924 17376
rect 17604 16288 17612 16352
rect 17676 16288 17692 16352
rect 17756 16288 17772 16352
rect 17836 16288 17852 16352
rect 17916 16288 17924 16352
rect 17604 15264 17924 16288
rect 17604 15200 17612 15264
rect 17676 15200 17692 15264
rect 17756 15200 17772 15264
rect 17836 15200 17852 15264
rect 17916 15200 17924 15264
rect 17604 14176 17924 15200
rect 17604 14112 17612 14176
rect 17676 14112 17692 14176
rect 17756 14112 17772 14176
rect 17836 14112 17852 14176
rect 17916 14112 17924 14176
rect 17604 13954 17924 14112
rect 17604 13718 17646 13954
rect 17882 13718 17924 13954
rect 17604 13088 17924 13718
rect 17604 13024 17612 13088
rect 17676 13024 17692 13088
rect 17756 13024 17772 13088
rect 17836 13024 17852 13088
rect 17916 13024 17924 13088
rect 17604 12000 17924 13024
rect 17604 11936 17612 12000
rect 17676 11936 17692 12000
rect 17756 11936 17772 12000
rect 17836 11936 17852 12000
rect 17916 11936 17924 12000
rect 17604 10912 17924 11936
rect 17604 10848 17612 10912
rect 17676 10848 17692 10912
rect 17756 10848 17772 10912
rect 17836 10848 17852 10912
rect 17916 10848 17924 10912
rect 17604 9824 17924 10848
rect 17604 9760 17612 9824
rect 17676 9760 17692 9824
rect 17756 9760 17772 9824
rect 17836 9760 17852 9824
rect 17916 9760 17924 9824
rect 17604 8954 17924 9760
rect 17604 8736 17646 8954
rect 17882 8736 17924 8954
rect 17604 8672 17612 8736
rect 17676 8672 17692 8718
rect 17756 8672 17772 8718
rect 17836 8672 17852 8718
rect 17916 8672 17924 8736
rect 17604 7648 17924 8672
rect 17604 7584 17612 7648
rect 17676 7584 17692 7648
rect 17756 7584 17772 7648
rect 17836 7584 17852 7648
rect 17916 7584 17924 7648
rect 17604 6560 17924 7584
rect 17604 6496 17612 6560
rect 17676 6496 17692 6560
rect 17756 6496 17772 6560
rect 17836 6496 17852 6560
rect 17916 6496 17924 6560
rect 17604 5472 17924 6496
rect 17604 5408 17612 5472
rect 17676 5408 17692 5472
rect 17756 5408 17772 5472
rect 17836 5408 17852 5472
rect 17916 5408 17924 5472
rect 17604 4384 17924 5408
rect 17604 4320 17612 4384
rect 17676 4320 17692 4384
rect 17756 4320 17772 4384
rect 17836 4320 17852 4384
rect 17916 4320 17924 4384
rect 17604 3954 17924 4320
rect 17604 3718 17646 3954
rect 17882 3718 17924 3954
rect 17604 3296 17924 3718
rect 17604 3232 17612 3296
rect 17676 3232 17692 3296
rect 17756 3232 17772 3296
rect 17836 3232 17852 3296
rect 17916 3232 17924 3296
rect 17604 2208 17924 3232
rect 17604 2144 17612 2208
rect 17676 2144 17692 2208
rect 17756 2144 17772 2208
rect 17836 2144 17852 2208
rect 17916 2144 17924 2208
rect 17604 2128 17924 2144
<< via4 >>
rect 1986 73058 2222 73294
rect 1986 68058 2222 68294
rect 1986 63058 2222 63294
rect 1986 58240 2222 58294
rect 1986 58176 2016 58240
rect 2016 58176 2032 58240
rect 2032 58176 2096 58240
rect 2096 58176 2112 58240
rect 2112 58176 2176 58240
rect 2176 58176 2192 58240
rect 2192 58176 2222 58240
rect 1986 58058 2222 58176
rect 1986 53058 2222 53294
rect 1986 48058 2222 48294
rect 1986 43058 2222 43294
rect 1986 38058 2222 38294
rect 1986 33216 2222 33294
rect 1986 33152 2016 33216
rect 2016 33152 2032 33216
rect 2032 33152 2096 33216
rect 2096 33152 2112 33216
rect 2112 33152 2176 33216
rect 2176 33152 2192 33216
rect 2192 33152 2222 33216
rect 1986 33058 2222 33152
rect 1986 28058 2222 28294
rect 1986 23058 2222 23294
rect 1986 18058 2222 18294
rect 1986 13058 2222 13294
rect 1986 8192 2222 8294
rect 1986 8128 2016 8192
rect 2016 8128 2032 8192
rect 2032 8128 2096 8192
rect 2096 8128 2112 8192
rect 2112 8128 2176 8192
rect 2176 8128 2192 8192
rect 2192 8128 2222 8192
rect 1986 8058 2222 8128
rect 1986 3058 2222 3294
rect 2646 73952 2676 73954
rect 2676 73952 2692 73954
rect 2692 73952 2756 73954
rect 2756 73952 2772 73954
rect 2772 73952 2836 73954
rect 2836 73952 2852 73954
rect 2852 73952 2882 73954
rect 2646 73718 2882 73952
rect 2646 68718 2882 68954
rect 2646 63718 2882 63954
rect 2646 58784 2882 58954
rect 2646 58720 2676 58784
rect 2676 58720 2692 58784
rect 2692 58720 2756 58784
rect 2756 58720 2772 58784
rect 2772 58720 2836 58784
rect 2836 58720 2852 58784
rect 2852 58720 2882 58784
rect 2646 58718 2882 58720
rect 2646 53718 2882 53954
rect 2646 48928 2676 48954
rect 2676 48928 2692 48954
rect 2692 48928 2756 48954
rect 2756 48928 2772 48954
rect 2772 48928 2836 48954
rect 2836 48928 2852 48954
rect 2852 48928 2882 48954
rect 2646 48718 2882 48928
rect 2646 43718 2882 43954
rect 2646 38718 2882 38954
rect 2646 33760 2882 33954
rect 2646 33718 2676 33760
rect 2676 33718 2692 33760
rect 2692 33718 2756 33760
rect 2756 33718 2772 33760
rect 2772 33718 2836 33760
rect 2836 33718 2852 33760
rect 2852 33718 2882 33760
rect 2646 28718 2882 28954
rect 2646 23904 2676 23954
rect 2676 23904 2692 23954
rect 2692 23904 2756 23954
rect 2756 23904 2772 23954
rect 2772 23904 2836 23954
rect 2836 23904 2852 23954
rect 2852 23904 2882 23954
rect 2646 23718 2882 23904
rect 2646 18718 2882 18954
rect 2646 13718 2882 13954
rect 2646 8736 2882 8954
rect 2646 8718 2676 8736
rect 2676 8718 2692 8736
rect 2692 8718 2756 8736
rect 2756 8718 2772 8736
rect 2772 8718 2836 8736
rect 2836 8718 2852 8736
rect 2852 8718 2882 8736
rect 6986 73058 7222 73294
rect 6986 68058 7222 68294
rect 6986 63058 7222 63294
rect 6986 58240 7222 58294
rect 6986 58176 7016 58240
rect 7016 58176 7032 58240
rect 7032 58176 7096 58240
rect 7096 58176 7112 58240
rect 7112 58176 7176 58240
rect 7176 58176 7192 58240
rect 7192 58176 7222 58240
rect 6986 58058 7222 58176
rect 6986 53058 7222 53294
rect 7646 73952 7676 73954
rect 7676 73952 7692 73954
rect 7692 73952 7756 73954
rect 7756 73952 7772 73954
rect 7772 73952 7836 73954
rect 7836 73952 7852 73954
rect 7852 73952 7882 73954
rect 7646 73718 7882 73952
rect 7646 68718 7882 68954
rect 7646 63718 7882 63954
rect 7646 58784 7882 58954
rect 7646 58720 7676 58784
rect 7676 58720 7692 58784
rect 7692 58720 7756 58784
rect 7756 58720 7772 58784
rect 7772 58720 7836 58784
rect 7836 58720 7852 58784
rect 7852 58720 7882 58784
rect 7646 58718 7882 58720
rect 7646 53718 7882 53954
rect 6986 48058 7222 48294
rect 7646 48928 7676 48954
rect 7676 48928 7692 48954
rect 7692 48928 7756 48954
rect 7756 48928 7772 48954
rect 7772 48928 7836 48954
rect 7836 48928 7852 48954
rect 7852 48928 7882 48954
rect 7646 48718 7882 48928
rect 7646 43718 7882 43954
rect 6986 43058 7222 43294
rect 6986 38058 7222 38294
rect 6986 33216 7222 33294
rect 6986 33152 7016 33216
rect 7016 33152 7032 33216
rect 7032 33152 7096 33216
rect 7096 33152 7112 33216
rect 7112 33152 7176 33216
rect 7176 33152 7192 33216
rect 7192 33152 7222 33216
rect 6986 33058 7222 33152
rect 6986 28058 7222 28294
rect 6986 23058 7222 23294
rect 6986 18058 7222 18294
rect 6986 13058 7222 13294
rect 6986 8192 7222 8294
rect 6986 8128 7016 8192
rect 7016 8128 7032 8192
rect 7032 8128 7096 8192
rect 7096 8128 7112 8192
rect 7112 8128 7176 8192
rect 7176 8128 7192 8192
rect 7192 8128 7222 8192
rect 6986 8058 7222 8128
rect 2646 3718 2882 3954
rect 6986 3058 7222 3294
rect 7646 38718 7882 38954
rect 7646 33760 7882 33954
rect 7646 33718 7676 33760
rect 7676 33718 7692 33760
rect 7692 33718 7756 33760
rect 7756 33718 7772 33760
rect 7772 33718 7836 33760
rect 7836 33718 7852 33760
rect 7852 33718 7882 33760
rect 7646 28718 7882 28954
rect 7646 23904 7676 23954
rect 7676 23904 7692 23954
rect 7692 23904 7756 23954
rect 7756 23904 7772 23954
rect 7772 23904 7836 23954
rect 7836 23904 7852 23954
rect 7852 23904 7882 23954
rect 7646 23718 7882 23904
rect 7646 18718 7882 18954
rect 7646 13718 7882 13954
rect 7646 8736 7882 8954
rect 7646 8718 7676 8736
rect 7676 8718 7692 8736
rect 7692 8718 7756 8736
rect 7756 8718 7772 8736
rect 7772 8718 7836 8736
rect 7836 8718 7852 8736
rect 7852 8718 7882 8736
rect 11986 73058 12222 73294
rect 11986 68058 12222 68294
rect 11986 63058 12222 63294
rect 11986 58240 12222 58294
rect 11986 58176 12016 58240
rect 12016 58176 12032 58240
rect 12032 58176 12096 58240
rect 12096 58176 12112 58240
rect 12112 58176 12176 58240
rect 12176 58176 12192 58240
rect 12192 58176 12222 58240
rect 11986 58058 12222 58176
rect 11986 53058 12222 53294
rect 11986 48058 12222 48294
rect 11986 43058 12222 43294
rect 11986 38058 12222 38294
rect 11986 33216 12222 33294
rect 11986 33152 12016 33216
rect 12016 33152 12032 33216
rect 12032 33152 12096 33216
rect 12096 33152 12112 33216
rect 12112 33152 12176 33216
rect 12176 33152 12192 33216
rect 12192 33152 12222 33216
rect 11986 33058 12222 33152
rect 11986 28058 12222 28294
rect 11986 23058 12222 23294
rect 11986 18058 12222 18294
rect 11986 13058 12222 13294
rect 11986 8192 12222 8294
rect 11986 8128 12016 8192
rect 12016 8128 12032 8192
rect 12032 8128 12096 8192
rect 12096 8128 12112 8192
rect 12112 8128 12176 8192
rect 12176 8128 12192 8192
rect 12192 8128 12222 8192
rect 11986 8058 12222 8128
rect 7646 3718 7882 3954
rect 11986 3058 12222 3294
rect 12646 73952 12676 73954
rect 12676 73952 12692 73954
rect 12692 73952 12756 73954
rect 12756 73952 12772 73954
rect 12772 73952 12836 73954
rect 12836 73952 12852 73954
rect 12852 73952 12882 73954
rect 12646 73718 12882 73952
rect 12646 68718 12882 68954
rect 12646 63718 12882 63954
rect 12646 58784 12882 58954
rect 12646 58720 12676 58784
rect 12676 58720 12692 58784
rect 12692 58720 12756 58784
rect 12756 58720 12772 58784
rect 12772 58720 12836 58784
rect 12836 58720 12852 58784
rect 12852 58720 12882 58784
rect 12646 58718 12882 58720
rect 12646 53718 12882 53954
rect 12646 48928 12676 48954
rect 12676 48928 12692 48954
rect 12692 48928 12756 48954
rect 12756 48928 12772 48954
rect 12772 48928 12836 48954
rect 12836 48928 12852 48954
rect 12852 48928 12882 48954
rect 12646 48718 12882 48928
rect 12646 43718 12882 43954
rect 12646 38718 12882 38954
rect 12646 33760 12882 33954
rect 12646 33718 12676 33760
rect 12676 33718 12692 33760
rect 12692 33718 12756 33760
rect 12756 33718 12772 33760
rect 12772 33718 12836 33760
rect 12836 33718 12852 33760
rect 12852 33718 12882 33760
rect 12646 28718 12882 28954
rect 12646 23904 12676 23954
rect 12676 23904 12692 23954
rect 12692 23904 12756 23954
rect 12756 23904 12772 23954
rect 12772 23904 12836 23954
rect 12836 23904 12852 23954
rect 12852 23904 12882 23954
rect 12646 23718 12882 23904
rect 12646 18718 12882 18954
rect 12646 13718 12882 13954
rect 12646 8736 12882 8954
rect 12646 8718 12676 8736
rect 12676 8718 12692 8736
rect 12692 8718 12756 8736
rect 12756 8718 12772 8736
rect 12772 8718 12836 8736
rect 12836 8718 12852 8736
rect 12852 8718 12882 8736
rect 16986 73058 17222 73294
rect 16986 68058 17222 68294
rect 16986 63058 17222 63294
rect 16986 58240 17222 58294
rect 16986 58176 17016 58240
rect 17016 58176 17032 58240
rect 17032 58176 17096 58240
rect 17096 58176 17112 58240
rect 17112 58176 17176 58240
rect 17176 58176 17192 58240
rect 17192 58176 17222 58240
rect 16986 58058 17222 58176
rect 16986 53058 17222 53294
rect 16986 48058 17222 48294
rect 16986 43058 17222 43294
rect 16986 38058 17222 38294
rect 16986 33216 17222 33294
rect 16986 33152 17016 33216
rect 17016 33152 17032 33216
rect 17032 33152 17096 33216
rect 17096 33152 17112 33216
rect 17112 33152 17176 33216
rect 17176 33152 17192 33216
rect 17192 33152 17222 33216
rect 16986 33058 17222 33152
rect 16986 28058 17222 28294
rect 16986 23058 17222 23294
rect 16986 18058 17222 18294
rect 16986 13058 17222 13294
rect 16986 8192 17222 8294
rect 16986 8128 17016 8192
rect 17016 8128 17032 8192
rect 17032 8128 17096 8192
rect 17096 8128 17112 8192
rect 17112 8128 17176 8192
rect 17176 8128 17192 8192
rect 17192 8128 17222 8192
rect 16986 8058 17222 8128
rect 12646 3718 12882 3954
rect 16986 3058 17222 3294
rect 17646 73952 17676 73954
rect 17676 73952 17692 73954
rect 17692 73952 17756 73954
rect 17756 73952 17772 73954
rect 17772 73952 17836 73954
rect 17836 73952 17852 73954
rect 17852 73952 17882 73954
rect 17646 73718 17882 73952
rect 17646 68718 17882 68954
rect 17646 63718 17882 63954
rect 17646 58784 17882 58954
rect 17646 58720 17676 58784
rect 17676 58720 17692 58784
rect 17692 58720 17756 58784
rect 17756 58720 17772 58784
rect 17772 58720 17836 58784
rect 17836 58720 17852 58784
rect 17852 58720 17882 58784
rect 17646 58718 17882 58720
rect 17646 53718 17882 53954
rect 17646 48928 17676 48954
rect 17676 48928 17692 48954
rect 17692 48928 17756 48954
rect 17756 48928 17772 48954
rect 17772 48928 17836 48954
rect 17836 48928 17852 48954
rect 17852 48928 17882 48954
rect 17646 48718 17882 48928
rect 17646 43718 17882 43954
rect 17646 38718 17882 38954
rect 17646 33760 17882 33954
rect 17646 33718 17676 33760
rect 17676 33718 17692 33760
rect 17692 33718 17756 33760
rect 17756 33718 17772 33760
rect 17772 33718 17836 33760
rect 17836 33718 17852 33760
rect 17852 33718 17882 33760
rect 17646 28718 17882 28954
rect 17646 23904 17676 23954
rect 17676 23904 17692 23954
rect 17692 23904 17756 23954
rect 17756 23904 17772 23954
rect 17772 23904 17836 23954
rect 17836 23904 17852 23954
rect 17852 23904 17882 23954
rect 17646 23718 17882 23904
rect 17646 18718 17882 18954
rect 17646 13718 17882 13954
rect 17646 8736 17882 8954
rect 17646 8718 17676 8736
rect 17676 8718 17692 8736
rect 17692 8718 17756 8736
rect 17756 8718 17772 8736
rect 17772 8718 17836 8736
rect 17836 8718 17852 8736
rect 17852 8718 17882 8736
rect 17646 3718 17882 3954
<< metal5 >>
rect 1056 73954 18908 73996
rect 1056 73718 2646 73954
rect 2882 73718 7646 73954
rect 7882 73718 12646 73954
rect 12882 73718 17646 73954
rect 17882 73718 18908 73954
rect 1056 73676 18908 73718
rect 1056 73294 18908 73336
rect 1056 73058 1986 73294
rect 2222 73058 6986 73294
rect 7222 73058 11986 73294
rect 12222 73058 16986 73294
rect 17222 73058 18908 73294
rect 1056 73016 18908 73058
rect 1056 68954 18908 68996
rect 1056 68718 2646 68954
rect 2882 68718 7646 68954
rect 7882 68718 12646 68954
rect 12882 68718 17646 68954
rect 17882 68718 18908 68954
rect 1056 68676 18908 68718
rect 1056 68294 18908 68336
rect 1056 68058 1986 68294
rect 2222 68058 6986 68294
rect 7222 68058 11986 68294
rect 12222 68058 16986 68294
rect 17222 68058 18908 68294
rect 1056 68016 18908 68058
rect 1056 63954 18908 63996
rect 1056 63718 2646 63954
rect 2882 63718 7646 63954
rect 7882 63718 12646 63954
rect 12882 63718 17646 63954
rect 17882 63718 18908 63954
rect 1056 63676 18908 63718
rect 1056 63294 18908 63336
rect 1056 63058 1986 63294
rect 2222 63058 6986 63294
rect 7222 63058 11986 63294
rect 12222 63058 16986 63294
rect 17222 63058 18908 63294
rect 1056 63016 18908 63058
rect 1056 58954 18908 58996
rect 1056 58718 2646 58954
rect 2882 58718 7646 58954
rect 7882 58718 12646 58954
rect 12882 58718 17646 58954
rect 17882 58718 18908 58954
rect 1056 58676 18908 58718
rect 1056 58294 18908 58336
rect 1056 58058 1986 58294
rect 2222 58058 6986 58294
rect 7222 58058 11986 58294
rect 12222 58058 16986 58294
rect 17222 58058 18908 58294
rect 1056 58016 18908 58058
rect 1056 53954 18908 53996
rect 1056 53718 2646 53954
rect 2882 53718 7646 53954
rect 7882 53718 12646 53954
rect 12882 53718 17646 53954
rect 17882 53718 18908 53954
rect 1056 53676 18908 53718
rect 1056 53294 18908 53336
rect 1056 53058 1986 53294
rect 2222 53058 6986 53294
rect 7222 53058 11986 53294
rect 12222 53058 16986 53294
rect 17222 53058 18908 53294
rect 1056 53016 18908 53058
rect 1056 48954 18908 48996
rect 1056 48718 2646 48954
rect 2882 48718 7646 48954
rect 7882 48718 12646 48954
rect 12882 48718 17646 48954
rect 17882 48718 18908 48954
rect 1056 48676 18908 48718
rect 1056 48294 18908 48336
rect 1056 48058 1986 48294
rect 2222 48058 6986 48294
rect 7222 48058 11986 48294
rect 12222 48058 16986 48294
rect 17222 48058 18908 48294
rect 1056 48016 18908 48058
rect 1056 43954 18908 43996
rect 1056 43718 2646 43954
rect 2882 43718 7646 43954
rect 7882 43718 12646 43954
rect 12882 43718 17646 43954
rect 17882 43718 18908 43954
rect 1056 43676 18908 43718
rect 1056 43294 18908 43336
rect 1056 43058 1986 43294
rect 2222 43058 6986 43294
rect 7222 43058 11986 43294
rect 12222 43058 16986 43294
rect 17222 43058 18908 43294
rect 1056 43016 18908 43058
rect 1056 38954 18908 38996
rect 1056 38718 2646 38954
rect 2882 38718 7646 38954
rect 7882 38718 12646 38954
rect 12882 38718 17646 38954
rect 17882 38718 18908 38954
rect 1056 38676 18908 38718
rect 1056 38294 18908 38336
rect 1056 38058 1986 38294
rect 2222 38058 6986 38294
rect 7222 38058 11986 38294
rect 12222 38058 16986 38294
rect 17222 38058 18908 38294
rect 1056 38016 18908 38058
rect 1056 33954 18908 33996
rect 1056 33718 2646 33954
rect 2882 33718 7646 33954
rect 7882 33718 12646 33954
rect 12882 33718 17646 33954
rect 17882 33718 18908 33954
rect 1056 33676 18908 33718
rect 1056 33294 18908 33336
rect 1056 33058 1986 33294
rect 2222 33058 6986 33294
rect 7222 33058 11986 33294
rect 12222 33058 16986 33294
rect 17222 33058 18908 33294
rect 1056 33016 18908 33058
rect 1056 28954 18908 28996
rect 1056 28718 2646 28954
rect 2882 28718 7646 28954
rect 7882 28718 12646 28954
rect 12882 28718 17646 28954
rect 17882 28718 18908 28954
rect 1056 28676 18908 28718
rect 1056 28294 18908 28336
rect 1056 28058 1986 28294
rect 2222 28058 6986 28294
rect 7222 28058 11986 28294
rect 12222 28058 16986 28294
rect 17222 28058 18908 28294
rect 1056 28016 18908 28058
rect 1056 23954 18908 23996
rect 1056 23718 2646 23954
rect 2882 23718 7646 23954
rect 7882 23718 12646 23954
rect 12882 23718 17646 23954
rect 17882 23718 18908 23954
rect 1056 23676 18908 23718
rect 1056 23294 18908 23336
rect 1056 23058 1986 23294
rect 2222 23058 6986 23294
rect 7222 23058 11986 23294
rect 12222 23058 16986 23294
rect 17222 23058 18908 23294
rect 1056 23016 18908 23058
rect 1056 18954 18908 18996
rect 1056 18718 2646 18954
rect 2882 18718 7646 18954
rect 7882 18718 12646 18954
rect 12882 18718 17646 18954
rect 17882 18718 18908 18954
rect 1056 18676 18908 18718
rect 1056 18294 18908 18336
rect 1056 18058 1986 18294
rect 2222 18058 6986 18294
rect 7222 18058 11986 18294
rect 12222 18058 16986 18294
rect 17222 18058 18908 18294
rect 1056 18016 18908 18058
rect 1056 13954 18908 13996
rect 1056 13718 2646 13954
rect 2882 13718 7646 13954
rect 7882 13718 12646 13954
rect 12882 13718 17646 13954
rect 17882 13718 18908 13954
rect 1056 13676 18908 13718
rect 1056 13294 18908 13336
rect 1056 13058 1986 13294
rect 2222 13058 6986 13294
rect 7222 13058 11986 13294
rect 12222 13058 16986 13294
rect 17222 13058 18908 13294
rect 1056 13016 18908 13058
rect 1056 8954 18908 8996
rect 1056 8718 2646 8954
rect 2882 8718 7646 8954
rect 7882 8718 12646 8954
rect 12882 8718 17646 8954
rect 17882 8718 18908 8954
rect 1056 8676 18908 8718
rect 1056 8294 18908 8336
rect 1056 8058 1986 8294
rect 2222 8058 6986 8294
rect 7222 8058 11986 8294
rect 12222 8058 16986 8294
rect 17222 8058 18908 8294
rect 1056 8016 18908 8058
rect 1056 3954 18908 3996
rect 1056 3718 2646 3954
rect 2882 3718 7646 3954
rect 7882 3718 12646 3954
rect 12882 3718 17646 3954
rect 17882 3718 18908 3954
rect 1056 3676 18908 3718
rect 1056 3294 18908 3336
rect 1056 3058 1986 3294
rect 2222 3058 6986 3294
rect 7222 3058 11986 3294
rect 12222 3058 16986 3294
rect 17222 3058 18908 3294
rect 1056 3016 18908 3058
use sky130_fd_sc_hd__buf_6  _168_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 12972 0 1 44608
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _169_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 9108 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _170_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 5336 0 1 28288
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  _171_
timestamp 1694700623
transform 1 0 6532 0 -1 47872
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _172_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 6532 0 -1 75072
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _173_
timestamp 1694700623
transform 1 0 12236 0 -1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _174_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 3220 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _175_
timestamp 1694700623
transform 1 0 12328 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _176_
timestamp 1694700623
transform 1 0 4968 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _177_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 17572 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _178_
timestamp 1694700623
transform 1 0 2300 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _179_
timestamp 1694700623
transform 1 0 17572 0 -1 67456
box -38 -48 866 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _180_
timestamp 1694700623
transform 1 0 15456 0 -1 40256
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  _181_
timestamp 1694700623
transform 1 0 5060 0 1 75072
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _182_
timestamp 1694700623
transform 1 0 14260 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_4  _183_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 11500 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _184_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 12236 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _185_
timestamp 1694700623
transform 1 0 7820 0 1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _186_
timestamp 1694700623
transform 1 0 10028 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _187_
timestamp 1694700623
transform 1 0 12328 0 1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _188_
timestamp 1694700623
transform 1 0 6532 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  _189_
timestamp 1694700623
transform 1 0 11408 0 1 55488
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _190_
timestamp 1694700623
transform 1 0 4692 0 -1 75072
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _191_
timestamp 1694700623
transform 1 0 15180 0 1 75072
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _192_
timestamp 1694700623
transform 1 0 8924 0 -1 60928
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _193_
timestamp 1694700623
transform 1 0 11868 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _194_
timestamp 1694700623
transform 1 0 3956 0 1 65280
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _195_
timestamp 1694700623
transform 1 0 7636 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _196_
timestamp 1694700623
transform 1 0 9108 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _197_
timestamp 1694700623
transform 1 0 12420 0 1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _198_
timestamp 1694700623
transform 1 0 2208 0 1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _199_
timestamp 1694700623
transform 1 0 15548 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _200_
timestamp 1694700623
transform 1 0 9384 0 -1 53312
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _201_
timestamp 1694700623
transform 1 0 8280 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _202_
timestamp 1694700623
transform 1 0 9844 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _203_
timestamp 1694700623
transform 1 0 1564 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _204_
timestamp 1694700623
transform 1 0 12972 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _205_
timestamp 1694700623
transform 1 0 17756 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_2  _206_
timestamp 1694700623
transform 1 0 16836 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _207_
timestamp 1694700623
transform 1 0 4140 0 1 62016
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _208_
timestamp 1694700623
transform 1 0 16836 0 -1 55488
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _209_
timestamp 1694700623
transform 1 0 14996 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  _210_
timestamp 1694700623
transform 1 0 17572 0 -1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _211_
timestamp 1694700623
transform 1 0 9108 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _212_
timestamp 1694700623
transform 1 0 5704 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _213_
timestamp 1694700623
transform 1 0 8096 0 -1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _214_
timestamp 1694700623
transform 1 0 7268 0 1 58752
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_2  _215_
timestamp 1694700623
transform 1 0 14720 0 1 58752
box -38 -48 866 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _216_
timestamp 1694700623
transform 1 0 9108 0 1 11968
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  _217_
timestamp 1694700623
transform 1 0 15640 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _218_
timestamp 1694700623
transform 1 0 2208 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _219_
timestamp 1694700623
transform 1 0 16100 0 1 59840
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _220_
timestamp 1694700623
transform 1 0 3956 0 1 69632
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _221_
timestamp 1694700623
transform 1 0 16928 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _222_
timestamp 1694700623
transform 1 0 4324 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _223_
timestamp 1694700623
transform 1 0 14260 0 -1 48960
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _224_
timestamp 1694700623
transform 1 0 16836 0 -1 75072
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _225_
timestamp 1694700623
transform 1 0 11868 0 -1 64192
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _226_
timestamp 1694700623
transform 1 0 6164 0 1 63104
box -38 -48 406 592
use sky130_fd_sc_hd__buf_6  _227_
timestamp 1694700623
transform 1 0 5060 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _228_
timestamp 1694700623
transform 1 0 6716 0 1 43520
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _229_
timestamp 1694700623
transform 1 0 11960 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _230_
timestamp 1694700623
transform 1 0 13708 0 -1 76160
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _231_
timestamp 1694700623
transform 1 0 16376 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _232_
timestamp 1694700623
transform 1 0 1564 0 -1 53312
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _233_
timestamp 1694700623
transform 1 0 8004 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _234_
timestamp 1694700623
transform 1 0 11684 0 -1 62016
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _235_
timestamp 1694700623
transform 1 0 16284 0 1 63104
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _236_
timestamp 1694700623
transform 1 0 1564 0 -1 44608
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _237_
timestamp 1694700623
transform 1 0 17940 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_2  _238_
timestamp 1694700623
transform 1 0 17388 0 -1 66368
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _239_
timestamp 1694700623
transform 1 0 8004 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _240_
timestamp 1694700623
transform 1 0 2668 0 1 50048
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _241_
timestamp 1694700623
transform 1 0 11684 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _242_
timestamp 1694700623
transform 1 0 12972 0 1 42432
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _243_
timestamp 1694700623
transform 1 0 4784 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _244_
timestamp 1694700623
transform 1 0 9108 0 -1 42432
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _245_
timestamp 1694700623
transform 1 0 8464 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_2  _246_
timestamp 1694700623
transform 1 0 6808 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _247_
timestamp 1694700623
transform 1 0 15824 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  _248_
timestamp 1694700623
transform 1 0 3128 0 -1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_2  _249_
timestamp 1694700623
transform 1 0 1932 0 1 69632
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _250_
timestamp 1694700623
transform 1 0 9660 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_2  _251_
timestamp 1694700623
transform 1 0 2668 0 1 46784
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _252_
timestamp 1694700623
transform 1 0 4140 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _253_
timestamp 1694700623
transform 1 0 15548 0 -1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _254_
timestamp 1694700623
transform 1 0 14352 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _255_
timestamp 1694700623
transform 1 0 6532 0 -1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _256_
timestamp 1694700623
transform 1 0 18032 0 -1 65280
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _257_
timestamp 1694700623
transform 1 0 12604 0 1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _258_
timestamp 1694700623
transform 1 0 17756 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_4  _259_
timestamp 1694700623
transform 1 0 6532 0 -1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_2  _260_
timestamp 1694700623
transform 1 0 14076 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _261_
timestamp 1694700623
transform 1 0 12972 0 1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _262_
timestamp 1694700623
transform 1 0 18032 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _263_
timestamp 1694700623
transform 1 0 14444 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _264_
timestamp 1694700623
transform 1 0 16100 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _265_
timestamp 1694700623
transform 1 0 6900 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _266_
timestamp 1694700623
transform 1 0 2944 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _267_
timestamp 1694700623
transform 1 0 12512 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _268_
timestamp 1694700623
transform 1 0 6992 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  _269_
timestamp 1694700623
transform 1 0 14904 0 1 69632
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _270_
timestamp 1694700623
transform 1 0 7912 0 -1 65280
box -38 -48 866 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _271_
timestamp 1694700623
transform 1 0 9108 0 1 69632
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_2  _272_
timestamp 1694700623
transform 1 0 1564 0 1 56576
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _273_
timestamp 1694700623
transform 1 0 9108 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_2  _274_
timestamp 1694700623
transform 1 0 9200 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _275_
timestamp 1694700623
transform 1 0 11500 0 1 76160
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_2  _276_
timestamp 1694700623
transform 1 0 1564 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _277_
timestamp 1694700623
transform 1 0 7912 0 -1 67456
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _278_
timestamp 1694700623
transform 1 0 11776 0 1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _279_
timestamp 1694700623
transform 1 0 2208 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_2  _280_
timestamp 1694700623
transform 1 0 1564 0 1 42432
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _281_
timestamp 1694700623
transform 1 0 16836 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _282_
timestamp 1694700623
transform 1 0 10304 0 -1 48960
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _283_
timestamp 1694700623
transform 1 0 10580 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _284_
timestamp 1694700623
transform 1 0 12052 0 1 73984
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _285_
timestamp 1694700623
transform 1 0 17020 0 1 71808
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _286_
timestamp 1694700623
transform 1 0 5428 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _287_
timestamp 1694700623
transform 1 0 9752 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _288_
timestamp 1694700623
transform 1 0 17112 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _289_
timestamp 1694700623
transform 1 0 12420 0 -1 56576
box -38 -48 958 592
use sky130_fd_sc_hd__buf_6  _290_
timestamp 1694700623
transform 1 0 14536 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _291_
timestamp 1694700623
transform 1 0 5704 0 1 41344
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _292_
timestamp 1694700623
transform 1 0 15272 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _293_
timestamp 1694700623
transform 1 0 9108 0 1 59840
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _294_
timestamp 1694700623
transform 1 0 11868 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _295_
timestamp 1694700623
transform 1 0 9568 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _296_
timestamp 1694700623
transform 1 0 2760 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _297_
timestamp 1694700623
transform 1 0 5704 0 1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _298_
timestamp 1694700623
transform 1 0 6624 0 1 25024
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  _299_
timestamp 1694700623
transform 1 0 10488 0 1 42432
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _300_
timestamp 1694700623
transform 1 0 16836 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_4  _301_
timestamp 1694700623
transform 1 0 14260 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_2  _302_
timestamp 1694700623
transform 1 0 8648 0 -1 76160
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _303_
timestamp 1694700623
transform 1 0 7544 0 1 59840
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _304_
timestamp 1694700623
transform 1 0 12236 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_2  _305_
timestamp 1694700623
transform 1 0 2300 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _306_
timestamp 1694700623
transform 1 0 8372 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _307_
timestamp 1694700623
transform 1 0 10120 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _308_
timestamp 1694700623
transform 1 0 12788 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _309_
timestamp 1694700623
transform 1 0 10212 0 -1 54400
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _310_
timestamp 1694700623
transform 1 0 7360 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _311_
timestamp 1694700623
transform 1 0 7820 0 -1 40256
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _312_
timestamp 1694700623
transform 1 0 3956 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _313_
timestamp 1694700623
transform 1 0 17572 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _314_
timestamp 1694700623
transform 1 0 14260 0 1 51136
box -38 -48 958 592
use sky130_fd_sc_hd__buf_6  _315_
timestamp 1694700623
transform 1 0 9936 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_2  _316_
timestamp 1694700623
transform 1 0 16008 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _317_
timestamp 1694700623
transform 1 0 7452 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _318_
timestamp 1694700623
transform 1 0 12788 0 -1 72896
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _319_
timestamp 1694700623
transform 1 0 2392 0 1 64192
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _320_
timestamp 1694700623
transform 1 0 7268 0 -1 73984
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _321_
timestamp 1694700623
transform 1 0 7544 0 1 75072
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _322_
timestamp 1694700623
transform 1 0 17296 0 -1 57664
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _323_
timestamp 1694700623
transform 1 0 14260 0 1 63104
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_4  _324_
timestamp 1694700623
transform 1 0 6624 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _325_
timestamp 1694700623
transform 1 0 17388 0 -1 77248
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  _326_
timestamp 1694700623
transform 1 0 6808 0 -1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _327_
timestamp 1694700623
transform 1 0 9016 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_4  _328_
timestamp 1694700623
transform 1 0 7452 0 1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_2  _329_
timestamp 1694700623
transform 1 0 2484 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _330_
timestamp 1694700623
transform 1 0 15364 0 -1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _331_
timestamp 1694700623
transform 1 0 5428 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_2  _332_
timestamp 1694700623
transform 1 0 2668 0 -1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _333_
timestamp 1694700623
transform 1 0 14352 0 -1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_2  _334_
timestamp 1694700623
transform 1 0 16744 0 1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _335_
timestamp 1694700623
transform 1 0 9752 0 -1 4352
box -38 -48 958 592
use sky130_fd_sc_hd__dfxtp_2  _336_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 2484 0 -1 3264
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _337_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 9568 0 -1 40256
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _338_
timestamp 1694700623
transform 1 0 15456 0 1 14144
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _339_
timestamp 1694700623
transform 1 0 15732 0 1 20672
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _340_
timestamp 1694700623
transform 1 0 4324 0 -1 44608
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _341_
timestamp 1694700623
transform 1 0 11776 0 1 64192
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_4  _342_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 14260 0 1 44608
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_2  _343_
timestamp 1694700623
transform 1 0 6532 0 -1 63104
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _344_
timestamp 1694700623
transform 1 0 3220 0 -1 59840
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _345_
timestamp 1694700623
transform 1 0 10764 0 1 11968
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _346_
timestamp 1694700623
transform 1 0 5980 0 1 70720
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _347_
timestamp 1694700623
transform 1 0 13248 0 -1 27200
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _348_
timestamp 1694700623
transform 1 0 7912 0 -1 23936
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _349_
timestamp 1694700623
transform 1 0 2208 0 -1 55488
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _350_
timestamp 1694700623
transform 1 0 14260 0 1 52224
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _351_
timestamp 1694700623
transform 1 0 9108 0 1 70720
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _352_
timestamp 1694700623
transform 1 0 8740 0 -1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _353_
timestamp 1694700623
transform 1 0 9108 0 1 68544
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _354_
timestamp 1694700623
transform 1 0 11684 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _355_
timestamp 1694700623
transform 1 0 8004 0 -1 50048
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _356_
timestamp 1694700623
transform 1 0 12236 0 1 3264
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _357_
timestamp 1694700623
transform 1 0 14536 0 -1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _358_
timestamp 1694700623
transform 1 0 1932 0 1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _359_
timestamp 1694700623
transform 1 0 14812 0 -1 75072
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _360_
timestamp 1694700623
transform 1 0 3128 0 -1 13056
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _361_
timestamp 1694700623
transform 1 0 7084 0 1 69632
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _362_
timestamp 1694700623
transform 1 0 6900 0 1 20672
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _363_
timestamp 1694700623
transform 1 0 16836 0 -1 31552
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _364_
timestamp 1694700623
transform 1 0 13892 0 -1 18496
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _365_
timestamp 1694700623
transform 1 0 5980 0 1 48960
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _366_
timestamp 1694700623
transform 1 0 14904 0 1 76160
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _367_
timestamp 1694700623
transform 1 0 14260 0 1 68544
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _368_
timestamp 1694700623
transform 1 0 12972 0 -1 65280
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _369_
timestamp 1694700623
transform 1 0 7728 0 -1 30464
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _370_
timestamp 1694700623
transform 1 0 14260 0 1 73984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _371_
timestamp 1694700623
transform 1 0 9108 0 1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _372_
timestamp 1694700623
transform 1 0 7084 0 1 16320
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _373_
timestamp 1694700623
transform 1 0 3956 0 1 51136
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _374_
timestamp 1694700623
transform 1 0 15456 0 1 70720
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _375_
timestamp 1694700623
transform 1 0 6624 0 1 72896
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _376_
timestamp 1694700623
transform 1 0 9568 0 -1 8704
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _377_
timestamp 1694700623
transform 1 0 11960 0 -1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _378_
timestamp 1694700623
transform 1 0 2760 0 -1 57664
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _379_
timestamp 1694700623
transform 1 0 3404 0 -1 48960
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _380_
timestamp 1694700623
transform 1 0 14260 0 1 59840
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _381_
timestamp 1694700623
transform 1 0 15548 0 1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _382_
timestamp 1694700623
transform 1 0 16836 0 1 15232
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _383_
timestamp 1694700623
transform 1 0 5060 0 1 5440
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _384_
timestamp 1694700623
transform 1 0 7268 0 -1 42432
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _385_
timestamp 1694700623
transform 1 0 15916 0 1 60928
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _386_
timestamp 1694700623
transform 1 0 3680 0 -1 39168
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _387_
timestamp 1694700623
transform 1 0 6532 0 -1 4352
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _388_
timestamp 1694700623
transform 1 0 3128 0 -1 56576
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _389_
timestamp 1694700623
transform 1 0 9016 0 -1 51136
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _390_
timestamp 1694700623
transform 1 0 1656 0 1 55488
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _391_
timestamp 1694700623
transform 1 0 3956 0 -1 76160
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _392_
timestamp 1694700623
transform 1 0 13340 0 -1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _393_
timestamp 1694700623
transform 1 0 16836 0 -1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _394_
timestamp 1694700623
transform 1 0 2024 0 1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _395_
timestamp 1694700623
transform 1 0 12880 0 -1 47872
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _396_
timestamp 1694700623
transform 1 0 4048 0 -1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _397_
timestamp 1694700623
transform 1 0 10396 0 1 51136
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _398_
timestamp 1694700623
transform 1 0 16836 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _399_
timestamp 1694700623
transform 1 0 5152 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _400_
timestamp 1694700623
transform 1 0 3036 0 -1 71808
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _401_
timestamp 1694700623
transform 1 0 3036 0 -1 50048
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _402_
timestamp 1694700623
transform 1 0 12236 0 -1 46784
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _403_
timestamp 1694700623
transform 1 0 13064 0 -1 35904
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _404_
timestamp 1694700623
transform 1 0 13524 0 -1 66368
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _405_
timestamp 1694700623
transform 1 0 10580 0 1 17408
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _406_
timestamp 1694700623
transform 1 0 9660 0 -1 69632
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _407_
timestamp 1694700623
transform 1 0 2116 0 -1 42432
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _408_
timestamp 1694700623
transform -1 0 4324 0 -1 9792
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_4  _409_
timestamp 1694700623
transform 1 0 2300 0 -1 8704
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_2  _410_
timestamp 1694700623
transform 1 0 12328 0 -1 53312
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _411_
timestamp 1694700623
transform 1 0 5980 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _412_
timestamp 1694700623
transform 1 0 6532 0 -1 60928
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_4  _413_
timestamp 1694700623
transform 1 0 11684 0 -1 5440
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_2  _414_
timestamp 1694700623
transform 1 0 3956 0 1 25024
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _415_
timestamp 1694700623
transform 1 0 5520 0 1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 9660 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp 1694700623
transform 1 0 10580 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_3
timestamp 1694700623
transform 1 0 2852 0 -1 59840
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_4
timestamp 1694700623
transform 1 0 4876 0 -1 59840
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_5
timestamp 1694700623
transform 1 0 4508 0 1 69632
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_6
timestamp 1694700623
transform 1 0 3312 0 1 69632
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_7
timestamp 1694700623
transform 1 0 4876 0 1 69632
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_8
timestamp 1694700623
transform 1 0 2944 0 1 69632
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_9
timestamp 1694700623
transform 1 0 2760 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_10
timestamp 1694700623
transform 1 0 4876 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_11
timestamp 1694700623
transform 1 0 2392 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_12
timestamp 1694700623
transform 1 0 5244 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_13
timestamp 1694700623
transform 1 0 6532 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_14
timestamp 1694700623
transform 1 0 6164 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_15
timestamp 1694700623
transform 1 0 12236 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_16
timestamp 1694700623
transform 1 0 11040 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_17
timestamp 1694700623
transform 1 0 12604 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_18
timestamp 1694700623
transform 1 0 15916 0 1 73984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_19
timestamp 1694700623
transform 1 0 13616 0 1 73984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_20
timestamp 1694700623
transform 1 0 16284 0 1 73984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_21
timestamp 1694700623
transform 1 0 4692 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_22
timestamp 1694700623
transform 1 0 5060 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_23
timestamp 1694700623
transform 1 0 3312 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_24
timestamp 1694700623
transform 1 0 5428 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_25
timestamp 1694700623
transform 1 0 2944 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_26
timestamp 1694700623
transform 1 0 6256 0 1 72896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_27
timestamp 1694700623
transform 1 0 8280 0 1 72896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_28
timestamp 1694700623
transform 1 0 5888 0 1 72896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_29
timestamp 1694700623
transform 1 0 5520 0 1 72896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_30
timestamp 1694700623
transform 1 0 9108 0 1 72896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_31
timestamp 1694700623
transform 1 0 13708 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_32
timestamp 1694700623
transform 1 0 3036 0 -1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_33
timestamp 1694700623
transform 1 0 8556 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_34
timestamp 1694700623
transform 1 0 9660 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_35
timestamp 1694700623
transform 1 0 15548 0 1 60928
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_36
timestamp 1694700623
transform 1 0 17572 0 1 60928
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_37
timestamp 1694700623
transform 1 0 1840 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_38
timestamp 1694700623
transform 1 0 2760 0 -1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_39
timestamp 1694700623
transform 1 0 17388 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_40
timestamp 1694700623
transform 1 0 8648 0 -1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_41
timestamp 1694700623
transform 1 0 4784 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_42
timestamp 1694700623
transform 1 0 7176 0 1 75072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_43
timestamp 1694700623
transform -1 0 2576 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_44
timestamp 1694700623
transform -1 0 4692 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_45
timestamp 1694700623
transform 1 0 1748 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_46
timestamp 1694700623
transform 1 0 3036 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_47
timestamp 1694700623
transform 1 0 1748 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_48
timestamp 1694700623
transform 1 0 8280 0 -1 60928
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_49
timestamp 1694700623
transform 1 0 5888 0 -1 60928
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_50
timestamp 1694700623
transform 1 0 8648 0 -1 60928
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_51
timestamp 1694700623
transform 1 0 5060 0 -1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_52
timestamp 1694700623
transform 1 0 4692 0 -1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_53
timestamp 1694700623
transform 1 0 13616 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_54
timestamp 1694700623
transform 1 0 11040 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_55
timestamp 1694700623
transform 1 0 11132 0 1 65280
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_56
timestamp 1694700623
transform 1 0 11868 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_57
timestamp 1694700623
transform 1 0 12052 0 1 67456
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_58
timestamp 1694700623
transform 1 0 14352 0 1 58752
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_59
timestamp 1694700623
transform 1 0 10212 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_60
timestamp 1694700623
transform 1 0 11132 0 1 76160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_61
timestamp 1694700623
transform 1 0 18216 0 1 76160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_62
timestamp 1694700623
transform 1 0 12880 0 -1 64192
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_63
timestamp 1694700623
transform 1 0 13248 0 -1 64192
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_64
timestamp 1694700623
transform 1 0 11040 0 -1 64192
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_65
timestamp 1694700623
transform 1 0 13616 0 -1 64192
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_66
timestamp 1694700623
transform 1 0 10672 0 -1 64192
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_67
timestamp 1694700623
transform 1 0 7084 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_68
timestamp 1694700623
transform 1 0 5888 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_69
timestamp 1694700623
transform 1 0 7452 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_70
timestamp 1694700623
transform 1 0 5520 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_71
timestamp 1694700623
transform 1 0 7820 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_72
timestamp 1694700623
transform 1 0 2576 0 1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_73
timestamp 1694700623
transform 1 0 2576 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_74
timestamp 1694700623
transform 1 0 11408 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_75
timestamp 1694700623
transform 1 0 2576 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_76
timestamp 1694700623
transform 1 0 9844 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_77
timestamp 1694700623
transform 1 0 11868 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_78
timestamp 1694700623
transform 1 0 12788 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_79
timestamp 1694700623
transform 1 0 11500 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_80
timestamp 1694700623
transform 1 0 13156 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_81
timestamp 1694700623
transform 1 0 8280 0 -1 63104
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_82
timestamp 1694700623
transform 1 0 5888 0 -1 63104
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_83
timestamp 1694700623
transform 1 0 8648 0 -1 63104
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_84
timestamp 1694700623
transform 1 0 5520 0 -1 63104
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_85
timestamp 1694700623
transform 1 0 9292 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_86
timestamp 1694700623
transform 1 0 2484 0 -1 59840
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_87
timestamp 1694700623
transform 1 0 8464 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_88
timestamp 1694700623
transform 1 0 10948 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_89
timestamp 1694700623
transform 1 0 2116 0 -1 59840
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_90
timestamp 1694700623
transform 1 0 5244 0 -1 59840
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_91
timestamp 1694700623
transform 1 0 7636 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_92
timestamp 1694700623
transform 1 0 8556 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_93
timestamp 1694700623
transform 1 0 7268 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_94
timestamp 1694700623
transform 1 0 8924 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_95
timestamp 1694700623
transform 1 0 6900 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_96
timestamp 1694700623
transform 1 0 14536 0 -1 77248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_97
timestamp 1694700623
transform 1 0 16836 0 1 77248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_98
timestamp 1694700623
transform 1 0 14168 0 -1 77248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_99
timestamp 1694700623
transform 1 0 17204 0 1 77248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_100
timestamp 1694700623
transform 1 0 13800 0 -1 77248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_101
timestamp 1694700623
transform 1 0 2392 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_102
timestamp 1694700623
transform 1 0 8280 0 -1 76160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_103
timestamp 1694700623
transform 1 0 9200 0 -1 76160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_104
timestamp 1694700623
transform 1 0 6808 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_105
timestamp 1694700623
transform 1 0 4416 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_106
timestamp 1694700623
transform 1 0 4048 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_107
timestamp 1694700623
transform 1 0 3312 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_108
timestamp 1694700623
transform 1 0 8096 0 1 75072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_109
timestamp 1694700623
transform -1 0 2208 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_110
timestamp 1694700623
transform 1 0 6808 0 1 75072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_111
timestamp 1694700623
transform -1 0 1840 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_112
timestamp 1694700623
transform -1 0 5060 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_113
timestamp 1694700623
transform 1 0 1932 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_114
timestamp 1694700623
transform 1 0 6532 0 -1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_115
timestamp 1694700623
transform 1 0 13984 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_116
timestamp 1694700623
transform 1 0 4324 0 -1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_117
timestamp 1694700623
transform 1 0 3956 0 -1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_118
timestamp 1694700623
transform 1 0 14352 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_119
timestamp 1694700623
transform 1 0 10672 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_120
timestamp 1694700623
transform 1 0 15732 0 1 58752
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_121
timestamp 1694700623
transform 1 0 8464 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_122
timestamp 1694700623
transform 1 0 13616 0 1 58752
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_123
timestamp 1694700623
transform 1 0 10580 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_124
timestamp 1694700623
transform 1 0 2116 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_125
timestamp 1694700623
transform 1 0 6072 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_126
timestamp 1694700623
transform 1 0 17204 0 -1 67456
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_127
timestamp 1694700623
transform 1 0 4876 0 1 75072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_128
timestamp 1694700623
transform 1 0 16928 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_129
timestamp 1694700623
transform 1 0 7084 0 1 76160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_130
timestamp 1694700623
transform 1 0 14996 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_131
timestamp 1694700623
transform 1 0 17664 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_132
timestamp 1694700623
transform 1 0 16192 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_133
timestamp 1694700623
transform 1 0 10672 0 -1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_134
timestamp 1694700623
transform 1 0 17756 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_135
timestamp 1694700623
transform 1 0 8280 0 -1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_136
timestamp 1694700623
transform 1 0 8464 0 1 75072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_137
timestamp 1694700623
transform -1 0 5428 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_138
timestamp 1694700623
transform 1 0 6440 0 1 75072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_139
timestamp 1694700623
transform 1 0 4784 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_140
timestamp 1694700623
transform -1 0 5796 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_141
timestamp 1694700623
transform 1 0 9108 0 1 75072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_142
timestamp 1694700623
transform 1 0 4416 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_143
timestamp 1694700623
transform 1 0 6072 0 1 75072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_144
timestamp 1694700623
transform 1 0 4048 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_145
timestamp 1694700623
transform -1 0 6716 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_146
timestamp 1694700623
transform 1 0 6256 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_147
timestamp 1694700623
transform 1 0 7912 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_148
timestamp 1694700623
transform 1 0 5888 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_149
timestamp 1694700623
transform 1 0 17020 0 -1 77248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_150
timestamp 1694700623
transform 1 0 16192 0 -1 77248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_151
timestamp 1694700623
transform 1 0 15824 0 -1 77248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_152
timestamp 1694700623
transform 1 0 17848 0 1 76160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_153
timestamp 1694700623
transform 1 0 17480 0 1 76160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_154
timestamp 1694700623
transform 1 0 17112 0 1 76160
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 1380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15
timestamp 1694700623
transform 1 0 2484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29
timestamp 1694700623
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 4876 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47
timestamp 1694700623
transform 1 0 5428 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_50 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 5704 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_54
timestamp 1694700623
transform 1 0 6072 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_57
timestamp 1694700623
transform 1 0 6348 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_63
timestamp 1694700623
transform 1 0 6900 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_67
timestamp 1694700623
transform 1 0 7268 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_71
timestamp 1694700623
transform 1 0 7636 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_75 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 8004 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_83
timestamp 1694700623
transform 1 0 8740 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85
timestamp 1694700623
transform 1 0 8924 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_101
timestamp 1694700623
transform 1 0 10396 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_109 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 11132 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113
timestamp 1694700623
transform 1 0 11500 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_125
timestamp 1694700623
transform 1 0 12604 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_137
timestamp 1694700623
transform 1 0 13708 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_141
timestamp 1694700623
transform 1 0 14076 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_149
timestamp 1694700623
transform 1 0 14812 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_161
timestamp 1694700623
transform 1 0 15916 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_167
timestamp 1694700623
transform 1 0 16468 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_169
timestamp 1694700623
transform 1 0 16652 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_181
timestamp 1694700623
transform 1 0 17756 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_188
timestamp 1694700623
transform 1 0 18400 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3
timestamp 1694700623
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_32
timestamp 1694700623
transform 1 0 4048 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_44
timestamp 1694700623
transform 1 0 5152 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_57
timestamp 1694700623
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_69
timestamp 1694700623
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_81
timestamp 1694700623
transform 1 0 8556 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_93
timestamp 1694700623
transform 1 0 9660 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_105
timestamp 1694700623
transform 1 0 10764 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_111
timestamp 1694700623
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_113
timestamp 1694700623
transform 1 0 11500 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_125
timestamp 1694700623
transform 1 0 12604 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_137
timestamp 1694700623
transform 1 0 13708 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_149
timestamp 1694700623
transform 1 0 14812 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_161
timestamp 1694700623
transform 1 0 15916 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_167
timestamp 1694700623
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_169
timestamp 1694700623
transform 1 0 16652 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_1_181
timestamp 1694700623
transform 1 0 17756 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_188
timestamp 1694700623
transform 1 0 18400 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3
timestamp 1694700623
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_15
timestamp 1694700623
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp 1694700623
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_29
timestamp 1694700623
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_41
timestamp 1694700623
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_53
timestamp 1694700623
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_65
timestamp 1694700623
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_77
timestamp 1694700623
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_83
timestamp 1694700623
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_85
timestamp 1694700623
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_97
timestamp 1694700623
transform 1 0 10028 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_109
timestamp 1694700623
transform 1 0 11132 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_2_138
timestamp 1694700623
transform 1 0 13800 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_2_141
timestamp 1694700623
transform 1 0 14076 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_153
timestamp 1694700623
transform 1 0 15180 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_165
timestamp 1694700623
transform 1 0 16284 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_177
timestamp 1694700623
transform 1 0 17388 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_189
timestamp 1694700623
transform 1 0 18492 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3
timestamp 1694700623
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_15
timestamp 1694700623
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_27
timestamp 1694700623
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_39
timestamp 1694700623
transform 1 0 4692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_51 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_55
timestamp 1694700623
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_57
timestamp 1694700623
transform 1 0 6348 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_3_76
timestamp 1694700623
transform 1 0 8096 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_88
timestamp 1694700623
transform 1 0 9200 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_3_104
timestamp 1694700623
transform 1 0 10672 0 -1 4352
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_3_113
timestamp 1694700623
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_125
timestamp 1694700623
transform 1 0 12604 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_137
timestamp 1694700623
transform 1 0 13708 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_149
timestamp 1694700623
transform 1 0 14812 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_161
timestamp 1694700623
transform 1 0 15916 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_167
timestamp 1694700623
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_169
timestamp 1694700623
transform 1 0 16652 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_181
timestamp 1694700623
transform 1 0 17756 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_189
timestamp 1694700623
transform 1 0 18492 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3
timestamp 1694700623
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_15
timestamp 1694700623
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 1694700623
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_29
timestamp 1694700623
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_41
timestamp 1694700623
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_53
timestamp 1694700623
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_65
timestamp 1694700623
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_77
timestamp 1694700623
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_83
timestamp 1694700623
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_85
timestamp 1694700623
transform 1 0 8924 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_4_93
timestamp 1694700623
transform 1 0 9660 0 1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_4_105
timestamp 1694700623
transform 1 0 10764 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_117
timestamp 1694700623
transform 1 0 11868 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_129
timestamp 1694700623
transform 1 0 12972 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_4_137
timestamp 1694700623
transform 1 0 13708 0 1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_4_141
timestamp 1694700623
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_153
timestamp 1694700623
transform 1 0 15180 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_165
timestamp 1694700623
transform 1 0 16284 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_177
timestamp 1694700623
transform 1 0 17388 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_189
timestamp 1694700623
transform 1 0 18492 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3
timestamp 1694700623
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_15
timestamp 1694700623
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_27
timestamp 1694700623
transform 1 0 3588 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_39
timestamp 1694700623
transform 1 0 4692 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_5_47
timestamp 1694700623
transform 1 0 5428 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_53
timestamp 1694700623
transform 1 0 5980 0 -1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_5_57
timestamp 1694700623
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_69
timestamp 1694700623
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_81
timestamp 1694700623
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_93
timestamp 1694700623
transform 1 0 9660 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_5_101
timestamp 1694700623
transform 1 0 10396 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_106
timestamp 1694700623
transform 1 0 10856 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_110
timestamp 1694700623
transform 1 0 11224 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_113
timestamp 1694700623
transform 1 0 11500 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_134
timestamp 1694700623
transform 1 0 13432 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_138
timestamp 1694700623
transform 1 0 13800 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_142
timestamp 1694700623
transform 1 0 14168 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_5_146
timestamp 1694700623
transform 1 0 14536 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_158
timestamp 1694700623
transform 1 0 15640 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_5_166
timestamp 1694700623
transform 1 0 16376 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_169
timestamp 1694700623
transform 1 0 16652 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_175
timestamp 1694700623
transform 1 0 17204 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_179
timestamp 1694700623
transform 1 0 17572 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_5_183
timestamp 1694700623
transform 1 0 17940 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_188
timestamp 1694700623
transform 1 0 18400 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3
timestamp 1694700623
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_15
timestamp 1694700623
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 1694700623
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_29
timestamp 1694700623
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_6_41
timestamp 1694700623
transform 1 0 4876 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_60
timestamp 1694700623
transform 1 0 6624 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_72
timestamp 1694700623
transform 1 0 7728 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_85
timestamp 1694700623
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_97
timestamp 1694700623
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_109
timestamp 1694700623
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_121
timestamp 1694700623
transform 1 0 12236 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_133
timestamp 1694700623
transform 1 0 13340 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_139
timestamp 1694700623
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_141
timestamp 1694700623
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_153
timestamp 1694700623
transform 1 0 15180 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_165
timestamp 1694700623
transform 1 0 16284 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_177
timestamp 1694700623
transform 1 0 17388 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_189
timestamp 1694700623
transform 1 0 18492 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3
timestamp 1694700623
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_15
timestamp 1694700623
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_27
timestamp 1694700623
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_39
timestamp 1694700623
transform 1 0 4692 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_51
timestamp 1694700623
transform 1 0 5796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_55
timestamp 1694700623
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_57
timestamp 1694700623
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_69
timestamp 1694700623
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_81
timestamp 1694700623
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_93
timestamp 1694700623
transform 1 0 9660 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_105
timestamp 1694700623
transform 1 0 10764 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_111
timestamp 1694700623
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_113
timestamp 1694700623
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_125
timestamp 1694700623
transform 1 0 12604 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_137
timestamp 1694700623
transform 1 0 13708 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_149
timestamp 1694700623
transform 1 0 14812 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_161
timestamp 1694700623
transform 1 0 15916 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_167
timestamp 1694700623
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_169
timestamp 1694700623
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_181
timestamp 1694700623
transform 1 0 17756 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_189
timestamp 1694700623
transform 1 0 18492 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3
timestamp 1694700623
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_15
timestamp 1694700623
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 1694700623
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_29
timestamp 1694700623
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_41
timestamp 1694700623
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_53
timestamp 1694700623
transform 1 0 5980 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_61
timestamp 1694700623
transform 1 0 6716 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_71
timestamp 1694700623
transform 1 0 7636 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp 1694700623
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_85
timestamp 1694700623
transform 1 0 8924 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_96
timestamp 1694700623
transform 1 0 9936 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_108
timestamp 1694700623
transform 1 0 11040 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_120
timestamp 1694700623
transform 1 0 12144 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_132
timestamp 1694700623
transform 1 0 13248 0 1 6528
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_8_141
timestamp 1694700623
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_153
timestamp 1694700623
transform 1 0 15180 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_165
timestamp 1694700623
transform 1 0 16284 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_177
timestamp 1694700623
transform 1 0 17388 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_183
timestamp 1694700623
transform 1 0 17940 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_188
timestamp 1694700623
transform 1 0 18400 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3
timestamp 1694700623
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_15
timestamp 1694700623
transform 1 0 2484 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_27
timestamp 1694700623
transform 1 0 3588 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_39
timestamp 1694700623
transform 1 0 4692 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_51
timestamp 1694700623
transform 1 0 5796 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_55
timestamp 1694700623
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_57
timestamp 1694700623
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_69
timestamp 1694700623
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_81
timestamp 1694700623
transform 1 0 8556 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_93
timestamp 1694700623
transform 1 0 9660 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_105
timestamp 1694700623
transform 1 0 10764 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_111
timestamp 1694700623
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_113
timestamp 1694700623
transform 1 0 11500 0 -1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_9_119
timestamp 1694700623
transform 1 0 12052 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_131
timestamp 1694700623
transform 1 0 13156 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_9_139
timestamp 1694700623
transform 1 0 13892 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_145
timestamp 1694700623
transform 1 0 14444 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_157
timestamp 1694700623
transform 1 0 15548 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_9_165
timestamp 1694700623
transform 1 0 16284 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_169
timestamp 1694700623
transform 1 0 16652 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_181
timestamp 1694700623
transform 1 0 17756 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_189
timestamp 1694700623
transform 1 0 18492 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3
timestamp 1694700623
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_15
timestamp 1694700623
transform 1 0 2484 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_19
timestamp 1694700623
transform 1 0 2852 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_22
timestamp 1694700623
transform 1 0 3128 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_26
timestamp 1694700623
transform 1 0 3496 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_29
timestamp 1694700623
transform 1 0 3772 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_37
timestamp 1694700623
transform 1 0 4508 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_41
timestamp 1694700623
transform 1 0 4876 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_45
timestamp 1694700623
transform 1 0 5244 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_49
timestamp 1694700623
transform 1 0 5612 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_61
timestamp 1694700623
transform 1 0 6716 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_73
timestamp 1694700623
transform 1 0 7820 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_10_81
timestamp 1694700623
transform 1 0 8556 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_85
timestamp 1694700623
transform 1 0 8924 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_96
timestamp 1694700623
transform 1 0 9936 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_108
timestamp 1694700623
transform 1 0 11040 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_112
timestamp 1694700623
transform 1 0 11408 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_115
timestamp 1694700623
transform 1 0 11684 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_119
timestamp 1694700623
transform 1 0 12052 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_125
timestamp 1694700623
transform 1 0 12604 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_129
timestamp 1694700623
transform 1 0 12972 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_10_133
timestamp 1694700623
transform 1 0 13340 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_139
timestamp 1694700623
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_141
timestamp 1694700623
transform 1 0 14076 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_153
timestamp 1694700623
transform 1 0 15180 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_165
timestamp 1694700623
transform 1 0 16284 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_177
timestamp 1694700623
transform 1 0 17388 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_189
timestamp 1694700623
transform 1 0 18492 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_11_3
timestamp 1694700623
transform 1 0 1380 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_11_11
timestamp 1694700623
transform 1 0 2116 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_11_32
timestamp 1694700623
transform 1 0 4048 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_44
timestamp 1694700623
transform 1 0 5152 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_57
timestamp 1694700623
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_69
timestamp 1694700623
transform 1 0 7452 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_81
timestamp 1694700623
transform 1 0 8556 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_11_89
timestamp 1694700623
transform 1 0 9292 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_109
timestamp 1694700623
transform 1 0 11132 0 -1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_11_113
timestamp 1694700623
transform 1 0 11500 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_125
timestamp 1694700623
transform 1 0 12604 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_137
timestamp 1694700623
transform 1 0 13708 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_143
timestamp 1694700623
transform 1 0 14260 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_154
timestamp 1694700623
transform 1 0 15272 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_11_166
timestamp 1694700623
transform 1 0 16376 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_11_169
timestamp 1694700623
transform 1 0 16652 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_185
timestamp 1694700623
transform 1 0 18124 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_189
timestamp 1694700623
transform 1 0 18492 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3
timestamp 1694700623
transform 1 0 1380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_15
timestamp 1694700623
transform 1 0 2484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_27
timestamp 1694700623
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_12_29
timestamp 1694700623
transform 1 0 3772 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_34
timestamp 1694700623
transform 1 0 4232 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_38
timestamp 1694700623
transform 1 0 4600 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_12_42
timestamp 1694700623
transform 1 0 4968 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_52
timestamp 1694700623
transform 1 0 5888 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_64
timestamp 1694700623
transform 1 0 6992 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_12_72
timestamp 1694700623
transform 1 0 7728 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_78
timestamp 1694700623
transform 1 0 8280 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_82
timestamp 1694700623
transform 1 0 8648 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_85
timestamp 1694700623
transform 1 0 8924 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_91
timestamp 1694700623
transform 1 0 9476 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_95
timestamp 1694700623
transform 1 0 9844 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_101
timestamp 1694700623
transform 1 0 10396 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_105
timestamp 1694700623
transform 1 0 10764 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_12_109
timestamp 1694700623
transform 1 0 11132 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_121
timestamp 1694700623
transform 1 0 12236 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_133
timestamp 1694700623
transform 1 0 13340 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_139
timestamp 1694700623
transform 1 0 13892 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_141
timestamp 1694700623
transform 1 0 14076 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_153
timestamp 1694700623
transform 1 0 15180 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_165
timestamp 1694700623
transform 1 0 16284 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_12_177
timestamp 1694700623
transform 1 0 17388 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_182
timestamp 1694700623
transform 1 0 17848 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_188
timestamp 1694700623
transform 1 0 18400 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_13_3
timestamp 1694700623
transform 1 0 1380 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_8
timestamp 1694700623
transform 1 0 1840 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_12
timestamp 1694700623
transform 1 0 2208 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_16
timestamp 1694700623
transform 1 0 2576 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_35
timestamp 1694700623
transform 1 0 4324 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_39
timestamp 1694700623
transform 1 0 4692 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_43
timestamp 1694700623
transform 1 0 5060 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_47
timestamp 1694700623
transform 1 0 5428 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_13_51
timestamp 1694700623
transform 1 0 5796 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_57
timestamp 1694700623
transform 1 0 6348 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_61
timestamp 1694700623
transform 1 0 6716 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_13_72
timestamp 1694700623
transform 1 0 7728 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_84
timestamp 1694700623
transform 1 0 8832 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_96
timestamp 1694700623
transform 1 0 9936 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_108
timestamp 1694700623
transform 1 0 11040 0 -1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_13_113
timestamp 1694700623
transform 1 0 11500 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_125
timestamp 1694700623
transform 1 0 12604 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_137
timestamp 1694700623
transform 1 0 13708 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_149
timestamp 1694700623
transform 1 0 14812 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_161
timestamp 1694700623
transform 1 0 15916 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_167
timestamp 1694700623
transform 1 0 16468 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_169
timestamp 1694700623
transform 1 0 16652 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_181
timestamp 1694700623
transform 1 0 17756 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_189
timestamp 1694700623
transform 1 0 18492 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_3
timestamp 1694700623
transform 1 0 1380 0 1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_14_9
timestamp 1694700623
transform 1 0 1932 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_21
timestamp 1694700623
transform 1 0 3036 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_27
timestamp 1694700623
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_29
timestamp 1694700623
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_41
timestamp 1694700623
transform 1 0 4876 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_14_45
timestamp 1694700623
transform 1 0 5244 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_51
timestamp 1694700623
transform 1 0 5796 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_54
timestamp 1694700623
transform 1 0 6072 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_58
timestamp 1694700623
transform 1 0 6440 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_72
timestamp 1694700623
transform 1 0 7728 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_14_76
timestamp 1694700623
transform 1 0 8096 0 1 9792
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_14_85
timestamp 1694700623
transform 1 0 8924 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_97
timestamp 1694700623
transform 1 0 10028 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_109
timestamp 1694700623
transform 1 0 11132 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_121
timestamp 1694700623
transform 1 0 12236 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_133
timestamp 1694700623
transform 1 0 13340 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_139
timestamp 1694700623
transform 1 0 13892 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_141
timestamp 1694700623
transform 1 0 14076 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_153
timestamp 1694700623
transform 1 0 15180 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_165
timestamp 1694700623
transform 1 0 16284 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_177
timestamp 1694700623
transform 1 0 17388 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_189
timestamp 1694700623
transform 1 0 18492 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_3
timestamp 1694700623
transform 1 0 1380 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_9
timestamp 1694700623
transform 1 0 1932 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_13
timestamp 1694700623
transform 1 0 2300 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_19
timestamp 1694700623
transform 1 0 2852 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_15_23
timestamp 1694700623
transform 1 0 3220 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_35
timestamp 1694700623
transform 1 0 4324 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_47
timestamp 1694700623
transform 1 0 5428 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_55
timestamp 1694700623
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_57
timestamp 1694700623
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_69
timestamp 1694700623
transform 1 0 7452 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_81
timestamp 1694700623
transform 1 0 8556 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_93
timestamp 1694700623
transform 1 0 9660 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_105
timestamp 1694700623
transform 1 0 10764 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_111
timestamp 1694700623
transform 1 0 11316 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_113
timestamp 1694700623
transform 1 0 11500 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_125
timestamp 1694700623
transform 1 0 12604 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_137
timestamp 1694700623
transform 1 0 13708 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_149
timestamp 1694700623
transform 1 0 14812 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_161
timestamp 1694700623
transform 1 0 15916 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_167
timestamp 1694700623
transform 1 0 16468 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_169
timestamp 1694700623
transform 1 0 16652 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_15_181
timestamp 1694700623
transform 1 0 17756 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_188
timestamp 1694700623
transform 1 0 18400 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_3
timestamp 1694700623
transform 1 0 1380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_15
timestamp 1694700623
transform 1 0 2484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_27
timestamp 1694700623
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_29
timestamp 1694700623
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_41
timestamp 1694700623
transform 1 0 4876 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_53
timestamp 1694700623
transform 1 0 5980 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_65
timestamp 1694700623
transform 1 0 7084 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_77
timestamp 1694700623
transform 1 0 8188 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_83
timestamp 1694700623
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_85
timestamp 1694700623
transform 1 0 8924 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_97
timestamp 1694700623
transform 1 0 10028 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_109
timestamp 1694700623
transform 1 0 11132 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_121
timestamp 1694700623
transform 1 0 12236 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_133
timestamp 1694700623
transform 1 0 13340 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_139
timestamp 1694700623
transform 1 0 13892 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_141
timestamp 1694700623
transform 1 0 14076 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_155
timestamp 1694700623
transform 1 0 15364 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_167
timestamp 1694700623
transform 1 0 16468 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_179
timestamp 1694700623
transform 1 0 17572 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_16_187
timestamp 1694700623
transform 1 0 18308 0 1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_17_3
timestamp 1694700623
transform 1 0 1380 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_15
timestamp 1694700623
transform 1 0 2484 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_27
timestamp 1694700623
transform 1 0 3588 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_39
timestamp 1694700623
transform 1 0 4692 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_51
timestamp 1694700623
transform 1 0 5796 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_55
timestamp 1694700623
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_57
timestamp 1694700623
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_69
timestamp 1694700623
transform 1 0 7452 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_81
timestamp 1694700623
transform 1 0 8556 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_93
timestamp 1694700623
transform 1 0 9660 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_105
timestamp 1694700623
transform 1 0 10764 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_111
timestamp 1694700623
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_113
timestamp 1694700623
transform 1 0 11500 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_125
timestamp 1694700623
transform 1 0 12604 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_137
timestamp 1694700623
transform 1 0 13708 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_149
timestamp 1694700623
transform 1 0 14812 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_161
timestamp 1694700623
transform 1 0 15916 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_167
timestamp 1694700623
transform 1 0 16468 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_169
timestamp 1694700623
transform 1 0 16652 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_181
timestamp 1694700623
transform 1 0 17756 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_189
timestamp 1694700623
transform 1 0 18492 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_3
timestamp 1694700623
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_15
timestamp 1694700623
transform 1 0 2484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp 1694700623
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_29
timestamp 1694700623
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_41
timestamp 1694700623
transform 1 0 4876 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_69
timestamp 1694700623
transform 1 0 7452 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_18_77
timestamp 1694700623
transform 1 0 8188 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_82
timestamp 1694700623
transform 1 0 8648 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_85
timestamp 1694700623
transform 1 0 8924 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_97
timestamp 1694700623
transform 1 0 10028 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_101
timestamp 1694700623
transform 1 0 10396 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_18_122
timestamp 1694700623
transform 1 0 12328 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_134
timestamp 1694700623
transform 1 0 13432 0 1 11968
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_18_141
timestamp 1694700623
transform 1 0 14076 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_153
timestamp 1694700623
transform 1 0 15180 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_165
timestamp 1694700623
transform 1 0 16284 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_177
timestamp 1694700623
transform 1 0 17388 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_183
timestamp 1694700623
transform 1 0 17940 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_188
timestamp 1694700623
transform 1 0 18400 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_19_3
timestamp 1694700623
transform 1 0 1380 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_19_11
timestamp 1694700623
transform 1 0 2116 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_16
timestamp 1694700623
transform 1 0 2576 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_20
timestamp 1694700623
transform 1 0 2944 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_39
timestamp 1694700623
transform 1 0 4692 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_43
timestamp 1694700623
transform 1 0 5060 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_19_47
timestamp 1694700623
transform 1 0 5428 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_55
timestamp 1694700623
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_57
timestamp 1694700623
transform 1 0 6348 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_69
timestamp 1694700623
transform 1 0 7452 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_81
timestamp 1694700623
transform 1 0 8556 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_93
timestamp 1694700623
transform 1 0 9660 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_105
timestamp 1694700623
transform 1 0 10764 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_111
timestamp 1694700623
transform 1 0 11316 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_113
timestamp 1694700623
transform 1 0 11500 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_125
timestamp 1694700623
transform 1 0 12604 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_137
timestamp 1694700623
transform 1 0 13708 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_149
timestamp 1694700623
transform 1 0 14812 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_161
timestamp 1694700623
transform 1 0 15916 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_167
timestamp 1694700623
transform 1 0 16468 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_169
timestamp 1694700623
transform 1 0 16652 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_187
timestamp 1694700623
transform 1 0 18308 0 -1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_20_3
timestamp 1694700623
transform 1 0 1380 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_15
timestamp 1694700623
transform 1 0 2484 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_27
timestamp 1694700623
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_29
timestamp 1694700623
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_41
timestamp 1694700623
transform 1 0 4876 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_53
timestamp 1694700623
transform 1 0 5980 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_65
timestamp 1694700623
transform 1 0 7084 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_77
timestamp 1694700623
transform 1 0 8188 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_83
timestamp 1694700623
transform 1 0 8740 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_85
timestamp 1694700623
transform 1 0 8924 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_97
timestamp 1694700623
transform 1 0 10028 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_109
timestamp 1694700623
transform 1 0 11132 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_121
timestamp 1694700623
transform 1 0 12236 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_133
timestamp 1694700623
transform 1 0 13340 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_139
timestamp 1694700623
transform 1 0 13892 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_141
timestamp 1694700623
transform 1 0 14076 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_153
timestamp 1694700623
transform 1 0 15180 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_161
timestamp 1694700623
transform 1 0 15916 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_171
timestamp 1694700623
transform 1 0 16836 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_183
timestamp 1694700623
transform 1 0 17940 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_189
timestamp 1694700623
transform 1 0 18492 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_3
timestamp 1694700623
transform 1 0 1380 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_15
timestamp 1694700623
transform 1 0 2484 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_27
timestamp 1694700623
transform 1 0 3588 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_39
timestamp 1694700623
transform 1 0 4692 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_51
timestamp 1694700623
transform 1 0 5796 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_55
timestamp 1694700623
transform 1 0 6164 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_57
timestamp 1694700623
transform 1 0 6348 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_21_62
timestamp 1694700623
transform 1 0 6808 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_74
timestamp 1694700623
transform 1 0 7912 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_86
timestamp 1694700623
transform 1 0 9016 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_98
timestamp 1694700623
transform 1 0 10120 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_21_110
timestamp 1694700623
transform 1 0 11224 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_21_113
timestamp 1694700623
transform 1 0 11500 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_125
timestamp 1694700623
transform 1 0 12604 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_137
timestamp 1694700623
transform 1 0 13708 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_149
timestamp 1694700623
transform 1 0 14812 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_161
timestamp 1694700623
transform 1 0 15916 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_167
timestamp 1694700623
transform 1 0 16468 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_169
timestamp 1694700623
transform 1 0 16652 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_181
timestamp 1694700623
transform 1 0 17756 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_189
timestamp 1694700623
transform 1 0 18492 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_3
timestamp 1694700623
transform 1 0 1380 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_15
timestamp 1694700623
transform 1 0 2484 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_27
timestamp 1694700623
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_29
timestamp 1694700623
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_41
timestamp 1694700623
transform 1 0 4876 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_53
timestamp 1694700623
transform 1 0 5980 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_65
timestamp 1694700623
transform 1 0 7084 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_22_74
timestamp 1694700623
transform 1 0 7912 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_82
timestamp 1694700623
transform 1 0 8648 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_22_85
timestamp 1694700623
transform 1 0 8924 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_97
timestamp 1694700623
transform 1 0 10028 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_109
timestamp 1694700623
transform 1 0 11132 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_121
timestamp 1694700623
transform 1 0 12236 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_133
timestamp 1694700623
transform 1 0 13340 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_139
timestamp 1694700623
transform 1 0 13892 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_141
timestamp 1694700623
transform 1 0 14076 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_22_153
timestamp 1694700623
transform 1 0 15180 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_22_173
timestamp 1694700623
transform 1 0 17020 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_22_181
timestamp 1694700623
transform 1 0 17756 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_188
timestamp 1694700623
transform 1 0 18400 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_3
timestamp 1694700623
transform 1 0 1380 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_7
timestamp 1694700623
transform 1 0 1748 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_10
timestamp 1694700623
transform 1 0 2024 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_23_16
timestamp 1694700623
transform 1 0 2576 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_28
timestamp 1694700623
transform 1 0 3680 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_40
timestamp 1694700623
transform 1 0 4784 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_52
timestamp 1694700623
transform 1 0 5888 0 -1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_23_57
timestamp 1694700623
transform 1 0 6348 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_69
timestamp 1694700623
transform 1 0 7452 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_81
timestamp 1694700623
transform 1 0 8556 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_93
timestamp 1694700623
transform 1 0 9660 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_105
timestamp 1694700623
transform 1 0 10764 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_111
timestamp 1694700623
transform 1 0 11316 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_113
timestamp 1694700623
transform 1 0 11500 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_125
timestamp 1694700623
transform 1 0 12604 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_137
timestamp 1694700623
transform 1 0 13708 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_149
timestamp 1694700623
transform 1 0 14812 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_161
timestamp 1694700623
transform 1 0 15916 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_167
timestamp 1694700623
transform 1 0 16468 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_169
timestamp 1694700623
transform 1 0 16652 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_177
timestamp 1694700623
transform 1 0 17388 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_188
timestamp 1694700623
transform 1 0 18400 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_3
timestamp 1694700623
transform 1 0 1380 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_15
timestamp 1694700623
transform 1 0 2484 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_27
timestamp 1694700623
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_29
timestamp 1694700623
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_41
timestamp 1694700623
transform 1 0 4876 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_53
timestamp 1694700623
transform 1 0 5980 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_65
timestamp 1694700623
transform 1 0 7084 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_77
timestamp 1694700623
transform 1 0 8188 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_83
timestamp 1694700623
transform 1 0 8740 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_85
timestamp 1694700623
transform 1 0 8924 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_97
timestamp 1694700623
transform 1 0 10028 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_109
timestamp 1694700623
transform 1 0 11132 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_24_120
timestamp 1694700623
transform 1 0 12144 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_24_133
timestamp 1694700623
transform 1 0 13340 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_139
timestamp 1694700623
transform 1 0 13892 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_141
timestamp 1694700623
transform 1 0 14076 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_153
timestamp 1694700623
transform 1 0 15180 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_165
timestamp 1694700623
transform 1 0 16284 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_24_188
timestamp 1694700623
transform 1 0 18400 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_25_3
timestamp 1694700623
transform 1 0 1380 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_15
timestamp 1694700623
transform 1 0 2484 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_27
timestamp 1694700623
transform 1 0 3588 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_39
timestamp 1694700623
transform 1 0 4692 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_51
timestamp 1694700623
transform 1 0 5796 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_55
timestamp 1694700623
transform 1 0 6164 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_25_57
timestamp 1694700623
transform 1 0 6348 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_25_65
timestamp 1694700623
transform 1 0 7084 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_69
timestamp 1694700623
transform 1 0 7452 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_73
timestamp 1694700623
transform 1 0 7820 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_79
timestamp 1694700623
transform 1 0 8372 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_83
timestamp 1694700623
transform 1 0 8740 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_91
timestamp 1694700623
transform 1 0 9476 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_25_95
timestamp 1694700623
transform 1 0 9844 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_107
timestamp 1694700623
transform 1 0 10948 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_111
timestamp 1694700623
transform 1 0 11316 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_113
timestamp 1694700623
transform 1 0 11500 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_125
timestamp 1694700623
transform 1 0 12604 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_137
timestamp 1694700623
transform 1 0 13708 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_149
timestamp 1694700623
transform 1 0 14812 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_161
timestamp 1694700623
transform 1 0 15916 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_167
timestamp 1694700623
transform 1 0 16468 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_169
timestamp 1694700623
transform 1 0 16652 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_25_181
timestamp 1694700623
transform 1 0 17756 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_25_188
timestamp 1694700623
transform 1 0 18400 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_26_3
timestamp 1694700623
transform 1 0 1380 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_15
timestamp 1694700623
transform 1 0 2484 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_27
timestamp 1694700623
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_29
timestamp 1694700623
transform 1 0 3772 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_41
timestamp 1694700623
transform 1 0 4876 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_26_56
timestamp 1694700623
transform 1 0 6256 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_64
timestamp 1694700623
transform 1 0 6992 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_82
timestamp 1694700623
transform 1 0 8648 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_26_85
timestamp 1694700623
transform 1 0 8924 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_97
timestamp 1694700623
transform 1 0 10028 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_109
timestamp 1694700623
transform 1 0 11132 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_121
timestamp 1694700623
transform 1 0 12236 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_133
timestamp 1694700623
transform 1 0 13340 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_139
timestamp 1694700623
transform 1 0 13892 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_141
timestamp 1694700623
transform 1 0 14076 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_153
timestamp 1694700623
transform 1 0 15180 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_165
timestamp 1694700623
transform 1 0 16284 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_177
timestamp 1694700623
transform 1 0 17388 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_185
timestamp 1694700623
transform 1 0 18124 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_189
timestamp 1694700623
transform 1 0 18492 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_3
timestamp 1694700623
transform 1 0 1380 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_15
timestamp 1694700623
transform 1 0 2484 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_27
timestamp 1694700623
transform 1 0 3588 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_39
timestamp 1694700623
transform 1 0 4692 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_51
timestamp 1694700623
transform 1 0 5796 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_55
timestamp 1694700623
transform 1 0 6164 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_57
timestamp 1694700623
transform 1 0 6348 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_69
timestamp 1694700623
transform 1 0 7452 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_81
timestamp 1694700623
transform 1 0 8556 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_93
timestamp 1694700623
transform 1 0 9660 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_101
timestamp 1694700623
transform 1 0 10396 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_107
timestamp 1694700623
transform 1 0 10948 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_111
timestamp 1694700623
transform 1 0 11316 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_113
timestamp 1694700623
transform 1 0 11500 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_125
timestamp 1694700623
transform 1 0 12604 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_137
timestamp 1694700623
transform 1 0 13708 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_149
timestamp 1694700623
transform 1 0 14812 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_161
timestamp 1694700623
transform 1 0 15916 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_167
timestamp 1694700623
transform 1 0 16468 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_169
timestamp 1694700623
transform 1 0 16652 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_181
timestamp 1694700623
transform 1 0 17756 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_189
timestamp 1694700623
transform 1 0 18492 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_3
timestamp 1694700623
transform 1 0 1380 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_15
timestamp 1694700623
transform 1 0 2484 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_27
timestamp 1694700623
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_29
timestamp 1694700623
transform 1 0 3772 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_41
timestamp 1694700623
transform 1 0 4876 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_53
timestamp 1694700623
transform 1 0 5980 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_65
timestamp 1694700623
transform 1 0 7084 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_77
timestamp 1694700623
transform 1 0 8188 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_83
timestamp 1694700623
transform 1 0 8740 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_85
timestamp 1694700623
transform 1 0 8924 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_97
timestamp 1694700623
transform 1 0 10028 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_28_120
timestamp 1694700623
transform 1 0 12144 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_128
timestamp 1694700623
transform 1 0 12880 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_138
timestamp 1694700623
transform 1 0 13800 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_28_141
timestamp 1694700623
transform 1 0 14076 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_153
timestamp 1694700623
transform 1 0 15180 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_165
timestamp 1694700623
transform 1 0 16284 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_177
timestamp 1694700623
transform 1 0 17388 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_189
timestamp 1694700623
transform 1 0 18492 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_3
timestamp 1694700623
transform 1 0 1380 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_15
timestamp 1694700623
transform 1 0 2484 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_27
timestamp 1694700623
transform 1 0 3588 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_39
timestamp 1694700623
transform 1 0 4692 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_51
timestamp 1694700623
transform 1 0 5796 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_55
timestamp 1694700623
transform 1 0 6164 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_57
timestamp 1694700623
transform 1 0 6348 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_69
timestamp 1694700623
transform 1 0 7452 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_81
timestamp 1694700623
transform 1 0 8556 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_93
timestamp 1694700623
transform 1 0 9660 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_105
timestamp 1694700623
transform 1 0 10764 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_111
timestamp 1694700623
transform 1 0 11316 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_113
timestamp 1694700623
transform 1 0 11500 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_125
timestamp 1694700623
transform 1 0 12604 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_29_137
timestamp 1694700623
transform 1 0 13708 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_29_156
timestamp 1694700623
transform 1 0 15456 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_169
timestamp 1694700623
transform 1 0 16652 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_29_181
timestamp 1694700623
transform 1 0 17756 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_29_188
timestamp 1694700623
transform 1 0 18400 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_30_3
timestamp 1694700623
transform 1 0 1380 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_15
timestamp 1694700623
transform 1 0 2484 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_27
timestamp 1694700623
transform 1 0 3588 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_29
timestamp 1694700623
transform 1 0 3772 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_41
timestamp 1694700623
transform 1 0 4876 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_53
timestamp 1694700623
transform 1 0 5980 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_65
timestamp 1694700623
transform 1 0 7084 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_77
timestamp 1694700623
transform 1 0 8188 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_83
timestamp 1694700623
transform 1 0 8740 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_85
timestamp 1694700623
transform 1 0 8924 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_97
timestamp 1694700623
transform 1 0 10028 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_109
timestamp 1694700623
transform 1 0 11132 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_121
timestamp 1694700623
transform 1 0 12236 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_133
timestamp 1694700623
transform 1 0 13340 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_139
timestamp 1694700623
transform 1 0 13892 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_141
timestamp 1694700623
transform 1 0 14076 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_153
timestamp 1694700623
transform 1 0 15180 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_165
timestamp 1694700623
transform 1 0 16284 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_177
timestamp 1694700623
transform 1 0 17388 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_189
timestamp 1694700623
transform 1 0 18492 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_3
timestamp 1694700623
transform 1 0 1380 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_15
timestamp 1694700623
transform 1 0 2484 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_27
timestamp 1694700623
transform 1 0 3588 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_39
timestamp 1694700623
transform 1 0 4692 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_51
timestamp 1694700623
transform 1 0 5796 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_55
timestamp 1694700623
transform 1 0 6164 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_57
timestamp 1694700623
transform 1 0 6348 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_69
timestamp 1694700623
transform 1 0 7452 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_81
timestamp 1694700623
transform 1 0 8556 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_93
timestamp 1694700623
transform 1 0 9660 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_105
timestamp 1694700623
transform 1 0 10764 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_111
timestamp 1694700623
transform 1 0 11316 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_113
timestamp 1694700623
transform 1 0 11500 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_117
timestamp 1694700623
transform 1 0 11868 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_121
timestamp 1694700623
transform 1 0 12236 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_133
timestamp 1694700623
transform 1 0 13340 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_145
timestamp 1694700623
transform 1 0 14444 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_157
timestamp 1694700623
transform 1 0 15548 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_31_165
timestamp 1694700623
transform 1 0 16284 0 -1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_31_169
timestamp 1694700623
transform 1 0 16652 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_181
timestamp 1694700623
transform 1 0 17756 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_31_189
timestamp 1694700623
transform 1 0 18492 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_3
timestamp 1694700623
transform 1 0 1380 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_15
timestamp 1694700623
transform 1 0 2484 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_27
timestamp 1694700623
transform 1 0 3588 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_29
timestamp 1694700623
transform 1 0 3772 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_41
timestamp 1694700623
transform 1 0 4876 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_53
timestamp 1694700623
transform 1 0 5980 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_65
timestamp 1694700623
transform 1 0 7084 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_77
timestamp 1694700623
transform 1 0 8188 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_83
timestamp 1694700623
transform 1 0 8740 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_85
timestamp 1694700623
transform 1 0 8924 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_97
timestamp 1694700623
transform 1 0 10028 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_109
timestamp 1694700623
transform 1 0 11132 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_121
timestamp 1694700623
transform 1 0 12236 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_133
timestamp 1694700623
transform 1 0 13340 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_139
timestamp 1694700623
transform 1 0 13892 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_141
timestamp 1694700623
transform 1 0 14076 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_153
timestamp 1694700623
transform 1 0 15180 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_165
timestamp 1694700623
transform 1 0 16284 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_177
timestamp 1694700623
transform 1 0 17388 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_183
timestamp 1694700623
transform 1 0 17940 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_188
timestamp 1694700623
transform 1 0 18400 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_3
timestamp 1694700623
transform 1 0 1380 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_14
timestamp 1694700623
transform 1 0 2392 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_33_18
timestamp 1694700623
transform 1 0 2760 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_30
timestamp 1694700623
transform 1 0 3864 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_42
timestamp 1694700623
transform 1 0 4968 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_33_54
timestamp 1694700623
transform 1 0 6072 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_33_57
timestamp 1694700623
transform 1 0 6348 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_69
timestamp 1694700623
transform 1 0 7452 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_81
timestamp 1694700623
transform 1 0 8556 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_93
timestamp 1694700623
transform 1 0 9660 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_105
timestamp 1694700623
transform 1 0 10764 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_111
timestamp 1694700623
transform 1 0 11316 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_113
timestamp 1694700623
transform 1 0 11500 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_33_131
timestamp 1694700623
transform 1 0 13156 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_33_143
timestamp 1694700623
transform 1 0 14260 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_33_154
timestamp 1694700623
transform 1 0 15272 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_33_166
timestamp 1694700623
transform 1 0 16376 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_33_169
timestamp 1694700623
transform 1 0 16652 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_33_181
timestamp 1694700623
transform 1 0 17756 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_33_189
timestamp 1694700623
transform 1 0 18492 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_3
timestamp 1694700623
transform 1 0 1380 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_15
timestamp 1694700623
transform 1 0 2484 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_27
timestamp 1694700623
transform 1 0 3588 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_29
timestamp 1694700623
transform 1 0 3772 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_41
timestamp 1694700623
transform 1 0 4876 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_34_53
timestamp 1694700623
transform 1 0 5980 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_57
timestamp 1694700623
transform 1 0 6348 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_61
timestamp 1694700623
transform 1 0 6716 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_80
timestamp 1694700623
transform 1 0 8464 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_85
timestamp 1694700623
transform 1 0 8924 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_34_96
timestamp 1694700623
transform 1 0 9936 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_108
timestamp 1694700623
transform 1 0 11040 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_120
timestamp 1694700623
transform 1 0 12144 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_132
timestamp 1694700623
transform 1 0 13248 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_34_141
timestamp 1694700623
transform 1 0 14076 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_145
timestamp 1694700623
transform 1 0 14444 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_155
timestamp 1694700623
transform 1 0 15364 0 1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_34_176
timestamp 1694700623
transform 1 0 17296 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_34_188
timestamp 1694700623
transform 1 0 18400 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_35_3
timestamp 1694700623
transform 1 0 1380 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_15
timestamp 1694700623
transform 1 0 2484 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_27
timestamp 1694700623
transform 1 0 3588 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_39
timestamp 1694700623
transform 1 0 4692 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_51
timestamp 1694700623
transform 1 0 5796 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_55
timestamp 1694700623
transform 1 0 6164 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_57
timestamp 1694700623
transform 1 0 6348 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_69
timestamp 1694700623
transform 1 0 7452 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_81
timestamp 1694700623
transform 1 0 8556 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_93
timestamp 1694700623
transform 1 0 9660 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_35_105
timestamp 1694700623
transform 1 0 10764 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_35_110
timestamp 1694700623
transform 1 0 11224 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_113
timestamp 1694700623
transform 1 0 11500 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_119
timestamp 1694700623
transform 1 0 12052 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_123
timestamp 1694700623
transform 1 0 12420 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_35_127
timestamp 1694700623
transform 1 0 12788 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_139
timestamp 1694700623
transform 1 0 13892 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_151
timestamp 1694700623
transform 1 0 14996 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_163
timestamp 1694700623
transform 1 0 16100 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_167
timestamp 1694700623
transform 1 0 16468 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_169
timestamp 1694700623
transform 1 0 16652 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_181
timestamp 1694700623
transform 1 0 17756 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_35_189
timestamp 1694700623
transform 1 0 18492 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_36_3
timestamp 1694700623
transform 1 0 1380 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_36_11
timestamp 1694700623
transform 1 0 2116 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_22
timestamp 1694700623
transform 1 0 3128 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_26
timestamp 1694700623
transform 1 0 3496 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_36_29
timestamp 1694700623
transform 1 0 3772 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_36_34
timestamp 1694700623
transform 1 0 4232 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_38
timestamp 1694700623
transform 1 0 4600 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_42
timestamp 1694700623
transform 1 0 4968 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_60
timestamp 1694700623
transform 1 0 6624 0 1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_36_67
timestamp 1694700623
transform 1 0 7268 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_36_79
timestamp 1694700623
transform 1 0 8372 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_83
timestamp 1694700623
transform 1 0 8740 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_85
timestamp 1694700623
transform 1 0 8924 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_97
timestamp 1694700623
transform 1 0 10028 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_109
timestamp 1694700623
transform 1 0 11132 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_121
timestamp 1694700623
transform 1 0 12236 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_133
timestamp 1694700623
transform 1 0 13340 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_139
timestamp 1694700623
transform 1 0 13892 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_36_141
timestamp 1694700623
transform 1 0 14076 0 1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_36_147
timestamp 1694700623
transform 1 0 14628 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_159
timestamp 1694700623
transform 1 0 15732 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_171
timestamp 1694700623
transform 1 0 16836 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_183
timestamp 1694700623
transform 1 0 17940 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_36_188
timestamp 1694700623
transform 1 0 18400 0 1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_37_3
timestamp 1694700623
transform 1 0 1380 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_15
timestamp 1694700623
transform 1 0 2484 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_27
timestamp 1694700623
transform 1 0 3588 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_39
timestamp 1694700623
transform 1 0 4692 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_51
timestamp 1694700623
transform 1 0 5796 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_55
timestamp 1694700623
transform 1 0 6164 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_57
timestamp 1694700623
transform 1 0 6348 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_69
timestamp 1694700623
transform 1 0 7452 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_81
timestamp 1694700623
transform 1 0 8556 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_93
timestamp 1694700623
transform 1 0 9660 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_105
timestamp 1694700623
transform 1 0 10764 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_111
timestamp 1694700623
transform 1 0 11316 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_113
timestamp 1694700623
transform 1 0 11500 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_125
timestamp 1694700623
transform 1 0 12604 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_137
timestamp 1694700623
transform 1 0 13708 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_149
timestamp 1694700623
transform 1 0 14812 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_161
timestamp 1694700623
transform 1 0 15916 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_167
timestamp 1694700623
transform 1 0 16468 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_169
timestamp 1694700623
transform 1 0 16652 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_173
timestamp 1694700623
transform 1 0 17020 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_37_183
timestamp 1694700623
transform 1 0 17940 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_189
timestamp 1694700623
transform 1 0 18492 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_3
timestamp 1694700623
transform 1 0 1380 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_15
timestamp 1694700623
transform 1 0 2484 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_38_27
timestamp 1694700623
transform 1 0 3588 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_29
timestamp 1694700623
transform 1 0 3772 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_41
timestamp 1694700623
transform 1 0 4876 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_53
timestamp 1694700623
transform 1 0 5980 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_65
timestamp 1694700623
transform 1 0 7084 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_77
timestamp 1694700623
transform 1 0 8188 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_83
timestamp 1694700623
transform 1 0 8740 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_85
timestamp 1694700623
transform 1 0 8924 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_97
timestamp 1694700623
transform 1 0 10028 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_109
timestamp 1694700623
transform 1 0 11132 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_121
timestamp 1694700623
transform 1 0 12236 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_133
timestamp 1694700623
transform 1 0 13340 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_139
timestamp 1694700623
transform 1 0 13892 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_141
timestamp 1694700623
transform 1 0 14076 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_153
timestamp 1694700623
transform 1 0 15180 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_165
timestamp 1694700623
transform 1 0 16284 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_177
timestamp 1694700623
transform 1 0 17388 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_38_189
timestamp 1694700623
transform 1 0 18492 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_3
timestamp 1694700623
transform 1 0 1380 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_15
timestamp 1694700623
transform 1 0 2484 0 -1 23936
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_39_26
timestamp 1694700623
transform 1 0 3496 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_38
timestamp 1694700623
transform 1 0 4600 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_50
timestamp 1694700623
transform 1 0 5704 0 -1 23936
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_39_57
timestamp 1694700623
transform 1 0 6348 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_69
timestamp 1694700623
transform 1 0 7452 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_73
timestamp 1694700623
transform 1 0 7820 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_91
timestamp 1694700623
transform 1 0 9476 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_103
timestamp 1694700623
transform 1 0 10580 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_39_111
timestamp 1694700623
transform 1 0 11316 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_113
timestamp 1694700623
transform 1 0 11500 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_125
timestamp 1694700623
transform 1 0 12604 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_137
timestamp 1694700623
transform 1 0 13708 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_149
timestamp 1694700623
transform 1 0 14812 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_161
timestamp 1694700623
transform 1 0 15916 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_167
timestamp 1694700623
transform 1 0 16468 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_39_169
timestamp 1694700623
transform 1 0 16652 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_39_180
timestamp 1694700623
transform 1 0 17664 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_39_188
timestamp 1694700623
transform 1 0 18400 0 -1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_40_3
timestamp 1694700623
transform 1 0 1380 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_15
timestamp 1694700623
transform 1 0 2484 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_27
timestamp 1694700623
transform 1 0 3588 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_29
timestamp 1694700623
transform 1 0 3772 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_41
timestamp 1694700623
transform 1 0 4876 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_53
timestamp 1694700623
transform 1 0 5980 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_65
timestamp 1694700623
transform 1 0 7084 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_77
timestamp 1694700623
transform 1 0 8188 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_83
timestamp 1694700623
transform 1 0 8740 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_85
timestamp 1694700623
transform 1 0 8924 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_97
timestamp 1694700623
transform 1 0 10028 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_109
timestamp 1694700623
transform 1 0 11132 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_121
timestamp 1694700623
transform 1 0 12236 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_133
timestamp 1694700623
transform 1 0 13340 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_139
timestamp 1694700623
transform 1 0 13892 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_141
timestamp 1694700623
transform 1 0 14076 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_153
timestamp 1694700623
transform 1 0 15180 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_165
timestamp 1694700623
transform 1 0 16284 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_177
timestamp 1694700623
transform 1 0 17388 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_183
timestamp 1694700623
transform 1 0 17940 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_40_188
timestamp 1694700623
transform 1 0 18400 0 1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_41_3
timestamp 1694700623
transform 1 0 1380 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_15
timestamp 1694700623
transform 1 0 2484 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_27
timestamp 1694700623
transform 1 0 3588 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_39
timestamp 1694700623
transform 1 0 4692 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_51
timestamp 1694700623
transform 1 0 5796 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_55
timestamp 1694700623
transform 1 0 6164 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_57
timestamp 1694700623
transform 1 0 6348 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_69
timestamp 1694700623
transform 1 0 7452 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_81
timestamp 1694700623
transform 1 0 8556 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_85
timestamp 1694700623
transform 1 0 8924 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_89
timestamp 1694700623
transform 1 0 9292 0 -1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_41_97
timestamp 1694700623
transform 1 0 10028 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_41_109
timestamp 1694700623
transform 1 0 11132 0 -1 25024
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_41_113
timestamp 1694700623
transform 1 0 11500 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_125
timestamp 1694700623
transform 1 0 12604 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_137
timestamp 1694700623
transform 1 0 13708 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_149
timestamp 1694700623
transform 1 0 14812 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_161
timestamp 1694700623
transform 1 0 15916 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_167
timestamp 1694700623
transform 1 0 16468 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_41_169
timestamp 1694700623
transform 1 0 16652 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_41_177
timestamp 1694700623
transform 1 0 17388 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_188
timestamp 1694700623
transform 1 0 18400 0 -1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_42_3
timestamp 1694700623
transform 1 0 1380 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_15
timestamp 1694700623
transform 1 0 2484 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_42_27
timestamp 1694700623
transform 1 0 3588 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_42_29
timestamp 1694700623
transform 1 0 3772 0 1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_42_48
timestamp 1694700623
transform 1 0 5520 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_70
timestamp 1694700623
transform 1 0 7544 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_42_82
timestamp 1694700623
transform 1 0 8648 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_42_85
timestamp 1694700623
transform 1 0 8924 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_42_93
timestamp 1694700623
transform 1 0 9660 0 1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_42_104
timestamp 1694700623
transform 1 0 10672 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_116
timestamp 1694700623
transform 1 0 11776 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_42_131
timestamp 1694700623
transform 1 0 13156 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_42_139
timestamp 1694700623
transform 1 0 13892 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_141
timestamp 1694700623
transform 1 0 14076 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_153
timestamp 1694700623
transform 1 0 15180 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_165
timestamp 1694700623
transform 1 0 16284 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_177
timestamp 1694700623
transform 1 0 17388 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_42_189
timestamp 1694700623
transform 1 0 18492 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_3
timestamp 1694700623
transform 1 0 1380 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_15
timestamp 1694700623
transform 1 0 2484 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_27
timestamp 1694700623
transform 1 0 3588 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_39
timestamp 1694700623
transform 1 0 4692 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_51
timestamp 1694700623
transform 1 0 5796 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_55
timestamp 1694700623
transform 1 0 6164 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_57
timestamp 1694700623
transform 1 0 6348 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_69
timestamp 1694700623
transform 1 0 7452 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_81
timestamp 1694700623
transform 1 0 8556 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_93
timestamp 1694700623
transform 1 0 9660 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_97
timestamp 1694700623
transform 1 0 10028 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_107
timestamp 1694700623
transform 1 0 10948 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_111
timestamp 1694700623
transform 1 0 11316 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_113
timestamp 1694700623
transform 1 0 11500 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_125
timestamp 1694700623
transform 1 0 12604 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_137
timestamp 1694700623
transform 1 0 13708 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_149
timestamp 1694700623
transform 1 0 14812 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_161
timestamp 1694700623
transform 1 0 15916 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_167
timestamp 1694700623
transform 1 0 16468 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_169
timestamp 1694700623
transform 1 0 16652 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_43_181
timestamp 1694700623
transform 1 0 17756 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_43_188
timestamp 1694700623
transform 1 0 18400 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_44_3
timestamp 1694700623
transform 1 0 1380 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_9
timestamp 1694700623
transform 1 0 1932 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_44_26
timestamp 1694700623
transform 1 0 3496 0 1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_44_29
timestamp 1694700623
transform 1 0 3772 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_41
timestamp 1694700623
transform 1 0 4876 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_47
timestamp 1694700623
transform 1 0 5428 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_64
timestamp 1694700623
transform 1 0 6992 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_76
timestamp 1694700623
transform 1 0 8096 0 1 26112
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_44_85
timestamp 1694700623
transform 1 0 8924 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_97
timestamp 1694700623
transform 1 0 10028 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_109
timestamp 1694700623
transform 1 0 11132 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_121
timestamp 1694700623
transform 1 0 12236 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_133
timestamp 1694700623
transform 1 0 13340 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_139
timestamp 1694700623
transform 1 0 13892 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_141
timestamp 1694700623
transform 1 0 14076 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_153
timestamp 1694700623
transform 1 0 15180 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_165
timestamp 1694700623
transform 1 0 16284 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_177
timestamp 1694700623
transform 1 0 17388 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_44_189
timestamp 1694700623
transform 1 0 18492 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_3
timestamp 1694700623
transform 1 0 1380 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_15
timestamp 1694700623
transform 1 0 2484 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_27
timestamp 1694700623
transform 1 0 3588 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_39
timestamp 1694700623
transform 1 0 4692 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_51
timestamp 1694700623
transform 1 0 5796 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_55
timestamp 1694700623
transform 1 0 6164 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_57
timestamp 1694700623
transform 1 0 6348 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_69
timestamp 1694700623
transform 1 0 7452 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_81
timestamp 1694700623
transform 1 0 8556 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_93
timestamp 1694700623
transform 1 0 9660 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_105
timestamp 1694700623
transform 1 0 10764 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_111
timestamp 1694700623
transform 1 0 11316 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_113
timestamp 1694700623
transform 1 0 11500 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_125
timestamp 1694700623
transform 1 0 12604 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_131
timestamp 1694700623
transform 1 0 13156 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_149
timestamp 1694700623
transform 1 0 14812 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_161
timestamp 1694700623
transform 1 0 15916 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_167
timestamp 1694700623
transform 1 0 16468 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_169
timestamp 1694700623
transform 1 0 16652 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_45_181
timestamp 1694700623
transform 1 0 17756 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_45_189
timestamp 1694700623
transform 1 0 18492 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_3
timestamp 1694700623
transform 1 0 1380 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_15
timestamp 1694700623
transform 1 0 2484 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_46_27
timestamp 1694700623
transform 1 0 3588 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_46_29
timestamp 1694700623
transform 1 0 3772 0 1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_46_35
timestamp 1694700623
transform 1 0 4324 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_47
timestamp 1694700623
transform 1 0 5428 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_59
timestamp 1694700623
transform 1 0 6532 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_71
timestamp 1694700623
transform 1 0 7636 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_46_83
timestamp 1694700623
transform 1 0 8740 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_85
timestamp 1694700623
transform 1 0 8924 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_97
timestamp 1694700623
transform 1 0 10028 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_109
timestamp 1694700623
transform 1 0 11132 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_121
timestamp 1694700623
transform 1 0 12236 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_133
timestamp 1694700623
transform 1 0 13340 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_139
timestamp 1694700623
transform 1 0 13892 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_141
timestamp 1694700623
transform 1 0 14076 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_153
timestamp 1694700623
transform 1 0 15180 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_165
timestamp 1694700623
transform 1 0 16284 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_177
timestamp 1694700623
transform 1 0 17388 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_46_187
timestamp 1694700623
transform 1 0 18308 0 1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_47_3
timestamp 1694700623
transform 1 0 1380 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_15
timestamp 1694700623
transform 1 0 2484 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_27
timestamp 1694700623
transform 1 0 3588 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_31
timestamp 1694700623
transform 1 0 3956 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_47_48
timestamp 1694700623
transform 1 0 5520 0 -1 28288
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_47_57
timestamp 1694700623
transform 1 0 6348 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_69
timestamp 1694700623
transform 1 0 7452 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_81
timestamp 1694700623
transform 1 0 8556 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_93
timestamp 1694700623
transform 1 0 9660 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_105
timestamp 1694700623
transform 1 0 10764 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_111
timestamp 1694700623
transform 1 0 11316 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_113
timestamp 1694700623
transform 1 0 11500 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_125
timestamp 1694700623
transform 1 0 12604 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_137
timestamp 1694700623
transform 1 0 13708 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_149
timestamp 1694700623
transform 1 0 14812 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_161
timestamp 1694700623
transform 1 0 15916 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_167
timestamp 1694700623
transform 1 0 16468 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_169
timestamp 1694700623
transform 1 0 16652 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_47_181
timestamp 1694700623
transform 1 0 17756 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_47_188
timestamp 1694700623
transform 1 0 18400 0 -1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_48_3
timestamp 1694700623
transform 1 0 1380 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_15
timestamp 1694700623
transform 1 0 2484 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_48_27
timestamp 1694700623
transform 1 0 3588 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_29
timestamp 1694700623
transform 1 0 3772 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_48_41
timestamp 1694700623
transform 1 0 4876 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_45
timestamp 1694700623
transform 1 0 5244 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_56
timestamp 1694700623
transform 1 0 6256 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_68
timestamp 1694700623
transform 1 0 7360 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_48_80
timestamp 1694700623
transform 1 0 8464 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_48_85
timestamp 1694700623
transform 1 0 8924 0 1 28288
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_48_97
timestamp 1694700623
transform 1 0 10028 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_109
timestamp 1694700623
transform 1 0 11132 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_121
timestamp 1694700623
transform 1 0 12236 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_133
timestamp 1694700623
transform 1 0 13340 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_139
timestamp 1694700623
transform 1 0 13892 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_141
timestamp 1694700623
transform 1 0 14076 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_153
timestamp 1694700623
transform 1 0 15180 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_165
timestamp 1694700623
transform 1 0 16284 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_177
timestamp 1694700623
transform 1 0 17388 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_48_189
timestamp 1694700623
transform 1 0 18492 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_3
timestamp 1694700623
transform 1 0 1380 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_15
timestamp 1694700623
transform 1 0 2484 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_27
timestamp 1694700623
transform 1 0 3588 0 -1 29376
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_49_39
timestamp 1694700623
transform 1 0 4692 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_51
timestamp 1694700623
transform 1 0 5796 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_55
timestamp 1694700623
transform 1 0 6164 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_57
timestamp 1694700623
transform 1 0 6348 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_69
timestamp 1694700623
transform 1 0 7452 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_81
timestamp 1694700623
transform 1 0 8556 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_49_89
timestamp 1694700623
transform 1 0 9292 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_49_101
timestamp 1694700623
transform 1 0 10396 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_49_109
timestamp 1694700623
transform 1 0 11132 0 -1 29376
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_49_113
timestamp 1694700623
transform 1 0 11500 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_125
timestamp 1694700623
transform 1 0 12604 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_137
timestamp 1694700623
transform 1 0 13708 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_149
timestamp 1694700623
transform 1 0 14812 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_161
timestamp 1694700623
transform 1 0 15916 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_167
timestamp 1694700623
transform 1 0 16468 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_169
timestamp 1694700623
transform 1 0 16652 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_181
timestamp 1694700623
transform 1 0 17756 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_49_189
timestamp 1694700623
transform 1 0 18492 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_3
timestamp 1694700623
transform 1 0 1380 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_15
timestamp 1694700623
transform 1 0 2484 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_50_27
timestamp 1694700623
transform 1 0 3588 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_29
timestamp 1694700623
transform 1 0 3772 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_41
timestamp 1694700623
transform 1 0 4876 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_53
timestamp 1694700623
transform 1 0 5980 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_65
timestamp 1694700623
transform 1 0 7084 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_77
timestamp 1694700623
transform 1 0 8188 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_83
timestamp 1694700623
transform 1 0 8740 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_85
timestamp 1694700623
transform 1 0 8924 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_97
timestamp 1694700623
transform 1 0 10028 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_109
timestamp 1694700623
transform 1 0 11132 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_121
timestamp 1694700623
transform 1 0 12236 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_133
timestamp 1694700623
transform 1 0 13340 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_139
timestamp 1694700623
transform 1 0 13892 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_141
timestamp 1694700623
transform 1 0 14076 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_50_153
timestamp 1694700623
transform 1 0 15180 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_157
timestamp 1694700623
transform 1 0 15548 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_167
timestamp 1694700623
transform 1 0 16468 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_50_179
timestamp 1694700623
transform 1 0 17572 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_183
timestamp 1694700623
transform 1 0 17940 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_50_188
timestamp 1694700623
transform 1 0 18400 0 1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_51_3
timestamp 1694700623
transform 1 0 1380 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_15
timestamp 1694700623
transform 1 0 2484 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_21
timestamp 1694700623
transform 1 0 3036 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_31
timestamp 1694700623
transform 1 0 3956 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_43
timestamp 1694700623
transform 1 0 5060 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_51_55
timestamp 1694700623
transform 1 0 6164 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_51_57
timestamp 1694700623
transform 1 0 6348 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_51_68
timestamp 1694700623
transform 1 0 7360 0 -1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_51_89
timestamp 1694700623
transform 1 0 9292 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_51_101
timestamp 1694700623
transform 1 0 10396 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_51_109
timestamp 1694700623
transform 1 0 11132 0 -1 30464
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_51_113
timestamp 1694700623
transform 1 0 11500 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_125
timestamp 1694700623
transform 1 0 12604 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_51_137
timestamp 1694700623
transform 1 0 13708 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_51_145
timestamp 1694700623
transform 1 0 14444 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_51_162
timestamp 1694700623
transform 1 0 16008 0 -1 30464
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_51_169
timestamp 1694700623
transform 1 0 16652 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_51_181
timestamp 1694700623
transform 1 0 17756 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_51_189
timestamp 1694700623
transform 1 0 18492 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_3
timestamp 1694700623
transform 1 0 1380 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_15
timestamp 1694700623
transform 1 0 2484 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_52_27
timestamp 1694700623
transform 1 0 3588 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_29
timestamp 1694700623
transform 1 0 3772 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_52_41
timestamp 1694700623
transform 1 0 4876 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_52_49
timestamp 1694700623
transform 1 0 5612 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_59
timestamp 1694700623
transform 1 0 6532 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_71
timestamp 1694700623
transform 1 0 7636 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_52_83
timestamp 1694700623
transform 1 0 8740 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_85
timestamp 1694700623
transform 1 0 8924 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_97
timestamp 1694700623
transform 1 0 10028 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_109
timestamp 1694700623
transform 1 0 11132 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_121
timestamp 1694700623
transform 1 0 12236 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_133
timestamp 1694700623
transform 1 0 13340 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_139
timestamp 1694700623
transform 1 0 13892 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_141
timestamp 1694700623
transform 1 0 14076 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_153
timestamp 1694700623
transform 1 0 15180 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_165
timestamp 1694700623
transform 1 0 16284 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_177
timestamp 1694700623
transform 1 0 17388 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_52_189
timestamp 1694700623
transform 1 0 18492 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_53_3
timestamp 1694700623
transform 1 0 1380 0 -1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_53_8
timestamp 1694700623
transform 1 0 1840 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_20
timestamp 1694700623
transform 1 0 2944 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_32
timestamp 1694700623
transform 1 0 4048 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_44
timestamp 1694700623
transform 1 0 5152 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_57
timestamp 1694700623
transform 1 0 6348 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_69
timestamp 1694700623
transform 1 0 7452 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_81
timestamp 1694700623
transform 1 0 8556 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_93
timestamp 1694700623
transform 1 0 9660 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_105
timestamp 1694700623
transform 1 0 10764 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_111
timestamp 1694700623
transform 1 0 11316 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_113
timestamp 1694700623
transform 1 0 11500 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_125
timestamp 1694700623
transform 1 0 12604 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_137
timestamp 1694700623
transform 1 0 13708 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_149
timestamp 1694700623
transform 1 0 14812 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_161
timestamp 1694700623
transform 1 0 15916 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_167
timestamp 1694700623
transform 1 0 16468 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_53_169
timestamp 1694700623
transform 1 0 16652 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_53_188
timestamp 1694700623
transform 1 0 18400 0 -1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_54_3
timestamp 1694700623
transform 1 0 1380 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_15
timestamp 1694700623
transform 1 0 2484 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_54_27
timestamp 1694700623
transform 1 0 3588 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_29
timestamp 1694700623
transform 1 0 3772 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_41
timestamp 1694700623
transform 1 0 4876 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_53
timestamp 1694700623
transform 1 0 5980 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_65
timestamp 1694700623
transform 1 0 7084 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_77
timestamp 1694700623
transform 1 0 8188 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_83
timestamp 1694700623
transform 1 0 8740 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_85
timestamp 1694700623
transform 1 0 8924 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_97
timestamp 1694700623
transform 1 0 10028 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_109
timestamp 1694700623
transform 1 0 11132 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_121
timestamp 1694700623
transform 1 0 12236 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_133
timestamp 1694700623
transform 1 0 13340 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_139
timestamp 1694700623
transform 1 0 13892 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_141
timestamp 1694700623
transform 1 0 14076 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_153
timestamp 1694700623
transform 1 0 15180 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_165
timestamp 1694700623
transform 1 0 16284 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_177
timestamp 1694700623
transform 1 0 17388 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_183
timestamp 1694700623
transform 1 0 17940 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_54_188
timestamp 1694700623
transform 1 0 18400 0 1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_55_3
timestamp 1694700623
transform 1 0 1380 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_15
timestamp 1694700623
transform 1 0 2484 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_27
timestamp 1694700623
transform 1 0 3588 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_39
timestamp 1694700623
transform 1 0 4692 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_51
timestamp 1694700623
transform 1 0 5796 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_55
timestamp 1694700623
transform 1 0 6164 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_57
timestamp 1694700623
transform 1 0 6348 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_61
timestamp 1694700623
transform 1 0 6716 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_71
timestamp 1694700623
transform 1 0 7636 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_83
timestamp 1694700623
transform 1 0 8740 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_95
timestamp 1694700623
transform 1 0 9844 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_107
timestamp 1694700623
transform 1 0 10948 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_111
timestamp 1694700623
transform 1 0 11316 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_113
timestamp 1694700623
transform 1 0 11500 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_117
timestamp 1694700623
transform 1 0 11868 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_134
timestamp 1694700623
transform 1 0 13432 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_146
timestamp 1694700623
transform 1 0 14536 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_55_158
timestamp 1694700623
transform 1 0 15640 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_55_166
timestamp 1694700623
transform 1 0 16376 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_169
timestamp 1694700623
transform 1 0 16652 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_55_187
timestamp 1694700623
transform 1 0 18308 0 -1 32640
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_56_3
timestamp 1694700623
transform 1 0 1380 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_15
timestamp 1694700623
transform 1 0 2484 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_56_27
timestamp 1694700623
transform 1 0 3588 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_29
timestamp 1694700623
transform 1 0 3772 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_41
timestamp 1694700623
transform 1 0 4876 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_53
timestamp 1694700623
transform 1 0 5980 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_65
timestamp 1694700623
transform 1 0 7084 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_77
timestamp 1694700623
transform 1 0 8188 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_83
timestamp 1694700623
transform 1 0 8740 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_85
timestamp 1694700623
transform 1 0 8924 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_97
timestamp 1694700623
transform 1 0 10028 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_109
timestamp 1694700623
transform 1 0 11132 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_121
timestamp 1694700623
transform 1 0 12236 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_133
timestamp 1694700623
transform 1 0 13340 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_139
timestamp 1694700623
transform 1 0 13892 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_141
timestamp 1694700623
transform 1 0 14076 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_56_153
timestamp 1694700623
transform 1 0 15180 0 1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_56_173
timestamp 1694700623
transform 1 0 17020 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_56_185
timestamp 1694700623
transform 1 0 18124 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_189
timestamp 1694700623
transform 1 0 18492 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_3
timestamp 1694700623
transform 1 0 1380 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_15
timestamp 1694700623
transform 1 0 2484 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_27
timestamp 1694700623
transform 1 0 3588 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_39
timestamp 1694700623
transform 1 0 4692 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_51
timestamp 1694700623
transform 1 0 5796 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_55
timestamp 1694700623
transform 1 0 6164 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_57
timestamp 1694700623
transform 1 0 6348 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_69
timestamp 1694700623
transform 1 0 7452 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_81
timestamp 1694700623
transform 1 0 8556 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_93
timestamp 1694700623
transform 1 0 9660 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_105
timestamp 1694700623
transform 1 0 10764 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_111
timestamp 1694700623
transform 1 0 11316 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_113
timestamp 1694700623
transform 1 0 11500 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_125
timestamp 1694700623
transform 1 0 12604 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_137
timestamp 1694700623
transform 1 0 13708 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_57_149
timestamp 1694700623
transform 1 0 14812 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_57_160
timestamp 1694700623
transform 1 0 15824 0 -1 33728
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_57_169
timestamp 1694700623
transform 1 0 16652 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_57_181
timestamp 1694700623
transform 1 0 17756 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_57_188
timestamp 1694700623
transform 1 0 18400 0 -1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_58_3
timestamp 1694700623
transform 1 0 1380 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_15
timestamp 1694700623
transform 1 0 2484 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_58_27
timestamp 1694700623
transform 1 0 3588 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_29
timestamp 1694700623
transform 1 0 3772 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_41
timestamp 1694700623
transform 1 0 4876 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_53
timestamp 1694700623
transform 1 0 5980 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_65
timestamp 1694700623
transform 1 0 7084 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_77
timestamp 1694700623
transform 1 0 8188 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_83
timestamp 1694700623
transform 1 0 8740 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_85
timestamp 1694700623
transform 1 0 8924 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_97
timestamp 1694700623
transform 1 0 10028 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_109
timestamp 1694700623
transform 1 0 11132 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_121
timestamp 1694700623
transform 1 0 12236 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_133
timestamp 1694700623
transform 1 0 13340 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_139
timestamp 1694700623
transform 1 0 13892 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_141
timestamp 1694700623
transform 1 0 14076 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_58_153
timestamp 1694700623
transform 1 0 15180 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_58_161
timestamp 1694700623
transform 1 0 15916 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_58_166
timestamp 1694700623
transform 1 0 16376 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_58_179
timestamp 1694700623
transform 1 0 17572 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_58_187
timestamp 1694700623
transform 1 0 18308 0 1 33728
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_59_3
timestamp 1694700623
transform 1 0 1380 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_59_15
timestamp 1694700623
transform 1 0 2484 0 -1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_59_26
timestamp 1694700623
transform 1 0 3496 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_38
timestamp 1694700623
transform 1 0 4600 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_50
timestamp 1694700623
transform 1 0 5704 0 -1 34816
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_59_57
timestamp 1694700623
transform 1 0 6348 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_69
timestamp 1694700623
transform 1 0 7452 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_59_81
timestamp 1694700623
transform 1 0 8556 0 -1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_59_99
timestamp 1694700623
transform 1 0 10212 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_59_111
timestamp 1694700623
transform 1 0 11316 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_59_113
timestamp 1694700623
transform 1 0 11500 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_59_130
timestamp 1694700623
transform 1 0 13064 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_59_149
timestamp 1694700623
transform 1 0 14812 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_59_153
timestamp 1694700623
transform 1 0 15180 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_59_164
timestamp 1694700623
transform 1 0 16192 0 -1 34816
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_59_169
timestamp 1694700623
transform 1 0 16652 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_59_181
timestamp 1694700623
transform 1 0 17756 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_59_189
timestamp 1694700623
transform 1 0 18492 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_3
timestamp 1694700623
transform 1 0 1380 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_15
timestamp 1694700623
transform 1 0 2484 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_60_27
timestamp 1694700623
transform 1 0 3588 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_29
timestamp 1694700623
transform 1 0 3772 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_41
timestamp 1694700623
transform 1 0 4876 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_53
timestamp 1694700623
transform 1 0 5980 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_60_65
timestamp 1694700623
transform 1 0 7084 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_60_82
timestamp 1694700623
transform 1 0 8648 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_60_85
timestamp 1694700623
transform 1 0 8924 0 1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_60_103
timestamp 1694700623
transform 1 0 10580 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_115
timestamp 1694700623
transform 1 0 11684 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_60_127
timestamp 1694700623
transform 1 0 12788 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_60_138
timestamp 1694700623
transform 1 0 13800 0 1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_60_141
timestamp 1694700623
transform 1 0 14076 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_153
timestamp 1694700623
transform 1 0 15180 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_165
timestamp 1694700623
transform 1 0 16284 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_177
timestamp 1694700623
transform 1 0 17388 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_60_189
timestamp 1694700623
transform 1 0 18492 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_3
timestamp 1694700623
transform 1 0 1380 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_15
timestamp 1694700623
transform 1 0 2484 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_27
timestamp 1694700623
transform 1 0 3588 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_39
timestamp 1694700623
transform 1 0 4692 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_61_51
timestamp 1694700623
transform 1 0 5796 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_55
timestamp 1694700623
transform 1 0 6164 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_57
timestamp 1694700623
transform 1 0 6348 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_69
timestamp 1694700623
transform 1 0 7452 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_81
timestamp 1694700623
transform 1 0 8556 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_93
timestamp 1694700623
transform 1 0 9660 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_105
timestamp 1694700623
transform 1 0 10764 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_111
timestamp 1694700623
transform 1 0 11316 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_61_113
timestamp 1694700623
transform 1 0 11500 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_61_125
timestamp 1694700623
transform 1 0 12604 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_129
timestamp 1694700623
transform 1 0 12972 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_147
timestamp 1694700623
transform 1 0 14628 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_61_159
timestamp 1694700623
transform 1 0 15732 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_61_167
timestamp 1694700623
transform 1 0 16468 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_169
timestamp 1694700623
transform 1 0 16652 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_61_181
timestamp 1694700623
transform 1 0 17756 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_61_188
timestamp 1694700623
transform 1 0 18400 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_62_3
timestamp 1694700623
transform 1 0 1380 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_62_11
timestamp 1694700623
transform 1 0 2116 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_62_21
timestamp 1694700623
transform 1 0 3036 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_27
timestamp 1694700623
transform 1 0 3588 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_29
timestamp 1694700623
transform 1 0 3772 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_41
timestamp 1694700623
transform 1 0 4876 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_53
timestamp 1694700623
transform 1 0 5980 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_65
timestamp 1694700623
transform 1 0 7084 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_77
timestamp 1694700623
transform 1 0 8188 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_83
timestamp 1694700623
transform 1 0 8740 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_85
timestamp 1694700623
transform 1 0 8924 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_97
timestamp 1694700623
transform 1 0 10028 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_62_109
timestamp 1694700623
transform 1 0 11132 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_62_114
timestamp 1694700623
transform 1 0 11592 0 1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_62_125
timestamp 1694700623
transform 1 0 12604 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_62_137
timestamp 1694700623
transform 1 0 13708 0 1 35904
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_62_141
timestamp 1694700623
transform 1 0 14076 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_153
timestamp 1694700623
transform 1 0 15180 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_165
timestamp 1694700623
transform 1 0 16284 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_177
timestamp 1694700623
transform 1 0 17388 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_62_189
timestamp 1694700623
transform 1 0 18492 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_3
timestamp 1694700623
transform 1 0 1380 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_15
timestamp 1694700623
transform 1 0 2484 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_27
timestamp 1694700623
transform 1 0 3588 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_39
timestamp 1694700623
transform 1 0 4692 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_51
timestamp 1694700623
transform 1 0 5796 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_55
timestamp 1694700623
transform 1 0 6164 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_57
timestamp 1694700623
transform 1 0 6348 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_69
timestamp 1694700623
transform 1 0 7452 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_75
timestamp 1694700623
transform 1 0 8004 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_85
timestamp 1694700623
transform 1 0 8924 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_97
timestamp 1694700623
transform 1 0 10028 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_63_109
timestamp 1694700623
transform 1 0 11132 0 -1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_63_113
timestamp 1694700623
transform 1 0 11500 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_125
timestamp 1694700623
transform 1 0 12604 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_137
timestamp 1694700623
transform 1 0 13708 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_149
timestamp 1694700623
transform 1 0 14812 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_161
timestamp 1694700623
transform 1 0 15916 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_167
timestamp 1694700623
transform 1 0 16468 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_169
timestamp 1694700623
transform 1 0 16652 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_63_181
timestamp 1694700623
transform 1 0 17756 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_63_189
timestamp 1694700623
transform 1 0 18492 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_64_3
timestamp 1694700623
transform 1 0 1380 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_64_25
timestamp 1694700623
transform 1 0 3404 0 1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_64_29
timestamp 1694700623
transform 1 0 3772 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_41
timestamp 1694700623
transform 1 0 4876 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_53
timestamp 1694700623
transform 1 0 5980 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_65
timestamp 1694700623
transform 1 0 7084 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_77
timestamp 1694700623
transform 1 0 8188 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_83
timestamp 1694700623
transform 1 0 8740 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_85
timestamp 1694700623
transform 1 0 8924 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_97
timestamp 1694700623
transform 1 0 10028 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_109
timestamp 1694700623
transform 1 0 11132 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_64_121
timestamp 1694700623
transform 1 0 12236 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_64_134
timestamp 1694700623
transform 1 0 13432 0 1 36992
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_64_141
timestamp 1694700623
transform 1 0 14076 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_153
timestamp 1694700623
transform 1 0 15180 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_165
timestamp 1694700623
transform 1 0 16284 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_177
timestamp 1694700623
transform 1 0 17388 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_183
timestamp 1694700623
transform 1 0 17940 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_64_188
timestamp 1694700623
transform 1 0 18400 0 1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_65_3
timestamp 1694700623
transform 1 0 1380 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_15
timestamp 1694700623
transform 1 0 2484 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_27
timestamp 1694700623
transform 1 0 3588 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_39
timestamp 1694700623
transform 1 0 4692 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_65_51
timestamp 1694700623
transform 1 0 5796 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_65_55
timestamp 1694700623
transform 1 0 6164 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_57
timestamp 1694700623
transform 1 0 6348 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_69
timestamp 1694700623
transform 1 0 7452 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_81
timestamp 1694700623
transform 1 0 8556 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_93
timestamp 1694700623
transform 1 0 9660 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_105
timestamp 1694700623
transform 1 0 10764 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_111
timestamp 1694700623
transform 1 0 11316 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_113
timestamp 1694700623
transform 1 0 11500 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_125
timestamp 1694700623
transform 1 0 12604 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_137
timestamp 1694700623
transform 1 0 13708 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_65_149
timestamp 1694700623
transform 1 0 14812 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_65_166
timestamp 1694700623
transform 1 0 16376 0 -1 38080
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_65_169
timestamp 1694700623
transform 1 0 16652 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_65_181
timestamp 1694700623
transform 1 0 17756 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_65_189
timestamp 1694700623
transform 1 0 18492 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_3
timestamp 1694700623
transform 1 0 1380 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_15
timestamp 1694700623
transform 1 0 2484 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_66_27
timestamp 1694700623
transform 1 0 3588 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_29
timestamp 1694700623
transform 1 0 3772 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_41
timestamp 1694700623
transform 1 0 4876 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_53
timestamp 1694700623
transform 1 0 5980 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_65
timestamp 1694700623
transform 1 0 7084 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_77
timestamp 1694700623
transform 1 0 8188 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_83
timestamp 1694700623
transform 1 0 8740 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_85
timestamp 1694700623
transform 1 0 8924 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_97
timestamp 1694700623
transform 1 0 10028 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_109
timestamp 1694700623
transform 1 0 11132 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_121
timestamp 1694700623
transform 1 0 12236 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_133
timestamp 1694700623
transform 1 0 13340 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_139
timestamp 1694700623
transform 1 0 13892 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_141
timestamp 1694700623
transform 1 0 14076 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_66_153
timestamp 1694700623
transform 1 0 15180 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_157
timestamp 1694700623
transform 1 0 15548 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_169
timestamp 1694700623
transform 1 0 16652 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_66_181
timestamp 1694700623
transform 1 0 17756 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_66_189
timestamp 1694700623
transform 1 0 18492 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_3
timestamp 1694700623
transform 1 0 1380 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_15
timestamp 1694700623
transform 1 0 2484 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_67_27
timestamp 1694700623
transform 1 0 3588 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_44
timestamp 1694700623
transform 1 0 5152 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_57
timestamp 1694700623
transform 1 0 6348 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_69
timestamp 1694700623
transform 1 0 7452 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_81
timestamp 1694700623
transform 1 0 8556 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_93
timestamp 1694700623
transform 1 0 9660 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_105
timestamp 1694700623
transform 1 0 10764 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_111
timestamp 1694700623
transform 1 0 11316 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_113
timestamp 1694700623
transform 1 0 11500 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_125
timestamp 1694700623
transform 1 0 12604 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_137
timestamp 1694700623
transform 1 0 13708 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_149
timestamp 1694700623
transform 1 0 14812 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_161
timestamp 1694700623
transform 1 0 15916 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_167
timestamp 1694700623
transform 1 0 16468 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_67_169
timestamp 1694700623
transform 1 0 16652 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_67_174
timestamp 1694700623
transform 1 0 17112 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_67_178
timestamp 1694700623
transform 1 0 17480 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_67_188
timestamp 1694700623
transform 1 0 18400 0 -1 39168
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_68_3
timestamp 1694700623
transform 1 0 1380 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_15
timestamp 1694700623
transform 1 0 2484 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_68_27
timestamp 1694700623
transform 1 0 3588 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_29
timestamp 1694700623
transform 1 0 3772 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_41
timestamp 1694700623
transform 1 0 4876 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_53
timestamp 1694700623
transform 1 0 5980 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_65
timestamp 1694700623
transform 1 0 7084 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_77
timestamp 1694700623
transform 1 0 8188 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_83
timestamp 1694700623
transform 1 0 8740 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_85
timestamp 1694700623
transform 1 0 8924 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_97
timestamp 1694700623
transform 1 0 10028 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_109
timestamp 1694700623
transform 1 0 11132 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_68_121
timestamp 1694700623
transform 1 0 12236 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_68_131
timestamp 1694700623
transform 1 0 13156 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_68_139
timestamp 1694700623
transform 1 0 13892 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_141
timestamp 1694700623
transform 1 0 14076 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_153
timestamp 1694700623
transform 1 0 15180 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_165
timestamp 1694700623
transform 1 0 16284 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_177
timestamp 1694700623
transform 1 0 17388 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_183
timestamp 1694700623
transform 1 0 17940 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_68_188
timestamp 1694700623
transform 1 0 18400 0 1 39168
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_69_3
timestamp 1694700623
transform 1 0 1380 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_15
timestamp 1694700623
transform 1 0 2484 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_27
timestamp 1694700623
transform 1 0 3588 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_39
timestamp 1694700623
transform 1 0 4692 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_69_51
timestamp 1694700623
transform 1 0 5796 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_69_55
timestamp 1694700623
transform 1 0 6164 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_57
timestamp 1694700623
transform 1 0 6348 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_69_69
timestamp 1694700623
transform 1 0 7452 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_69_82
timestamp 1694700623
transform 1 0 8648 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_69_90
timestamp 1694700623
transform 1 0 9384 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_69_108
timestamp 1694700623
transform 1 0 11040 0 -1 40256
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_69_113
timestamp 1694700623
transform 1 0 11500 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_125
timestamp 1694700623
transform 1 0 12604 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_137
timestamp 1694700623
transform 1 0 13708 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_149
timestamp 1694700623
transform 1 0 14812 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_155
timestamp 1694700623
transform 1 0 15364 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_69_166
timestamp 1694700623
transform 1 0 16376 0 -1 40256
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_69_169
timestamp 1694700623
transform 1 0 16652 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_69_181
timestamp 1694700623
transform 1 0 17756 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_69_189
timestamp 1694700623
transform 1 0 18492 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_3
timestamp 1694700623
transform 1 0 1380 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_15
timestamp 1694700623
transform 1 0 2484 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_70_27
timestamp 1694700623
transform 1 0 3588 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_29
timestamp 1694700623
transform 1 0 3772 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_41
timestamp 1694700623
transform 1 0 4876 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_53
timestamp 1694700623
transform 1 0 5980 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_65
timestamp 1694700623
transform 1 0 7084 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_77
timestamp 1694700623
transform 1 0 8188 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_83
timestamp 1694700623
transform 1 0 8740 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_85
timestamp 1694700623
transform 1 0 8924 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_97
timestamp 1694700623
transform 1 0 10028 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_109
timestamp 1694700623
transform 1 0 11132 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_121
timestamp 1694700623
transform 1 0 12236 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_133
timestamp 1694700623
transform 1 0 13340 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_139
timestamp 1694700623
transform 1 0 13892 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_141
timestamp 1694700623
transform 1 0 14076 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_153
timestamp 1694700623
transform 1 0 15180 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_165
timestamp 1694700623
transform 1 0 16284 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_177
timestamp 1694700623
transform 1 0 17388 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_70_189
timestamp 1694700623
transform 1 0 18492 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_3
timestamp 1694700623
transform 1 0 1380 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_15
timestamp 1694700623
transform 1 0 2484 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_27
timestamp 1694700623
transform 1 0 3588 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_39
timestamp 1694700623
transform 1 0 4692 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_71_51
timestamp 1694700623
transform 1 0 5796 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_71_55
timestamp 1694700623
transform 1 0 6164 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_57
timestamp 1694700623
transform 1 0 6348 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_69
timestamp 1694700623
transform 1 0 7452 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_81
timestamp 1694700623
transform 1 0 8556 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_93
timestamp 1694700623
transform 1 0 9660 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_105
timestamp 1694700623
transform 1 0 10764 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_111
timestamp 1694700623
transform 1 0 11316 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_113
timestamp 1694700623
transform 1 0 11500 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_125
timestamp 1694700623
transform 1 0 12604 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_137
timestamp 1694700623
transform 1 0 13708 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_149
timestamp 1694700623
transform 1 0 14812 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_161
timestamp 1694700623
transform 1 0 15916 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_167
timestamp 1694700623
transform 1 0 16468 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_169
timestamp 1694700623
transform 1 0 16652 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_71_181
timestamp 1694700623
transform 1 0 17756 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_71_188
timestamp 1694700623
transform 1 0 18400 0 -1 41344
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_72_3
timestamp 1694700623
transform 1 0 1380 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_15
timestamp 1694700623
transform 1 0 2484 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_72_27
timestamp 1694700623
transform 1 0 3588 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_29
timestamp 1694700623
transform 1 0 3772 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_72_41
timestamp 1694700623
transform 1 0 4876 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_72_49
timestamp 1694700623
transform 1 0 5612 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_59
timestamp 1694700623
transform 1 0 6532 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_71
timestamp 1694700623
transform 1 0 7636 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_72_83
timestamp 1694700623
transform 1 0 8740 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_85
timestamp 1694700623
transform 1 0 8924 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_97
timestamp 1694700623
transform 1 0 10028 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_109
timestamp 1694700623
transform 1 0 11132 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_121
timestamp 1694700623
transform 1 0 12236 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_133
timestamp 1694700623
transform 1 0 13340 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_139
timestamp 1694700623
transform 1 0 13892 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_141
timestamp 1694700623
transform 1 0 14076 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_153
timestamp 1694700623
transform 1 0 15180 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_165
timestamp 1694700623
transform 1 0 16284 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_177
timestamp 1694700623
transform 1 0 17388 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_72_189
timestamp 1694700623
transform 1 0 18492 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_73_3
timestamp 1694700623
transform 1 0 1380 0 -1 42432
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_73_28
timestamp 1694700623
transform 1 0 3680 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_40
timestamp 1694700623
transform 1 0 4784 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_73_52
timestamp 1694700623
transform 1 0 5888 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_73_57
timestamp 1694700623
transform 1 0 6348 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_73_65
timestamp 1694700623
transform 1 0 7084 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_73_83
timestamp 1694700623
transform 1 0 8740 0 -1 42432
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_73_96
timestamp 1694700623
transform 1 0 9936 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_73_108
timestamp 1694700623
transform 1 0 11040 0 -1 42432
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_73_113
timestamp 1694700623
transform 1 0 11500 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_125
timestamp 1694700623
transform 1 0 12604 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_137
timestamp 1694700623
transform 1 0 13708 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_149
timestamp 1694700623
transform 1 0 14812 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_161
timestamp 1694700623
transform 1 0 15916 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_167
timestamp 1694700623
transform 1 0 16468 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_169
timestamp 1694700623
transform 1 0 16652 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_73_181
timestamp 1694700623
transform 1 0 17756 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_73_189
timestamp 1694700623
transform 1 0 18492 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_74_3
timestamp 1694700623
transform 1 0 1380 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_74_14
timestamp 1694700623
transform 1 0 2392 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_74_21
timestamp 1694700623
transform 1 0 3036 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_27
timestamp 1694700623
transform 1 0 3588 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_29
timestamp 1694700623
transform 1 0 3772 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_41
timestamp 1694700623
transform 1 0 4876 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_53
timestamp 1694700623
transform 1 0 5980 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_65
timestamp 1694700623
transform 1 0 7084 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_77
timestamp 1694700623
transform 1 0 8188 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_83
timestamp 1694700623
transform 1 0 8740 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_74_85
timestamp 1694700623
transform 1 0 8924 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_74_93
timestamp 1694700623
transform 1 0 9660 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_74_97
timestamp 1694700623
transform 1 0 10028 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_74_101
timestamp 1694700623
transform 1 0 10396 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_111
timestamp 1694700623
transform 1 0 11316 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_123
timestamp 1694700623
transform 1 0 12420 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_74_138
timestamp 1694700623
transform 1 0 13800 0 1 42432
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_74_141
timestamp 1694700623
transform 1 0 14076 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_153
timestamp 1694700623
transform 1 0 15180 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_165
timestamp 1694700623
transform 1 0 16284 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_177
timestamp 1694700623
transform 1 0 17388 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_74_189
timestamp 1694700623
transform 1 0 18492 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_3
timestamp 1694700623
transform 1 0 1380 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_15
timestamp 1694700623
transform 1 0 2484 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_27
timestamp 1694700623
transform 1 0 3588 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_39
timestamp 1694700623
transform 1 0 4692 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_75_51
timestamp 1694700623
transform 1 0 5796 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_75_55
timestamp 1694700623
transform 1 0 6164 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_57
timestamp 1694700623
transform 1 0 6348 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_69
timestamp 1694700623
transform 1 0 7452 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_81
timestamp 1694700623
transform 1 0 8556 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_93
timestamp 1694700623
transform 1 0 9660 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_105
timestamp 1694700623
transform 1 0 10764 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_111
timestamp 1694700623
transform 1 0 11316 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_113
timestamp 1694700623
transform 1 0 11500 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_125
timestamp 1694700623
transform 1 0 12604 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_137
timestamp 1694700623
transform 1 0 13708 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_149
timestamp 1694700623
transform 1 0 14812 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_161
timestamp 1694700623
transform 1 0 15916 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_167
timestamp 1694700623
transform 1 0 16468 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_169
timestamp 1694700623
transform 1 0 16652 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_75_181
timestamp 1694700623
transform 1 0 17756 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_75_188
timestamp 1694700623
transform 1 0 18400 0 -1 43520
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_76_3
timestamp 1694700623
transform 1 0 1380 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_15
timestamp 1694700623
transform 1 0 2484 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_76_27
timestamp 1694700623
transform 1 0 3588 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_29
timestamp 1694700623
transform 1 0 3772 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_41
timestamp 1694700623
transform 1 0 4876 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_76_53
timestamp 1694700623
transform 1 0 5980 0 1 43520
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_76_70
timestamp 1694700623
transform 1 0 7544 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_76_82
timestamp 1694700623
transform 1 0 8648 0 1 43520
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_76_85
timestamp 1694700623
transform 1 0 8924 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_97
timestamp 1694700623
transform 1 0 10028 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_109
timestamp 1694700623
transform 1 0 11132 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_121
timestamp 1694700623
transform 1 0 12236 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_133
timestamp 1694700623
transform 1 0 13340 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_139
timestamp 1694700623
transform 1 0 13892 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_141
timestamp 1694700623
transform 1 0 14076 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_153
timestamp 1694700623
transform 1 0 15180 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_165
timestamp 1694700623
transform 1 0 16284 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_177
timestamp 1694700623
transform 1 0 17388 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_76_189
timestamp 1694700623
transform 1 0 18492 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_77_3
timestamp 1694700623
transform 1 0 1380 0 -1 44608
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_77_14
timestamp 1694700623
transform 1 0 2392 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_77_26
timestamp 1694700623
transform 1 0 3496 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_77_34
timestamp 1694700623
transform 1 0 4232 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_77_52
timestamp 1694700623
transform 1 0 5888 0 -1 44608
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_77_57
timestamp 1694700623
transform 1 0 6348 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_69
timestamp 1694700623
transform 1 0 7452 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_81
timestamp 1694700623
transform 1 0 8556 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_93
timestamp 1694700623
transform 1 0 9660 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_105
timestamp 1694700623
transform 1 0 10764 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_111
timestamp 1694700623
transform 1 0 11316 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_113
timestamp 1694700623
transform 1 0 11500 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_125
timestamp 1694700623
transform 1 0 12604 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_137
timestamp 1694700623
transform 1 0 13708 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_149
timestamp 1694700623
transform 1 0 14812 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_161
timestamp 1694700623
transform 1 0 15916 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_167
timestamp 1694700623
transform 1 0 16468 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_169
timestamp 1694700623
transform 1 0 16652 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_77_181
timestamp 1694700623
transform 1 0 17756 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_77_189
timestamp 1694700623
transform 1 0 18492 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_3
timestamp 1694700623
transform 1 0 1380 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_15
timestamp 1694700623
transform 1 0 2484 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_78_27
timestamp 1694700623
transform 1 0 3588 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_29
timestamp 1694700623
transform 1 0 3772 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_41
timestamp 1694700623
transform 1 0 4876 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_53
timestamp 1694700623
transform 1 0 5980 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_65
timestamp 1694700623
transform 1 0 7084 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_77
timestamp 1694700623
transform 1 0 8188 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_83
timestamp 1694700623
transform 1 0 8740 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_85
timestamp 1694700623
transform 1 0 8924 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_97
timestamp 1694700623
transform 1 0 10028 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_109
timestamp 1694700623
transform 1 0 11132 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_78_121
timestamp 1694700623
transform 1 0 12236 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_78_138
timestamp 1694700623
transform 1 0 13800 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_78_141
timestamp 1694700623
transform 1 0 14076 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_78_162
timestamp 1694700623
transform 1 0 16008 0 1 44608
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_78_169
timestamp 1694700623
transform 1 0 16652 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_78_181
timestamp 1694700623
transform 1 0 17756 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_78_188
timestamp 1694700623
transform 1 0 18400 0 1 44608
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_79_3
timestamp 1694700623
transform 1 0 1380 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_15
timestamp 1694700623
transform 1 0 2484 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_27
timestamp 1694700623
transform 1 0 3588 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_39
timestamp 1694700623
transform 1 0 4692 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_79_51
timestamp 1694700623
transform 1 0 5796 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_79_55
timestamp 1694700623
transform 1 0 6164 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_57
timestamp 1694700623
transform 1 0 6348 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_69
timestamp 1694700623
transform 1 0 7452 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_81
timestamp 1694700623
transform 1 0 8556 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_93
timestamp 1694700623
transform 1 0 9660 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_105
timestamp 1694700623
transform 1 0 10764 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_111
timestamp 1694700623
transform 1 0 11316 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_113
timestamp 1694700623
transform 1 0 11500 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_125
timestamp 1694700623
transform 1 0 12604 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_137
timestamp 1694700623
transform 1 0 13708 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_149
timestamp 1694700623
transform 1 0 14812 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_161
timestamp 1694700623
transform 1 0 15916 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_167
timestamp 1694700623
transform 1 0 16468 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_169
timestamp 1694700623
transform 1 0 16652 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_79_181
timestamp 1694700623
transform 1 0 17756 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_79_189
timestamp 1694700623
transform 1 0 18492 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_3
timestamp 1694700623
transform 1 0 1380 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_15
timestamp 1694700623
transform 1 0 2484 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_80_27
timestamp 1694700623
transform 1 0 3588 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_29
timestamp 1694700623
transform 1 0 3772 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_41
timestamp 1694700623
transform 1 0 4876 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_53
timestamp 1694700623
transform 1 0 5980 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_65
timestamp 1694700623
transform 1 0 7084 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_77
timestamp 1694700623
transform 1 0 8188 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_83
timestamp 1694700623
transform 1 0 8740 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_85
timestamp 1694700623
transform 1 0 8924 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_97
timestamp 1694700623
transform 1 0 10028 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_109
timestamp 1694700623
transform 1 0 11132 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_121
timestamp 1694700623
transform 1 0 12236 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_133
timestamp 1694700623
transform 1 0 13340 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_139
timestamp 1694700623
transform 1 0 13892 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_141
timestamp 1694700623
transform 1 0 14076 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_153
timestamp 1694700623
transform 1 0 15180 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_165
timestamp 1694700623
transform 1 0 16284 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_177
timestamp 1694700623
transform 1 0 17388 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_80_189
timestamp 1694700623
transform 1 0 18492 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_3
timestamp 1694700623
transform 1 0 1380 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_15
timestamp 1694700623
transform 1 0 2484 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_27
timestamp 1694700623
transform 1 0 3588 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_39
timestamp 1694700623
transform 1 0 4692 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_81_51
timestamp 1694700623
transform 1 0 5796 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_81_55
timestamp 1694700623
transform 1 0 6164 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_57
timestamp 1694700623
transform 1 0 6348 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_69
timestamp 1694700623
transform 1 0 7452 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_81
timestamp 1694700623
transform 1 0 8556 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_93
timestamp 1694700623
transform 1 0 9660 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_105
timestamp 1694700623
transform 1 0 10764 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_111
timestamp 1694700623
transform 1 0 11316 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_81_113
timestamp 1694700623
transform 1 0 11500 0 -1 46784
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_81_138
timestamp 1694700623
transform 1 0 13800 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_150
timestamp 1694700623
transform 1 0 14904 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_162
timestamp 1694700623
transform 1 0 16008 0 -1 46784
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_81_169
timestamp 1694700623
transform 1 0 16652 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_81_181
timestamp 1694700623
transform 1 0 17756 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_81_189
timestamp 1694700623
transform 1 0 18492 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_3
timestamp 1694700623
transform 1 0 1380 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_82_15
timestamp 1694700623
transform 1 0 2484 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_82_26
timestamp 1694700623
transform 1 0 3496 0 1 46784
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_82_29
timestamp 1694700623
transform 1 0 3772 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_41
timestamp 1694700623
transform 1 0 4876 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_53
timestamp 1694700623
transform 1 0 5980 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_82_65
timestamp 1694700623
transform 1 0 7084 0 1 46784
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_82_71
timestamp 1694700623
transform 1 0 7636 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_82_83
timestamp 1694700623
transform 1 0 8740 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_85
timestamp 1694700623
transform 1 0 8924 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_97
timestamp 1694700623
transform 1 0 10028 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_109
timestamp 1694700623
transform 1 0 11132 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_121
timestamp 1694700623
transform 1 0 12236 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_133
timestamp 1694700623
transform 1 0 13340 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_139
timestamp 1694700623
transform 1 0 13892 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_141
timestamp 1694700623
transform 1 0 14076 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_153
timestamp 1694700623
transform 1 0 15180 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_165
timestamp 1694700623
transform 1 0 16284 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_177
timestamp 1694700623
transform 1 0 17388 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_183
timestamp 1694700623
transform 1 0 17940 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_82_188
timestamp 1694700623
transform 1 0 18400 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_83_3
timestamp 1694700623
transform 1 0 1380 0 -1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_83_11
timestamp 1694700623
transform 1 0 2116 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_83_16
timestamp 1694700623
transform 1 0 2576 0 -1 47872
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_83_24
timestamp 1694700623
transform 1 0 3312 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_83_36
timestamp 1694700623
transform 1 0 4416 0 -1 47872
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_83_43
timestamp 1694700623
transform 1 0 5060 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_83_55
timestamp 1694700623
transform 1 0 6164 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_83_57
timestamp 1694700623
transform 1 0 6348 0 -1 47872
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_83_68
timestamp 1694700623
transform 1 0 7360 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_80
timestamp 1694700623
transform 1 0 8464 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_92
timestamp 1694700623
transform 1 0 9568 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_83_104
timestamp 1694700623
transform 1 0 10672 0 -1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_83_113
timestamp 1694700623
transform 1 0 11500 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_83_120
timestamp 1694700623
transform 1 0 12144 0 -1 47872
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_83_145
timestamp 1694700623
transform 1 0 14444 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_83_157
timestamp 1694700623
transform 1 0 15548 0 -1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_83_165
timestamp 1694700623
transform 1 0 16284 0 -1 47872
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_83_169
timestamp 1694700623
transform 1 0 16652 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_83_181
timestamp 1694700623
transform 1 0 17756 0 -1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_83_189
timestamp 1694700623
transform 1 0 18492 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_3
timestamp 1694700623
transform 1 0 1380 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_15
timestamp 1694700623
transform 1 0 2484 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_84_27
timestamp 1694700623
transform 1 0 3588 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_29
timestamp 1694700623
transform 1 0 3772 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_41
timestamp 1694700623
transform 1 0 4876 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_53
timestamp 1694700623
transform 1 0 5980 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_65
timestamp 1694700623
transform 1 0 7084 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_77
timestamp 1694700623
transform 1 0 8188 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_83
timestamp 1694700623
transform 1 0 8740 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_85
timestamp 1694700623
transform 1 0 8924 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_97
timestamp 1694700623
transform 1 0 10028 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_109
timestamp 1694700623
transform 1 0 11132 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_121
timestamp 1694700623
transform 1 0 12236 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_133
timestamp 1694700623
transform 1 0 13340 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_139
timestamp 1694700623
transform 1 0 13892 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_141
timestamp 1694700623
transform 1 0 14076 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_153
timestamp 1694700623
transform 1 0 15180 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_165
timestamp 1694700623
transform 1 0 16284 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_177
timestamp 1694700623
transform 1 0 17388 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_84_189
timestamp 1694700623
transform 1 0 18492 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_3
timestamp 1694700623
transform 1 0 1380 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_15
timestamp 1694700623
transform 1 0 2484 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_85_23
timestamp 1694700623
transform 1 0 3220 0 -1 48960
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_85_41
timestamp 1694700623
transform 1 0 4876 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_85_53
timestamp 1694700623
transform 1 0 5980 0 -1 48960
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_85_57
timestamp 1694700623
transform 1 0 6348 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_72
timestamp 1694700623
transform 1 0 7728 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_84
timestamp 1694700623
transform 1 0 8832 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_85_96
timestamp 1694700623
transform 1 0 9936 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_85_109
timestamp 1694700623
transform 1 0 11132 0 -1 48960
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_85_113
timestamp 1694700623
transform 1 0 11500 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_125
timestamp 1694700623
transform 1 0 12604 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_137
timestamp 1694700623
transform 1 0 13708 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_85_152
timestamp 1694700623
transform 1 0 15088 0 -1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_85_163
timestamp 1694700623
transform 1 0 16100 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_85_167
timestamp 1694700623
transform 1 0 16468 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_169
timestamp 1694700623
transform 1 0 16652 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_85_181
timestamp 1694700623
transform 1 0 17756 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_85_188
timestamp 1694700623
transform 1 0 18400 0 -1 48960
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_86_3
timestamp 1694700623
transform 1 0 1380 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_15
timestamp 1694700623
transform 1 0 2484 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_86_27
timestamp 1694700623
transform 1 0 3588 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_29
timestamp 1694700623
transform 1 0 3772 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_41
timestamp 1694700623
transform 1 0 4876 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_69
timestamp 1694700623
transform 1 0 7452 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_86_81
timestamp 1694700623
transform 1 0 8556 0 1 48960
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_86_85
timestamp 1694700623
transform 1 0 8924 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_97
timestamp 1694700623
transform 1 0 10028 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_109
timestamp 1694700623
transform 1 0 11132 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_121
timestamp 1694700623
transform 1 0 12236 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_133
timestamp 1694700623
transform 1 0 13340 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_139
timestamp 1694700623
transform 1 0 13892 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_141
timestamp 1694700623
transform 1 0 14076 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_153
timestamp 1694700623
transform 1 0 15180 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_165
timestamp 1694700623
transform 1 0 16284 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_177
timestamp 1694700623
transform 1 0 17388 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_86_189
timestamp 1694700623
transform 1 0 18492 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_3
timestamp 1694700623
transform 1 0 1380 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_15
timestamp 1694700623
transform 1 0 2484 0 -1 50048
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_87_38
timestamp 1694700623
transform 1 0 4600 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_50
timestamp 1694700623
transform 1 0 5704 0 -1 50048
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_87_57
timestamp 1694700623
transform 1 0 6348 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_69
timestamp 1694700623
transform 1 0 7452 0 -1 50048
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_87_92
timestamp 1694700623
transform 1 0 9568 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_87_104
timestamp 1694700623
transform 1 0 10672 0 -1 50048
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_87_113
timestamp 1694700623
transform 1 0 11500 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_125
timestamp 1694700623
transform 1 0 12604 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_137
timestamp 1694700623
transform 1 0 13708 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_149
timestamp 1694700623
transform 1 0 14812 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_161
timestamp 1694700623
transform 1 0 15916 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_167
timestamp 1694700623
transform 1 0 16468 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_169
timestamp 1694700623
transform 1 0 16652 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_87_181
timestamp 1694700623
transform 1 0 17756 0 -1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_87_189
timestamp 1694700623
transform 1 0 18492 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_3
timestamp 1694700623
transform 1 0 1380 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_88_15
timestamp 1694700623
transform 1 0 2484 0 1 50048
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_88_26
timestamp 1694700623
transform 1 0 3496 0 1 50048
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_88_29
timestamp 1694700623
transform 1 0 3772 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_41
timestamp 1694700623
transform 1 0 4876 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_53
timestamp 1694700623
transform 1 0 5980 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_65
timestamp 1694700623
transform 1 0 7084 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_77
timestamp 1694700623
transform 1 0 8188 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_83
timestamp 1694700623
transform 1 0 8740 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_85
timestamp 1694700623
transform 1 0 8924 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_97
timestamp 1694700623
transform 1 0 10028 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_109
timestamp 1694700623
transform 1 0 11132 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_121
timestamp 1694700623
transform 1 0 12236 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_133
timestamp 1694700623
transform 1 0 13340 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_139
timestamp 1694700623
transform 1 0 13892 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_88_141
timestamp 1694700623
transform 1 0 14076 0 1 50048
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_88_146
timestamp 1694700623
transform 1 0 14536 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_158
timestamp 1694700623
transform 1 0 15640 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_170
timestamp 1694700623
transform 1 0 16744 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_88_182
timestamp 1694700623
transform 1 0 17848 0 1 50048
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_89_3
timestamp 1694700623
transform 1 0 1380 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_15
timestamp 1694700623
transform 1 0 2484 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_27
timestamp 1694700623
transform 1 0 3588 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_39
timestamp 1694700623
transform 1 0 4692 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_89_51
timestamp 1694700623
transform 1 0 5796 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_89_55
timestamp 1694700623
transform 1 0 6164 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_57
timestamp 1694700623
transform 1 0 6348 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_89_69
timestamp 1694700623
transform 1 0 7452 0 -1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_89_77
timestamp 1694700623
transform 1 0 8188 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_89_80
timestamp 1694700623
transform 1 0 8464 0 -1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_89_84
timestamp 1694700623
transform 1 0 8832 0 -1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_89_102
timestamp 1694700623
transform 1 0 10488 0 -1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_89_106
timestamp 1694700623
transform 1 0 10856 0 -1 51136
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_89_113
timestamp 1694700623
transform 1 0 11500 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_125
timestamp 1694700623
transform 1 0 12604 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_137
timestamp 1694700623
transform 1 0 13708 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_149
timestamp 1694700623
transform 1 0 14812 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_161
timestamp 1694700623
transform 1 0 15916 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_167
timestamp 1694700623
transform 1 0 16468 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_169
timestamp 1694700623
transform 1 0 16652 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_89_181
timestamp 1694700623
transform 1 0 17756 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_89_188
timestamp 1694700623
transform 1 0 18400 0 -1 51136
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_90_3
timestamp 1694700623
transform 1 0 1380 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_15
timestamp 1694700623
transform 1 0 2484 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_90_27
timestamp 1694700623
transform 1 0 3588 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_90_29
timestamp 1694700623
transform 1 0 3772 0 1 51136
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_90_48
timestamp 1694700623
transform 1 0 5520 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_60
timestamp 1694700623
transform 1 0 6624 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_72
timestamp 1694700623
transform 1 0 7728 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_78
timestamp 1694700623
transform 1 0 8280 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_90_82
timestamp 1694700623
transform 1 0 8648 0 1 51136
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_90_85
timestamp 1694700623
transform 1 0 8924 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_90_97
timestamp 1694700623
transform 1 0 10028 0 1 51136
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_90_118
timestamp 1694700623
transform 1 0 11960 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_90_130
timestamp 1694700623
transform 1 0 13064 0 1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_90_138
timestamp 1694700623
transform 1 0 13800 0 1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_90_141
timestamp 1694700623
transform 1 0 14076 0 1 51136
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_90_153
timestamp 1694700623
transform 1 0 15180 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_165
timestamp 1694700623
transform 1 0 16284 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_177
timestamp 1694700623
transform 1 0 17388 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_90_189
timestamp 1694700623
transform 1 0 18492 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_3
timestamp 1694700623
transform 1 0 1380 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_15
timestamp 1694700623
transform 1 0 2484 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_27
timestamp 1694700623
transform 1 0 3588 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_39
timestamp 1694700623
transform 1 0 4692 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_91_51
timestamp 1694700623
transform 1 0 5796 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_91_55
timestamp 1694700623
transform 1 0 6164 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_57
timestamp 1694700623
transform 1 0 6348 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_69
timestamp 1694700623
transform 1 0 7452 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_81
timestamp 1694700623
transform 1 0 8556 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_93
timestamp 1694700623
transform 1 0 9660 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_105
timestamp 1694700623
transform 1 0 10764 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_111
timestamp 1694700623
transform 1 0 11316 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_113
timestamp 1694700623
transform 1 0 11500 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_125
timestamp 1694700623
transform 1 0 12604 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_137
timestamp 1694700623
transform 1 0 13708 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_149
timestamp 1694700623
transform 1 0 14812 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_161
timestamp 1694700623
transform 1 0 15916 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_167
timestamp 1694700623
transform 1 0 16468 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_169
timestamp 1694700623
transform 1 0 16652 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_91_181
timestamp 1694700623
transform 1 0 17756 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_91_187
timestamp 1694700623
transform 1 0 18308 0 -1 52224
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_92_3
timestamp 1694700623
transform 1 0 1380 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_15
timestamp 1694700623
transform 1 0 2484 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_92_27
timestamp 1694700623
transform 1 0 3588 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_29
timestamp 1694700623
transform 1 0 3772 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_41
timestamp 1694700623
transform 1 0 4876 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_53
timestamp 1694700623
transform 1 0 5980 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_65
timestamp 1694700623
transform 1 0 7084 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_77
timestamp 1694700623
transform 1 0 8188 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_83
timestamp 1694700623
transform 1 0 8740 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_85
timestamp 1694700623
transform 1 0 8924 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_97
timestamp 1694700623
transform 1 0 10028 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_109
timestamp 1694700623
transform 1 0 11132 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_121
timestamp 1694700623
transform 1 0 12236 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_133
timestamp 1694700623
transform 1 0 13340 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_139
timestamp 1694700623
transform 1 0 13892 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_92_141
timestamp 1694700623
transform 1 0 14076 0 1 52224
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_92_160
timestamp 1694700623
transform 1 0 15824 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_172
timestamp 1694700623
transform 1 0 16928 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_92_188
timestamp 1694700623
transform 1 0 18400 0 1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_93_3
timestamp 1694700623
transform 1 0 1380 0 -1 53312
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_93_14
timestamp 1694700623
transform 1 0 2392 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_26
timestamp 1694700623
transform 1 0 3496 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_38
timestamp 1694700623
transform 1 0 4600 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_50
timestamp 1694700623
transform 1 0 5704 0 -1 53312
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_93_57
timestamp 1694700623
transform 1 0 6348 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_93_69
timestamp 1694700623
transform 1 0 7452 0 -1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_93_77
timestamp 1694700623
transform 1 0 8188 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_93_84
timestamp 1694700623
transform 1 0 8832 0 -1 53312
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_93_99
timestamp 1694700623
transform 1 0 10212 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_93_111
timestamp 1694700623
transform 1 0 11316 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_93_113
timestamp 1694700623
transform 1 0 11500 0 -1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_93_121
timestamp 1694700623
transform 1 0 12236 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_139
timestamp 1694700623
transform 1 0 13892 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_151
timestamp 1694700623
transform 1 0 14996 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_93_163
timestamp 1694700623
transform 1 0 16100 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_93_167
timestamp 1694700623
transform 1 0 16468 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_169
timestamp 1694700623
transform 1 0 16652 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_93_181
timestamp 1694700623
transform 1 0 17756 0 -1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_93_189
timestamp 1694700623
transform 1 0 18492 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_3
timestamp 1694700623
transform 1 0 1380 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_15
timestamp 1694700623
transform 1 0 2484 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_94_27
timestamp 1694700623
transform 1 0 3588 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_29
timestamp 1694700623
transform 1 0 3772 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_41
timestamp 1694700623
transform 1 0 4876 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_53
timestamp 1694700623
transform 1 0 5980 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_65
timestamp 1694700623
transform 1 0 7084 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_77
timestamp 1694700623
transform 1 0 8188 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_83
timestamp 1694700623
transform 1 0 8740 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_85
timestamp 1694700623
transform 1 0 8924 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_97
timestamp 1694700623
transform 1 0 10028 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_109
timestamp 1694700623
transform 1 0 11132 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_121
timestamp 1694700623
transform 1 0 12236 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_133
timestamp 1694700623
transform 1 0 13340 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_139
timestamp 1694700623
transform 1 0 13892 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_141
timestamp 1694700623
transform 1 0 14076 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_153
timestamp 1694700623
transform 1 0 15180 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_165
timestamp 1694700623
transform 1 0 16284 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_177
timestamp 1694700623
transform 1 0 17388 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_94_189
timestamp 1694700623
transform 1 0 18492 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_3
timestamp 1694700623
transform 1 0 1380 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_15
timestamp 1694700623
transform 1 0 2484 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_27
timestamp 1694700623
transform 1 0 3588 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_39
timestamp 1694700623
transform 1 0 4692 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_95_51
timestamp 1694700623
transform 1 0 5796 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_95_55
timestamp 1694700623
transform 1 0 6164 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_57
timestamp 1694700623
transform 1 0 6348 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_69
timestamp 1694700623
transform 1 0 7452 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_81
timestamp 1694700623
transform 1 0 8556 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_95_93
timestamp 1694700623
transform 1 0 9660 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_95_97
timestamp 1694700623
transform 1 0 10028 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_95_108
timestamp 1694700623
transform 1 0 11040 0 -1 54400
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_95_113
timestamp 1694700623
transform 1 0 11500 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_95_125
timestamp 1694700623
transform 1 0 12604 0 -1 54400
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_95_130
timestamp 1694700623
transform 1 0 13064 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_142
timestamp 1694700623
transform 1 0 14168 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_154
timestamp 1694700623
transform 1 0 15272 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_95_166
timestamp 1694700623
transform 1 0 16376 0 -1 54400
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_95_169
timestamp 1694700623
transform 1 0 16652 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_95_181
timestamp 1694700623
transform 1 0 17756 0 -1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_95_189
timestamp 1694700623
transform 1 0 18492 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_3
timestamp 1694700623
transform 1 0 1380 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_15
timestamp 1694700623
transform 1 0 2484 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_96_27
timestamp 1694700623
transform 1 0 3588 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_29
timestamp 1694700623
transform 1 0 3772 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_41
timestamp 1694700623
transform 1 0 4876 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_53
timestamp 1694700623
transform 1 0 5980 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_65
timestamp 1694700623
transform 1 0 7084 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_77
timestamp 1694700623
transform 1 0 8188 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_83
timestamp 1694700623
transform 1 0 8740 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_85
timestamp 1694700623
transform 1 0 8924 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_97
timestamp 1694700623
transform 1 0 10028 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_109
timestamp 1694700623
transform 1 0 11132 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_121
timestamp 1694700623
transform 1 0 12236 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_133
timestamp 1694700623
transform 1 0 13340 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_139
timestamp 1694700623
transform 1 0 13892 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_141
timestamp 1694700623
transform 1 0 14076 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_153
timestamp 1694700623
transform 1 0 15180 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_165
timestamp 1694700623
transform 1 0 16284 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_177
timestamp 1694700623
transform 1 0 17388 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_183
timestamp 1694700623
transform 1 0 17940 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_96_188
timestamp 1694700623
transform 1 0 18400 0 1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_97_3
timestamp 1694700623
transform 1 0 1380 0 -1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_97_11
timestamp 1694700623
transform 1 0 2116 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_97_29
timestamp 1694700623
transform 1 0 3772 0 -1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_97_33
timestamp 1694700623
transform 1 0 4140 0 -1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_97_37
timestamp 1694700623
transform 1 0 4508 0 -1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_97_41
timestamp 1694700623
transform 1 0 4876 0 -1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_97_45
timestamp 1694700623
transform 1 0 5244 0 -1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_97_51
timestamp 1694700623
transform 1 0 5796 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_97_55
timestamp 1694700623
transform 1 0 6164 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_97_57
timestamp 1694700623
transform 1 0 6348 0 -1 55488
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_97_61
timestamp 1694700623
transform 1 0 6716 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_73
timestamp 1694700623
transform 1 0 7820 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_85
timestamp 1694700623
transform 1 0 8924 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_97
timestamp 1694700623
transform 1 0 10028 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_97_109
timestamp 1694700623
transform 1 0 11132 0 -1 55488
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_97_113
timestamp 1694700623
transform 1 0 11500 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_125
timestamp 1694700623
transform 1 0 12604 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_137
timestamp 1694700623
transform 1 0 13708 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_149
timestamp 1694700623
transform 1 0 14812 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_161
timestamp 1694700623
transform 1 0 15916 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_167
timestamp 1694700623
transform 1 0 16468 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_97_169
timestamp 1694700623
transform 1 0 16652 0 -1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_97_180
timestamp 1694700623
transform 1 0 17664 0 -1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_97_188
timestamp 1694700623
transform 1 0 18400 0 -1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_98_3
timestamp 1694700623
transform 1 0 1380 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_98_22
timestamp 1694700623
transform 1 0 3128 0 1 55488
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_98_29
timestamp 1694700623
transform 1 0 3772 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_41
timestamp 1694700623
transform 1 0 4876 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_53
timestamp 1694700623
transform 1 0 5980 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_65
timestamp 1694700623
transform 1 0 7084 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_77
timestamp 1694700623
transform 1 0 8188 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_83
timestamp 1694700623
transform 1 0 8740 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_85
timestamp 1694700623
transform 1 0 8924 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_97
timestamp 1694700623
transform 1 0 10028 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_98_109
timestamp 1694700623
transform 1 0 11132 0 1 55488
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_98_121
timestamp 1694700623
transform 1 0 12236 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_133
timestamp 1694700623
transform 1 0 13340 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_139
timestamp 1694700623
transform 1 0 13892 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_141
timestamp 1694700623
transform 1 0 14076 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_153
timestamp 1694700623
transform 1 0 15180 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_165
timestamp 1694700623
transform 1 0 16284 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_177
timestamp 1694700623
transform 1 0 17388 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_98_189
timestamp 1694700623
transform 1 0 18492 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_99_3
timestamp 1694700623
transform 1 0 1380 0 -1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_99_11
timestamp 1694700623
transform 1 0 2116 0 -1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_99_16
timestamp 1694700623
transform 1 0 2576 0 -1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_99_20
timestamp 1694700623
transform 1 0 2944 0 -1 56576
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_99_38
timestamp 1694700623
transform 1 0 4600 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_50
timestamp 1694700623
transform 1 0 5704 0 -1 56576
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_99_57
timestamp 1694700623
transform 1 0 6348 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_69
timestamp 1694700623
transform 1 0 7452 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_81
timestamp 1694700623
transform 1 0 8556 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_93
timestamp 1694700623
transform 1 0 9660 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_105
timestamp 1694700623
transform 1 0 10764 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_111
timestamp 1694700623
transform 1 0 11316 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_99_113
timestamp 1694700623
transform 1 0 11500 0 -1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_99_121
timestamp 1694700623
transform 1 0 12236 0 -1 56576
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_99_133
timestamp 1694700623
transform 1 0 13340 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_145
timestamp 1694700623
transform 1 0 14444 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_99_157
timestamp 1694700623
transform 1 0 15548 0 -1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_99_165
timestamp 1694700623
transform 1 0 16284 0 -1 56576
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_99_169
timestamp 1694700623
transform 1 0 16652 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_99_181
timestamp 1694700623
transform 1 0 17756 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_99_188
timestamp 1694700623
transform 1 0 18400 0 -1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_100_3
timestamp 1694700623
transform 1 0 1380 0 1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_100_14
timestamp 1694700623
transform 1 0 2392 0 1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_100_18
timestamp 1694700623
transform 1 0 2760 0 1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_100_26
timestamp 1694700623
transform 1 0 3496 0 1 56576
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_100_29
timestamp 1694700623
transform 1 0 3772 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_41
timestamp 1694700623
transform 1 0 4876 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_53
timestamp 1694700623
transform 1 0 5980 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_65
timestamp 1694700623
transform 1 0 7084 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_77
timestamp 1694700623
transform 1 0 8188 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_83
timestamp 1694700623
transform 1 0 8740 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_85
timestamp 1694700623
transform 1 0 8924 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_97
timestamp 1694700623
transform 1 0 10028 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_109
timestamp 1694700623
transform 1 0 11132 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_121
timestamp 1694700623
transform 1 0 12236 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_133
timestamp 1694700623
transform 1 0 13340 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_139
timestamp 1694700623
transform 1 0 13892 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_141
timestamp 1694700623
transform 1 0 14076 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_153
timestamp 1694700623
transform 1 0 15180 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_165
timestamp 1694700623
transform 1 0 16284 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_177
timestamp 1694700623
transform 1 0 17388 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_100_189
timestamp 1694700623
transform 1 0 18492 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_101_3
timestamp 1694700623
transform 1 0 1380 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_101_11
timestamp 1694700623
transform 1 0 2116 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_101_16
timestamp 1694700623
transform 1 0 2576 0 -1 57664
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_101_34
timestamp 1694700623
transform 1 0 4232 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_101_46
timestamp 1694700623
transform 1 0 5336 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_101_54
timestamp 1694700623
transform 1 0 6072 0 -1 57664
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_101_57
timestamp 1694700623
transform 1 0 6348 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_69
timestamp 1694700623
transform 1 0 7452 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_81
timestamp 1694700623
transform 1 0 8556 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_93
timestamp 1694700623
transform 1 0 9660 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_101_105
timestamp 1694700623
transform 1 0 10764 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_101_111
timestamp 1694700623
transform 1 0 11316 0 -1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_101_113
timestamp 1694700623
transform 1 0 11500 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_125
timestamp 1694700623
transform 1 0 12604 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_137
timestamp 1694700623
transform 1 0 13708 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_101_149
timestamp 1694700623
transform 1 0 14812 0 -1 57664
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_101_154
timestamp 1694700623
transform 1 0 15272 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_101_166
timestamp 1694700623
transform 1 0 16376 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_101_169
timestamp 1694700623
transform 1 0 16652 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_101_174
timestamp 1694700623
transform 1 0 17112 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_101_185
timestamp 1694700623
transform 1 0 18124 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_101_189
timestamp 1694700623
transform 1 0 18492 0 -1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_102_3
timestamp 1694700623
transform 1 0 1380 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_15
timestamp 1694700623
transform 1 0 2484 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_102_27
timestamp 1694700623
transform 1 0 3588 0 1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_102_29
timestamp 1694700623
transform 1 0 3772 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_41
timestamp 1694700623
transform 1 0 4876 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_53
timestamp 1694700623
transform 1 0 5980 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_65
timestamp 1694700623
transform 1 0 7084 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_102_77
timestamp 1694700623
transform 1 0 8188 0 1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_102_83
timestamp 1694700623
transform 1 0 8740 0 1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_102_85
timestamp 1694700623
transform 1 0 8924 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_97
timestamp 1694700623
transform 1 0 10028 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_109
timestamp 1694700623
transform 1 0 11132 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_121
timestamp 1694700623
transform 1 0 12236 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_102_133
timestamp 1694700623
transform 1 0 13340 0 1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_102_139
timestamp 1694700623
transform 1 0 13892 0 1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_102_141
timestamp 1694700623
transform 1 0 14076 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_153
timestamp 1694700623
transform 1 0 15180 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_165
timestamp 1694700623
transform 1 0 16284 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_177
timestamp 1694700623
transform 1 0 17388 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_102_189
timestamp 1694700623
transform 1 0 18492 0 1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_103_3
timestamp 1694700623
transform 1 0 1380 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_15
timestamp 1694700623
transform 1 0 2484 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_27
timestamp 1694700623
transform 1 0 3588 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_39
timestamp 1694700623
transform 1 0 4692 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_103_51
timestamp 1694700623
transform 1 0 5796 0 -1 58752
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_103_55
timestamp 1694700623
transform 1 0 6164 0 -1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_103_57
timestamp 1694700623
transform 1 0 6348 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_69
timestamp 1694700623
transform 1 0 7452 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_81
timestamp 1694700623
transform 1 0 8556 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_93
timestamp 1694700623
transform 1 0 9660 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_103_105
timestamp 1694700623
transform 1 0 10764 0 -1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_103_111
timestamp 1694700623
transform 1 0 11316 0 -1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_103_113
timestamp 1694700623
transform 1 0 11500 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_125
timestamp 1694700623
transform 1 0 12604 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_137
timestamp 1694700623
transform 1 0 13708 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_149
timestamp 1694700623
transform 1 0 14812 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_103_161
timestamp 1694700623
transform 1 0 15916 0 -1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_103_167
timestamp 1694700623
transform 1 0 16468 0 -1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_103_169
timestamp 1694700623
transform 1 0 16652 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_103_181
timestamp 1694700623
transform 1 0 17756 0 -1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_103_188
timestamp 1694700623
transform 1 0 18400 0 -1 58752
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_104_3
timestamp 1694700623
transform 1 0 1380 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_15
timestamp 1694700623
transform 1 0 2484 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_104_27
timestamp 1694700623
transform 1 0 3588 0 1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_104_29
timestamp 1694700623
transform 1 0 3772 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_41
timestamp 1694700623
transform 1 0 4876 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_53
timestamp 1694700623
transform 1 0 5980 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_104_65
timestamp 1694700623
transform 1 0 7084 0 1 58752
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_104_77
timestamp 1694700623
transform 1 0 8188 0 1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_104_83
timestamp 1694700623
transform 1 0 8740 0 1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_104_85
timestamp 1694700623
transform 1 0 8924 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_97
timestamp 1694700623
transform 1 0 10028 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_109
timestamp 1694700623
transform 1 0 11132 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_121
timestamp 1694700623
transform 1 0 12236 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_104_133
timestamp 1694700623
transform 1 0 13340 0 1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_104_138
timestamp 1694700623
transform 1 0 13800 0 1 58752
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_104_141
timestamp 1694700623
transform 1 0 14076 0 1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_104_146
timestamp 1694700623
transform 1 0 14536 0 1 58752
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_104_157
timestamp 1694700623
transform 1 0 15548 0 1 58752
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_104_161
timestamp 1694700623
transform 1 0 15916 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_173
timestamp 1694700623
transform 1 0 17020 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_104_185
timestamp 1694700623
transform 1 0 18124 0 1 58752
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_104_189
timestamp 1694700623
transform 1 0 18492 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_105_3
timestamp 1694700623
transform 1 0 1380 0 -1 59840
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_105_13
timestamp 1694700623
transform 1 0 2300 0 -1 59840
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_105_17
timestamp 1694700623
transform 1 0 2668 0 -1 59840
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_105_21
timestamp 1694700623
transform 1 0 3036 0 -1 59840
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_105_39
timestamp 1694700623
transform 1 0 4692 0 -1 59840
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_105_43
timestamp 1694700623
transform 1 0 5060 0 -1 59840
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_105_47
timestamp 1694700623
transform 1 0 5428 0 -1 59840
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_105_55
timestamp 1694700623
transform 1 0 6164 0 -1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_105_57
timestamp 1694700623
transform 1 0 6348 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_69
timestamp 1694700623
transform 1 0 7452 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_81
timestamp 1694700623
transform 1 0 8556 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_93
timestamp 1694700623
transform 1 0 9660 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_105_105
timestamp 1694700623
transform 1 0 10764 0 -1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_105_111
timestamp 1694700623
transform 1 0 11316 0 -1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_105_113
timestamp 1694700623
transform 1 0 11500 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_125
timestamp 1694700623
transform 1 0 12604 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_137
timestamp 1694700623
transform 1 0 13708 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_149
timestamp 1694700623
transform 1 0 14812 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_105_161
timestamp 1694700623
transform 1 0 15916 0 -1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_105_167
timestamp 1694700623
transform 1 0 16468 0 -1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_105_169
timestamp 1694700623
transform 1 0 16652 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_105_181
timestamp 1694700623
transform 1 0 17756 0 -1 59840
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_105_189
timestamp 1694700623
transform 1 0 18492 0 -1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_106_3
timestamp 1694700623
transform 1 0 1380 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_15
timestamp 1694700623
transform 1 0 2484 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_106_27
timestamp 1694700623
transform 1 0 3588 0 1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_106_29
timestamp 1694700623
transform 1 0 3772 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_41
timestamp 1694700623
transform 1 0 4876 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_53
timestamp 1694700623
transform 1 0 5980 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_106_65
timestamp 1694700623
transform 1 0 7084 0 1 59840
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_106_69
timestamp 1694700623
transform 1 0 7452 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_106_79
timestamp 1694700623
transform 1 0 8372 0 1 59840
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_106_83
timestamp 1694700623
transform 1 0 8740 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_106_85
timestamp 1694700623
transform 1 0 8924 0 1 59840
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_106_96
timestamp 1694700623
transform 1 0 9936 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_108
timestamp 1694700623
transform 1 0 11040 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_120
timestamp 1694700623
transform 1 0 12144 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_106_132
timestamp 1694700623
transform 1 0 13248 0 1 59840
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_106_141
timestamp 1694700623
transform 1 0 14076 0 1 59840
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_106_159
timestamp 1694700623
transform 1 0 15732 0 1 59840
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_106_172
timestamp 1694700623
transform 1 0 16928 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_106_188
timestamp 1694700623
transform 1 0 18400 0 1 59840
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_107_3
timestamp 1694700623
transform 1 0 1380 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_15
timestamp 1694700623
transform 1 0 2484 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_27
timestamp 1694700623
transform 1 0 3588 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_39
timestamp 1694700623
transform 1 0 4692 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_107_51
timestamp 1694700623
transform 1 0 5796 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_107_54
timestamp 1694700623
transform 1 0 6072 0 -1 60928
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_107_57
timestamp 1694700623
transform 1 0 6348 0 -1 60928
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_107_76
timestamp 1694700623
transform 1 0 8096 0 -1 60928
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_107_80
timestamp 1694700623
transform 1 0 8464 0 -1 60928
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_107_84
timestamp 1694700623
transform 1 0 8832 0 -1 60928
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_107_94
timestamp 1694700623
transform 1 0 9752 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_107_106
timestamp 1694700623
transform 1 0 10856 0 -1 60928
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_107_113
timestamp 1694700623
transform 1 0 11500 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_125
timestamp 1694700623
transform 1 0 12604 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_137
timestamp 1694700623
transform 1 0 13708 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_149
timestamp 1694700623
transform 1 0 14812 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_107_161
timestamp 1694700623
transform 1 0 15916 0 -1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_107_167
timestamp 1694700623
transform 1 0 16468 0 -1 60928
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_107_169
timestamp 1694700623
transform 1 0 16652 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_107_181
timestamp 1694700623
transform 1 0 17756 0 -1 60928
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_107_189
timestamp 1694700623
transform 1 0 18492 0 -1 60928
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_108_3
timestamp 1694700623
transform 1 0 1380 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_108_15
timestamp 1694700623
transform 1 0 2484 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_108_27
timestamp 1694700623
transform 1 0 3588 0 1 60928
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_108_29
timestamp 1694700623
transform 1 0 3772 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_108_41
timestamp 1694700623
transform 1 0 4876 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_108_53
timestamp 1694700623
transform 1 0 5980 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_108_65
timestamp 1694700623
transform 1 0 7084 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_108_77
timestamp 1694700623
transform 1 0 8188 0 1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_108_83
timestamp 1694700623
transform 1 0 8740 0 1 60928
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_108_85
timestamp 1694700623
transform 1 0 8924 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_108_97
timestamp 1694700623
transform 1 0 10028 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_108_109
timestamp 1694700623
transform 1 0 11132 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_108_121
timestamp 1694700623
transform 1 0 12236 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_108_133
timestamp 1694700623
transform 1 0 13340 0 1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_108_139
timestamp 1694700623
transform 1 0 13892 0 1 60928
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_108_141
timestamp 1694700623
transform 1 0 14076 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_108_153
timestamp 1694700623
transform 1 0 15180 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_108_159
timestamp 1694700623
transform 1 0 15732 0 1 60928
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_108_177
timestamp 1694700623
transform 1 0 17388 0 1 60928
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_108_181
timestamp 1694700623
transform 1 0 17756 0 1 60928
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_108_189
timestamp 1694700623
transform 1 0 18492 0 1 60928
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_109_3
timestamp 1694700623
transform 1 0 1380 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_109_15
timestamp 1694700623
transform 1 0 2484 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_109_27
timestamp 1694700623
transform 1 0 3588 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_109_39
timestamp 1694700623
transform 1 0 4692 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_109_51
timestamp 1694700623
transform 1 0 5796 0 -1 62016
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_109_55
timestamp 1694700623
transform 1 0 6164 0 -1 62016
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_109_57
timestamp 1694700623
transform 1 0 6348 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_109_69
timestamp 1694700623
transform 1 0 7452 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_109_81
timestamp 1694700623
transform 1 0 8556 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_109_93
timestamp 1694700623
transform 1 0 9660 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_109_105
timestamp 1694700623
transform 1 0 10764 0 -1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_109_111
timestamp 1694700623
transform 1 0 11316 0 -1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_109_113
timestamp 1694700623
transform 1 0 11500 0 -1 62016
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_109_124
timestamp 1694700623
transform 1 0 12512 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_109_136
timestamp 1694700623
transform 1 0 13616 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_109_148
timestamp 1694700623
transform 1 0 14720 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_109_160
timestamp 1694700623
transform 1 0 15824 0 -1 62016
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_109_169
timestamp 1694700623
transform 1 0 16652 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_109_181
timestamp 1694700623
transform 1 0 17756 0 -1 62016
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_109_189
timestamp 1694700623
transform 1 0 18492 0 -1 62016
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_110_3
timestamp 1694700623
transform 1 0 1380 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_110_15
timestamp 1694700623
transform 1 0 2484 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_110_27
timestamp 1694700623
transform 1 0 3588 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_110_29
timestamp 1694700623
transform 1 0 3772 0 1 62016
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_110_37
timestamp 1694700623
transform 1 0 4508 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_110_49
timestamp 1694700623
transform 1 0 5612 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_110_61
timestamp 1694700623
transform 1 0 6716 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_110_73
timestamp 1694700623
transform 1 0 7820 0 1 62016
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_110_81
timestamp 1694700623
transform 1 0 8556 0 1 62016
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_110_85
timestamp 1694700623
transform 1 0 8924 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_110_97
timestamp 1694700623
transform 1 0 10028 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_110_109
timestamp 1694700623
transform 1 0 11132 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_110_121
timestamp 1694700623
transform 1 0 12236 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_110_133
timestamp 1694700623
transform 1 0 13340 0 1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_110_139
timestamp 1694700623
transform 1 0 13892 0 1 62016
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_110_141
timestamp 1694700623
transform 1 0 14076 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_110_153
timestamp 1694700623
transform 1 0 15180 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_110_165
timestamp 1694700623
transform 1 0 16284 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_110_177
timestamp 1694700623
transform 1 0 17388 0 1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_110_183
timestamp 1694700623
transform 1 0 17940 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_110_188
timestamp 1694700623
transform 1 0 18400 0 1 62016
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_111_3
timestamp 1694700623
transform 1 0 1380 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_111_15
timestamp 1694700623
transform 1 0 2484 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_111_27
timestamp 1694700623
transform 1 0 3588 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_111_39
timestamp 1694700623
transform 1 0 4692 0 -1 63104
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_111_47
timestamp 1694700623
transform 1 0 5428 0 -1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_111_50
timestamp 1694700623
transform 1 0 5704 0 -1 63104
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_111_54
timestamp 1694700623
transform 1 0 6072 0 -1 63104
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_111_57
timestamp 1694700623
transform 1 0 6348 0 -1 63104
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_111_76
timestamp 1694700623
transform 1 0 8096 0 -1 63104
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_111_80
timestamp 1694700623
transform 1 0 8464 0 -1 63104
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_111_84
timestamp 1694700623
transform 1 0 8832 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_111_96
timestamp 1694700623
transform 1 0 9936 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_111_108
timestamp 1694700623
transform 1 0 11040 0 -1 63104
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_111_113
timestamp 1694700623
transform 1 0 11500 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_111_125
timestamp 1694700623
transform 1 0 12604 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_111_137
timestamp 1694700623
transform 1 0 13708 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_111_149
timestamp 1694700623
transform 1 0 14812 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_111_161
timestamp 1694700623
transform 1 0 15916 0 -1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_111_167
timestamp 1694700623
transform 1 0 16468 0 -1 63104
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_111_169
timestamp 1694700623
transform 1 0 16652 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_111_181
timestamp 1694700623
transform 1 0 17756 0 -1 63104
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_111_189
timestamp 1694700623
transform 1 0 18492 0 -1 63104
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_112_3
timestamp 1694700623
transform 1 0 1380 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_112_15
timestamp 1694700623
transform 1 0 2484 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_112_27
timestamp 1694700623
transform 1 0 3588 0 1 63104
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_112_29
timestamp 1694700623
transform 1 0 3772 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_112_41
timestamp 1694700623
transform 1 0 4876 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_112_53
timestamp 1694700623
transform 1 0 5980 0 1 63104
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_112_59
timestamp 1694700623
transform 1 0 6532 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_112_71
timestamp 1694700623
transform 1 0 7636 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_112_83
timestamp 1694700623
transform 1 0 8740 0 1 63104
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_112_85
timestamp 1694700623
transform 1 0 8924 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_112_97
timestamp 1694700623
transform 1 0 10028 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_112_109
timestamp 1694700623
transform 1 0 11132 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_112_121
timestamp 1694700623
transform 1 0 12236 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_112_133
timestamp 1694700623
transform 1 0 13340 0 1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_112_139
timestamp 1694700623
transform 1 0 13892 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_112_141
timestamp 1694700623
transform 1 0 14076 0 1 63104
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_112_147
timestamp 1694700623
transform 1 0 14628 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_112_159
timestamp 1694700623
transform 1 0 15732 0 1 63104
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_112_168
timestamp 1694700623
transform 1 0 16560 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_112_180
timestamp 1694700623
transform 1 0 17664 0 1 63104
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_112_188
timestamp 1694700623
transform 1 0 18400 0 1 63104
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_113_3
timestamp 1694700623
transform 1 0 1380 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_113_15
timestamp 1694700623
transform 1 0 2484 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_113_27
timestamp 1694700623
transform 1 0 3588 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_113_39
timestamp 1694700623
transform 1 0 4692 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_113_51
timestamp 1694700623
transform 1 0 5796 0 -1 64192
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_113_55
timestamp 1694700623
transform 1 0 6164 0 -1 64192
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_113_57
timestamp 1694700623
transform 1 0 6348 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_113_69
timestamp 1694700623
transform 1 0 7452 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_113_81
timestamp 1694700623
transform 1 0 8556 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_113_93
timestamp 1694700623
transform 1 0 9660 0 -1 64192
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_113_101
timestamp 1694700623
transform 1 0 10396 0 -1 64192
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_113_106
timestamp 1694700623
transform 1 0 10856 0 -1 64192
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_113_110
timestamp 1694700623
transform 1 0 11224 0 -1 64192
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_113_113
timestamp 1694700623
transform 1 0 11500 0 -1 64192
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_113_126
timestamp 1694700623
transform 1 0 12696 0 -1 64192
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_113_130
timestamp 1694700623
transform 1 0 13064 0 -1 64192
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_113_134
timestamp 1694700623
transform 1 0 13432 0 -1 64192
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_113_138
timestamp 1694700623
transform 1 0 13800 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_113_150
timestamp 1694700623
transform 1 0 14904 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_113_162
timestamp 1694700623
transform 1 0 16008 0 -1 64192
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_113_169
timestamp 1694700623
transform 1 0 16652 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_113_181
timestamp 1694700623
transform 1 0 17756 0 -1 64192
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_113_188
timestamp 1694700623
transform 1 0 18400 0 -1 64192
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_114_3
timestamp 1694700623
transform 1 0 1380 0 1 64192
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_114_11
timestamp 1694700623
transform 1 0 2116 0 1 64192
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_114_17
timestamp 1694700623
transform 1 0 2668 0 1 64192
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_114_25
timestamp 1694700623
transform 1 0 3404 0 1 64192
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_114_29
timestamp 1694700623
transform 1 0 3772 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_114_41
timestamp 1694700623
transform 1 0 4876 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_114_53
timestamp 1694700623
transform 1 0 5980 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_114_65
timestamp 1694700623
transform 1 0 7084 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_114_77
timestamp 1694700623
transform 1 0 8188 0 1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_114_83
timestamp 1694700623
transform 1 0 8740 0 1 64192
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_114_85
timestamp 1694700623
transform 1 0 8924 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_114_97
timestamp 1694700623
transform 1 0 10028 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_114_109
timestamp 1694700623
transform 1 0 11132 0 1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_114_115
timestamp 1694700623
transform 1 0 11684 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_114_133
timestamp 1694700623
transform 1 0 13340 0 1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_114_139
timestamp 1694700623
transform 1 0 13892 0 1 64192
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_114_141
timestamp 1694700623
transform 1 0 14076 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_114_153
timestamp 1694700623
transform 1 0 15180 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_114_165
timestamp 1694700623
transform 1 0 16284 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_114_177
timestamp 1694700623
transform 1 0 17388 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_114_189
timestamp 1694700623
transform 1 0 18492 0 1 64192
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_115_3
timestamp 1694700623
transform 1 0 1380 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_115_15
timestamp 1694700623
transform 1 0 2484 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_115_27
timestamp 1694700623
transform 1 0 3588 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_115_39
timestamp 1694700623
transform 1 0 4692 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_115_51
timestamp 1694700623
transform 1 0 5796 0 -1 65280
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_115_55
timestamp 1694700623
transform 1 0 6164 0 -1 65280
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_115_57
timestamp 1694700623
transform 1 0 6348 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_115_69
timestamp 1694700623
transform 1 0 7452 0 -1 65280
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_115_73
timestamp 1694700623
transform 1 0 7820 0 -1 65280
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_115_83
timestamp 1694700623
transform 1 0 8740 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_115_95
timestamp 1694700623
transform 1 0 9844 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_115_107
timestamp 1694700623
transform 1 0 10948 0 -1 65280
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_115_111
timestamp 1694700623
transform 1 0 11316 0 -1 65280
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_115_113
timestamp 1694700623
transform 1 0 11500 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_115_125
timestamp 1694700623
transform 1 0 12604 0 -1 65280
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_115_145
timestamp 1694700623
transform 1 0 14444 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_115_157
timestamp 1694700623
transform 1 0 15548 0 -1 65280
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_115_165
timestamp 1694700623
transform 1 0 16284 0 -1 65280
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_115_169
timestamp 1694700623
transform 1 0 16652 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_115_181
timestamp 1694700623
transform 1 0 17756 0 -1 65280
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_115_188
timestamp 1694700623
transform 1 0 18400 0 -1 65280
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_116_3
timestamp 1694700623
transform 1 0 1380 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_116_15
timestamp 1694700623
transform 1 0 2484 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_116_27
timestamp 1694700623
transform 1 0 3588 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_116_29
timestamp 1694700623
transform 1 0 3772 0 1 65280
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_116_40
timestamp 1694700623
transform 1 0 4784 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_116_52
timestamp 1694700623
transform 1 0 5888 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_116_64
timestamp 1694700623
transform 1 0 6992 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_116_76
timestamp 1694700623
transform 1 0 8096 0 1 65280
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_116_85
timestamp 1694700623
transform 1 0 8924 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_116_97
timestamp 1694700623
transform 1 0 10028 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_116_111
timestamp 1694700623
transform 1 0 11316 0 1 65280
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_116_125
timestamp 1694700623
transform 1 0 12604 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_116_137
timestamp 1694700623
transform 1 0 13708 0 1 65280
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_116_141
timestamp 1694700623
transform 1 0 14076 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_116_153
timestamp 1694700623
transform 1 0 15180 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_116_165
timestamp 1694700623
transform 1 0 16284 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_116_177
timestamp 1694700623
transform 1 0 17388 0 1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_116_183
timestamp 1694700623
transform 1 0 17940 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_116_188
timestamp 1694700623
transform 1 0 18400 0 1 65280
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_117_3
timestamp 1694700623
transform 1 0 1380 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_15
timestamp 1694700623
transform 1 0 2484 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_27
timestamp 1694700623
transform 1 0 3588 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_39
timestamp 1694700623
transform 1 0 4692 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_117_51
timestamp 1694700623
transform 1 0 5796 0 -1 66368
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_117_55
timestamp 1694700623
transform 1 0 6164 0 -1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_117_57
timestamp 1694700623
transform 1 0 6348 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_69
timestamp 1694700623
transform 1 0 7452 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_81
timestamp 1694700623
transform 1 0 8556 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_93
timestamp 1694700623
transform 1 0 9660 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_117_105
timestamp 1694700623
transform 1 0 10764 0 -1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_117_111
timestamp 1694700623
transform 1 0 11316 0 -1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_117_113
timestamp 1694700623
transform 1 0 11500 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_117_125
timestamp 1694700623
transform 1 0 12604 0 -1 66368
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_117_133
timestamp 1694700623
transform 1 0 13340 0 -1 66368
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_117_152
timestamp 1694700623
transform 1 0 15088 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_117_164
timestamp 1694700623
transform 1 0 16192 0 -1 66368
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_117_169
timestamp 1694700623
transform 1 0 16652 0 -1 66368
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_117_186
timestamp 1694700623
transform 1 0 18216 0 -1 66368
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_118_3
timestamp 1694700623
transform 1 0 1380 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_15
timestamp 1694700623
transform 1 0 2484 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_118_27
timestamp 1694700623
transform 1 0 3588 0 1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_118_29
timestamp 1694700623
transform 1 0 3772 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_41
timestamp 1694700623
transform 1 0 4876 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_53
timestamp 1694700623
transform 1 0 5980 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_65
timestamp 1694700623
transform 1 0 7084 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_118_77
timestamp 1694700623
transform 1 0 8188 0 1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_118_83
timestamp 1694700623
transform 1 0 8740 0 1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_118_85
timestamp 1694700623
transform 1 0 8924 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_97
timestamp 1694700623
transform 1 0 10028 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_109
timestamp 1694700623
transform 1 0 11132 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_121
timestamp 1694700623
transform 1 0 12236 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_118_133
timestamp 1694700623
transform 1 0 13340 0 1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_118_139
timestamp 1694700623
transform 1 0 13892 0 1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_118_141
timestamp 1694700623
transform 1 0 14076 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_153
timestamp 1694700623
transform 1 0 15180 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_165
timestamp 1694700623
transform 1 0 16284 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_177
timestamp 1694700623
transform 1 0 17388 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_118_189
timestamp 1694700623
transform 1 0 18492 0 1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_119_3
timestamp 1694700623
transform 1 0 1380 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_15
timestamp 1694700623
transform 1 0 2484 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_27
timestamp 1694700623
transform 1 0 3588 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_39
timestamp 1694700623
transform 1 0 4692 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_119_51
timestamp 1694700623
transform 1 0 5796 0 -1 67456
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_119_55
timestamp 1694700623
transform 1 0 6164 0 -1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_119_57
timestamp 1694700623
transform 1 0 6348 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_119_69
timestamp 1694700623
transform 1 0 7452 0 -1 67456
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_119_73
timestamp 1694700623
transform 1 0 7820 0 -1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_119_78
timestamp 1694700623
transform 1 0 8280 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_90
timestamp 1694700623
transform 1 0 9384 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_119_102
timestamp 1694700623
transform 1 0 10488 0 -1 67456
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_119_110
timestamp 1694700623
transform 1 0 11224 0 -1 67456
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_119_113
timestamp 1694700623
transform 1 0 11500 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_125
timestamp 1694700623
transform 1 0 12604 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_137
timestamp 1694700623
transform 1 0 13708 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_149
timestamp 1694700623
transform 1 0 14812 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_119_161
timestamp 1694700623
transform 1 0 15916 0 -1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_119_167
timestamp 1694700623
transform 1 0 16468 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_119_169
timestamp 1694700623
transform 1 0 16652 0 -1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_119_177
timestamp 1694700623
transform 1 0 17388 0 -1 67456
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_119_188
timestamp 1694700623
transform 1 0 18400 0 -1 67456
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_120_3
timestamp 1694700623
transform 1 0 1380 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_15
timestamp 1694700623
transform 1 0 2484 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_120_27
timestamp 1694700623
transform 1 0 3588 0 1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_120_29
timestamp 1694700623
transform 1 0 3772 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_41
timestamp 1694700623
transform 1 0 4876 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_53
timestamp 1694700623
transform 1 0 5980 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_65
timestamp 1694700623
transform 1 0 7084 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_120_77
timestamp 1694700623
transform 1 0 8188 0 1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_120_83
timestamp 1694700623
transform 1 0 8740 0 1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_120_85
timestamp 1694700623
transform 1 0 8924 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_97
timestamp 1694700623
transform 1 0 10028 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_120_109
timestamp 1694700623
transform 1 0 11132 0 1 67456
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_120_117
timestamp 1694700623
transform 1 0 11868 0 1 67456
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_120_121
timestamp 1694700623
transform 1 0 12236 0 1 67456
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_120_126
timestamp 1694700623
transform 1 0 12696 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_120_138
timestamp 1694700623
transform 1 0 13800 0 1 67456
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_120_141
timestamp 1694700623
transform 1 0 14076 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_153
timestamp 1694700623
transform 1 0 15180 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_165
timestamp 1694700623
transform 1 0 16284 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_120_177
timestamp 1694700623
transform 1 0 17388 0 1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_120_183
timestamp 1694700623
transform 1 0 17940 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_120_188
timestamp 1694700623
transform 1 0 18400 0 1 67456
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_121_3
timestamp 1694700623
transform 1 0 1380 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_15
timestamp 1694700623
transform 1 0 2484 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_27
timestamp 1694700623
transform 1 0 3588 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_39
timestamp 1694700623
transform 1 0 4692 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_121_51
timestamp 1694700623
transform 1 0 5796 0 -1 68544
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_121_55
timestamp 1694700623
transform 1 0 6164 0 -1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_121_57
timestamp 1694700623
transform 1 0 6348 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_69
timestamp 1694700623
transform 1 0 7452 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_81
timestamp 1694700623
transform 1 0 8556 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_93
timestamp 1694700623
transform 1 0 9660 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_121_105
timestamp 1694700623
transform 1 0 10764 0 -1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_121_111
timestamp 1694700623
transform 1 0 11316 0 -1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_121_113
timestamp 1694700623
transform 1 0 11500 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_125
timestamp 1694700623
transform 1 0 12604 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_137
timestamp 1694700623
transform 1 0 13708 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_149
timestamp 1694700623
transform 1 0 14812 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_121_161
timestamp 1694700623
transform 1 0 15916 0 -1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_121_167
timestamp 1694700623
transform 1 0 16468 0 -1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_121_169
timestamp 1694700623
transform 1 0 16652 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_121_181
timestamp 1694700623
transform 1 0 17756 0 -1 68544
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_121_189
timestamp 1694700623
transform 1 0 18492 0 -1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_122_3
timestamp 1694700623
transform 1 0 1380 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_15
timestamp 1694700623
transform 1 0 2484 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_122_27
timestamp 1694700623
transform 1 0 3588 0 1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_122_29
timestamp 1694700623
transform 1 0 3772 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_41
timestamp 1694700623
transform 1 0 4876 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_53
timestamp 1694700623
transform 1 0 5980 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_65
timestamp 1694700623
transform 1 0 7084 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_122_77
timestamp 1694700623
transform 1 0 8188 0 1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_122_83
timestamp 1694700623
transform 1 0 8740 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_122_85
timestamp 1694700623
transform 1 0 8924 0 1 68544
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_122_104
timestamp 1694700623
transform 1 0 10672 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_116
timestamp 1694700623
transform 1 0 11776 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_128
timestamp 1694700623
transform 1 0 12880 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_122_141
timestamp 1694700623
transform 1 0 14076 0 1 68544
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_122_159
timestamp 1694700623
transform 1 0 15732 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_171
timestamp 1694700623
transform 1 0 16836 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_122_183
timestamp 1694700623
transform 1 0 17940 0 1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_122_189
timestamp 1694700623
transform 1 0 18492 0 1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_123_3
timestamp 1694700623
transform 1 0 1380 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_15
timestamp 1694700623
transform 1 0 2484 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_27
timestamp 1694700623
transform 1 0 3588 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_39
timestamp 1694700623
transform 1 0 4692 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_123_51
timestamp 1694700623
transform 1 0 5796 0 -1 69632
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_123_55
timestamp 1694700623
transform 1 0 6164 0 -1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_123_57
timestamp 1694700623
transform 1 0 6348 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_69
timestamp 1694700623
transform 1 0 7452 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_81
timestamp 1694700623
transform 1 0 8556 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_123_110
timestamp 1694700623
transform 1 0 11224 0 -1 69632
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_123_113
timestamp 1694700623
transform 1 0 11500 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_125
timestamp 1694700623
transform 1 0 12604 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_137
timestamp 1694700623
transform 1 0 13708 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_149
timestamp 1694700623
transform 1 0 14812 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_123_161
timestamp 1694700623
transform 1 0 15916 0 -1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_123_167
timestamp 1694700623
transform 1 0 16468 0 -1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_123_169
timestamp 1694700623
transform 1 0 16652 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_123_181
timestamp 1694700623
transform 1 0 17756 0 -1 69632
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_123_189
timestamp 1694700623
transform 1 0 18492 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_124_3
timestamp 1694700623
transform 1 0 1380 0 1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_124_18
timestamp 1694700623
transform 1 0 2760 0 1 69632
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_124_22
timestamp 1694700623
transform 1 0 3128 0 1 69632
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_124_26
timestamp 1694700623
transform 1 0 3496 0 1 69632
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_124_29
timestamp 1694700623
transform 1 0 3772 0 1 69632
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_124_35
timestamp 1694700623
transform 1 0 4324 0 1 69632
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_124_39
timestamp 1694700623
transform 1 0 4692 0 1 69632
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_124_43
timestamp 1694700623
transform 1 0 5060 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_124_55
timestamp 1694700623
transform 1 0 6164 0 1 69632
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_124_63
timestamp 1694700623
transform 1 0 6900 0 1 69632
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_124_82
timestamp 1694700623
transform 1 0 8648 0 1 69632
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_124_85
timestamp 1694700623
transform 1 0 8924 0 1 69632
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_124_97
timestamp 1694700623
transform 1 0 10028 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_109
timestamp 1694700623
transform 1 0 11132 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_121
timestamp 1694700623
transform 1 0 12236 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_124_133
timestamp 1694700623
transform 1 0 13340 0 1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_124_139
timestamp 1694700623
transform 1 0 13892 0 1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_124_141
timestamp 1694700623
transform 1 0 14076 0 1 69632
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_124_149
timestamp 1694700623
transform 1 0 14812 0 1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_124_159
timestamp 1694700623
transform 1 0 15732 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_171
timestamp 1694700623
transform 1 0 16836 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_124_183
timestamp 1694700623
transform 1 0 17940 0 1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_124_188
timestamp 1694700623
transform 1 0 18400 0 1 69632
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_125_3
timestamp 1694700623
transform 1 0 1380 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_15
timestamp 1694700623
transform 1 0 2484 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_27
timestamp 1694700623
transform 1 0 3588 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_39
timestamp 1694700623
transform 1 0 4692 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_125_51
timestamp 1694700623
transform 1 0 5796 0 -1 70720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_125_55
timestamp 1694700623
transform 1 0 6164 0 -1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_125_57
timestamp 1694700623
transform 1 0 6348 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_69
timestamp 1694700623
transform 1 0 7452 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_81
timestamp 1694700623
transform 1 0 8556 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_93
timestamp 1694700623
transform 1 0 9660 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_125_105
timestamp 1694700623
transform 1 0 10764 0 -1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_125_111
timestamp 1694700623
transform 1 0 11316 0 -1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_125_113
timestamp 1694700623
transform 1 0 11500 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_125
timestamp 1694700623
transform 1 0 12604 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_137
timestamp 1694700623
transform 1 0 13708 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_149
timestamp 1694700623
transform 1 0 14812 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_125_161
timestamp 1694700623
transform 1 0 15916 0 -1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_125_167
timestamp 1694700623
transform 1 0 16468 0 -1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_125_169
timestamp 1694700623
transform 1 0 16652 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_125_181
timestamp 1694700623
transform 1 0 17756 0 -1 70720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_125_189
timestamp 1694700623
transform 1 0 18492 0 -1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_126_3
timestamp 1694700623
transform 1 0 1380 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_15
timestamp 1694700623
transform 1 0 2484 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_126_27
timestamp 1694700623
transform 1 0 3588 0 1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_126_29
timestamp 1694700623
transform 1 0 3772 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_41
timestamp 1694700623
transform 1 0 4876 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_70
timestamp 1694700623
transform 1 0 7544 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_126_82
timestamp 1694700623
transform 1 0 8648 0 1 70720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_126_85
timestamp 1694700623
transform 1 0 8924 0 1 70720
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_126_104
timestamp 1694700623
transform 1 0 10672 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_116
timestamp 1694700623
transform 1 0 11776 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_128
timestamp 1694700623
transform 1 0 12880 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_141
timestamp 1694700623
transform 1 0 14076 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_126_153
timestamp 1694700623
transform 1 0 15180 0 1 70720
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_126_172
timestamp 1694700623
transform 1 0 16928 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_126_184
timestamp 1694700623
transform 1 0 18032 0 1 70720
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_127_3
timestamp 1694700623
transform 1 0 1380 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_127_15
timestamp 1694700623
transform 1 0 2484 0 -1 71808
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_127_38
timestamp 1694700623
transform 1 0 4600 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_127_50
timestamp 1694700623
transform 1 0 5704 0 -1 71808
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_127_57
timestamp 1694700623
transform 1 0 6348 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_69
timestamp 1694700623
transform 1 0 7452 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_81
timestamp 1694700623
transform 1 0 8556 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_93
timestamp 1694700623
transform 1 0 9660 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_127_105
timestamp 1694700623
transform 1 0 10764 0 -1 71808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_127_111
timestamp 1694700623
transform 1 0 11316 0 -1 71808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_127_113
timestamp 1694700623
transform 1 0 11500 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_125
timestamp 1694700623
transform 1 0 12604 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_137
timestamp 1694700623
transform 1 0 13708 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_149
timestamp 1694700623
transform 1 0 14812 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_127_161
timestamp 1694700623
transform 1 0 15916 0 -1 71808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_127_167
timestamp 1694700623
transform 1 0 16468 0 -1 71808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_127_169
timestamp 1694700623
transform 1 0 16652 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_127_181
timestamp 1694700623
transform 1 0 17756 0 -1 71808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_127_188
timestamp 1694700623
transform 1 0 18400 0 -1 71808
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_128_3
timestamp 1694700623
transform 1 0 1380 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_15
timestamp 1694700623
transform 1 0 2484 0 1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_128_27
timestamp 1694700623
transform 1 0 3588 0 1 71808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_128_29
timestamp 1694700623
transform 1 0 3772 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_41
timestamp 1694700623
transform 1 0 4876 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_53
timestamp 1694700623
transform 1 0 5980 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_65
timestamp 1694700623
transform 1 0 7084 0 1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_128_77
timestamp 1694700623
transform 1 0 8188 0 1 71808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_128_83
timestamp 1694700623
transform 1 0 8740 0 1 71808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_128_85
timestamp 1694700623
transform 1 0 8924 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_97
timestamp 1694700623
transform 1 0 10028 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_109
timestamp 1694700623
transform 1 0 11132 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_121
timestamp 1694700623
transform 1 0 12236 0 1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_128_133
timestamp 1694700623
transform 1 0 13340 0 1 71808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_128_139
timestamp 1694700623
transform 1 0 13892 0 1 71808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_128_141
timestamp 1694700623
transform 1 0 14076 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_153
timestamp 1694700623
transform 1 0 15180 0 1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_128_165
timestamp 1694700623
transform 1 0 16284 0 1 71808
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_128_176
timestamp 1694700623
transform 1 0 17296 0 1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_128_188
timestamp 1694700623
transform 1 0 18400 0 1 71808
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_129_3
timestamp 1694700623
transform 1 0 1380 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_15
timestamp 1694700623
transform 1 0 2484 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_27
timestamp 1694700623
transform 1 0 3588 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_39
timestamp 1694700623
transform 1 0 4692 0 -1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_129_51
timestamp 1694700623
transform 1 0 5796 0 -1 72896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_129_55
timestamp 1694700623
transform 1 0 6164 0 -1 72896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_129_57
timestamp 1694700623
transform 1 0 6348 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_69
timestamp 1694700623
transform 1 0 7452 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_81
timestamp 1694700623
transform 1 0 8556 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_93
timestamp 1694700623
transform 1 0 9660 0 -1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_129_105
timestamp 1694700623
transform 1 0 10764 0 -1 72896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_129_111
timestamp 1694700623
transform 1 0 11316 0 -1 72896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_129_113
timestamp 1694700623
transform 1 0 11500 0 -1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_129_125
timestamp 1694700623
transform 1 0 12604 0 -1 72896
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_129_136
timestamp 1694700623
transform 1 0 13616 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_148
timestamp 1694700623
transform 1 0 14720 0 -1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_129_160
timestamp 1694700623
transform 1 0 15824 0 -1 72896
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_129_169
timestamp 1694700623
transform 1 0 16652 0 -1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_129_181
timestamp 1694700623
transform 1 0 17756 0 -1 72896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_129_189
timestamp 1694700623
transform 1 0 18492 0 -1 72896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_130_3
timestamp 1694700623
transform 1 0 1380 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_15
timestamp 1694700623
transform 1 0 2484 0 1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_130_27
timestamp 1694700623
transform 1 0 3588 0 1 72896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_130_29
timestamp 1694700623
transform 1 0 3772 0 1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_130_41
timestamp 1694700623
transform 1 0 4876 0 1 72896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_130_47
timestamp 1694700623
transform 1 0 5428 0 1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_130_50
timestamp 1694700623
transform 1 0 5704 0 1 72896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_130_54
timestamp 1694700623
transform 1 0 6072 0 1 72896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_130_58
timestamp 1694700623
transform 1 0 6440 0 1 72896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_130_76
timestamp 1694700623
transform 1 0 8096 0 1 72896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_130_80
timestamp 1694700623
transform 1 0 8464 0 1 72896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_130_85
timestamp 1694700623
transform 1 0 8924 0 1 72896
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_130_89
timestamp 1694700623
transform 1 0 9292 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_101
timestamp 1694700623
transform 1 0 10396 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_113
timestamp 1694700623
transform 1 0 11500 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_125
timestamp 1694700623
transform 1 0 12604 0 1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_130_137
timestamp 1694700623
transform 1 0 13708 0 1 72896
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_130_141
timestamp 1694700623
transform 1 0 14076 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_153
timestamp 1694700623
transform 1 0 15180 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_165
timestamp 1694700623
transform 1 0 16284 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_177
timestamp 1694700623
transform 1 0 17388 0 1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_130_189
timestamp 1694700623
transform 1 0 18492 0 1 72896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_131_3
timestamp 1694700623
transform 1 0 1380 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_15
timestamp 1694700623
transform 1 0 2484 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_27
timestamp 1694700623
transform 1 0 3588 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_39
timestamp 1694700623
transform 1 0 4692 0 -1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_131_51
timestamp 1694700623
transform 1 0 5796 0 -1 73984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_131_55
timestamp 1694700623
transform 1 0 6164 0 -1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_131_57
timestamp 1694700623
transform 1 0 6348 0 -1 73984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_131_65
timestamp 1694700623
transform 1 0 7084 0 -1 73984
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_131_76
timestamp 1694700623
transform 1 0 8096 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_88
timestamp 1694700623
transform 1 0 9200 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_100
timestamp 1694700623
transform 1 0 10304 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_113
timestamp 1694700623
transform 1 0 11500 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_125
timestamp 1694700623
transform 1 0 12604 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_137
timestamp 1694700623
transform 1 0 13708 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_149
timestamp 1694700623
transform 1 0 14812 0 -1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_131_161
timestamp 1694700623
transform 1 0 15916 0 -1 73984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_131_167
timestamp 1694700623
transform 1 0 16468 0 -1 73984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_131_169
timestamp 1694700623
transform 1 0 16652 0 -1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_131_181
timestamp 1694700623
transform 1 0 17756 0 -1 73984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_131_188
timestamp 1694700623
transform 1 0 18400 0 -1 73984
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_132_3
timestamp 1694700623
transform 1 0 1380 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_15
timestamp 1694700623
transform 1 0 2484 0 1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_132_27
timestamp 1694700623
transform 1 0 3588 0 1 73984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_132_29
timestamp 1694700623
transform 1 0 3772 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_41
timestamp 1694700623
transform 1 0 4876 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_53
timestamp 1694700623
transform 1 0 5980 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_65
timestamp 1694700623
transform 1 0 7084 0 1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_132_77
timestamp 1694700623
transform 1 0 8188 0 1 73984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_132_83
timestamp 1694700623
transform 1 0 8740 0 1 73984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_132_85
timestamp 1694700623
transform 1 0 8924 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_97
timestamp 1694700623
transform 1 0 10028 0 1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_132_109
timestamp 1694700623
transform 1 0 11132 0 1 73984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_132_117
timestamp 1694700623
transform 1 0 11868 0 1 73984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_132_128
timestamp 1694700623
transform 1 0 12880 0 1 73984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_132_138
timestamp 1694700623
transform 1 0 13800 0 1 73984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_132_141
timestamp 1694700623
transform 1 0 14076 0 1 73984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_132_159
timestamp 1694700623
transform 1 0 15732 0 1 73984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_132_163
timestamp 1694700623
transform 1 0 16100 0 1 73984
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_132_167
timestamp 1694700623
transform 1 0 16468 0 1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_132_179
timestamp 1694700623
transform 1 0 17572 0 1 73984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_132_187
timestamp 1694700623
transform 1 0 18308 0 1 73984
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_133_3
timestamp 1694700623
transform 1 0 1380 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_15
timestamp 1694700623
transform 1 0 2484 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_27
timestamp 1694700623
transform 1 0 3588 0 -1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_133_48
timestamp 1694700623
transform 1 0 5520 0 -1 75072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_133_57
timestamp 1694700623
transform 1 0 6348 0 -1 75072
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_133_63
timestamp 1694700623
transform 1 0 6900 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_75
timestamp 1694700623
transform 1 0 8004 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_87
timestamp 1694700623
transform 1 0 9108 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_99
timestamp 1694700623
transform 1 0 10212 0 -1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_133_111
timestamp 1694700623
transform 1 0 11316 0 -1 75072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_133_113
timestamp 1694700623
transform 1 0 11500 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_125
timestamp 1694700623
transform 1 0 12604 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_137
timestamp 1694700623
transform 1 0 13708 0 -1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_133_166
timestamp 1694700623
transform 1 0 16376 0 -1 75072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_133_169
timestamp 1694700623
transform 1 0 16652 0 -1 75072
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_133_175
timestamp 1694700623
transform 1 0 17204 0 -1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_133_187
timestamp 1694700623
transform 1 0 18308 0 -1 75072
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_134_3
timestamp 1694700623
transform 1 0 1380 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_15
timestamp 1694700623
transform 1 0 2484 0 1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_134_27
timestamp 1694700623
transform 1 0 3588 0 1 75072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_134_29
timestamp 1694700623
transform 1 0 3772 0 1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_134_52
timestamp 1694700623
transform 1 0 5888 0 1 75072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_134_56
timestamp 1694700623
transform 1 0 6256 0 1 75072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_134_60
timestamp 1694700623
transform 1 0 6624 0 1 75072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_134_64
timestamp 1694700623
transform 1 0 6992 0 1 75072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_134_68
timestamp 1694700623
transform 1 0 7360 0 1 75072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_134_74
timestamp 1694700623
transform 1 0 7912 0 1 75072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_134_78
timestamp 1694700623
transform 1 0 8280 0 1 75072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_134_82
timestamp 1694700623
transform 1 0 8648 0 1 75072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_134_85
timestamp 1694700623
transform 1 0 8924 0 1 75072
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_134_89
timestamp 1694700623
transform 1 0 9292 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_101
timestamp 1694700623
transform 1 0 10396 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_113
timestamp 1694700623
transform 1 0 11500 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_125
timestamp 1694700623
transform 1 0 12604 0 1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_134_137
timestamp 1694700623
transform 1 0 13708 0 1 75072
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_134_141
timestamp 1694700623
transform 1 0 14076 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_156
timestamp 1694700623
transform 1 0 15456 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_168
timestamp 1694700623
transform 1 0 16560 0 1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_134_180
timestamp 1694700623
transform 1 0 17664 0 1 75072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_134_188
timestamp 1694700623
transform 1 0 18400 0 1 75072
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_135_3
timestamp 1694700623
transform 1 0 1380 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_15
timestamp 1694700623
transform 1 0 2484 0 -1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_135_27
timestamp 1694700623
transform 1 0 3588 0 -1 76160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_135_48
timestamp 1694700623
transform 1 0 5520 0 -1 76160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_135_57
timestamp 1694700623
transform 1 0 6348 0 -1 76160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_135_71
timestamp 1694700623
transform 1 0 7636 0 -1 76160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_135_77
timestamp 1694700623
transform 1 0 8188 0 -1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_135_80
timestamp 1694700623
transform 1 0 8464 0 -1 76160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_135_86
timestamp 1694700623
transform 1 0 9016 0 -1 76160
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_135_90
timestamp 1694700623
transform 1 0 9384 0 -1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_135_102
timestamp 1694700623
transform 1 0 10488 0 -1 76160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_135_110
timestamp 1694700623
transform 1 0 11224 0 -1 76160
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_135_113
timestamp 1694700623
transform 1 0 11500 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_125
timestamp 1694700623
transform 1 0 12604 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_146
timestamp 1694700623
transform 1 0 14536 0 -1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_135_158
timestamp 1694700623
transform 1 0 15640 0 -1 76160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_135_166
timestamp 1694700623
transform 1 0 16376 0 -1 76160
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_135_169
timestamp 1694700623
transform 1 0 16652 0 -1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_135_181
timestamp 1694700623
transform 1 0 17756 0 -1 76160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_135_189
timestamp 1694700623
transform 1 0 18492 0 -1 76160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_136_3
timestamp 1694700623
transform 1 0 1380 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_15
timestamp 1694700623
transform 1 0 2484 0 1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_136_27
timestamp 1694700623
transform 1 0 3588 0 1 76160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_136_29
timestamp 1694700623
transform 1 0 3772 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_41
timestamp 1694700623
transform 1 0 4876 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_53
timestamp 1694700623
transform 1 0 5980 0 1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_136_67
timestamp 1694700623
transform 1 0 7268 0 1 76160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_136_81
timestamp 1694700623
transform 1 0 8556 0 1 76160
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_136_85
timestamp 1694700623
transform 1 0 8924 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_97
timestamp 1694700623
transform 1 0 10028 0 1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_136_111
timestamp 1694700623
transform 1 0 11316 0 1 76160
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_136_117
timestamp 1694700623
transform 1 0 11868 0 1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_136_129
timestamp 1694700623
transform 1 0 12972 0 1 76160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_136_137
timestamp 1694700623
transform 1 0 13708 0 1 76160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_136_141
timestamp 1694700623
transform 1 0 14076 0 1 76160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_136_149
timestamp 1694700623
transform 1 0 14812 0 1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_136_166
timestamp 1694700623
transform 1 0 16376 0 1 76160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_136_176
timestamp 1694700623
transform 1 0 17296 0 1 76160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_136_180
timestamp 1694700623
transform 1 0 17664 0 1 76160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_136_184
timestamp 1694700623
transform 1 0 18032 0 1 76160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_136_188
timestamp 1694700623
transform 1 0 18400 0 1 76160
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_137_3
timestamp 1694700623
transform 1 0 1380 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_15
timestamp 1694700623
transform 1 0 2484 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_27
timestamp 1694700623
transform 1 0 3588 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_39
timestamp 1694700623
transform 1 0 4692 0 -1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_137_51
timestamp 1694700623
transform 1 0 5796 0 -1 77248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_137_55
timestamp 1694700623
transform 1 0 6164 0 -1 77248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_137_57
timestamp 1694700623
transform 1 0 6348 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_69
timestamp 1694700623
transform 1 0 7452 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_81
timestamp 1694700623
transform 1 0 8556 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_93
timestamp 1694700623
transform 1 0 9660 0 -1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_137_105
timestamp 1694700623
transform 1 0 10764 0 -1 77248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_137_111
timestamp 1694700623
transform 1 0 11316 0 -1 77248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_137_113
timestamp 1694700623
transform 1 0 11500 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_125
timestamp 1694700623
transform 1 0 12604 0 -1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_137_137
timestamp 1694700623
transform 1 0 13708 0 -1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_137_140
timestamp 1694700623
transform 1 0 13984 0 -1 77248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_137_144
timestamp 1694700623
transform 1 0 14352 0 -1 77248
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_137_148
timestamp 1694700623
transform 1 0 14720 0 -1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_137_162
timestamp 1694700623
transform 1 0 16008 0 -1 77248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_137_166
timestamp 1694700623
transform 1 0 16376 0 -1 77248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_137_169
timestamp 1694700623
transform 1 0 16652 0 -1 77248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_137_175
timestamp 1694700623
transform 1 0 17204 0 -1 77248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_137_187
timestamp 1694700623
transform 1 0 18308 0 -1 77248
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_138_3
timestamp 1694700623
transform 1 0 1380 0 1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_138_15
timestamp 1694700623
transform 1 0 2484 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_138_27
timestamp 1694700623
transform 1 0 3588 0 1 77248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_138_29
timestamp 1694700623
transform 1 0 3772 0 1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_138_41
timestamp 1694700623
transform 1 0 4876 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_138_53
timestamp 1694700623
transform 1 0 5980 0 1 77248
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_138_57
timestamp 1694700623
transform 1 0 6348 0 1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_138_69
timestamp 1694700623
transform 1 0 7452 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_138_81
timestamp 1694700623
transform 1 0 8556 0 1 77248
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_138_85
timestamp 1694700623
transform 1 0 8924 0 1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_138_97
timestamp 1694700623
transform 1 0 10028 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_138_109
timestamp 1694700623
transform 1 0 11132 0 1 77248
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_138_113
timestamp 1694700623
transform 1 0 11500 0 1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_138_125
timestamp 1694700623
transform 1 0 12604 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_138_137
timestamp 1694700623
transform 1 0 13708 0 1 77248
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_138_141
timestamp 1694700623
transform 1 0 14076 0 1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_138_153
timestamp 1694700623
transform 1 0 15180 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_138_165
timestamp 1694700623
transform 1 0 16284 0 1 77248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_138_169
timestamp 1694700623
transform 1 0 16652 0 1 77248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_138_173
timestamp 1694700623
transform 1 0 17020 0 1 77248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_138_177
timestamp 1694700623
transform 1 0 17388 0 1 77248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_138_183
timestamp 1694700623
transform 1 0 17940 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_138_188
timestamp 1694700623
transform 1 0 18400 0 1 77248
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  input1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 17848 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input2
timestamp 1694700623
transform 1 0 6532 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 14260 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output4
timestamp 1694700623
transform 1 0 18032 0 1 77248
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output5
timestamp 1694700623
transform 1 0 18032 0 -1 58752
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output6
timestamp 1694700623
transform 1 0 18032 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output7
timestamp 1694700623
transform 1 0 18032 0 1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output8
timestamp 1694700623
transform 1 0 18032 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output9
timestamp 1694700623
transform 1 0 18032 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output10
timestamp 1694700623
transform 1 0 18032 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output11
timestamp 1694700623
transform 1 0 18032 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output12
timestamp 1694700623
transform 1 0 18032 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output13
timestamp 1694700623
transform 1 0 18032 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output14
timestamp 1694700623
transform 1 0 18032 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output15
timestamp 1694700623
transform 1 0 18032 0 1 75072
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output16
timestamp 1694700623
transform 1 0 18032 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output17
timestamp 1694700623
transform 1 0 18032 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output18
timestamp 1694700623
transform 1 0 18032 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output19
timestamp 1694700623
transform 1 0 18032 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output20
timestamp 1694700623
transform 1 0 18032 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output21
timestamp 1694700623
transform 1 0 18032 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output22
timestamp 1694700623
transform 1 0 18032 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output23
timestamp 1694700623
transform 1 0 18032 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output24
timestamp 1694700623
transform 1 0 18032 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output25
timestamp 1694700623
transform 1 0 18032 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output26
timestamp 1694700623
transform 1 0 18032 0 -1 73984
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output27
timestamp 1694700623
transform 1 0 18032 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output28
timestamp 1694700623
transform 1 0 18032 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output29
timestamp 1694700623
transform 1 0 18032 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output30
timestamp 1694700623
transform 1 0 18032 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output31
timestamp 1694700623
transform 1 0 18032 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output32
timestamp 1694700623
transform 1 0 18032 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output33
timestamp 1694700623
transform 1 0 18032 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output34
timestamp 1694700623
transform 1 0 18032 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output35
timestamp 1694700623
transform 1 0 18032 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output36
timestamp 1694700623
transform 1 0 18032 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output37
timestamp 1694700623
transform 1 0 18032 0 -1 71808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output38
timestamp 1694700623
transform 1 0 18032 0 1 69632
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output39
timestamp 1694700623
transform 1 0 18032 0 1 67456
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output40
timestamp 1694700623
transform 1 0 18032 0 1 65280
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output41
timestamp 1694700623
transform 1 0 18032 0 -1 64192
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output42
timestamp 1694700623
transform 1 0 18032 0 1 62016
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output43
timestamp 1694700623
transform 1 0 18032 0 1 59840
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output44
timestamp 1694700623
transform 1 0 10028 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1694700623
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1694700623
transform -1 0 18860 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1694700623
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1694700623
transform -1 0 18860 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1694700623
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1694700623
transform -1 0 18860 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1694700623
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1694700623
transform -1 0 18860 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1694700623
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1694700623
transform -1 0 18860 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1694700623
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1694700623
transform -1 0 18860 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1694700623
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1694700623
transform -1 0 18860 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1694700623
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1694700623
transform -1 0 18860 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1694700623
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1694700623
transform -1 0 18860 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1694700623
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1694700623
transform -1 0 18860 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1694700623
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1694700623
transform -1 0 18860 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1694700623
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1694700623
transform -1 0 18860 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1694700623
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1694700623
transform -1 0 18860 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1694700623
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1694700623
transform -1 0 18860 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1694700623
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1694700623
transform -1 0 18860 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1694700623
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1694700623
transform -1 0 18860 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1694700623
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1694700623
transform -1 0 18860 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1694700623
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1694700623
transform -1 0 18860 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1694700623
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1694700623
transform -1 0 18860 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1694700623
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1694700623
transform -1 0 18860 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1694700623
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1694700623
transform -1 0 18860 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1694700623
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1694700623
transform -1 0 18860 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1694700623
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1694700623
transform -1 0 18860 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1694700623
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1694700623
transform -1 0 18860 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1694700623
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1694700623
transform -1 0 18860 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1694700623
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1694700623
transform -1 0 18860 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1694700623
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1694700623
transform -1 0 18860 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1694700623
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1694700623
transform -1 0 18860 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1694700623
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1694700623
transform -1 0 18860 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1694700623
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1694700623
transform -1 0 18860 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1694700623
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1694700623
transform -1 0 18860 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1694700623
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1694700623
transform -1 0 18860 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1694700623
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1694700623
transform -1 0 18860 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1694700623
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1694700623
transform -1 0 18860 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1694700623
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1694700623
transform -1 0 18860 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1694700623
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1694700623
transform -1 0 18860 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1694700623
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1694700623
transform -1 0 18860 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1694700623
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1694700623
transform -1 0 18860 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1694700623
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1694700623
transform -1 0 18860 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1694700623
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1694700623
transform -1 0 18860 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1694700623
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1694700623
transform -1 0 18860 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1694700623
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1694700623
transform -1 0 18860 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1694700623
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1694700623
transform -1 0 18860 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1694700623
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1694700623
transform -1 0 18860 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1694700623
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1694700623
transform -1 0 18860 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1694700623
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1694700623
transform -1 0 18860 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1694700623
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1694700623
transform -1 0 18860 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1694700623
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1694700623
transform -1 0 18860 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1694700623
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1694700623
transform -1 0 18860 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1694700623
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1694700623
transform -1 0 18860 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1694700623
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1694700623
transform -1 0 18860 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1694700623
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1694700623
transform -1 0 18860 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1694700623
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1694700623
transform -1 0 18860 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1694700623
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1694700623
transform -1 0 18860 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1694700623
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1694700623
transform -1 0 18860 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1694700623
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1694700623
transform -1 0 18860 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1694700623
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1694700623
transform -1 0 18860 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1694700623
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1694700623
transform -1 0 18860 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1694700623
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1694700623
transform -1 0 18860 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1694700623
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1694700623
transform -1 0 18860 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1694700623
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1694700623
transform -1 0 18860 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1694700623
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1694700623
transform -1 0 18860 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1694700623
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1694700623
transform -1 0 18860 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 1694700623
transform 1 0 1104 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 1694700623
transform -1 0 18860 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 1694700623
transform 1 0 1104 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 1694700623
transform -1 0 18860 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_130
timestamp 1694700623
transform 1 0 1104 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_131
timestamp 1694700623
transform -1 0 18860 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_132
timestamp 1694700623
transform 1 0 1104 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_133
timestamp 1694700623
transform -1 0 18860 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_134
timestamp 1694700623
transform 1 0 1104 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_135
timestamp 1694700623
transform -1 0 18860 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_136
timestamp 1694700623
transform 1 0 1104 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_137
timestamp 1694700623
transform -1 0 18860 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_138
timestamp 1694700623
transform 1 0 1104 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_139
timestamp 1694700623
transform -1 0 18860 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_140
timestamp 1694700623
transform 1 0 1104 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_141
timestamp 1694700623
transform -1 0 18860 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_142
timestamp 1694700623
transform 1 0 1104 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_143
timestamp 1694700623
transform -1 0 18860 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_144
timestamp 1694700623
transform 1 0 1104 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_145
timestamp 1694700623
transform -1 0 18860 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_146
timestamp 1694700623
transform 1 0 1104 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_147
timestamp 1694700623
transform -1 0 18860 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_148
timestamp 1694700623
transform 1 0 1104 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_149
timestamp 1694700623
transform -1 0 18860 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_150
timestamp 1694700623
transform 1 0 1104 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_151
timestamp 1694700623
transform -1 0 18860 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_152
timestamp 1694700623
transform 1 0 1104 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_153
timestamp 1694700623
transform -1 0 18860 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_154
timestamp 1694700623
transform 1 0 1104 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_155
timestamp 1694700623
transform -1 0 18860 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_156
timestamp 1694700623
transform 1 0 1104 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_157
timestamp 1694700623
transform -1 0 18860 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_158
timestamp 1694700623
transform 1 0 1104 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_159
timestamp 1694700623
transform -1 0 18860 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_160
timestamp 1694700623
transform 1 0 1104 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_161
timestamp 1694700623
transform -1 0 18860 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_162
timestamp 1694700623
transform 1 0 1104 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_163
timestamp 1694700623
transform -1 0 18860 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_164
timestamp 1694700623
transform 1 0 1104 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_165
timestamp 1694700623
transform -1 0 18860 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_166
timestamp 1694700623
transform 1 0 1104 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_167
timestamp 1694700623
transform -1 0 18860 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_168
timestamp 1694700623
transform 1 0 1104 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_169
timestamp 1694700623
transform -1 0 18860 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_170
timestamp 1694700623
transform 1 0 1104 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_171
timestamp 1694700623
transform -1 0 18860 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_172
timestamp 1694700623
transform 1 0 1104 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_173
timestamp 1694700623
transform -1 0 18860 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_174
timestamp 1694700623
transform 1 0 1104 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_175
timestamp 1694700623
transform -1 0 18860 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_176
timestamp 1694700623
transform 1 0 1104 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_177
timestamp 1694700623
transform -1 0 18860 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_178
timestamp 1694700623
transform 1 0 1104 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_179
timestamp 1694700623
transform -1 0 18860 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_180
timestamp 1694700623
transform 1 0 1104 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_181
timestamp 1694700623
transform -1 0 18860 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_182
timestamp 1694700623
transform 1 0 1104 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_183
timestamp 1694700623
transform -1 0 18860 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_184
timestamp 1694700623
transform 1 0 1104 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_185
timestamp 1694700623
transform -1 0 18860 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_186
timestamp 1694700623
transform 1 0 1104 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_187
timestamp 1694700623
transform -1 0 18860 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_188
timestamp 1694700623
transform 1 0 1104 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_189
timestamp 1694700623
transform -1 0 18860 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_190
timestamp 1694700623
transform 1 0 1104 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_191
timestamp 1694700623
transform -1 0 18860 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_192
timestamp 1694700623
transform 1 0 1104 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_193
timestamp 1694700623
transform -1 0 18860 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_194
timestamp 1694700623
transform 1 0 1104 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_195
timestamp 1694700623
transform -1 0 18860 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_196
timestamp 1694700623
transform 1 0 1104 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_197
timestamp 1694700623
transform -1 0 18860 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_198
timestamp 1694700623
transform 1 0 1104 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_199
timestamp 1694700623
transform -1 0 18860 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_200
timestamp 1694700623
transform 1 0 1104 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_201
timestamp 1694700623
transform -1 0 18860 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_202
timestamp 1694700623
transform 1 0 1104 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_203
timestamp 1694700623
transform -1 0 18860 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_204
timestamp 1694700623
transform 1 0 1104 0 1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_205
timestamp 1694700623
transform -1 0 18860 0 1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_206
timestamp 1694700623
transform 1 0 1104 0 -1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_207
timestamp 1694700623
transform -1 0 18860 0 -1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_208
timestamp 1694700623
transform 1 0 1104 0 1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_209
timestamp 1694700623
transform -1 0 18860 0 1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_210
timestamp 1694700623
transform 1 0 1104 0 -1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_211
timestamp 1694700623
transform -1 0 18860 0 -1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_212
timestamp 1694700623
transform 1 0 1104 0 1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_213
timestamp 1694700623
transform -1 0 18860 0 1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_214
timestamp 1694700623
transform 1 0 1104 0 -1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_215
timestamp 1694700623
transform -1 0 18860 0 -1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_216
timestamp 1694700623
transform 1 0 1104 0 1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_217
timestamp 1694700623
transform -1 0 18860 0 1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_218
timestamp 1694700623
transform 1 0 1104 0 -1 62016
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_219
timestamp 1694700623
transform -1 0 18860 0 -1 62016
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_220
timestamp 1694700623
transform 1 0 1104 0 1 62016
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_221
timestamp 1694700623
transform -1 0 18860 0 1 62016
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_222
timestamp 1694700623
transform 1 0 1104 0 -1 63104
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_223
timestamp 1694700623
transform -1 0 18860 0 -1 63104
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_224
timestamp 1694700623
transform 1 0 1104 0 1 63104
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_225
timestamp 1694700623
transform -1 0 18860 0 1 63104
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_226
timestamp 1694700623
transform 1 0 1104 0 -1 64192
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_227
timestamp 1694700623
transform -1 0 18860 0 -1 64192
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_228
timestamp 1694700623
transform 1 0 1104 0 1 64192
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_229
timestamp 1694700623
transform -1 0 18860 0 1 64192
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_230
timestamp 1694700623
transform 1 0 1104 0 -1 65280
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_231
timestamp 1694700623
transform -1 0 18860 0 -1 65280
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_232
timestamp 1694700623
transform 1 0 1104 0 1 65280
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_233
timestamp 1694700623
transform -1 0 18860 0 1 65280
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_234
timestamp 1694700623
transform 1 0 1104 0 -1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_235
timestamp 1694700623
transform -1 0 18860 0 -1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_236
timestamp 1694700623
transform 1 0 1104 0 1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_237
timestamp 1694700623
transform -1 0 18860 0 1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_238
timestamp 1694700623
transform 1 0 1104 0 -1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_239
timestamp 1694700623
transform -1 0 18860 0 -1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_240
timestamp 1694700623
transform 1 0 1104 0 1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_241
timestamp 1694700623
transform -1 0 18860 0 1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_242
timestamp 1694700623
transform 1 0 1104 0 -1 68544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_243
timestamp 1694700623
transform -1 0 18860 0 -1 68544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_244
timestamp 1694700623
transform 1 0 1104 0 1 68544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_245
timestamp 1694700623
transform -1 0 18860 0 1 68544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_246
timestamp 1694700623
transform 1 0 1104 0 -1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_247
timestamp 1694700623
transform -1 0 18860 0 -1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_248
timestamp 1694700623
transform 1 0 1104 0 1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_249
timestamp 1694700623
transform -1 0 18860 0 1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_250
timestamp 1694700623
transform 1 0 1104 0 -1 70720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_251
timestamp 1694700623
transform -1 0 18860 0 -1 70720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_252
timestamp 1694700623
transform 1 0 1104 0 1 70720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_253
timestamp 1694700623
transform -1 0 18860 0 1 70720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_254
timestamp 1694700623
transform 1 0 1104 0 -1 71808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_255
timestamp 1694700623
transform -1 0 18860 0 -1 71808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_256
timestamp 1694700623
transform 1 0 1104 0 1 71808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_257
timestamp 1694700623
transform -1 0 18860 0 1 71808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_258
timestamp 1694700623
transform 1 0 1104 0 -1 72896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_259
timestamp 1694700623
transform -1 0 18860 0 -1 72896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_260
timestamp 1694700623
transform 1 0 1104 0 1 72896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_261
timestamp 1694700623
transform -1 0 18860 0 1 72896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_262
timestamp 1694700623
transform 1 0 1104 0 -1 73984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_263
timestamp 1694700623
transform -1 0 18860 0 -1 73984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_264
timestamp 1694700623
transform 1 0 1104 0 1 73984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_265
timestamp 1694700623
transform -1 0 18860 0 1 73984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_266
timestamp 1694700623
transform 1 0 1104 0 -1 75072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_267
timestamp 1694700623
transform -1 0 18860 0 -1 75072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_268
timestamp 1694700623
transform 1 0 1104 0 1 75072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_269
timestamp 1694700623
transform -1 0 18860 0 1 75072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_270
timestamp 1694700623
transform 1 0 1104 0 -1 76160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_271
timestamp 1694700623
transform -1 0 18860 0 -1 76160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_272
timestamp 1694700623
transform 1 0 1104 0 1 76160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_273
timestamp 1694700623
transform -1 0 18860 0 1 76160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_274
timestamp 1694700623
transform 1 0 1104 0 -1 77248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_275
timestamp 1694700623
transform -1 0 18860 0 -1 77248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_276
timestamp 1694700623
transform 1 0 1104 0 1 77248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_277
timestamp 1694700623
transform -1 0 18860 0 1 77248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1694700623
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1694700623
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1694700623
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1694700623
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1694700623
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1694700623
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1694700623
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1694700623
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1694700623
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1694700623
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1694700623
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1694700623
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1694700623
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1694700623
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1694700623
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1694700623
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1694700623
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1694700623
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1694700623
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1694700623
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1694700623
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1694700623
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1694700623
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1694700623
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1694700623
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1694700623
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1694700623
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1694700623
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1694700623
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1694700623
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1694700623
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1694700623
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1694700623
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1694700623
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1694700623
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1694700623
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1694700623
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1694700623
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1694700623
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1694700623
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1694700623
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1694700623
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1694700623
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1694700623
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1694700623
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1694700623
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1694700623
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1694700623
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1694700623
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1694700623
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1694700623
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1694700623
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1694700623
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1694700623
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1694700623
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1694700623
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1694700623
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1694700623
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1694700623
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1694700623
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1694700623
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1694700623
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1694700623
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1694700623
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1694700623
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1694700623
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1694700623
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1694700623
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1694700623
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1694700623
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1694700623
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1694700623
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1694700623
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1694700623
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1694700623
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1694700623
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1694700623
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1694700623
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1694700623
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1694700623
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1694700623
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1694700623
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1694700623
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1694700623
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1694700623
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1694700623
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1694700623
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1694700623
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1694700623
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1694700623
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1694700623
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1694700623
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1694700623
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1694700623
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1694700623
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1694700623
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1694700623
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1694700623
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1694700623
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1694700623
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1694700623
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1694700623
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1694700623
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1694700623
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1694700623
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1694700623
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1694700623
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1694700623
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1694700623
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1694700623
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1694700623
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1694700623
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1694700623
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1694700623
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1694700623
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1694700623
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1694700623
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1694700623
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1694700623
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1694700623
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1694700623
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1694700623
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1694700623
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1694700623
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1694700623
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1694700623
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1694700623
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1694700623
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1694700623
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1694700623
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1694700623
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1694700623
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1694700623
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1694700623
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1694700623
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1694700623
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1694700623
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1694700623
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1694700623
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1694700623
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1694700623
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1694700623
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1694700623
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1694700623
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1694700623
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1694700623
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1694700623
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1694700623
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1694700623
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1694700623
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1694700623
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1694700623
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1694700623
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1694700623
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1694700623
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1694700623
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1694700623
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1694700623
transform 1 0 16560 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 1694700623
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 1694700623
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 1694700623
transform 1 0 13984 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 1694700623
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 1694700623
transform 1 0 11408 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 1694700623
transform 1 0 16560 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 1694700623
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 1694700623
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 1694700623
transform 1 0 13984 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 1694700623
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 1694700623
transform 1 0 11408 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 1694700623
transform 1 0 16560 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 1694700623
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 1694700623
transform 1 0 8832 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 1694700623
transform 1 0 13984 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 1694700623
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 1694700623
transform 1 0 11408 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 1694700623
transform 1 0 16560 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 1694700623
transform 1 0 3680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 1694700623
transform 1 0 8832 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 1694700623
transform 1 0 13984 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 1694700623
transform 1 0 6256 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 1694700623
transform 1 0 11408 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 1694700623
transform 1 0 16560 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 1694700623
transform 1 0 3680 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 1694700623
transform 1 0 8832 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 1694700623
transform 1 0 13984 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 1694700623
transform 1 0 6256 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 1694700623
transform 1 0 11408 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 1694700623
transform 1 0 16560 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 1694700623
transform 1 0 3680 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 1694700623
transform 1 0 8832 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_469
timestamp 1694700623
transform 1 0 13984 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_470
timestamp 1694700623
transform 1 0 6256 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_471
timestamp 1694700623
transform 1 0 11408 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_472
timestamp 1694700623
transform 1 0 16560 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_473
timestamp 1694700623
transform 1 0 3680 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_474
timestamp 1694700623
transform 1 0 8832 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_475
timestamp 1694700623
transform 1 0 13984 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_476
timestamp 1694700623
transform 1 0 6256 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_477
timestamp 1694700623
transform 1 0 11408 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_478
timestamp 1694700623
transform 1 0 16560 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_479
timestamp 1694700623
transform 1 0 3680 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_480
timestamp 1694700623
transform 1 0 8832 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_481
timestamp 1694700623
transform 1 0 13984 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_482
timestamp 1694700623
transform 1 0 6256 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_483
timestamp 1694700623
transform 1 0 11408 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_484
timestamp 1694700623
transform 1 0 16560 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_485
timestamp 1694700623
transform 1 0 3680 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_486
timestamp 1694700623
transform 1 0 8832 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_487
timestamp 1694700623
transform 1 0 13984 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_488
timestamp 1694700623
transform 1 0 6256 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_489
timestamp 1694700623
transform 1 0 11408 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_490
timestamp 1694700623
transform 1 0 16560 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_491
timestamp 1694700623
transform 1 0 3680 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_492
timestamp 1694700623
transform 1 0 8832 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_493
timestamp 1694700623
transform 1 0 13984 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_494
timestamp 1694700623
transform 1 0 6256 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_495
timestamp 1694700623
transform 1 0 11408 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_496
timestamp 1694700623
transform 1 0 16560 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_497
timestamp 1694700623
transform 1 0 3680 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_498
timestamp 1694700623
transform 1 0 8832 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_499
timestamp 1694700623
transform 1 0 13984 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_500
timestamp 1694700623
transform 1 0 6256 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_501
timestamp 1694700623
transform 1 0 11408 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_502
timestamp 1694700623
transform 1 0 16560 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_503
timestamp 1694700623
transform 1 0 3680 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_504
timestamp 1694700623
transform 1 0 8832 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_505
timestamp 1694700623
transform 1 0 13984 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_506
timestamp 1694700623
transform 1 0 6256 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_507
timestamp 1694700623
transform 1 0 11408 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_508
timestamp 1694700623
transform 1 0 16560 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_509
timestamp 1694700623
transform 1 0 3680 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_510
timestamp 1694700623
transform 1 0 8832 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_511
timestamp 1694700623
transform 1 0 13984 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_512
timestamp 1694700623
transform 1 0 6256 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_513
timestamp 1694700623
transform 1 0 11408 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_514
timestamp 1694700623
transform 1 0 16560 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_515
timestamp 1694700623
transform 1 0 3680 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_516
timestamp 1694700623
transform 1 0 8832 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_517
timestamp 1694700623
transform 1 0 13984 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_518
timestamp 1694700623
transform 1 0 6256 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_519
timestamp 1694700623
transform 1 0 11408 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_520
timestamp 1694700623
transform 1 0 16560 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_521
timestamp 1694700623
transform 1 0 3680 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_522
timestamp 1694700623
transform 1 0 8832 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_523
timestamp 1694700623
transform 1 0 13984 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_524
timestamp 1694700623
transform 1 0 6256 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_525
timestamp 1694700623
transform 1 0 11408 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_526
timestamp 1694700623
transform 1 0 16560 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_527
timestamp 1694700623
transform 1 0 3680 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_528
timestamp 1694700623
transform 1 0 8832 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_529
timestamp 1694700623
transform 1 0 13984 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_530
timestamp 1694700623
transform 1 0 6256 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_531
timestamp 1694700623
transform 1 0 11408 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_532
timestamp 1694700623
transform 1 0 16560 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_533
timestamp 1694700623
transform 1 0 3680 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_534
timestamp 1694700623
transform 1 0 8832 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_535
timestamp 1694700623
transform 1 0 13984 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_536
timestamp 1694700623
transform 1 0 6256 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_537
timestamp 1694700623
transform 1 0 11408 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_538
timestamp 1694700623
transform 1 0 16560 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_539
timestamp 1694700623
transform 1 0 3680 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_540
timestamp 1694700623
transform 1 0 8832 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_541
timestamp 1694700623
transform 1 0 13984 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_542
timestamp 1694700623
transform 1 0 6256 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_543
timestamp 1694700623
transform 1 0 11408 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_544
timestamp 1694700623
transform 1 0 16560 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_545
timestamp 1694700623
transform 1 0 3680 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_546
timestamp 1694700623
transform 1 0 8832 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_547
timestamp 1694700623
transform 1 0 13984 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_548
timestamp 1694700623
transform 1 0 6256 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_549
timestamp 1694700623
transform 1 0 11408 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_550
timestamp 1694700623
transform 1 0 16560 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_551
timestamp 1694700623
transform 1 0 3680 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_552
timestamp 1694700623
transform 1 0 8832 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_553
timestamp 1694700623
transform 1 0 13984 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_554
timestamp 1694700623
transform 1 0 6256 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_555
timestamp 1694700623
transform 1 0 11408 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_556
timestamp 1694700623
transform 1 0 16560 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_557
timestamp 1694700623
transform 1 0 3680 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_558
timestamp 1694700623
transform 1 0 8832 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_559
timestamp 1694700623
transform 1 0 13984 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_560
timestamp 1694700623
transform 1 0 6256 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_561
timestamp 1694700623
transform 1 0 11408 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_562
timestamp 1694700623
transform 1 0 16560 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_563
timestamp 1694700623
transform 1 0 3680 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_564
timestamp 1694700623
transform 1 0 8832 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_565
timestamp 1694700623
transform 1 0 13984 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_566
timestamp 1694700623
transform 1 0 6256 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_567
timestamp 1694700623
transform 1 0 11408 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_568
timestamp 1694700623
transform 1 0 16560 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_569
timestamp 1694700623
transform 1 0 3680 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_570
timestamp 1694700623
transform 1 0 8832 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_571
timestamp 1694700623
transform 1 0 13984 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_572
timestamp 1694700623
transform 1 0 6256 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_573
timestamp 1694700623
transform 1 0 11408 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_574
timestamp 1694700623
transform 1 0 16560 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_575
timestamp 1694700623
transform 1 0 3680 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_576
timestamp 1694700623
transform 1 0 8832 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_577
timestamp 1694700623
transform 1 0 13984 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_578
timestamp 1694700623
transform 1 0 6256 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_579
timestamp 1694700623
transform 1 0 11408 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_580
timestamp 1694700623
transform 1 0 16560 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_581
timestamp 1694700623
transform 1 0 3680 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_582
timestamp 1694700623
transform 1 0 8832 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_583
timestamp 1694700623
transform 1 0 13984 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_584
timestamp 1694700623
transform 1 0 6256 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_585
timestamp 1694700623
transform 1 0 11408 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_586
timestamp 1694700623
transform 1 0 16560 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_587
timestamp 1694700623
transform 1 0 3680 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_588
timestamp 1694700623
transform 1 0 8832 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_589
timestamp 1694700623
transform 1 0 13984 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_590
timestamp 1694700623
transform 1 0 6256 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_591
timestamp 1694700623
transform 1 0 11408 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_592
timestamp 1694700623
transform 1 0 16560 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_593
timestamp 1694700623
transform 1 0 3680 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_594
timestamp 1694700623
transform 1 0 8832 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_595
timestamp 1694700623
transform 1 0 13984 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_596
timestamp 1694700623
transform 1 0 6256 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_597
timestamp 1694700623
transform 1 0 11408 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_598
timestamp 1694700623
transform 1 0 16560 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_599
timestamp 1694700623
transform 1 0 3680 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_600
timestamp 1694700623
transform 1 0 8832 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_601
timestamp 1694700623
transform 1 0 13984 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_602
timestamp 1694700623
transform 1 0 6256 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_603
timestamp 1694700623
transform 1 0 11408 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_604
timestamp 1694700623
transform 1 0 16560 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_605
timestamp 1694700623
transform 1 0 3680 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_606
timestamp 1694700623
transform 1 0 8832 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_607
timestamp 1694700623
transform 1 0 13984 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_608
timestamp 1694700623
transform 1 0 6256 0 -1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_609
timestamp 1694700623
transform 1 0 11408 0 -1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_610
timestamp 1694700623
transform 1 0 16560 0 -1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_611
timestamp 1694700623
transform 1 0 3680 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_612
timestamp 1694700623
transform 1 0 8832 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_613
timestamp 1694700623
transform 1 0 13984 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_614
timestamp 1694700623
transform 1 0 6256 0 -1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_615
timestamp 1694700623
transform 1 0 11408 0 -1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_616
timestamp 1694700623
transform 1 0 16560 0 -1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_617
timestamp 1694700623
transform 1 0 3680 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_618
timestamp 1694700623
transform 1 0 8832 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_619
timestamp 1694700623
transform 1 0 13984 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_620
timestamp 1694700623
transform 1 0 6256 0 -1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_621
timestamp 1694700623
transform 1 0 11408 0 -1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_622
timestamp 1694700623
transform 1 0 16560 0 -1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_623
timestamp 1694700623
transform 1 0 3680 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_624
timestamp 1694700623
transform 1 0 8832 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_625
timestamp 1694700623
transform 1 0 13984 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_626
timestamp 1694700623
transform 1 0 6256 0 -1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_627
timestamp 1694700623
transform 1 0 11408 0 -1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_628
timestamp 1694700623
transform 1 0 16560 0 -1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_629
timestamp 1694700623
transform 1 0 3680 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_630
timestamp 1694700623
transform 1 0 8832 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_631
timestamp 1694700623
transform 1 0 13984 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_632
timestamp 1694700623
transform 1 0 6256 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_633
timestamp 1694700623
transform 1 0 11408 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_634
timestamp 1694700623
transform 1 0 16560 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_635
timestamp 1694700623
transform 1 0 3680 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_636
timestamp 1694700623
transform 1 0 8832 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_637
timestamp 1694700623
transform 1 0 13984 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_638
timestamp 1694700623
transform 1 0 6256 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_639
timestamp 1694700623
transform 1 0 11408 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_640
timestamp 1694700623
transform 1 0 16560 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_641
timestamp 1694700623
transform 1 0 3680 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_642
timestamp 1694700623
transform 1 0 8832 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_643
timestamp 1694700623
transform 1 0 13984 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_644
timestamp 1694700623
transform 1 0 6256 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_645
timestamp 1694700623
transform 1 0 11408 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_646
timestamp 1694700623
transform 1 0 16560 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_647
timestamp 1694700623
transform 1 0 3680 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_648
timestamp 1694700623
transform 1 0 8832 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_649
timestamp 1694700623
transform 1 0 13984 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_650
timestamp 1694700623
transform 1 0 6256 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_651
timestamp 1694700623
transform 1 0 11408 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_652
timestamp 1694700623
transform 1 0 16560 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_653
timestamp 1694700623
transform 1 0 3680 0 1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_654
timestamp 1694700623
transform 1 0 8832 0 1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_655
timestamp 1694700623
transform 1 0 13984 0 1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_656
timestamp 1694700623
transform 1 0 6256 0 -1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_657
timestamp 1694700623
transform 1 0 11408 0 -1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_658
timestamp 1694700623
transform 1 0 16560 0 -1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_659
timestamp 1694700623
transform 1 0 3680 0 1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_660
timestamp 1694700623
transform 1 0 8832 0 1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_661
timestamp 1694700623
transform 1 0 13984 0 1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_662
timestamp 1694700623
transform 1 0 6256 0 -1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_663
timestamp 1694700623
transform 1 0 11408 0 -1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_664
timestamp 1694700623
transform 1 0 16560 0 -1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_665
timestamp 1694700623
transform 1 0 3680 0 1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_666
timestamp 1694700623
transform 1 0 8832 0 1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_667
timestamp 1694700623
transform 1 0 13984 0 1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_668
timestamp 1694700623
transform 1 0 6256 0 -1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_669
timestamp 1694700623
transform 1 0 11408 0 -1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_670
timestamp 1694700623
transform 1 0 16560 0 -1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_671
timestamp 1694700623
transform 1 0 3680 0 1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_672
timestamp 1694700623
transform 1 0 8832 0 1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_673
timestamp 1694700623
transform 1 0 13984 0 1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_674
timestamp 1694700623
transform 1 0 6256 0 -1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_675
timestamp 1694700623
transform 1 0 11408 0 -1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_676
timestamp 1694700623
transform 1 0 16560 0 -1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_677
timestamp 1694700623
transform 1 0 3680 0 1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_678
timestamp 1694700623
transform 1 0 8832 0 1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_679
timestamp 1694700623
transform 1 0 13984 0 1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_680
timestamp 1694700623
transform 1 0 6256 0 -1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_681
timestamp 1694700623
transform 1 0 11408 0 -1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_682
timestamp 1694700623
transform 1 0 16560 0 -1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_683
timestamp 1694700623
transform 1 0 3680 0 1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_684
timestamp 1694700623
transform 1 0 8832 0 1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_685
timestamp 1694700623
transform 1 0 13984 0 1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_686
timestamp 1694700623
transform 1 0 6256 0 -1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_687
timestamp 1694700623
transform 1 0 11408 0 -1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_688
timestamp 1694700623
transform 1 0 16560 0 -1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_689
timestamp 1694700623
transform 1 0 3680 0 1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_690
timestamp 1694700623
transform 1 0 8832 0 1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_691
timestamp 1694700623
transform 1 0 13984 0 1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_692
timestamp 1694700623
transform 1 0 6256 0 -1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_693
timestamp 1694700623
transform 1 0 11408 0 -1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_694
timestamp 1694700623
transform 1 0 16560 0 -1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_695
timestamp 1694700623
transform 1 0 3680 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_696
timestamp 1694700623
transform 1 0 6256 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_697
timestamp 1694700623
transform 1 0 8832 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_698
timestamp 1694700623
transform 1 0 11408 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_699
timestamp 1694700623
transform 1 0 13984 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_700
timestamp 1694700623
transform 1 0 16560 0 1 77248
box -38 -48 130 592
<< labels >>
flabel metal4 s 2604 2128 2924 77840 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 7604 2128 7924 77840 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 12604 2128 12924 77840 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 17604 2128 17924 77840 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal5 s 1056 3676 18908 3996 0 FreeSans 2560 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal5 s 1056 8676 18908 8996 0 FreeSans 2560 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal5 s 1056 13676 18908 13996 0 FreeSans 2560 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal5 s 1056 18676 18908 18996 0 FreeSans 2560 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal5 s 1056 23676 18908 23996 0 FreeSans 2560 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal5 s 1056 28676 18908 28996 0 FreeSans 2560 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal5 s 1056 33676 18908 33996 0 FreeSans 2560 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal5 s 1056 38676 18908 38996 0 FreeSans 2560 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal5 s 1056 43676 18908 43996 0 FreeSans 2560 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal5 s 1056 48676 18908 48996 0 FreeSans 2560 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal5 s 1056 53676 18908 53996 0 FreeSans 2560 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal5 s 1056 58676 18908 58996 0 FreeSans 2560 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal5 s 1056 63676 18908 63996 0 FreeSans 2560 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal5 s 1056 68676 18908 68996 0 FreeSans 2560 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal5 s 1056 73676 18908 73996 0 FreeSans 2560 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 1944 2128 2264 77840 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 6944 2128 7264 77840 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 11944 2128 12264 77840 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 16944 2128 17264 77840 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal5 s 1056 3016 18908 3336 0 FreeSans 2560 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal5 s 1056 8016 18908 8336 0 FreeSans 2560 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal5 s 1056 13016 18908 13336 0 FreeSans 2560 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal5 s 1056 18016 18908 18336 0 FreeSans 2560 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal5 s 1056 23016 18908 23336 0 FreeSans 2560 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal5 s 1056 28016 18908 28336 0 FreeSans 2560 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal5 s 1056 33016 18908 33336 0 FreeSans 2560 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal5 s 1056 38016 18908 38336 0 FreeSans 2560 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal5 s 1056 43016 18908 43336 0 FreeSans 2560 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal5 s 1056 48016 18908 48336 0 FreeSans 2560 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal5 s 1056 53016 18908 53336 0 FreeSans 2560 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal5 s 1056 58016 18908 58336 0 FreeSans 2560 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal5 s 1056 63016 18908 63336 0 FreeSans 2560 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal5 s 1056 68016 18908 68336 0 FreeSans 2560 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal5 s 1056 73016 18908 73336 0 FreeSans 2560 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal2 s 2042 0 2098 800 0 FreeSans 224 90 0 0 clk
port 2 nsew signal input
flabel metal3 s 19200 76984 20000 77104 0 FreeSans 480 0 0 0 data_reg[0]
port 3 nsew signal tristate
flabel metal3 s 19200 57944 20000 58064 0 FreeSans 480 0 0 0 data_reg[10]
port 4 nsew signal tristate
flabel metal3 s 19200 56040 20000 56160 0 FreeSans 480 0 0 0 data_reg[11]
port 5 nsew signal tristate
flabel metal3 s 19200 54136 20000 54256 0 FreeSans 480 0 0 0 data_reg[12]
port 6 nsew signal tristate
flabel metal3 s 19200 52232 20000 52352 0 FreeSans 480 0 0 0 data_reg[13]
port 7 nsew signal tristate
flabel metal3 s 19200 50328 20000 50448 0 FreeSans 480 0 0 0 data_reg[14]
port 8 nsew signal tristate
flabel metal3 s 19200 48424 20000 48544 0 FreeSans 480 0 0 0 data_reg[15]
port 9 nsew signal tristate
flabel metal3 s 19200 46520 20000 46640 0 FreeSans 480 0 0 0 data_reg[16]
port 10 nsew signal tristate
flabel metal3 s 19200 44616 20000 44736 0 FreeSans 480 0 0 0 data_reg[17]
port 11 nsew signal tristate
flabel metal3 s 19200 42712 20000 42832 0 FreeSans 480 0 0 0 data_reg[18]
port 12 nsew signal tristate
flabel metal3 s 19200 40808 20000 40928 0 FreeSans 480 0 0 0 data_reg[19]
port 13 nsew signal tristate
flabel metal3 s 19200 75080 20000 75200 0 FreeSans 480 0 0 0 data_reg[1]
port 14 nsew signal tristate
flabel metal3 s 19200 38904 20000 39024 0 FreeSans 480 0 0 0 data_reg[20]
port 15 nsew signal tristate
flabel metal3 s 19200 37000 20000 37120 0 FreeSans 480 0 0 0 data_reg[21]
port 16 nsew signal tristate
flabel metal3 s 19200 35096 20000 35216 0 FreeSans 480 0 0 0 data_reg[22]
port 17 nsew signal tristate
flabel metal3 s 19200 33192 20000 33312 0 FreeSans 480 0 0 0 data_reg[23]
port 18 nsew signal tristate
flabel metal3 s 19200 31288 20000 31408 0 FreeSans 480 0 0 0 data_reg[24]
port 19 nsew signal tristate
flabel metal3 s 19200 29384 20000 29504 0 FreeSans 480 0 0 0 data_reg[25]
port 20 nsew signal tristate
flabel metal3 s 19200 27480 20000 27600 0 FreeSans 480 0 0 0 data_reg[26]
port 21 nsew signal tristate
flabel metal3 s 19200 25576 20000 25696 0 FreeSans 480 0 0 0 data_reg[27]
port 22 nsew signal tristate
flabel metal3 s 19200 23672 20000 23792 0 FreeSans 480 0 0 0 data_reg[28]
port 23 nsew signal tristate
flabel metal3 s 19200 21768 20000 21888 0 FreeSans 480 0 0 0 data_reg[29]
port 24 nsew signal tristate
flabel metal3 s 19200 73176 20000 73296 0 FreeSans 480 0 0 0 data_reg[2]
port 25 nsew signal tristate
flabel metal3 s 19200 19864 20000 19984 0 FreeSans 480 0 0 0 data_reg[30]
port 26 nsew signal tristate
flabel metal3 s 19200 17960 20000 18080 0 FreeSans 480 0 0 0 data_reg[31]
port 27 nsew signal tristate
flabel metal3 s 19200 16056 20000 16176 0 FreeSans 480 0 0 0 data_reg[32]
port 28 nsew signal tristate
flabel metal3 s 19200 14152 20000 14272 0 FreeSans 480 0 0 0 data_reg[33]
port 29 nsew signal tristate
flabel metal3 s 19200 12248 20000 12368 0 FreeSans 480 0 0 0 data_reg[34]
port 30 nsew signal tristate
flabel metal3 s 19200 10344 20000 10464 0 FreeSans 480 0 0 0 data_reg[35]
port 31 nsew signal tristate
flabel metal3 s 19200 8440 20000 8560 0 FreeSans 480 0 0 0 data_reg[36]
port 32 nsew signal tristate
flabel metal3 s 19200 6536 20000 6656 0 FreeSans 480 0 0 0 data_reg[37]
port 33 nsew signal tristate
flabel metal3 s 19200 4632 20000 4752 0 FreeSans 480 0 0 0 data_reg[38]
port 34 nsew signal tristate
flabel metal3 s 19200 2728 20000 2848 0 FreeSans 480 0 0 0 data_reg[39]
port 35 nsew signal tristate
flabel metal3 s 19200 71272 20000 71392 0 FreeSans 480 0 0 0 data_reg[3]
port 36 nsew signal tristate
flabel metal3 s 19200 69368 20000 69488 0 FreeSans 480 0 0 0 data_reg[4]
port 37 nsew signal tristate
flabel metal3 s 19200 67464 20000 67584 0 FreeSans 480 0 0 0 data_reg[5]
port 38 nsew signal tristate
flabel metal3 s 19200 65560 20000 65680 0 FreeSans 480 0 0 0 data_reg[6]
port 39 nsew signal tristate
flabel metal3 s 19200 63656 20000 63776 0 FreeSans 480 0 0 0 data_reg[7]
port 40 nsew signal tristate
flabel metal3 s 19200 61752 20000 61872 0 FreeSans 480 0 0 0 data_reg[8]
port 41 nsew signal tristate
flabel metal3 s 19200 59848 20000 59968 0 FreeSans 480 0 0 0 data_reg[9]
port 42 nsew signal tristate
flabel metal2 s 17866 0 17922 800 0 FreeSans 224 90 0 0 load
port 43 nsew signal input
flabel metal2 s 5998 0 6054 800 0 FreeSans 224 90 0 0 serial_in
port 44 nsew signal input
flabel metal2 s 9954 0 10010 800 0 FreeSans 224 90 0 0 serial_out
port 45 nsew signal tristate
flabel metal2 s 13910 0 13966 800 0 FreeSans 224 90 0 0 shift_enable
port 46 nsew signal input
rlabel metal1 9982 77248 9982 77248 0 VGND
rlabel metal1 9982 77792 9982 77792 0 VPWR
rlabel metal1 4227 3094 4227 3094 0 _000_
rlabel metal1 8362 40018 8362 40018 0 _001_
rlabel metal1 13554 14314 13554 14314 0 _002_
rlabel metal1 5014 9928 5014 9928 0 _003_
rlabel metal1 2484 50694 2484 50694 0 _004_
rlabel metal1 11714 64362 11714 64362 0 _005_
rlabel metal1 14444 50150 14444 50150 0 _006_
rlabel metal1 5796 62798 5796 62798 0 _007_
rlabel metal1 5244 59398 5244 59398 0 _008_
rlabel via1 11081 12206 11081 12206 0 _009_
rlabel metal2 15226 73304 15226 73304 0 _010_
rlabel metal1 13386 26928 13386 26928 0 _011_
rlabel metal1 7544 14586 7544 14586 0 _012_
rlabel metal1 3910 55284 3910 55284 0 _013_
rlabel metal1 15083 52462 15083 52462 0 _014_
rlabel metal2 1150 42670 1150 42670 0 _015_
rlabel metal1 8546 34578 8546 34578 0 _016_
rlabel metal1 14352 62798 14352 62798 0 _017_
rlabel metal2 4370 41344 4370 41344 0 _018_
rlabel metal1 11684 57222 11684 57222 0 _019_
rlabel metal2 8142 4250 8142 4250 0 _020_
rlabel metal1 13248 58990 13248 58990 0 _021_
rlabel metal1 2054 37162 2054 37162 0 _022_
rlabel via1 15129 74834 15129 74834 0 _023_
rlabel metal1 5152 69734 5152 69734 0 _024_
rlabel metal2 6624 64860 6624 64860 0 _025_
rlabel metal1 17940 74630 17940 74630 0 _026_
rlabel metal1 11760 31382 11760 31382 0 _027_
rlabel via1 14209 18326 14209 18326 0 _028_
rlabel metal2 16422 47090 16422 47090 0 _029_
rlabel metal1 17112 77350 17112 77350 0 _030_
rlabel metal1 15456 63478 15456 63478 0 _031_
rlabel metal1 16233 65110 16233 65110 0 _032_
rlabel metal1 8096 9146 8096 9146 0 _033_
rlabel metal2 13524 44948 13524 44948 0 _034_
rlabel metal1 7114 34986 7114 34986 0 _035_
rlabel metal1 4784 52938 4784 52938 0 _036_
rlabel metal1 14996 48858 14996 48858 0 _037_
rlabel via1 15773 70890 15773 70890 0 _038_
rlabel metal1 2162 8058 2162 8058 0 _039_
rlabel metal1 14260 21862 14260 21862 0 _040_
rlabel metal1 18400 64906 18400 64906 0 _041_
rlabel via1 3077 57426 3077 57426 0 _042_
rlabel via2 13846 7259 13846 7259 0 _043_
rlabel via1 14577 60010 14577 60010 0 _044_
rlabel metal1 16003 32810 16003 32810 0 _045_
rlabel metal1 16866 15402 16866 15402 0 _046_
rlabel metal1 5791 5678 5791 5678 0 _047_
rlabel metal1 9062 52462 9062 52462 0 _048_
rlabel via1 16233 61098 16233 61098 0 _049_
rlabel metal1 8326 55862 8326 55862 0 _050_
rlabel metal1 3956 4046 3956 4046 0 _051_
rlabel metal1 1886 56202 1886 56202 0 _052_
rlabel via2 16238 5219 16238 5219 0 _053_
rlabel metal1 1410 55658 1410 55658 0 _054_
rlabel metal1 16882 72250 16882 72250 0 _055_
rlabel metal2 13294 34748 13294 34748 0 _056_
rlabel metal1 12880 56270 12880 56270 0 _057_
rlabel metal1 11454 31994 11454 31994 0 _058_
rlabel metal1 12795 47702 12795 47702 0 _059_
rlabel metal1 3848 28118 3848 28118 0 _060_
rlabel metal1 10672 51238 10672 51238 0 _061_
rlabel metal1 17245 12886 17245 12886 0 _062_
rlabel metal1 7038 21862 7038 21862 0 _063_
rlabel metal2 12466 35513 12466 35513 0 _064_
rlabel metal1 6302 51238 6302 51238 0 _065_
rlabel via1 12553 46614 12553 46614 0 _066_
rlabel metal1 12404 35734 12404 35734 0 _067_
rlabel metal2 4232 57324 4232 57324 0 _068_
rlabel metal1 13662 42806 13662 42806 0 _069_
rlabel metal1 8724 69462 8724 69462 0 _070_
rlabel metal1 1840 42738 1840 42738 0 _071_
rlabel via2 6670 9571 6670 9571 0 _072_
rlabel metal1 2576 8398 2576 8398 0 _073_
rlabel metal2 17526 75820 17526 75820 0 _074_
rlabel metal1 6596 12138 6596 12138 0 _075_
rlabel metal1 6670 60656 6670 60656 0 _076_
rlabel metal1 6164 55250 6164 55250 0 _077_
rlabel metal1 13110 8466 13110 8466 0 _078_
rlabel metal2 8234 5202 8234 5202 0 _079_
rlabel metal1 18170 67218 18170 67218 0 _080_
rlabel metal1 7268 28594 7268 28594 0 _081_
rlabel metal1 6578 74834 6578 74834 0 _082_
rlabel metal1 12282 34680 12282 34680 0 _083_
rlabel metal1 5198 10064 5198 10064 0 _084_
rlabel metal3 1633 55692 1633 55692 0 _085_
rlabel metal1 17066 42534 17066 42534 0 _086_
rlabel metal2 5106 62730 5106 62730 0 _087_
rlabel metal3 13041 55828 13041 55828 0 _088_
rlabel metal1 9108 8874 9108 8874 0 _089_
rlabel metal1 11822 21862 11822 21862 0 _090_
rlabel metal2 4646 63036 4646 63036 0 _091_
rlabel metal1 6440 74970 6440 74970 0 _092_
rlabel metal2 8050 60384 8050 60384 0 _093_
rlabel metal3 4025 65212 4025 65212 0 _094_
rlabel metal1 9798 6834 9798 6834 0 _095_
rlabel metal2 14030 35054 14030 35054 0 _096_
rlabel metal3 9039 52564 9039 52564 0 _097_
rlabel metal2 1794 28390 1794 28390 0 _098_
rlabel metal1 13800 17782 13800 17782 0 _099_
rlabel via3 4301 62220 4301 62220 0 _100_
rlabel metal2 16882 56406 16882 56406 0 _101_
rlabel metal1 17894 20366 17894 20366 0 _102_
rlabel metal1 7544 5202 7544 5202 0 _103_
rlabel metal1 5704 58990 5704 58990 0 _104_
rlabel via2 13754 58837 13754 58837 0 _105_
rlabel metal1 15410 36550 15410 36550 0 _106_
rlabel metal2 4002 69666 4002 69666 0 _107_
rlabel metal1 8234 20230 8234 20230 0 _108_
rlabel metal2 16744 58412 16744 58412 0 _109_
rlabel metal2 9706 63546 9706 63546 0 _110_
rlabel metal1 2806 53006 2806 53006 0 _111_
rlabel metal3 9361 19924 9361 19924 0 _112_
rlabel metal1 15180 44846 15180 44846 0 _113_
rlabel metal3 1679 40596 1679 40596 0 _114_
rlabel metal1 14122 61914 14122 61914 0 _115_
rlabel metal1 18124 27438 18124 27438 0 _116_
rlabel metal2 17526 65501 17526 65501 0 _117_
rlabel metal1 7498 21522 7498 21522 0 _118_
rlabel metal1 13018 42806 13018 42806 0 _119_
rlabel metal1 8878 53074 8878 53074 0 _120_
rlabel metal3 7659 6732 7659 6732 0 _121_
rlabel metal1 3220 69802 3220 69802 0 _122_
rlabel metal3 1909 69292 1909 69292 0 _123_
rlabel metal1 3588 7854 3588 7854 0 _124_
rlabel metal1 14904 21998 14904 21998 0 _125_
rlabel metal1 18768 65042 18768 65042 0 _126_
rlabel metal1 15686 16558 15686 16558 0 _127_
rlabel via3 14237 8228 14237 8228 0 _128_
rlabel metal1 18492 51986 18492 51986 0 _129_
rlabel metal1 15410 20298 15410 20298 0 _130_
rlabel metal2 7038 9707 7038 9707 0 _131_
rlabel metal2 9522 18802 9522 18802 0 _132_
rlabel metal1 1886 42670 1886 42670 0 _133_
rlabel metal1 8142 65178 8142 65178 0 _134_
rlabel metal1 2622 56950 2622 56950 0 _135_
rlabel via2 11270 76245 11270 76245 0 _136_
rlabel metal1 1794 20298 1794 20298 0 _137_
rlabel metal2 2346 18571 2346 18571 0 _138_
rlabel via1 1697 42534 1697 42534 0 _139_
rlabel metal2 1564 40732 1564 40732 0 _140_
rlabel metal2 16882 73236 16882 73236 0 _141_
rlabel metal2 690 29002 690 29002 0 _142_
rlabel metal3 13455 55692 13455 55692 0 _143_
rlabel metal1 14950 20842 14950 20842 0 _144_
rlabel metal1 15364 38318 15364 38318 0 _145_
rlabel metal1 9844 60214 9844 60214 0 _146_
rlabel metal1 7544 29274 7544 29274 0 _147_
rlabel metal1 6210 25330 6210 25330 0 _148_
rlabel metal1 17204 38930 17204 38930 0 _149_
rlabel via2 15318 11203 15318 11203 0 _150_
rlabel metal1 7452 59942 7452 59942 0 _151_
rlabel metal1 1932 22066 1932 22066 0 _152_
rlabel metal3 11339 54060 11339 54060 0 _153_
rlabel metal1 8832 54026 8832 54026 0 _154_
rlabel metal1 6486 40154 6486 40154 0 _155_
rlabel metal1 15962 24650 15962 24650 0 _156_
rlabel metal2 17480 42636 17480 42636 0 _157_
rlabel metal1 12374 13498 12374 13498 0 _158_
rlabel metal1 4761 64430 4761 64430 0 _159_
rlabel metal2 7314 74596 7314 74596 0 _160_
rlabel metal2 15594 60452 15594 60452 0 _161_
rlabel metal1 17296 76942 17296 76942 0 _162_
rlabel metal1 6808 32198 6808 32198 0 _163_
rlabel via2 2622 10693 2622 10693 0 _164_
rlabel metal2 15410 36312 15410 36312 0 _165_
rlabel metal2 14398 9418 14398 9418 0 _166_
rlabel metal1 16606 31824 16606 31824 0 _167_
rlabel metal1 2438 2958 2438 2958 0 clk
rlabel metal2 18262 77197 18262 77197 0 data_reg[0]
rlabel metal2 18262 58157 18262 58157 0 data_reg[10]
rlabel via2 18262 56117 18262 56117 0 data_reg[11]
rlabel metal2 18262 54349 18262 54349 0 data_reg[12]
rlabel metal2 18262 52445 18262 52445 0 data_reg[13]
rlabel metal2 18262 50541 18262 50541 0 data_reg[14]
rlabel via2 18262 48501 18262 48501 0 data_reg[15]
rlabel metal2 18262 46733 18262 46733 0 data_reg[16]
rlabel via2 18262 44693 18262 44693 0 data_reg[17]
rlabel metal2 18262 42925 18262 42925 0 data_reg[18]
rlabel via2 18262 40885 18262 40885 0 data_reg[19]
rlabel via2 18262 75157 18262 75157 0 data_reg[1]
rlabel metal2 18262 39117 18262 39117 0 data_reg[20]
rlabel via2 18262 37077 18262 37077 0 data_reg[21]
rlabel metal2 18262 35309 18262 35309 0 data_reg[22]
rlabel via2 18262 33269 18262 33269 0 data_reg[23]
rlabel metal2 18262 31501 18262 31501 0 data_reg[24]
rlabel via2 18262 29461 18262 29461 0 data_reg[25]
rlabel metal1 18078 27846 18078 27846 0 data_reg[26]
rlabel via2 18262 25653 18262 25653 0 data_reg[27]
rlabel metal2 18262 23885 18262 23885 0 data_reg[28]
rlabel via2 18262 21845 18262 21845 0 data_reg[29]
rlabel metal2 18262 73389 18262 73389 0 data_reg[2]
rlabel via2 18262 19941 18262 19941 0 data_reg[30]
rlabel via2 18262 18037 18262 18037 0 data_reg[31]
rlabel metal2 18262 16167 18262 16167 0 data_reg[32]
rlabel via2 18262 14229 18262 14229 0 data_reg[33]
rlabel via2 18262 12325 18262 12325 0 data_reg[34]
rlabel via2 18262 10421 18262 10421 0 data_reg[35]
rlabel metal2 18262 8653 18262 8653 0 data_reg[36]
rlabel via2 18262 6613 18262 6613 0 data_reg[37]
rlabel metal2 18262 4845 18262 4845 0 data_reg[38]
rlabel via2 18262 2805 18262 2805 0 data_reg[39]
rlabel via2 18262 71349 18262 71349 0 data_reg[3]
rlabel metal2 18262 69581 18262 69581 0 data_reg[4]
rlabel metal2 18262 67677 18262 67677 0 data_reg[5]
rlabel via2 18262 65637 18262 65637 0 data_reg[6]
rlabel via2 18262 63733 18262 63733 0 data_reg[7]
rlabel metal2 18262 61965 18262 61965 0 data_reg[8]
rlabel via2 18262 59925 18262 59925 0 data_reg[9]
rlabel metal2 17894 1367 17894 1367 0 load
rlabel metal1 14444 20910 14444 20910 0 net1
rlabel metal1 6578 60010 6578 60010 0 net10
rlabel metal1 16100 60214 16100 60214 0 net11
rlabel metal1 18814 44846 18814 44846 0 net12
rlabel metal1 18308 43282 18308 43282 0 net13
rlabel metal1 18170 15368 18170 15368 0 net14
rlabel metal1 17319 75310 17319 75310 0 net15
rlabel metal1 8510 65042 8510 65042 0 net16
rlabel metal1 2346 56814 2346 56814 0 net17
rlabel metal1 13018 35632 13018 35632 0 net18
rlabel metal1 2162 20332 2162 20332 0 net19
rlabel metal1 5796 2278 5796 2278 0 net2
rlabel metal2 18078 33932 18078 33932 0 net20
rlabel metal1 2438 42738 2438 42738 0 net21
rlabel metal1 6670 55590 6670 55590 0 net22
rlabel metal2 12466 72896 12466 72896 0 net23
rlabel metal1 14950 34714 14950 34714 0 net24
rlabel metal1 18354 32198 18354 32198 0 net25
rlabel metal2 1978 53278 1978 53278 0 net26
rlabel metal1 12052 19822 12052 19822 0 net27
rlabel metal1 18676 18258 18676 18258 0 net28
rlabel metal1 14536 16082 14536 16082 0 net29
rlabel metal1 13846 44778 13846 44778 0 net3
rlabel metal1 18814 14382 18814 14382 0 net30
rlabel metal2 18078 12580 18078 12580 0 net31
rlabel metal1 9545 11118 9545 11118 0 net32
rlabel metal1 8050 60010 8050 60010 0 net33
rlabel metal1 5566 11798 5566 11798 0 net34
rlabel metal1 17802 5202 17802 5202 0 net35
rlabel metal2 10626 53295 10626 53295 0 net36
rlabel metal1 13892 61846 13892 61846 0 net37
rlabel metal1 1978 44472 1978 44472 0 net38
rlabel metal1 17526 42534 17526 42534 0 net39
rlabel metal1 18630 44370 18630 44370 0 net4
rlabel metal1 10534 61370 10534 61370 0 net40
rlabel metal1 18308 63954 18308 63954 0 net41
rlabel metal1 18354 62254 18354 62254 0 net42
rlabel metal1 18676 60078 18676 60078 0 net43
rlabel metal1 9476 2414 9476 2414 0 net44
rlabel metal1 17388 58514 17388 58514 0 net5
rlabel metal1 8280 57562 8280 57562 0 net6
rlabel metal2 18262 44268 18262 44268 0 net7
rlabel metal1 18032 52462 18032 52462 0 net8
rlabel metal2 4186 57120 4186 57120 0 net9
rlabel metal2 6026 1588 6026 1588 0 serial_in
rlabel metal2 9982 1520 9982 1520 0 serial_out
rlabel metal2 13938 1554 13938 1554 0 shift_enable
rlabel metal2 2484 50388 2484 50388 0 shift_reg\[10\]
rlabel metal2 6900 31892 6900 31892 0 shift_reg\[11\]
rlabel metal1 6624 3162 6624 3162 0 shift_reg\[12\]
rlabel metal1 9522 20978 9522 20978 0 shift_reg\[13\]
rlabel metal1 15042 14586 15042 14586 0 shift_reg\[14\]
rlabel metal1 15088 21114 15088 21114 0 shift_reg\[15\]
rlabel metal1 16928 15062 16928 15062 0 shift_reg\[16\]
rlabel metal1 14444 63546 14444 63546 0 shift_reg\[17\]
rlabel metal2 16836 58276 16836 58276 0 shift_reg\[18\]
rlabel metal1 11500 62390 11500 62390 0 shift_reg\[19\]
rlabel metal2 14214 57766 14214 57766 0 shift_reg\[1\]
rlabel metal1 5773 59738 5773 59738 0 shift_reg\[20\]
rlabel metal2 2300 44404 2300 44404 0 shift_reg\[21\]
rlabel metal1 9844 39338 9844 39338 0 shift_reg\[22\]
rlabel metal1 5290 20502 5290 20502 0 shift_reg\[23\]
rlabel metal1 9016 60758 9016 60758 0 shift_reg\[24\]
rlabel metal1 4094 65382 4094 65382 0 shift_reg\[25\]
rlabel via2 9706 6715 9706 6715 0 shift_reg\[26\]
rlabel metal1 6302 36142 6302 36142 0 shift_reg\[27\]
rlabel metal1 10074 53142 10074 53142 0 shift_reg\[28\]
rlabel metal3 10465 67660 10465 67660 0 shift_reg\[29\]
rlabel metal1 11270 54298 11270 54298 0 shift_reg\[2\]
rlabel metal1 13294 17714 13294 17714 0 shift_reg\[30\]
rlabel metal1 17066 55250 17066 55250 0 shift_reg\[31\]
rlabel metal1 16974 55318 16974 55318 0 shift_reg\[32\]
rlabel metal1 9200 7922 9200 7922 0 shift_reg\[33\]
rlabel metal2 15226 50864 15226 50864 0 shift_reg\[34\]
rlabel metal1 15410 58922 15410 58922 0 shift_reg\[35\]
rlabel metal1 15042 59942 15042 59942 0 shift_reg\[36\]
rlabel metal2 16422 60095 16422 60095 0 shift_reg\[37\]
rlabel metal2 16882 20162 16882 20162 0 shift_reg\[38\]
rlabel metal1 11776 63954 11776 63954 0 shift_reg\[39\]
rlabel metal2 16606 13209 16606 13209 0 shift_reg\[3\]
rlabel metal2 2162 44574 2162 44574 0 shift_reg\[4\]
rlabel metal1 16790 57494 16790 57494 0 shift_reg\[5\]
rlabel metal2 6854 51680 6854 51680 0 shift_reg\[6\]
rlabel metal2 13202 42432 13202 42432 0 shift_reg\[7\]
rlabel metal2 7958 60333 7958 60333 0 shift_reg\[8\]
rlabel metal2 12558 42307 12558 42307 0 shift_reg\[9\]
<< properties >>
string FIXED_BBOX 0 0 20000 80000
<< end >>
