magic
tech sky130A
magscale 1 2
timestamp 1699972208
<< metal1 >>
rect 23396 117265 23541 120592
rect 23390 117120 23396 117265
rect 23541 117120 23547 117265
rect 23395 112070 23558 112697
rect 23389 111907 23395 112070
rect 23558 111907 23564 112070
rect 23353 104222 23507 104791
rect 23353 104102 23370 104222
rect 23490 104102 23507 104222
rect 23353 104085 23507 104102
rect 23377 99887 23523 100185
rect 23371 99741 23377 99887
rect 23523 99741 23529 99887
rect 23370 96825 23527 97196
rect 23364 96668 23370 96825
rect 23527 96668 23533 96825
rect 23383 93901 23525 94183
rect 23377 93759 23383 93901
rect 23525 93759 23531 93901
rect 23396 66484 23402 66604
rect 23522 66484 23528 66604
rect 23402 66238 23522 66484
rect 23416 63362 23422 63482
rect 23542 63362 23548 63482
rect 23422 63264 23542 63362
rect 23414 60500 23420 60620
rect 23540 60500 23546 60620
rect 23420 60400 23540 60500
rect 23414 60282 23540 60400
rect 23420 60280 23540 60282
rect 23396 55710 23402 55830
rect 23522 55710 23528 55830
rect 23402 55624 23522 55710
rect 36146 55216 36266 55222
rect 32476 55096 36146 55216
rect 36146 55090 36266 55096
rect 36402 50998 36522 51004
rect 32462 50878 36402 50998
rect 36402 50872 36522 50878
rect 36626 48828 36746 48834
rect 32482 48708 36626 48828
rect 36626 48702 36746 48708
rect 23408 47906 23414 48026
rect 23534 47906 23540 48026
rect 23414 47770 23534 47906
rect 36864 47670 36984 47676
rect 32462 47550 36864 47670
rect 36864 47544 36984 47550
rect 37068 46644 37188 46650
rect 32462 46524 37068 46644
rect 37068 46518 37188 46524
rect 37308 45640 37428 45646
rect 32462 45520 37308 45640
rect 37308 45514 37428 45520
rect 23420 40002 23426 40122
rect 23546 40002 23552 40122
rect 23426 39916 23546 40002
<< via1 >>
rect 23396 117120 23541 117265
rect 23395 111907 23558 112070
rect 23370 104102 23490 104222
rect 23377 99741 23523 99887
rect 23370 96668 23527 96825
rect 23383 93759 23525 93901
rect 23402 66484 23522 66604
rect 23422 63362 23542 63482
rect 23420 60500 23540 60620
rect 23402 55710 23522 55830
rect 36146 55096 36266 55216
rect 36402 50878 36522 50998
rect 36626 48708 36746 48828
rect 23414 47906 23534 48026
rect 36864 47550 36984 47670
rect 37068 46524 37188 46644
rect 37308 45520 37428 45640
rect 23426 40002 23546 40122
<< metal2 >>
rect 41279 121449 41288 122419
rect 42258 121449 42267 122419
rect 45288 122379 46258 122388
rect 41288 119602 42258 121449
rect 45288 119602 46258 121409
rect 49279 121403 49288 122373
rect 50258 121403 50267 122373
rect 49288 119602 50258 121403
rect 53279 121315 53288 122285
rect 54258 121315 54267 122285
rect 53288 119602 54258 121315
rect 57279 121189 57288 122159
rect 58258 121189 58267 122159
rect 57288 119602 58258 121189
rect 41712 119180 41768 119602
rect 45668 119180 45724 119602
rect 49624 119180 49680 119602
rect 53580 119180 53636 119602
rect 57536 119180 57592 119602
rect 23396 117265 23541 117271
rect 39441 117252 39551 117256
rect 23541 117247 39556 117252
rect 23541 117137 39441 117247
rect 39551 117137 39556 117247
rect 23541 117132 39556 117137
rect 39441 117128 39551 117132
rect 23396 117114 23541 117120
rect 39349 115348 39459 115352
rect 30314 115343 39464 115348
rect 30314 115233 39349 115343
rect 39459 115233 39464 115343
rect 30314 115228 39464 115233
rect 23395 112070 23558 112076
rect 30314 112048 30434 115228
rect 39349 115224 39459 115228
rect 39357 113444 39467 113448
rect 23558 111928 30434 112048
rect 30646 113439 39472 113444
rect 30646 113329 39357 113439
rect 39467 113329 39472 113439
rect 30646 113324 39472 113329
rect 23395 111901 23558 111907
rect 23370 104222 23490 104228
rect 30646 104222 30766 113324
rect 39357 113320 39467 113324
rect 39311 111540 39421 111544
rect 23490 104102 30766 104222
rect 30928 111535 39426 111540
rect 30928 111425 39311 111535
rect 39421 111425 39426 111535
rect 30928 111420 39426 111425
rect 23370 104096 23490 104102
rect 23377 99887 23523 99893
rect 30928 99874 31048 111420
rect 39311 111416 39421 111420
rect 39321 109636 39431 109640
rect 23523 99754 31048 99874
rect 31240 109631 39436 109636
rect 31240 109521 39321 109631
rect 39431 109521 39436 109631
rect 31240 109516 39436 109521
rect 23377 99735 23523 99741
rect 23370 96825 23527 96831
rect 31240 96806 31360 109516
rect 39321 109512 39431 109516
rect 39293 107732 39403 107736
rect 23527 96686 31360 96806
rect 31504 107727 39408 107732
rect 31504 107617 39293 107727
rect 39403 107617 39408 107727
rect 31504 107612 39408 107617
rect 23370 96662 23527 96668
rect 23383 93901 23525 93907
rect 31504 93890 31624 107612
rect 39293 107608 39403 107612
rect 37760 94399 37880 94404
rect 37756 94289 37765 94399
rect 37875 94289 37884 94399
rect 23525 93770 31624 93890
rect 23383 93753 23525 93759
rect 37760 81944 37880 94289
rect 38026 92495 38146 92500
rect 38022 92385 38031 92495
rect 38141 92385 38150 92495
rect 31660 81824 37880 81944
rect 31660 79000 31780 81824
rect 38026 81670 38146 92385
rect 38232 90591 38352 90596
rect 38228 90481 38237 90591
rect 38347 90481 38356 90591
rect 31651 78880 31660 79000
rect 31761 78880 31780 79000
rect 31892 81550 38146 81670
rect 31892 78806 32012 81550
rect 38232 81420 38352 90481
rect 38488 88687 38608 88692
rect 38484 88577 38493 88687
rect 38603 88577 38612 88687
rect 31883 78686 31892 78806
rect 31992 78686 32012 78806
rect 32072 81300 38352 81420
rect 32072 78614 32192 81300
rect 38488 81180 38608 88577
rect 38752 86792 38848 86800
rect 38749 86783 38859 86792
rect 38749 86664 38859 86673
rect 32306 81060 38608 81180
rect 32063 78494 32072 78614
rect 32192 78494 32201 78614
rect 32306 78426 32426 81060
rect 32563 80930 32649 80934
rect 38752 80930 38848 86664
rect 38910 84767 38919 84902
rect 39054 84767 39063 84902
rect 32558 80925 38848 80930
rect 32558 80839 32563 80925
rect 32649 80839 38848 80925
rect 32558 80834 38848 80839
rect 32563 80830 32649 80834
rect 32759 80742 32845 80746
rect 38938 80742 39034 84767
rect 39115 82860 39124 83024
rect 39288 82860 39297 83024
rect 32754 80737 39034 80742
rect 32754 80651 32759 80737
rect 32845 80651 39034 80737
rect 32754 80646 39034 80651
rect 32759 80642 32845 80646
rect 32571 80526 32657 80530
rect 39158 80526 39254 82860
rect 39362 81071 39458 81084
rect 39346 80961 39355 81071
rect 39465 80961 39474 81071
rect 32566 80521 39254 80526
rect 32566 80435 32571 80521
rect 32657 80435 39254 80521
rect 32566 80430 39254 80435
rect 32571 80426 32657 80430
rect 32837 80346 32923 80350
rect 39362 80346 39458 80961
rect 32832 80341 39458 80346
rect 32832 80255 32837 80341
rect 32923 80255 39458 80341
rect 32832 80250 39458 80255
rect 32837 80246 32923 80250
rect 32297 78306 32306 78426
rect 32426 78306 32435 78426
rect 15846 76408 15966 76418
rect 15846 76309 16629 76408
rect 24688 76310 25296 76406
rect 30200 76310 30742 76406
rect 15846 73572 15966 76309
rect 16084 76261 16204 76272
rect 16084 76164 16642 76261
rect 24742 76166 25122 76262
rect 16084 74315 16204 76164
rect 16080 74205 16089 74315
rect 16199 74205 16208 74315
rect 16084 74200 16204 74205
rect 25026 73790 25122 76166
rect 25200 73970 25296 76310
rect 30202 76166 30602 76262
rect 30506 74470 30602 76166
rect 30646 74650 30742 76310
rect 30637 74554 30646 74650
rect 30742 74554 30751 74650
rect 30497 74374 30506 74470
rect 30602 74374 30611 74470
rect 25200 73874 28328 73970
rect 25026 73694 28134 73790
rect 28232 73746 28328 73874
rect 25829 73572 25939 73576
rect 15846 73567 25944 73572
rect 15846 73457 25829 73567
rect 25939 73457 25944 73567
rect 28038 73560 28134 73694
rect 28223 73650 28232 73746
rect 28328 73650 28337 73746
rect 28029 73464 28038 73560
rect 28134 73464 28143 73560
rect 15846 73452 25944 73457
rect 25829 73448 25939 73452
rect 23402 66604 23522 66610
rect 30585 66606 30695 66610
rect 28796 66604 30700 66606
rect 23522 66601 30700 66604
rect 23522 66491 30585 66601
rect 30695 66491 30700 66601
rect 23522 66486 30700 66491
rect 23522 66484 29500 66486
rect 23402 66478 23522 66484
rect 30585 66482 30695 66486
rect 32624 66019 32633 66129
rect 32743 66019 32752 66129
rect 32644 65474 32733 66019
rect 33218 65729 33227 65839
rect 33337 65729 33346 65839
rect 33236 65476 33329 65729
rect 23422 63482 23542 63488
rect 30297 63482 30407 63486
rect 23542 63477 30412 63482
rect 23542 63367 30297 63477
rect 30407 63367 30412 63477
rect 23542 63362 30412 63367
rect 23422 63356 23542 63362
rect 30297 63358 30407 63362
rect 23420 60620 23540 60626
rect 23540 60500 30556 60620
rect 23420 60494 23540 60500
rect 23402 55830 23522 55836
rect 29808 55830 29928 55840
rect 23522 55710 30186 55830
rect 23402 55704 23522 55710
rect 23408 48064 29484 48184
rect 23408 48032 23528 48064
rect 23408 48026 23534 48032
rect 23408 47906 23414 48026
rect 23408 47902 23534 47906
rect 23414 47900 23534 47902
rect 29364 40434 29484 48064
rect 29808 40700 29928 55710
rect 30436 40955 30556 60500
rect 36151 55216 36261 55220
rect 36140 55096 36146 55216
rect 36266 55096 36272 55216
rect 36151 55092 36261 55096
rect 36407 50998 36517 51002
rect 36396 50878 36402 50998
rect 36522 50878 36528 50998
rect 36407 50874 36517 50878
rect 36631 48828 36741 48832
rect 36620 48708 36626 48828
rect 36746 48708 36752 48828
rect 36631 48704 36741 48708
rect 36869 47670 36979 47674
rect 36858 47550 36864 47670
rect 36984 47550 36990 47670
rect 36869 47546 36979 47550
rect 37073 46644 37183 46648
rect 37062 46524 37068 46644
rect 37188 46524 37194 46644
rect 37073 46520 37183 46524
rect 37313 45640 37423 45644
rect 37302 45520 37308 45640
rect 37428 45520 37434 45640
rect 37313 45516 37423 45520
rect 30432 40845 30441 40955
rect 30551 40845 30560 40955
rect 30436 40840 30556 40845
rect 30247 40700 30357 40704
rect 29808 40695 30362 40700
rect 29808 40585 30247 40695
rect 30357 40585 30362 40695
rect 29808 40580 30362 40585
rect 30247 40576 30357 40580
rect 30463 40434 30573 40438
rect 29364 40429 30578 40434
rect 29364 40319 30463 40429
rect 30573 40319 30578 40429
rect 29364 40314 30578 40319
rect 30463 40310 30573 40314
rect 23426 40122 23546 40128
rect 23546 40117 30392 40122
rect 23546 40007 30277 40117
rect 30387 40007 30396 40117
rect 23546 40002 30392 40007
rect 23426 39996 23546 40002
<< via2 >>
rect 41288 121449 42258 122419
rect 45288 121409 46258 122379
rect 49288 121403 50258 122373
rect 53288 121315 54258 122285
rect 57288 121189 58258 122159
rect 39441 117137 39551 117247
rect 39349 115233 39459 115343
rect 39357 113329 39467 113439
rect 39311 111425 39421 111535
rect 39321 109521 39431 109631
rect 39293 107617 39403 107727
rect 37765 94289 37875 94399
rect 38031 92385 38141 92495
rect 38237 90481 38347 90591
rect 31660 78880 31761 79000
rect 38493 88577 38603 88687
rect 31892 78686 31992 78806
rect 38749 86673 38859 86783
rect 32072 78494 32192 78614
rect 38919 84767 39054 84902
rect 32563 80839 32649 80925
rect 39124 82860 39288 83024
rect 32759 80651 32845 80737
rect 39355 80961 39465 81071
rect 32571 80435 32657 80521
rect 32837 80255 32923 80341
rect 32306 78306 32426 78426
rect 16089 74205 16199 74315
rect 30646 74554 30742 74650
rect 30506 74374 30602 74470
rect 25829 73457 25939 73567
rect 28232 73650 28328 73746
rect 28038 73464 28134 73560
rect 30585 66491 30695 66601
rect 32633 66019 32743 66129
rect 33227 65729 33337 65839
rect 30297 63367 30407 63477
rect 36151 55101 36261 55211
rect 36407 50883 36517 50993
rect 36631 48713 36741 48823
rect 36869 47555 36979 47665
rect 37073 46529 37183 46639
rect 37313 45525 37423 45635
rect 30441 40845 30551 40955
rect 30247 40585 30357 40695
rect 30463 40319 30573 40429
rect 30277 40007 30387 40117
<< metal3 >>
rect -8704 459120 -4244 461120
rect -9044 456660 -4244 459120
rect -8704 399284 -4244 456660
rect -8704 396674 -8426 399284
rect -4476 396674 -4244 399284
rect -8704 396452 -4244 396674
rect 956 459120 5416 461120
rect 956 456660 5756 459120
rect 956 399298 5416 456660
rect 127517 427426 128487 460073
rect 127517 426458 127518 427426
rect 128486 426458 128487 427426
rect 127517 426457 128487 426458
rect 127518 426452 128486 426457
rect 170925 421880 171895 460071
rect 170925 420912 170926 421880
rect 171894 420912 171895 421880
rect 170925 420911 171895 420912
rect 170926 420906 171894 420911
rect 213771 414686 214741 460049
rect 213771 413718 213772 414686
rect 214740 413718 214741 414686
rect 213771 413717 214741 413718
rect 213772 413712 214740 413717
rect 257093 410356 258063 460067
rect 257093 409388 257094 410356
rect 258062 409388 258063 410356
rect 257093 409387 258063 409388
rect 257094 409382 258062 409387
rect 300471 406092 301441 459983
rect 300471 405124 300472 406092
rect 301440 405124 301441 406092
rect 300471 405123 301441 405124
rect 300472 405118 301440 405123
rect 956 396688 1170 399298
rect 5120 396688 5416 399298
rect 956 396468 5416 396688
rect 41277 121454 41283 122424
rect 42263 121454 42269 122424
rect 45283 122384 46253 122390
rect 46253 122379 46263 122384
rect 41283 121449 41288 121454
rect 42258 121449 42263 121454
rect 41283 121444 42263 121449
rect 46258 121409 46263 122379
rect 46253 121404 46263 121409
rect 49277 121408 49283 122378
rect 50263 121408 50269 122378
rect 45283 121398 46253 121404
rect 49283 121403 49288 121408
rect 50258 121403 50263 121408
rect 49283 121398 50263 121403
rect 53277 121320 53283 122290
rect 54263 121320 54269 122290
rect 53283 121315 53288 121320
rect 54258 121315 54263 121320
rect 53283 121310 54263 121315
rect 57277 121194 57283 122164
rect 58263 121194 58269 122164
rect 57283 121189 57288 121194
rect 58258 121189 58263 121194
rect 57283 121184 58263 121189
rect 39408 117247 39818 117252
rect 39408 117137 39441 117247
rect 39551 117137 39818 117247
rect 39408 117132 39818 117137
rect 39344 115343 40212 115348
rect 39344 115233 39349 115343
rect 39459 115233 40212 115343
rect 39344 115228 40212 115233
rect 39352 113439 40222 113444
rect 39352 113329 39357 113439
rect 39467 113329 40222 113439
rect 39352 113324 40222 113329
rect 39306 111535 40152 111540
rect 39306 111425 39311 111535
rect 39421 111425 40152 111535
rect 39306 111420 40152 111425
rect 39316 109631 40122 109636
rect 39316 109521 39321 109631
rect 39431 109521 40122 109631
rect 39316 109516 40122 109521
rect 39288 107727 40138 107732
rect 39288 107617 39293 107727
rect 39403 107617 40138 107727
rect 39288 107612 40138 107617
rect 37760 94399 40052 94404
rect 37760 94289 37765 94399
rect 37875 94289 40052 94399
rect 37760 94284 40052 94289
rect 38026 92495 40222 92500
rect 38026 92385 38031 92495
rect 38141 92385 40222 92495
rect 38026 92380 40222 92385
rect 38232 90591 40254 90596
rect 38232 90481 38237 90591
rect 38347 90481 40254 90591
rect 38232 90476 40254 90481
rect 38488 88687 39754 88692
rect 38488 88577 38493 88687
rect 38603 88577 39754 88687
rect 38488 88572 39754 88577
rect 38744 86783 39754 86788
rect 38744 86673 38749 86783
rect 38859 86673 39754 86783
rect 38744 86668 39754 86673
rect 38914 84902 39059 84907
rect 38914 84767 38919 84902
rect 39054 84767 39897 84902
rect 38914 84762 39059 84767
rect 39119 83024 39293 83029
rect 39119 82860 39124 83024
rect 39288 82860 39766 83024
rect 39119 82855 39293 82860
rect 39350 81071 39754 81076
rect 39350 80961 39355 81071
rect 39465 80961 39754 81071
rect 39350 80956 39754 80961
rect 26490 80925 32654 80930
rect 26490 80839 32563 80925
rect 32649 80839 32654 80925
rect 26490 80834 32654 80839
rect 26490 78986 26586 80834
rect 24950 78890 26586 78986
rect 26666 80737 32850 80742
rect 26666 80651 32759 80737
rect 32845 80651 32850 80737
rect 26666 80646 32850 80651
rect 26666 78794 26762 80646
rect 24868 78698 26762 78794
rect 26878 80521 32662 80526
rect 26878 80435 32571 80521
rect 32657 80435 32662 80521
rect 26878 80430 32662 80435
rect 26878 78602 26974 80430
rect 24630 78506 26974 78602
rect 27062 80341 32928 80346
rect 27062 80255 32837 80341
rect 32923 80255 32928 80341
rect 27062 80250 32928 80255
rect 27062 78410 27158 80250
rect 38734 79150 39754 79172
rect 38732 79052 39754 79150
rect 31649 78875 31655 79005
rect 31756 79000 31766 79005
rect 31761 78880 31766 79000
rect 31756 78875 31766 78880
rect 31881 78681 31887 78811
rect 31987 78806 31997 78811
rect 31992 78686 31997 78806
rect 31987 78681 31997 78686
rect 32061 78489 32067 78619
rect 32187 78614 32197 78619
rect 32192 78494 32197 78614
rect 32187 78489 32197 78494
rect 24854 78314 27158 78410
rect 32295 78301 32301 78431
rect 32421 78426 32431 78431
rect 32426 78306 32431 78426
rect 32421 78301 32431 78306
rect 30641 74650 30747 74655
rect 38732 74650 38828 79052
rect 38930 77268 39026 77286
rect 38926 77148 39764 77268
rect 30641 74554 30646 74650
rect 30742 74554 38828 74650
rect 30641 74549 30747 74554
rect 30501 74470 30607 74475
rect 38930 74470 39026 77148
rect 39190 75244 39756 75364
rect 30501 74374 30506 74470
rect 30602 74374 39026 74470
rect 30501 74369 30607 74374
rect 16084 74315 21872 74320
rect 16084 74205 16089 74315
rect 16199 74205 21872 74315
rect 39194 74230 39290 75244
rect 16084 74200 21872 74205
rect 21752 74054 21872 74200
rect 31536 74134 39290 74230
rect 21752 73934 24748 74054
rect 24628 73808 24748 73934
rect 27760 73808 27880 73812
rect 24628 73688 27880 73808
rect 25824 73567 27626 73572
rect 25824 73457 25829 73567
rect 25939 73457 27626 73567
rect 25824 73452 27626 73457
rect 27506 72990 27626 73452
rect 27760 73254 27880 73688
rect 28227 73746 28333 73751
rect 31536 73746 31632 74134
rect 28227 73650 28232 73746
rect 28328 73650 31632 73746
rect 28227 73645 28333 73650
rect 28033 73560 28139 73565
rect 28033 73464 28038 73560
rect 28134 73464 36704 73560
rect 28033 73459 28139 73464
rect 36608 73460 36704 73464
rect 36608 73340 39788 73460
rect 27760 73134 36414 73254
rect 27506 72870 36126 72990
rect 36006 69652 36126 72870
rect 36294 71556 36414 73134
rect 36294 71436 40048 71556
rect 36006 69532 39988 69652
rect 39282 67628 39996 67748
rect 30580 66601 30700 66606
rect 30580 66491 30585 66601
rect 30695 66491 30700 66601
rect 30292 63477 30412 63482
rect 30292 63367 30297 63477
rect 30407 63367 30412 63477
rect 30292 41170 30412 63367
rect 30580 41394 30700 66491
rect 39282 66134 39402 67628
rect 32628 66129 39402 66134
rect 32628 66019 32633 66129
rect 32743 66019 39402 66129
rect 32628 66014 39402 66019
rect 33222 65839 39904 65844
rect 33222 65729 33227 65839
rect 33337 65729 39904 65839
rect 33222 65724 39904 65729
rect 36146 63820 40074 63940
rect 36146 55211 36266 63820
rect 36146 55101 36151 55211
rect 36261 55101 36266 55211
rect 36146 55096 36266 55101
rect 36402 61916 40082 62036
rect 36402 50993 36522 61916
rect 36402 50883 36407 50993
rect 36517 50883 36522 50993
rect 36402 50878 36522 50883
rect 36626 60012 39884 60132
rect 36626 48823 36746 60012
rect 36626 48713 36631 48823
rect 36741 48713 36746 48823
rect 36626 48708 36746 48713
rect 36864 58108 39878 58228
rect 36864 47665 36984 58108
rect 36864 47555 36869 47665
rect 36979 47555 36984 47665
rect 36864 47550 36984 47555
rect 37068 56204 40082 56324
rect 37068 46639 37188 56204
rect 37068 46529 37073 46639
rect 37183 46529 37188 46639
rect 37068 46524 37188 46529
rect 37308 54300 40254 54420
rect 37308 45635 37428 54300
rect 37308 45525 37313 45635
rect 37423 45525 37428 45635
rect 37308 45520 37428 45525
rect 37624 52396 40152 52516
rect 30580 41274 31428 41394
rect 30292 41050 31176 41170
rect 30436 40955 30970 40960
rect 30436 40845 30441 40955
rect 30551 40845 30970 40955
rect 30436 40840 30970 40845
rect 30242 40695 30784 40700
rect 30242 40585 30247 40695
rect 30357 40585 30784 40695
rect 30242 40580 30784 40585
rect 30458 40429 30578 40434
rect 30458 40319 30463 40429
rect 30573 40319 30578 40429
rect 30272 40117 30392 40122
rect 30272 40007 30277 40117
rect 30387 40007 30392 40117
rect 30272 37528 30392 40007
rect 30458 37738 30578 40319
rect 30664 37996 30784 40580
rect 30850 38254 30970 40840
rect 31056 38512 31176 41050
rect 31308 38758 31428 41274
rect 37624 38758 37744 52396
rect 31308 38638 37744 38758
rect 38028 50492 40434 50612
rect 38028 38512 38148 50492
rect 31056 38392 38148 38512
rect 38336 48588 39844 48708
rect 38336 38254 38456 48588
rect 30850 38134 38456 38254
rect 38704 46684 40128 46804
rect 38704 37996 38824 46684
rect 30664 37876 38824 37996
rect 39122 44780 40004 44900
rect 39122 37738 39242 44780
rect 30458 37618 39242 37738
rect 39332 42876 39776 42996
rect 39332 37528 39452 42876
rect 30272 37408 39452 37528
rect 84236 -122680 89036 -110420
rect 94236 -122480 99036 -110420
<< via3 >>
rect -8426 396674 -4476 399284
rect 127518 426458 128486 427426
rect 170926 420912 171894 421880
rect 213772 413718 214740 414686
rect 257094 409388 258062 410356
rect 300472 405124 301440 406092
rect 1170 396688 5120 399298
rect 41283 122419 42263 122424
rect 41283 121454 41288 122419
rect 41288 121454 42258 122419
rect 42258 121454 42263 122419
rect 45283 122379 46253 122384
rect 45283 121409 45288 122379
rect 45288 121409 46253 122379
rect 45283 121404 46253 121409
rect 49283 122373 50263 122378
rect 49283 121408 49288 122373
rect 49288 121408 50258 122373
rect 50258 121408 50263 122373
rect 53283 122285 54263 122290
rect 53283 121320 53288 122285
rect 53288 121320 54258 122285
rect 54258 121320 54263 122285
rect 57283 122159 58263 122164
rect 57283 121194 57288 122159
rect 57288 121194 58258 122159
rect 58258 121194 58263 122159
rect 31655 79000 31756 79005
rect 31655 78880 31660 79000
rect 31660 78880 31756 79000
rect 31655 78875 31756 78880
rect 31887 78806 31987 78811
rect 31887 78686 31892 78806
rect 31892 78686 31987 78806
rect 31887 78681 31987 78686
rect 32067 78614 32187 78619
rect 32067 78494 32072 78614
rect 32072 78494 32187 78614
rect 32067 78489 32187 78494
rect 32301 78426 32421 78431
rect 32301 78306 32306 78426
rect 32306 78306 32421 78426
rect 32301 78301 32421 78306
<< metal4 >>
rect 127517 427426 128487 427427
rect 127517 426458 127518 427426
rect 128486 426458 128487 427426
rect 127517 426457 128487 426458
rect 170925 421880 171895 421881
rect 170925 420912 170926 421880
rect 171894 420912 171895 421880
rect 170925 420911 171895 420912
rect 213771 414686 214741 414687
rect 213771 413718 213772 414686
rect 214740 413718 214741 414686
rect 213771 413717 214741 413718
rect 257093 410356 258063 410357
rect 257093 409388 257094 410356
rect 258062 409388 258063 410356
rect 257093 409387 258063 409388
rect 300471 406092 301441 406093
rect 300471 405124 300472 406092
rect 301440 405124 301441 406092
rect 300471 405123 301441 405124
rect -10290 399496 85976 399520
rect -10290 399298 82932 399496
rect -10290 399284 1170 399298
rect -10290 396674 -8426 399284
rect -4476 396688 1170 399284
rect 5120 396688 82932 399298
rect -4476 396674 82932 396688
rect -10290 396476 82932 396674
rect 85952 396476 85976 399496
rect -10290 396452 85976 396476
rect 41282 121454 41283 121455
rect 42263 121454 42264 121455
rect 41282 121453 42264 121454
rect 46252 122384 46254 122385
rect 46253 121404 46254 122384
rect 49282 121408 49283 121409
rect 50263 121408 50264 121409
rect 49282 121407 50264 121408
rect 46252 121403 46254 121404
rect 53282 121320 53283 121321
rect 54263 121320 54264 121321
rect 53282 121319 54264 121320
rect 57282 121194 57283 121195
rect 58263 121194 58264 121195
rect 57282 121193 58264 121194
rect 31654 79005 31757 79006
rect 31654 78991 31655 79005
rect 30510 78890 31655 78991
rect 31654 78875 31655 78890
rect 31756 78875 31757 79005
rect 31654 78874 31757 78875
rect 31886 78811 31988 78812
rect 31886 78796 31887 78811
rect 30498 78696 31887 78796
rect 31886 78681 31887 78696
rect 31987 78681 31988 78811
rect 31886 78680 31988 78681
rect 32066 78619 32188 78620
rect 32066 78603 32067 78619
rect 30496 78506 32067 78603
rect 32066 78489 32067 78506
rect 32187 78489 32188 78619
rect 32066 78488 32188 78489
rect 32300 78431 32422 78432
rect 32300 78418 32301 78431
rect 30389 78315 32301 78418
rect 32300 78301 32301 78315
rect 32421 78301 32422 78431
rect 32300 78300 32422 78301
rect 32115 66220 38565 66277
rect 32115 65852 37716 66220
rect 38450 65852 38565 66220
rect 32115 65797 38565 65852
rect 31132 40750 40272 40778
rect 31132 40748 39902 40750
rect 31132 40508 31162 40748
rect 31582 40508 39902 40748
rect 31132 40504 39902 40508
rect 40246 40504 40272 40750
rect 31132 40478 40272 40504
<< via4 >>
rect 127541 426481 128463 427403
rect 170949 420935 171871 421857
rect 213795 413741 214717 414663
rect 257117 409411 258039 410333
rect 300495 405147 301417 406069
rect 82932 396476 85952 399496
rect 41282 122424 42264 122425
rect 41282 121455 41283 122424
rect 41283 121455 42263 122424
rect 42263 121455 42264 122424
rect 45282 122384 46252 122385
rect 45282 121404 45283 122384
rect 45283 121404 46252 122384
rect 49282 122378 50264 122379
rect 49282 121409 49283 122378
rect 49283 121409 50263 122378
rect 50263 121409 50264 122378
rect 53282 122290 54264 122291
rect 45282 121403 46252 121404
rect 53282 121321 53283 122290
rect 53283 121321 54263 122290
rect 54263 121321 54264 122290
rect 57282 122164 58264 122165
rect 57282 121195 57283 122164
rect 57283 121195 58263 122164
rect 58263 121195 58264 122164
rect 37716 65852 38450 66220
rect 31162 40508 31582 40748
rect 39902 40504 40246 40750
<< metal5 >>
rect 37391 427403 128487 427427
rect 37391 426481 127541 427403
rect 128463 426481 128487 427403
rect 37391 426457 128487 426481
rect 37391 122425 38361 426457
rect 43149 421857 171895 421881
rect 43149 420935 170949 421857
rect 171871 420935 171895 421857
rect 43149 420911 171895 420935
rect 41258 122425 42288 122449
rect 37391 121455 41282 122425
rect 42264 121455 42288 122425
rect 41258 121431 42288 121455
rect 43149 122379 44119 420911
rect 49288 414663 214741 414687
rect 49288 413741 213795 414663
rect 214717 413741 214741 414663
rect 49288 413717 214741 413741
rect 45258 122385 46276 122409
rect 49288 122403 50258 413717
rect 53288 410333 258063 410357
rect 53288 409411 257117 410333
rect 258039 409411 258063 410333
rect 53288 409387 258063 409411
rect 45258 122379 45282 122385
rect 43149 121409 45282 122379
rect 45258 121403 45282 121409
rect 46252 121403 46276 122385
rect 45258 121379 46276 121403
rect 49258 122379 50288 122403
rect 49258 121409 49282 122379
rect 50264 121409 50288 122379
rect 53288 122315 54258 409387
rect 57288 406069 301441 406093
rect 57288 405147 300495 406069
rect 301417 405147 301441 406069
rect 57288 405123 301441 405147
rect 49258 121385 50288 121409
rect 53258 122291 54288 122315
rect 53258 121321 53282 122291
rect 54264 121321 54288 122291
rect 57288 122189 58258 405123
rect 82908 399496 85976 399520
rect 82908 396476 82932 399496
rect 85952 396476 85976 399496
rect 53258 121297 54288 121321
rect 57258 122165 58288 122189
rect 57258 121195 57282 122165
rect 58264 121195 58288 122165
rect 57258 121171 58288 121195
rect -41400 111217 15839 111537
rect -43144 109536 14753 109873
rect -44878 108216 13771 108536
rect 37648 66644 42412 66964
rect 55648 66644 62412 66964
rect 37648 66220 38566 66644
rect 37648 65852 37716 66220
rect 38450 65852 38566 66220
rect 37648 65798 38566 65852
rect 59344 63982 62412 66644
rect 82908 63982 85976 396476
rect 59344 60914 85976 63982
rect 39872 45984 43752 46304
rect 39874 40750 40272 45984
rect 39874 40504 39902 40750
rect 40246 40504 40272 40750
rect 39874 40478 40272 40504
rect -56662 21296 854 25934
rect -56900 7514 542 12152
rect -50943 -15355 5189 -11352
rect -44867 -28019 48454 -20496
rect -26953 -40398 58454 -32868
use shiftreg  shiftreg_0
timestamp 1699972208
transform -1 0 59634 0 -1 119980
box 658 0 20000 77840
use uwb_transmitter  uwb_transmitter_0
timestamp 1699972208
transform 1 0 13102 0 1 113100
box -78304 -228320 86125 331063
<< labels >>
flabel metal5 -56662 21296 854 25934 0 FreeSans 1600 0 0 0 rfoutn
port 4 nsew
flabel metal5 -56900 7514 542 12152 0 FreeSans 1600 0 0 0 rfoutp
port 5 nsew
flabel metal5 -50943 -15355 5189 -11352 0 FreeSans 1600 0 0 0 utrig
port 1 nsew
flabel metal5 -44867 -28019 48454 -20496 0 FreeSans 1600 0 0 0 avdd
port 2 nsew
flabel metal5 -26953 -40398 58454 -32868 0 FreeSans 1600 0 0 0 vss
port 0 nsew
flabel metal5 -43144 109536 14753 109873 0 FreeSans 1600 0 0 0 pat1ext
port 8 nsew
flabel metal2 45668 119180 45724 119980 0 FreeSans 1600 0 0 0 sen
port 10 nsew
flabel metal2 49624 119180 49680 119980 0 FreeSans 1600 0 0 0 sdo
port 12 nsew
flabel metal2 53580 119180 53636 119980 0 FreeSans 1600 0 0 0 sdi
port 13 nsew
flabel metal2 57536 119180 57592 119980 0 FreeSans 1600 0 0 0 sclk
port 14 nsew
flabel metal2 41712 119180 41768 119980 0 FreeSans 1600 0 0 0 sload
port 15 nsew
flabel metal5 -41400 111217 15839 111537 0 FreeSans 1600 0 0 0 osct1ext
port 16 nsew
flabel metal5 -44878 108216 13771 108536 0 FreeSans 1600 0 0 0 osct2ext
port 17 nsew
flabel metal4 32115 65797 37716 66277 0 FreeSans 1600 0 0 0 dvdd
port 18 nsew
<< end >>
