magic
tech sky130A
magscale 1 2
timestamp 1696931086
<< error_p >>
rect -172 -147 -114 -141
rect 115 -147 173 -141
rect -172 -181 -160 -147
rect 115 -181 127 -147
rect -172 -187 -114 -181
rect 115 -187 173 -181
<< nwell >>
rect -455 -319 455 319
<< pmos >>
rect -255 -100 -225 100
rect -159 -100 -129 100
rect -63 -100 -33 100
rect 33 -100 63 100
rect 129 -100 159 100
rect 225 -100 255 100
<< pdiff >>
rect -317 88 -255 100
rect -317 -88 -305 88
rect -271 -88 -255 88
rect -317 -100 -255 -88
rect -225 88 -159 100
rect -225 -88 -209 88
rect -175 -88 -159 88
rect -225 -100 -159 -88
rect -129 88 -63 100
rect -129 -88 -113 88
rect -79 -88 -63 88
rect -129 -100 -63 -88
rect -33 88 33 100
rect -33 -88 -17 88
rect 17 -88 33 88
rect -33 -100 33 -88
rect 63 88 129 100
rect 63 -88 79 88
rect 113 -88 129 88
rect 63 -100 129 -88
rect 159 88 225 100
rect 159 -88 175 88
rect 209 -88 225 88
rect 159 -100 225 -88
rect 255 88 317 100
rect 255 -88 271 88
rect 305 -88 317 88
rect 255 -100 317 -88
<< pdiffc >>
rect -305 -88 -271 88
rect -209 -88 -175 88
rect -113 -88 -79 88
rect -17 -88 17 88
rect 79 -88 113 88
rect 175 -88 209 88
rect 271 -88 305 88
<< nsubdiff >>
rect -419 249 -323 283
rect 323 249 419 283
rect -419 187 -385 249
rect 385 187 419 249
rect -419 -249 -385 -187
rect 385 -249 419 -187
rect -419 -283 -323 -249
rect 323 -283 419 -249
<< nsubdiffcont >>
rect -323 249 323 283
rect -419 -187 -385 187
rect 385 -187 419 187
rect -323 -283 323 -249
<< poly >>
rect -255 100 -225 126
rect -159 100 -129 126
rect -63 100 -33 126
rect 33 100 63 126
rect 129 100 159 126
rect 225 100 255 126
rect -255 -131 -225 -100
rect -159 -131 -129 -100
rect -63 -131 -33 -100
rect 33 -131 63 -100
rect 129 -131 159 -100
rect 225 -131 255 -100
rect -291 -147 -225 -131
rect -291 -181 -275 -147
rect -241 -181 -225 -147
rect -291 -197 -225 -181
rect -176 -147 -110 -131
rect -176 -181 -160 -147
rect -126 -181 -110 -147
rect -176 -197 -110 -181
rect -63 -147 63 -131
rect -63 -181 -47 -147
rect 47 -181 63 -147
rect -63 -197 63 -181
rect 111 -147 177 -131
rect 111 -181 127 -147
rect 161 -181 177 -147
rect 111 -197 177 -181
rect 225 -147 291 -131
rect 225 -181 241 -147
rect 275 -181 291 -147
rect 225 -197 291 -181
<< polycont >>
rect -275 -181 -241 -147
rect -160 -181 -126 -147
rect -47 -181 47 -147
rect 127 -181 161 -147
rect 241 -181 275 -147
<< locali >>
rect -419 249 -323 283
rect 323 249 419 283
rect -419 187 -385 249
rect 385 187 419 249
rect -305 88 -271 104
rect -305 -104 -271 -88
rect -209 88 -175 104
rect -209 -104 -175 -88
rect -113 88 -79 104
rect -113 -104 -79 -88
rect -17 88 17 104
rect -17 -104 17 -88
rect 79 88 113 104
rect 79 -104 113 -88
rect 175 88 209 104
rect 175 -104 209 -88
rect 271 88 305 104
rect 271 -104 305 -88
rect -291 -181 -275 -147
rect -241 -181 -225 -147
rect -176 -181 -160 -147
rect -126 -181 -110 -147
rect -63 -181 -47 -147
rect 47 -181 63 -147
rect 111 -181 127 -147
rect 161 -181 177 -147
rect 225 -181 241 -147
rect 275 -181 291 -147
rect -419 -249 -385 -187
rect 385 -249 419 -187
rect -419 -283 -323 -249
rect 323 -283 419 -249
<< viali >>
rect -305 -88 -271 88
rect -209 -88 -175 88
rect -113 -88 -79 88
rect -17 -88 17 88
rect 79 -88 113 88
rect 175 -88 209 88
rect 271 -88 305 88
rect -160 -181 -126 -147
rect -47 -181 47 -147
rect 127 -181 161 -147
<< metal1 >>
rect -311 88 -265 100
rect -311 -88 -305 88
rect -271 -88 -265 88
rect -311 -100 -265 -88
rect -215 88 -169 100
rect -215 -88 -209 88
rect -175 -88 -169 88
rect -215 -100 -169 -88
rect -119 88 -73 100
rect -119 -88 -113 88
rect -79 -88 -73 88
rect -119 -100 -73 -88
rect -23 88 23 100
rect -23 -88 -17 88
rect 17 -88 23 88
rect -23 -100 23 -88
rect 73 88 119 100
rect 73 -88 79 88
rect 113 -88 119 88
rect 73 -100 119 -88
rect 169 88 215 100
rect 169 -88 175 88
rect 209 -88 215 88
rect 169 -100 215 -88
rect 265 88 311 100
rect 265 -88 271 88
rect 305 -88 311 88
rect 265 -100 311 -88
rect -172 -147 -114 -141
rect -172 -181 -160 -147
rect -126 -181 -114 -147
rect -172 -187 -114 -181
rect -59 -147 59 -141
rect -59 -181 -47 -147
rect 47 -181 59 -147
rect -59 -187 59 -181
rect 115 -147 173 -141
rect 115 -181 127 -147
rect 161 -181 173 -147
rect 115 -187 173 -181
<< properties >>
string FIXED_BBOX -402 -266 402 266
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 1 l 0.15 m 1 nf 6 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
