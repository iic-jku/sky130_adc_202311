magic
tech sky130A
magscale 1 2
timestamp 1515178157
<< checkpaint >>
rect -1260 -1258 35460 13226
<< viali >>
rect 29929 11305 29963 11339
rect 27813 11237 27847 11271
rect 1915 11203 1949 11237
rect 4813 11203 4847 11237
rect 9091 11203 9125 11237
rect 11759 11203 11793 11237
rect 14565 11203 14599 11237
rect 17417 11203 17451 11237
rect 20269 11203 20303 11237
rect 21695 11203 21729 11237
rect 3709 11169 3743 11203
rect 6469 11169 6503 11203
rect 7297 11169 7331 11203
rect 9965 11169 9999 11203
rect 12817 11169 12851 11203
rect 15669 11169 15703 11203
rect 18521 11169 18555 11203
rect 23397 11169 23431 11203
rect 24409 11169 24443 11203
rect 25237 11169 25271 11203
rect 25329 11169 25363 11203
rect 26065 11169 26099 11203
rect 27261 11169 27295 11203
rect 27905 11169 27939 11203
rect 28917 11169 28951 11203
rect 24593 11101 24627 11135
rect 26249 11101 26283 11135
rect 28365 11101 28399 11135
rect 25053 11033 25087 11067
rect 27169 11033 27203 11067
rect 24225 10965 24259 10999
rect 25881 10965 25915 10999
rect 30205 10761 30239 10795
rect 30757 10761 30791 10795
rect 1593 10557 1627 10591
rect 4721 10557 4755 10591
rect 9413 10557 9447 10591
rect 10517 10557 10551 10591
rect 15025 10557 15059 10591
rect 18061 10557 18095 10591
rect 18521 10557 18555 10591
rect 21373 10557 21407 10591
rect 23949 10557 23983 10591
rect 27721 10557 27755 10591
rect 3387 10523 3421 10557
rect 6469 10523 6503 10557
rect 7665 10523 7699 10557
rect 12219 10523 12253 10557
rect 13369 10523 13403 10557
rect 16313 10523 16347 10557
rect 20315 10523 20349 10557
rect 23121 10523 23155 10557
rect 25697 10523 25731 10557
rect 29423 10523 29457 10557
rect 27077 10421 27111 10455
rect 23305 10217 23339 10251
rect 18797 10149 18831 10183
rect 22845 10149 22879 10183
rect 2237 10115 2271 10149
rect 6239 10115 6273 10149
rect 9367 10115 9401 10149
rect 11897 10115 11931 10149
rect 15025 10115 15059 10149
rect 17647 10115 17681 10149
rect 21603 10115 21637 10149
rect 25973 10115 26007 10149
rect 28549 10115 28583 10149
rect 31723 10115 31757 10149
rect 3985 10081 4019 10115
rect 4445 10081 4479 10115
rect 7573 10081 7607 10115
rect 10149 10081 10183 10115
rect 13277 10081 13311 10115
rect 15945 10081 15979 10115
rect 18889 10081 18923 10115
rect 19901 10081 19935 10115
rect 23489 10081 23523 10115
rect 24225 10081 24259 10115
rect 26801 10081 26835 10115
rect 29929 10081 29963 10115
rect 18705 10013 18739 10047
rect 22385 10013 22419 10047
rect 23673 10013 23707 10047
rect 22477 9945 22511 9979
rect 19257 9877 19291 9911
rect 19717 9605 19751 9639
rect 19901 9605 19935 9639
rect 15853 9537 15887 9571
rect 3709 9469 3743 9503
rect 4721 9469 4755 9503
rect 7297 9469 7331 9503
rect 10425 9469 10459 9503
rect 13093 9469 13127 9503
rect 17233 9469 17267 9503
rect 20637 9469 20671 9503
rect 20729 9469 20763 9503
rect 21465 9469 21499 9503
rect 24501 9469 24535 9503
rect 29193 9469 29227 9503
rect 29653 9469 29687 9503
rect 1961 9435 1995 9469
rect 6515 9435 6549 9469
rect 9091 9435 9125 9469
rect 12173 9435 12207 9469
rect 14795 9435 14829 9469
rect 18889 9435 18923 9469
rect 23121 9435 23155 9469
rect 26203 9435 26237 9469
rect 27445 9435 27479 9469
rect 31401 9435 31435 9469
rect 16037 9401 16071 9435
rect 20177 9401 20211 9435
rect 15945 9333 15979 9367
rect 16405 9333 16439 9367
rect 7389 9129 7423 9163
rect 8677 9129 8711 9163
rect 12173 9129 12207 9163
rect 27721 9061 27755 9095
rect 28917 9061 28951 9095
rect 1915 9027 1949 9061
rect 4721 9027 4755 9061
rect 11345 9027 11379 9061
rect 15025 9027 15059 9061
rect 16221 9027 16255 9061
rect 20545 9027 20579 9061
rect 23351 9027 23385 9061
rect 26847 9027 26881 9061
rect 31723 9027 31757 9061
rect 3709 8993 3743 9027
rect 6469 8993 6503 9027
rect 7481 8993 7515 9027
rect 9597 8993 9631 9027
rect 13277 8993 13311 9027
rect 17877 8993 17911 9027
rect 18797 8993 18831 9027
rect 21649 8993 21683 9027
rect 24409 8993 24443 9027
rect 25053 8993 25087 9027
rect 27813 8993 27847 9027
rect 28457 8993 28491 9027
rect 30021 8993 30055 9027
rect 7297 8925 7331 8959
rect 8493 8925 8527 8959
rect 8585 8925 8619 8959
rect 24225 8925 24259 8959
rect 7849 8857 7883 8891
rect 9045 8857 9079 8891
rect 24593 8789 24627 8823
rect 28365 8789 28399 8823
rect 3709 8381 3743 8415
rect 4721 8381 4755 8415
rect 7297 8381 7331 8415
rect 10517 8381 10551 8415
rect 15025 8381 15059 8415
rect 15945 8381 15979 8415
rect 18613 8381 18647 8415
rect 21465 8381 21499 8415
rect 23949 8381 23983 8415
rect 27169 8381 27203 8415
rect 32137 8381 32171 8415
rect 1915 8347 1949 8381
rect 6515 8347 6549 8381
rect 9091 8347 9125 8381
rect 12173 8347 12207 8381
rect 13369 8347 13403 8381
rect 17693 8347 17727 8381
rect 20269 8347 20303 8381
rect 23167 8347 23201 8381
rect 25743 8347 25777 8381
rect 28825 8347 28859 8381
rect 30435 8347 30469 8381
rect 17509 8041 17543 8075
rect 26893 8041 26927 8075
rect 28549 8041 28583 8075
rect 11897 7973 11931 8007
rect 13277 7973 13311 8007
rect 16773 7973 16807 8007
rect 2099 7939 2133 7973
rect 6147 7939 6181 7973
rect 11115 7939 11149 7973
rect 15485 7939 15519 7973
rect 21603 7939 21637 7973
rect 24593 7939 24627 7973
rect 30711 7939 30745 7973
rect 3893 7905 3927 7939
rect 4353 7905 4387 7939
rect 7389 7905 7423 7939
rect 7481 7905 7515 7939
rect 9413 7905 9447 7939
rect 12081 7905 12115 7939
rect 13829 7905 13863 7939
rect 16681 7905 16715 7939
rect 19901 7905 19935 7939
rect 22569 7905 22603 7939
rect 23397 7905 23431 7939
rect 26249 7905 26283 7939
rect 26985 7905 27019 7939
rect 27997 7905 28031 7939
rect 32413 7905 32447 7939
rect 7297 7837 7331 7871
rect 8769 7837 8803 7871
rect 12265 7837 12299 7871
rect 16957 7837 16991 7871
rect 17969 7837 18003 7871
rect 18981 7837 19015 7871
rect 22753 7837 22787 7871
rect 23581 7837 23615 7871
rect 27537 7837 27571 7871
rect 8309 7769 8343 7803
rect 8401 7769 8435 7803
rect 12909 7769 12943 7803
rect 17601 7769 17635 7803
rect 18521 7769 18555 7803
rect 18613 7769 18647 7803
rect 29101 7769 29135 7803
rect 7849 7701 7883 7735
rect 12817 7701 12851 7735
rect 16313 7701 16347 7735
rect 22385 7701 22419 7735
rect 23213 7701 23247 7735
rect 25145 7497 25179 7531
rect 27077 7497 27111 7531
rect 28181 7497 28215 7531
rect 30941 7497 30975 7531
rect 10425 7429 10459 7463
rect 19625 7429 19659 7463
rect 19717 7429 19751 7463
rect 21465 7429 21499 7463
rect 3065 7361 3099 7395
rect 10149 7361 10183 7395
rect 10609 7361 10643 7395
rect 11253 7361 11287 7395
rect 14933 7361 14967 7395
rect 20085 7361 20119 7395
rect 21373 7361 21407 7395
rect 21833 7361 21867 7395
rect 26065 7361 26099 7395
rect 27629 7361 27663 7395
rect 1777 7293 1811 7327
rect 2421 7293 2455 7327
rect 6837 7293 6871 7327
rect 7297 7293 7331 7327
rect 12265 7293 12299 7327
rect 14841 7293 14875 7327
rect 15669 7293 15703 7327
rect 15945 7293 15979 7327
rect 17141 7293 17175 7327
rect 20545 7293 20579 7327
rect 24593 7293 24627 7327
rect 25329 7293 25363 7327
rect 25421 7293 25455 7327
rect 26157 7293 26191 7327
rect 29837 7293 29871 7327
rect 5089 7259 5123 7293
rect 9091 7259 9125 7293
rect 14013 7259 14047 7293
rect 18797 7259 18831 7293
rect 22891 7259 22925 7293
rect 1961 7225 1995 7259
rect 11345 7225 11379 7259
rect 11437 7225 11471 7259
rect 30389 7225 30423 7259
rect 1593 7157 1627 7191
rect 11805 7157 11839 7191
rect 20729 7157 20763 7191
rect 28733 7157 28767 7191
rect 29285 7157 29319 7191
rect 2421 6953 2455 6987
rect 3985 6953 4019 6987
rect 25145 6953 25179 6987
rect 29929 6953 29963 6987
rect 3617 6885 3651 6919
rect 24225 6885 24259 6919
rect 27445 6885 27479 6919
rect 4813 6851 4847 6885
rect 8861 6851 8895 6885
rect 10471 6851 10505 6885
rect 14565 6851 14599 6885
rect 17141 6851 17175 6885
rect 20315 6851 20349 6885
rect 22845 6851 22879 6885
rect 2329 6817 2363 6851
rect 6561 6817 6595 6851
rect 7113 6817 7147 6851
rect 12265 6817 12299 6851
rect 12909 6817 12943 6851
rect 15485 6817 15519 6851
rect 18613 6817 18647 6851
rect 21097 6817 21131 6851
rect 24409 6817 24443 6851
rect 25237 6817 25271 6851
rect 25881 6817 25915 6851
rect 28549 6817 28583 6851
rect 2237 6749 2271 6783
rect 3433 6749 3467 6783
rect 3525 6749 3559 6783
rect 24593 6749 24627 6783
rect 27997 6749 28031 6783
rect 26341 6681 26375 6715
rect 29101 6681 29135 6715
rect 2789 6613 2823 6647
rect 25789 6613 25823 6647
rect 26893 6613 26927 6647
rect 20637 6409 20671 6443
rect 30665 6409 30699 6443
rect 2513 6341 2547 6375
rect 15761 6341 15795 6375
rect 16681 6341 16715 6375
rect 1961 6273 1995 6307
rect 3617 6273 3651 6307
rect 27169 6273 27203 6307
rect 2145 6205 2179 6239
rect 6377 6205 6411 6239
rect 7297 6205 7331 6239
rect 10425 6205 10459 6239
rect 13093 6205 13127 6239
rect 16129 6205 16163 6239
rect 17049 6205 17083 6239
rect 17969 6205 18003 6239
rect 20729 6205 20763 6239
rect 21465 6205 21499 6239
rect 24409 6205 24443 6239
rect 28089 6205 28123 6239
rect 4629 6171 4663 6205
rect 9091 6171 9125 6205
rect 12219 6171 12253 6205
rect 14795 6171 14829 6205
rect 19717 6171 19751 6205
rect 23167 6171 23201 6205
rect 26203 6171 26237 6205
rect 29837 6171 29871 6205
rect 2053 6137 2087 6171
rect 2973 6069 3007 6103
rect 3341 6069 3375 6103
rect 3433 6069 3467 6103
rect 15669 6069 15703 6103
rect 16589 6069 16623 6103
rect 3617 5865 3651 5899
rect 3985 5865 4019 5899
rect 4813 5763 4847 5797
rect 9091 5763 9125 5797
rect 11943 5763 11977 5797
rect 14565 5763 14599 5797
rect 17647 5763 17681 5797
rect 21235 5763 21269 5797
rect 25973 5763 26007 5797
rect 28595 5763 28629 5797
rect 31723 5763 31757 5797
rect 2421 5729 2455 5763
rect 6561 5729 6595 5763
rect 7297 5729 7331 5763
rect 10241 5729 10275 5763
rect 12817 5729 12851 5763
rect 15853 5729 15887 5763
rect 18521 5729 18555 5763
rect 19533 5729 19567 5763
rect 22477 5729 22511 5763
rect 23121 5729 23155 5763
rect 23213 5729 23247 5763
rect 24225 5729 24259 5763
rect 26801 5729 26835 5763
rect 29929 5729 29963 5763
rect 2237 5661 2271 5695
rect 2329 5661 2363 5695
rect 3433 5661 3467 5695
rect 3525 5661 3559 5695
rect 18705 5661 18739 5695
rect 22293 5661 22327 5695
rect 22937 5593 22971 5627
rect 2789 5525 2823 5559
rect 16865 5321 16899 5355
rect 20453 5321 20487 5355
rect 9137 5253 9171 5287
rect 16957 5253 16991 5287
rect 1961 5185 1995 5219
rect 4537 5185 4571 5219
rect 8585 5185 8619 5219
rect 16221 5185 16255 5219
rect 20821 5185 20855 5219
rect 1593 5117 1627 5151
rect 1777 5117 1811 5151
rect 3709 5117 3743 5151
rect 4721 5117 4755 5151
rect 7941 5117 7975 5151
rect 9965 5117 9999 5151
rect 13001 5117 13035 5151
rect 16037 5117 16071 5151
rect 17969 5117 18003 5151
rect 20637 5117 20671 5151
rect 21465 5117 21499 5151
rect 25973 5117 26007 5151
rect 29101 5117 29135 5151
rect 32137 5117 32171 5151
rect 6193 5083 6227 5117
rect 11759 5083 11793 5117
rect 14749 5083 14783 5117
rect 19625 5083 19659 5117
rect 23167 5083 23201 5117
rect 24317 5083 24351 5117
rect 27445 5083 27479 5117
rect 30435 5083 30469 5117
rect 2421 5049 2455 5083
rect 8769 5049 8803 5083
rect 16129 5049 16163 5083
rect 17325 5049 17359 5083
rect 4629 4981 4663 5015
rect 5089 4981 5123 5015
rect 8677 4981 8711 5015
rect 15669 4981 15703 5015
rect 23673 4777 23707 4811
rect 2237 4675 2271 4709
rect 6193 4675 6227 4709
rect 9321 4675 9355 4709
rect 11943 4675 11977 4709
rect 15025 4675 15059 4709
rect 17647 4675 17681 4709
rect 21695 4675 21729 4709
rect 25973 4675 26007 4709
rect 28549 4675 28583 4709
rect 31723 4675 31757 4709
rect 3985 4641 4019 4675
rect 4445 4641 4479 4675
rect 7665 4641 7699 4675
rect 10241 4641 10275 4675
rect 13277 4641 13311 4675
rect 15945 4641 15979 4675
rect 19993 4641 20027 4675
rect 22661 4641 22695 4675
rect 22753 4641 22787 4675
rect 23305 4641 23339 4675
rect 23489 4641 23523 4675
rect 24225 4641 24259 4675
rect 26801 4641 26835 4675
rect 29929 4641 29963 4675
rect 18981 4573 19015 4607
rect 18613 4505 18647 4539
rect 18521 4437 18555 4471
rect 22477 4437 22511 4471
rect 4997 4233 5031 4267
rect 4445 4097 4479 4131
rect 5733 4097 5767 4131
rect 3709 4029 3743 4063
rect 4537 4029 4571 4063
rect 6745 4029 6779 4063
rect 9965 4029 9999 4063
rect 15025 4029 15059 4063
rect 16129 4029 16163 4063
rect 18797 4029 18831 4063
rect 21465 4029 21499 4063
rect 25973 4029 26007 4063
rect 27169 4029 27203 4063
rect 31677 4029 31711 4063
rect 1961 3995 1995 4029
rect 8493 3995 8527 4029
rect 11759 3995 11793 4029
rect 13369 3995 13403 4029
rect 17877 3995 17911 4029
rect 20453 3995 20487 4029
rect 23167 3995 23201 4029
rect 24317 3995 24351 4029
rect 28871 3995 28905 4029
rect 30021 3995 30055 4029
rect 5917 3961 5951 3995
rect 4629 3893 4663 3927
rect 5825 3893 5859 3927
rect 6285 3893 6319 3927
rect 9413 3893 9447 3927
rect 21097 3689 21131 3723
rect 22293 3689 22327 3723
rect 1777 3621 1811 3655
rect 12173 3621 12207 3655
rect 27169 3621 27203 3655
rect 4813 3587 4847 3621
rect 16681 3587 16715 3621
rect 20315 3587 20349 3621
rect 26295 3587 26329 3621
rect 3985 3553 4019 3587
rect 6561 3553 6595 3587
rect 7297 3553 7331 3587
rect 8125 3553 8159 3587
rect 9137 3553 9171 3587
rect 14105 3553 14139 3587
rect 14933 3553 14967 3587
rect 18521 3553 18555 3587
rect 21281 3553 21315 3587
rect 22109 3553 22143 3587
rect 22937 3553 22971 3587
rect 23029 3553 23063 3587
rect 24501 3553 24535 3587
rect 2789 3485 2823 3519
rect 8217 3485 8251 3519
rect 8309 3485 8343 3519
rect 11713 3485 11747 3519
rect 13461 3485 13495 3519
rect 17969 3485 18003 3519
rect 21465 3485 21499 3519
rect 21925 3485 21959 3519
rect 2145 3417 2179 3451
rect 7113 3417 7147 3451
rect 7757 3417 7791 3451
rect 10819 3417 10853 3451
rect 11897 3417 11931 3451
rect 17601 3417 17635 3451
rect 2237 3349 2271 3383
rect 17509 3349 17543 3383
rect 22753 3349 22787 3383
rect 23673 3349 23707 3383
rect 27629 3349 27663 3383
rect 16405 3145 16439 3179
rect 23213 3145 23247 3179
rect 20085 3077 20119 3111
rect 27077 3077 27111 3111
rect 15853 3009 15887 3043
rect 20453 3009 20487 3043
rect 25605 3009 25639 3043
rect 1685 2941 1719 2975
rect 6745 2941 6779 2975
rect 7297 2941 7331 2975
rect 12449 2941 12483 2975
rect 13093 2941 13127 2975
rect 15945 2941 15979 2975
rect 17509 2941 17543 2975
rect 21373 2941 21407 2975
rect 22293 2941 22327 2975
rect 22477 2941 22511 2975
rect 22661 2941 22695 2975
rect 23305 2941 23339 2975
rect 23857 2941 23891 2975
rect 23949 2941 23983 2975
rect 24593 2941 24627 2975
rect 26249 2941 26283 2975
rect 3387 2907 3421 2941
rect 5089 2907 5123 2941
rect 9045 2907 9079 2941
rect 10747 2907 10781 2941
rect 14795 2907 14829 2941
rect 19165 2907 19199 2941
rect 16037 2873 16071 2907
rect 16865 2873 16899 2907
rect 21649 2873 21683 2907
rect 24501 2873 24535 2907
rect 19993 2805 20027 2839
rect 25145 2805 25179 2839
rect 27629 2805 27663 2839
rect 24777 2601 24811 2635
rect 22017 2533 22051 2567
rect 23581 2533 23615 2567
rect 25881 2533 25915 2567
rect 26985 2533 27019 2567
rect 2007 2499 2041 2533
rect 4813 2499 4847 2533
rect 9367 2499 9401 2533
rect 11943 2499 11977 2533
rect 14565 2499 14599 2533
rect 17371 2499 17405 2533
rect 18889 2499 18923 2533
rect 3801 2465 3835 2499
rect 6561 2465 6595 2499
rect 7573 2465 7607 2499
rect 10149 2465 10183 2499
rect 12817 2465 12851 2499
rect 15577 2465 15611 2499
rect 20637 2465 20671 2499
rect 22201 2465 22235 2499
rect 22385 2465 22419 2499
rect 22845 2465 22879 2499
rect 23673 2465 23707 2499
rect 25329 2465 25363 2499
rect 21557 2397 21591 2431
rect 21281 2329 21315 2363
rect 26433 2329 26467 2363
rect 21097 2261 21131 2295
rect 22937 2261 22971 2295
rect 24225 2261 24259 2295
rect 15669 2057 15703 2091
rect 22109 2057 22143 2091
rect 22661 2057 22695 2091
rect 25513 2057 25547 2091
rect 26065 2057 26099 2091
rect 15761 1989 15795 2023
rect 16773 1989 16807 2023
rect 20821 1989 20855 2023
rect 21465 1989 21499 2023
rect 23305 1989 23339 2023
rect 17049 1921 17083 1955
rect 24409 1921 24443 1955
rect 1685 1853 1719 1887
rect 6745 1853 6779 1887
rect 9413 1853 9447 1887
rect 10425 1853 10459 1887
rect 15117 1853 15151 1887
rect 17969 1853 18003 1887
rect 20453 1853 20487 1887
rect 20637 1853 20671 1887
rect 21373 1853 21407 1887
rect 22017 1853 22051 1887
rect 22845 1853 22879 1887
rect 24961 1853 24995 1887
rect 3341 1819 3375 1853
rect 5043 1819 5077 1853
rect 7665 1819 7699 1853
rect 12219 1819 12253 1853
rect 13369 1819 13403 1853
rect 19671 1819 19705 1853
rect 16129 1785 16163 1819
rect 16589 1717 16623 1751
rect 23949 1717 23983 1751
rect 21649 1513 21683 1547
rect 22845 1513 22879 1547
rect 3663 1411 3697 1445
rect 6239 1411 6273 1445
rect 9367 1411 9401 1445
rect 10517 1411 10551 1445
rect 14795 1411 14829 1445
rect 17647 1411 17681 1445
rect 19303 1411 19337 1445
rect 1961 1377 1995 1411
rect 4537 1377 4571 1411
rect 7573 1377 7607 1411
rect 12265 1377 12299 1411
rect 13001 1377 13035 1411
rect 15945 1377 15979 1411
rect 21005 1377 21039 1411
rect 21741 1377 21775 1411
rect 24225 1309 24259 1343
rect 24869 1309 24903 1343
rect 22293 1241 22327 1275
rect 23397 1241 23431 1275
rect 20269 969 20303 1003
rect 25329 969 25363 1003
rect 14105 901 14139 935
rect 21465 901 21499 935
rect 13001 833 13035 867
rect 13093 833 13127 867
rect 18889 833 18923 867
rect 19349 833 19383 867
rect 22109 833 22143 867
rect 22661 833 22695 867
rect 24869 833 24903 867
rect 3617 765 3651 799
rect 4445 765 4479 799
rect 7297 765 7331 799
rect 10149 765 10183 799
rect 14933 765 14967 799
rect 15669 765 15703 799
rect 18705 765 18739 799
rect 19533 765 19567 799
rect 20177 765 20211 799
rect 21533 765 21567 799
rect 24225 765 24259 799
rect 1961 731 1995 765
rect 6239 731 6273 765
rect 9091 731 9125 765
rect 11943 731 11977 765
rect 17417 731 17451 765
rect 14473 697 14507 731
rect 23121 697 23155 731
rect 13185 629 13219 663
rect 13553 629 13587 663
rect 14013 629 14047 663
rect 15025 629 15059 663
rect 18521 629 18555 663
rect 19717 629 19751 663
<< metal1 >>
rect 4154 11908 4160 11960
rect 4212 11948 4218 11960
rect 22370 11948 22376 11960
rect 4212 11920 22376 11948
rect 4212 11908 4218 11920
rect 22370 11908 22376 11920
rect 22428 11948 22434 11960
rect 30190 11948 30196 11960
rect 22428 11920 30196 11948
rect 22428 11908 22434 11920
rect 30190 11908 30196 11920
rect 30248 11908 30254 11960
rect 3694 11840 3700 11892
rect 3752 11880 3758 11892
rect 12434 11880 12440 11892
rect 3752 11852 12440 11880
rect 3752 11840 3758 11852
rect 12434 11840 12440 11852
rect 12492 11840 12498 11892
rect 12526 11840 12532 11892
rect 12584 11880 12590 11892
rect 20438 11880 20444 11892
rect 12584 11852 20444 11880
rect 12584 11840 12590 11852
rect 20438 11840 20444 11852
rect 20496 11840 20502 11892
rect 30742 11880 30748 11892
rect 28966 11852 30748 11880
rect 3786 11812 3792 11824
rect 2746 11784 3792 11812
rect 1026 11704 1032 11756
rect 1084 11744 1090 11756
rect 2746 11744 2774 11784
rect 3786 11772 3792 11784
rect 3844 11772 3850 11824
rect 3970 11772 3976 11824
rect 4028 11812 4034 11824
rect 20622 11812 20628 11824
rect 4028 11784 20628 11812
rect 4028 11772 4034 11784
rect 20622 11772 20628 11784
rect 20680 11772 20686 11824
rect 12894 11744 12900 11756
rect 1084 11716 2774 11744
rect 3620 11716 12900 11744
rect 1084 11704 1090 11716
rect 2130 11636 2136 11688
rect 2188 11676 2194 11688
rect 3620 11676 3648 11716
rect 12894 11704 12900 11716
rect 12952 11704 12958 11756
rect 12986 11704 12992 11756
rect 13044 11744 13050 11756
rect 14918 11744 14924 11756
rect 13044 11716 14924 11744
rect 13044 11704 13050 11716
rect 14918 11704 14924 11716
rect 14976 11704 14982 11756
rect 21910 11744 21916 11756
rect 15120 11716 21916 11744
rect 2188 11648 3648 11676
rect 2188 11636 2194 11648
rect 3878 11636 3884 11688
rect 3936 11676 3942 11688
rect 15120 11676 15148 11716
rect 21910 11704 21916 11716
rect 21968 11704 21974 11756
rect 28966 11744 28994 11852
rect 30742 11840 30748 11852
rect 30800 11840 30806 11892
rect 22848 11716 28994 11744
rect 3936 11648 15148 11676
rect 3936 11636 3942 11648
rect 15194 11636 15200 11688
rect 15252 11676 15258 11688
rect 22848 11676 22876 11716
rect 15252 11648 22876 11676
rect 15252 11636 15258 11648
rect 22922 11636 22928 11688
rect 22980 11676 22986 11688
rect 29914 11676 29920 11688
rect 22980 11648 29920 11676
rect 22980 11636 22986 11648
rect 29914 11636 29920 11648
rect 29972 11636 29978 11688
rect 934 11568 940 11620
rect 992 11608 998 11620
rect 3050 11608 3056 11620
rect 992 11580 3056 11608
rect 992 11568 998 11580
rect 3050 11568 3056 11580
rect 3108 11568 3114 11620
rect 4062 11568 4068 11620
rect 4120 11608 4126 11620
rect 12342 11608 12348 11620
rect 4120 11580 12348 11608
rect 4120 11568 4126 11580
rect 12342 11568 12348 11580
rect 12400 11568 12406 11620
rect 12434 11568 12440 11620
rect 12492 11608 12498 11620
rect 21450 11608 21456 11620
rect 12492 11580 21456 11608
rect 12492 11568 12498 11580
rect 21450 11568 21456 11580
rect 21508 11568 21514 11620
rect 21818 11568 21824 11620
rect 21876 11608 21882 11620
rect 25682 11608 25688 11620
rect 21876 11580 25688 11608
rect 21876 11568 21882 11580
rect 25682 11568 25688 11580
rect 25740 11568 25746 11620
rect 2774 11500 2780 11552
rect 2832 11540 2838 11552
rect 4706 11540 4712 11552
rect 2832 11512 4712 11540
rect 2832 11500 2838 11512
rect 4706 11500 4712 11512
rect 4764 11500 4770 11552
rect 4798 11500 4804 11552
rect 4856 11540 4862 11552
rect 7282 11540 7288 11552
rect 4856 11512 7288 11540
rect 4856 11500 4862 11512
rect 7282 11500 7288 11512
rect 7340 11500 7346 11552
rect 9674 11500 9680 11552
rect 9732 11540 9738 11552
rect 12066 11540 12072 11552
rect 9732 11512 12072 11540
rect 9732 11500 9738 11512
rect 12066 11500 12072 11512
rect 12124 11500 12130 11552
rect 12158 11500 12164 11552
rect 12216 11540 12222 11552
rect 12986 11540 12992 11552
rect 12216 11512 12992 11540
rect 12216 11500 12222 11512
rect 12986 11500 12992 11512
rect 13044 11500 13050 11552
rect 13078 11500 13084 11552
rect 13136 11540 13142 11552
rect 14550 11540 14556 11552
rect 13136 11512 14556 11540
rect 13136 11500 13142 11512
rect 14550 11500 14556 11512
rect 14608 11500 14614 11552
rect 15930 11500 15936 11552
rect 15988 11540 15994 11552
rect 17402 11540 17408 11552
rect 15988 11512 17408 11540
rect 15988 11500 15994 11512
rect 17402 11500 17408 11512
rect 17460 11500 17466 11552
rect 18046 11500 18052 11552
rect 18104 11540 18110 11552
rect 20254 11540 20260 11552
rect 18104 11512 20260 11540
rect 18104 11500 18110 11512
rect 20254 11500 20260 11512
rect 20312 11500 20318 11552
rect 21358 11500 21364 11552
rect 21416 11540 21422 11552
rect 23934 11540 23940 11552
rect 21416 11512 23940 11540
rect 21416 11500 21422 11512
rect 23934 11500 23940 11512
rect 23992 11500 23998 11552
rect 1104 11450 33028 11472
rect 1104 11398 11610 11450
rect 11662 11398 11674 11450
rect 11726 11398 11738 11450
rect 11790 11398 11802 11450
rect 11854 11398 11866 11450
rect 11918 11398 21610 11450
rect 21662 11398 21674 11450
rect 21726 11398 21738 11450
rect 21790 11398 21802 11450
rect 21854 11398 21866 11450
rect 21918 11398 31610 11450
rect 31662 11398 31674 11450
rect 31726 11398 31738 11450
rect 31790 11398 31802 11450
rect 31854 11398 31866 11450
rect 31918 11398 33028 11450
rect 1104 11376 33028 11398
rect 24118 11296 24124 11348
rect 24176 11336 24182 11348
rect 27706 11336 27712 11348
rect 24176 11308 27712 11336
rect 24176 11296 24182 11308
rect 27706 11296 27712 11308
rect 27764 11296 27770 11348
rect 29914 11296 29920 11348
rect 29972 11296 29978 11348
rect 1903 11237 1961 11243
rect 1903 11234 1915 11237
rect 1596 11212 1915 11234
rect 1578 11160 1584 11212
rect 1636 11206 1915 11212
rect 1636 11160 1642 11206
rect 1903 11203 1915 11206
rect 1949 11203 1961 11237
rect 1903 11197 1961 11203
rect 3694 11160 3700 11212
rect 3752 11160 3758 11212
rect 4798 11194 4804 11246
rect 4856 11194 4862 11246
rect 9079 11237 9137 11243
rect 6454 11160 6460 11212
rect 6512 11160 6518 11212
rect 7282 11160 7288 11212
rect 7340 11160 7346 11212
rect 9079 11203 9091 11237
rect 9125 11234 9137 11237
rect 11747 11237 11805 11243
rect 9125 11212 9398 11234
rect 9125 11206 9404 11212
rect 9125 11203 9137 11206
rect 9079 11197 9137 11203
rect 9370 11172 9404 11206
rect 9398 11160 9404 11172
rect 9456 11160 9462 11212
rect 9950 11160 9956 11212
rect 10008 11160 10014 11212
rect 11747 11203 11759 11237
rect 11793 11234 11805 11237
rect 12066 11234 12072 11280
rect 11793 11228 12072 11234
rect 12124 11228 12130 11280
rect 11793 11206 12112 11228
rect 11793 11203 11805 11206
rect 11747 11197 11805 11203
rect 12158 11160 12164 11212
rect 12216 11200 12222 11212
rect 12805 11203 12863 11209
rect 12805 11200 12817 11203
rect 12216 11172 12817 11200
rect 12216 11160 12222 11172
rect 12805 11169 12817 11172
rect 12851 11169 12863 11203
rect 14550 11194 14556 11246
rect 14608 11194 14614 11246
rect 12805 11163 12863 11169
rect 15654 11160 15660 11212
rect 15712 11160 15718 11212
rect 17402 11194 17408 11246
rect 17460 11194 17466 11246
rect 17770 11160 17776 11212
rect 17828 11200 17834 11212
rect 18509 11203 18567 11209
rect 18509 11200 18521 11203
rect 17828 11172 18521 11200
rect 17828 11160 17834 11172
rect 18509 11169 18521 11172
rect 18555 11169 18567 11203
rect 20254 11194 20260 11246
rect 20312 11194 20318 11246
rect 21358 11228 21364 11280
rect 21416 11234 21422 11280
rect 27801 11271 27859 11277
rect 27801 11268 27813 11271
rect 21683 11237 21741 11243
rect 21683 11234 21695 11237
rect 21416 11228 21695 11234
rect 21376 11206 21695 11228
rect 21683 11203 21695 11206
rect 21729 11203 21741 11237
rect 24412 11240 26004 11268
rect 21683 11197 21741 11203
rect 18509 11163 18567 11169
rect 23106 11160 23112 11212
rect 23164 11200 23170 11212
rect 24412 11209 24440 11240
rect 23385 11203 23443 11209
rect 23385 11200 23397 11203
rect 23164 11172 23397 11200
rect 23164 11160 23170 11172
rect 23385 11169 23397 11172
rect 23431 11169 23443 11203
rect 23385 11163 23443 11169
rect 24397 11203 24455 11209
rect 24397 11169 24409 11203
rect 24443 11169 24455 11203
rect 24397 11163 24455 11169
rect 25225 11203 25283 11209
rect 25225 11169 25237 11203
rect 25271 11169 25283 11203
rect 25225 11163 25283 11169
rect 24026 11092 24032 11144
rect 24084 11132 24090 11144
rect 24581 11135 24639 11141
rect 24581 11132 24593 11135
rect 24084 11104 24593 11132
rect 24084 11092 24090 11104
rect 24581 11101 24593 11104
rect 24627 11132 24639 11135
rect 25130 11132 25136 11144
rect 24627 11104 25136 11132
rect 24627 11101 24639 11104
rect 24581 11095 24639 11101
rect 25130 11092 25136 11104
rect 25188 11092 25194 11144
rect 25240 11132 25268 11163
rect 25314 11160 25320 11212
rect 25372 11200 25378 11212
rect 25866 11200 25872 11212
rect 25372 11172 25872 11200
rect 25372 11160 25378 11172
rect 25866 11160 25872 11172
rect 25924 11160 25930 11212
rect 25976 11132 26004 11240
rect 26068 11240 27813 11268
rect 26068 11209 26096 11240
rect 27801 11237 27813 11240
rect 27847 11237 27859 11271
rect 27801 11231 27859 11237
rect 26053 11203 26111 11209
rect 26053 11169 26065 11203
rect 26099 11169 26111 11203
rect 26878 11200 26884 11212
rect 26053 11163 26111 11169
rect 26160 11172 26884 11200
rect 26160 11132 26188 11172
rect 26878 11160 26884 11172
rect 26936 11160 26942 11212
rect 27246 11160 27252 11212
rect 27304 11160 27310 11212
rect 27890 11160 27896 11212
rect 27948 11200 27954 11212
rect 28905 11203 28963 11209
rect 28905 11200 28917 11203
rect 27948 11172 28917 11200
rect 27948 11160 27954 11172
rect 28905 11169 28917 11172
rect 28951 11169 28963 11203
rect 28905 11163 28963 11169
rect 25240 11104 25360 11132
rect 25976 11104 26188 11132
rect 23382 11024 23388 11076
rect 23440 11064 23446 11076
rect 25041 11067 25099 11073
rect 25041 11064 25053 11067
rect 23440 11036 25053 11064
rect 23440 11024 23446 11036
rect 25041 11033 25053 11036
rect 25087 11033 25099 11067
rect 25332 11064 25360 11104
rect 26234 11092 26240 11144
rect 26292 11092 26298 11144
rect 27264 11132 27292 11160
rect 28353 11135 28411 11141
rect 28353 11132 28365 11135
rect 27264 11104 28365 11132
rect 28353 11101 28365 11104
rect 28399 11101 28411 11135
rect 28353 11095 28411 11101
rect 27157 11067 27215 11073
rect 27157 11064 27169 11067
rect 25332 11036 27169 11064
rect 25041 11027 25099 11033
rect 27157 11033 27169 11036
rect 27203 11033 27215 11067
rect 27157 11027 27215 11033
rect 23474 10956 23480 11008
rect 23532 10996 23538 11008
rect 24213 10999 24271 11005
rect 24213 10996 24225 10999
rect 23532 10968 24225 10996
rect 23532 10956 23538 10968
rect 24213 10965 24225 10968
rect 24259 10965 24271 10999
rect 24213 10959 24271 10965
rect 24302 10956 24308 11008
rect 24360 10996 24366 11008
rect 25869 10999 25927 11005
rect 25869 10996 25881 10999
rect 24360 10968 25881 10996
rect 24360 10956 24366 10968
rect 25869 10965 25881 10968
rect 25915 10965 25927 10999
rect 25869 10959 25927 10965
rect 1104 10906 33028 10928
rect 1104 10854 10950 10906
rect 11002 10854 11014 10906
rect 11066 10854 11078 10906
rect 11130 10854 11142 10906
rect 11194 10854 11206 10906
rect 11258 10854 20950 10906
rect 21002 10854 21014 10906
rect 21066 10854 21078 10906
rect 21130 10854 21142 10906
rect 21194 10854 21206 10906
rect 21258 10854 30950 10906
rect 31002 10854 31014 10906
rect 31066 10854 31078 10906
rect 31130 10854 31142 10906
rect 31194 10854 31206 10906
rect 31258 10854 33028 10906
rect 1104 10832 33028 10854
rect 30190 10752 30196 10804
rect 30248 10752 30254 10804
rect 30742 10752 30748 10804
rect 30800 10752 30806 10804
rect 17586 10616 17592 10668
rect 17644 10656 17650 10668
rect 17644 10628 18552 10656
rect 17644 10616 17650 10628
rect 1578 10548 1584 10600
rect 1636 10548 1642 10600
rect 4709 10591 4767 10597
rect 4709 10588 4721 10591
rect 3375 10557 3433 10563
rect 3375 10523 3387 10557
rect 3421 10554 3433 10557
rect 3712 10560 4721 10588
rect 3712 10554 3740 10560
rect 3421 10526 3740 10554
rect 4709 10557 4721 10560
rect 4755 10557 4767 10591
rect 4709 10551 4767 10557
rect 3421 10523 3433 10526
rect 3375 10517 3433 10523
rect 6454 10514 6460 10566
rect 6512 10514 6518 10566
rect 7650 10514 7656 10566
rect 7708 10514 7714 10566
rect 9398 10548 9404 10600
rect 9456 10548 9462 10600
rect 10505 10591 10563 10597
rect 10505 10557 10517 10591
rect 10551 10588 10563 10591
rect 10778 10588 10784 10600
rect 10551 10560 10784 10588
rect 10551 10557 10563 10560
rect 10505 10551 10563 10557
rect 10778 10548 10784 10560
rect 10836 10548 10842 10600
rect 12207 10557 12265 10563
rect 12207 10523 12219 10557
rect 12253 10554 12265 10557
rect 12253 10532 12572 10554
rect 12253 10526 12532 10532
rect 12253 10523 12265 10526
rect 12207 10517 12265 10523
rect 12526 10480 12532 10526
rect 12584 10480 12590 10532
rect 13354 10514 13360 10566
rect 13412 10514 13418 10566
rect 15010 10548 15016 10600
rect 15068 10548 15074 10600
rect 16298 10514 16304 10566
rect 16356 10514 16362 10566
rect 18046 10548 18052 10600
rect 18104 10548 18110 10600
rect 18524 10597 18552 10628
rect 20714 10616 20720 10668
rect 20772 10656 20778 10668
rect 20772 10628 21864 10656
rect 20772 10616 20778 10628
rect 18509 10591 18567 10597
rect 18509 10557 18521 10591
rect 18555 10557 18567 10591
rect 21361 10591 21419 10597
rect 21361 10588 21373 10591
rect 18509 10551 18567 10557
rect 20303 10557 20361 10563
rect 20303 10523 20315 10557
rect 20349 10554 20361 10557
rect 20640 10560 21373 10588
rect 20640 10554 20668 10560
rect 20349 10526 20668 10554
rect 21361 10557 21373 10560
rect 21407 10557 21419 10591
rect 21361 10551 21419 10557
rect 20349 10523 20361 10526
rect 20303 10517 20361 10523
rect 21836 10452 21864 10628
rect 23106 10514 23112 10566
rect 23164 10514 23170 10566
rect 23934 10548 23940 10600
rect 23992 10548 23998 10600
rect 27709 10591 27767 10597
rect 25682 10514 25688 10566
rect 25740 10514 25746 10566
rect 27709 10557 27721 10591
rect 27755 10588 27767 10591
rect 27755 10560 28120 10588
rect 27755 10557 27767 10560
rect 27709 10551 27767 10557
rect 22002 10452 22008 10464
rect 21836 10424 22008 10452
rect 22002 10412 22008 10424
rect 22060 10412 22066 10464
rect 26050 10412 26056 10464
rect 26108 10452 26114 10464
rect 27065 10455 27123 10461
rect 27065 10452 27077 10455
rect 26108 10424 27077 10452
rect 26108 10412 26114 10424
rect 27065 10421 27077 10424
rect 27111 10421 27123 10455
rect 28092 10452 28120 10560
rect 29411 10557 29469 10563
rect 29411 10523 29423 10557
rect 29457 10554 29469 10557
rect 29457 10526 29776 10554
rect 29457 10523 29469 10526
rect 29411 10517 29469 10523
rect 29748 10520 29776 10526
rect 29914 10520 29920 10532
rect 29748 10492 29920 10520
rect 29914 10480 29920 10492
rect 29972 10480 29978 10532
rect 28350 10452 28356 10464
rect 28092 10424 28356 10452
rect 27065 10415 27123 10421
rect 28350 10412 28356 10424
rect 28408 10412 28414 10464
rect 1104 10362 33028 10384
rect 1104 10310 11610 10362
rect 11662 10310 11674 10362
rect 11726 10310 11738 10362
rect 11790 10310 11802 10362
rect 11854 10310 11866 10362
rect 11918 10310 21610 10362
rect 21662 10310 21674 10362
rect 21726 10310 21738 10362
rect 21790 10310 21802 10362
rect 21854 10310 21866 10362
rect 21918 10310 31610 10362
rect 31662 10310 31674 10362
rect 31726 10310 31738 10362
rect 31790 10310 31802 10362
rect 31854 10310 31866 10362
rect 31918 10310 33028 10362
rect 1104 10288 33028 10310
rect 17954 10208 17960 10260
rect 18012 10248 18018 10260
rect 19058 10248 19064 10260
rect 18012 10220 19064 10248
rect 18012 10208 18018 10220
rect 19058 10208 19064 10220
rect 19116 10208 19122 10260
rect 20530 10248 20536 10260
rect 20180 10220 20536 10248
rect 9950 10180 9956 10192
rect 2222 10106 2228 10158
rect 2280 10106 2286 10158
rect 6227 10149 6285 10155
rect 3973 10115 4031 10121
rect 3973 10081 3985 10115
rect 4019 10112 4031 10115
rect 4154 10112 4160 10124
rect 4019 10084 4160 10112
rect 4019 10081 4031 10084
rect 3973 10075 4031 10081
rect 4154 10072 4160 10084
rect 4212 10072 4218 10124
rect 4433 10115 4491 10121
rect 4433 10081 4445 10115
rect 4479 10081 4491 10115
rect 6227 10115 6239 10149
rect 6273 10146 6285 10149
rect 9355 10149 9413 10155
rect 6273 10118 6592 10146
rect 6273 10115 6285 10118
rect 6227 10109 6285 10115
rect 6564 10112 6592 10118
rect 6822 10112 6828 10124
rect 6564 10084 6828 10112
rect 4433 10075 4491 10081
rect 3510 10004 3516 10056
rect 3568 10044 3574 10056
rect 4448 10044 4476 10075
rect 6822 10072 6828 10084
rect 6880 10072 6886 10124
rect 7190 10072 7196 10124
rect 7248 10112 7254 10124
rect 7561 10115 7619 10121
rect 7561 10112 7573 10115
rect 7248 10084 7573 10112
rect 7248 10072 7254 10084
rect 7561 10081 7573 10084
rect 7607 10081 7619 10115
rect 9355 10115 9367 10149
rect 9401 10146 9413 10149
rect 9692 10152 9956 10180
rect 9692 10146 9720 10152
rect 9401 10118 9720 10146
rect 9950 10140 9956 10152
rect 10008 10140 10014 10192
rect 11885 10149 11943 10155
rect 9401 10115 9413 10118
rect 9355 10109 9413 10115
rect 7561 10075 7619 10081
rect 9766 10072 9772 10124
rect 9824 10112 9830 10124
rect 10137 10115 10195 10121
rect 10137 10112 10149 10115
rect 9824 10084 10149 10112
rect 9824 10072 9830 10084
rect 10137 10081 10149 10084
rect 10183 10081 10195 10115
rect 11885 10115 11897 10149
rect 11931 10146 11943 10149
rect 11974 10146 11980 10158
rect 11931 10118 11980 10146
rect 11931 10115 11943 10118
rect 11885 10109 11943 10115
rect 11974 10106 11980 10118
rect 12032 10106 12038 10158
rect 10137 10075 10195 10081
rect 12526 10072 12532 10124
rect 12584 10112 12590 10124
rect 13265 10115 13323 10121
rect 13265 10112 13277 10115
rect 12584 10084 13277 10112
rect 12584 10072 12590 10084
rect 13265 10081 13277 10084
rect 13311 10081 13323 10115
rect 15010 10106 15016 10158
rect 15068 10106 15074 10158
rect 17635 10149 17693 10155
rect 13265 10075 13323 10081
rect 15930 10072 15936 10124
rect 15988 10072 15994 10124
rect 17635 10115 17647 10149
rect 17681 10146 17693 10149
rect 17681 10118 18000 10146
rect 18046 10140 18052 10192
rect 18104 10180 18110 10192
rect 18785 10183 18843 10189
rect 18785 10180 18797 10183
rect 18104 10152 18797 10180
rect 18104 10140 18110 10152
rect 18785 10149 18797 10152
rect 18831 10180 18843 10183
rect 18831 10152 19748 10180
rect 18831 10149 18843 10152
rect 18785 10143 18843 10149
rect 17681 10115 17693 10118
rect 17635 10109 17693 10115
rect 17972 10112 18000 10118
rect 18877 10115 18935 10121
rect 18877 10112 18889 10115
rect 17972 10084 18889 10112
rect 18877 10081 18889 10084
rect 18923 10081 18935 10115
rect 19720 10112 19748 10152
rect 19794 10112 19800 10124
rect 19720 10084 19800 10112
rect 18877 10075 18935 10081
rect 19794 10072 19800 10084
rect 19852 10072 19858 10124
rect 19889 10115 19947 10121
rect 19889 10081 19901 10115
rect 19935 10112 19947 10115
rect 20180 10112 20208 10220
rect 20530 10208 20536 10220
rect 20588 10208 20594 10260
rect 22002 10208 22008 10260
rect 22060 10248 22066 10260
rect 23293 10251 23351 10257
rect 23293 10248 23305 10251
rect 22060 10220 23305 10248
rect 22060 10208 22066 10220
rect 23293 10217 23305 10220
rect 23339 10217 23351 10251
rect 23293 10211 23351 10217
rect 19935 10084 20208 10112
rect 21591 10149 21649 10155
rect 21591 10115 21603 10149
rect 21637 10146 21649 10149
rect 21637 10118 21956 10146
rect 22094 10140 22100 10192
rect 22152 10180 22158 10192
rect 22833 10183 22891 10189
rect 22833 10180 22845 10183
rect 22152 10152 22845 10180
rect 22152 10140 22158 10152
rect 22833 10149 22845 10152
rect 22879 10180 22891 10183
rect 23382 10180 23388 10192
rect 22879 10152 23388 10180
rect 22879 10149 22891 10152
rect 22833 10143 22891 10149
rect 23382 10140 23388 10152
rect 23440 10140 23446 10192
rect 21637 10115 21649 10118
rect 21591 10109 21649 10115
rect 21928 10112 21956 10118
rect 22002 10112 22008 10124
rect 21928 10084 22008 10112
rect 19935 10081 19947 10084
rect 19889 10075 19947 10081
rect 22002 10072 22008 10084
rect 22060 10072 22066 10124
rect 23477 10115 23535 10121
rect 23477 10081 23489 10115
rect 23523 10112 23535 10115
rect 24118 10112 24124 10124
rect 23523 10084 24124 10112
rect 23523 10081 23535 10084
rect 23477 10075 23535 10081
rect 24118 10072 24124 10084
rect 24176 10072 24182 10124
rect 24210 10072 24216 10124
rect 24268 10072 24274 10124
rect 25958 10106 25964 10158
rect 26016 10106 26022 10158
rect 26786 10072 26792 10124
rect 26844 10072 26850 10124
rect 28534 10106 28540 10158
rect 28592 10106 28598 10158
rect 31711 10149 31769 10155
rect 29914 10072 29920 10124
rect 29972 10072 29978 10124
rect 31711 10115 31723 10149
rect 31757 10146 31769 10149
rect 31757 10124 32076 10146
rect 31757 10118 32036 10124
rect 31757 10115 31769 10118
rect 31711 10109 31769 10115
rect 32030 10072 32036 10118
rect 32088 10072 32094 10124
rect 3568 10016 4476 10044
rect 18693 10047 18751 10053
rect 3568 10004 3574 10016
rect 18693 10013 18705 10047
rect 18739 10013 18751 10047
rect 20254 10044 20260 10056
rect 18693 10007 18751 10013
rect 18892 10016 20260 10044
rect 18708 9976 18736 10007
rect 18892 9976 18920 10016
rect 20254 10004 20260 10016
rect 20312 10004 20318 10056
rect 22370 10004 22376 10056
rect 22428 10004 22434 10056
rect 23661 10047 23719 10053
rect 23661 10013 23673 10047
rect 23707 10013 23719 10047
rect 23661 10007 23719 10013
rect 18708 9948 18920 9976
rect 22094 9936 22100 9988
rect 22152 9976 22158 9988
rect 22465 9979 22523 9985
rect 22465 9976 22477 9979
rect 22152 9948 22477 9976
rect 22152 9936 22158 9948
rect 22465 9945 22477 9948
rect 22511 9945 22523 9979
rect 23676 9976 23704 10007
rect 24118 9976 24124 9988
rect 23676 9948 24124 9976
rect 22465 9939 22523 9945
rect 24118 9936 24124 9948
rect 24176 9936 24182 9988
rect 18046 9868 18052 9920
rect 18104 9908 18110 9920
rect 18966 9908 18972 9920
rect 18104 9880 18972 9908
rect 18104 9868 18110 9880
rect 18966 9868 18972 9880
rect 19024 9868 19030 9920
rect 19150 9868 19156 9920
rect 19208 9908 19214 9920
rect 19245 9911 19303 9917
rect 19245 9908 19257 9911
rect 19208 9880 19257 9908
rect 19208 9868 19214 9880
rect 19245 9877 19257 9880
rect 19291 9877 19303 9911
rect 19245 9871 19303 9877
rect 1104 9818 33028 9840
rect 1104 9766 10950 9818
rect 11002 9766 11014 9818
rect 11066 9766 11078 9818
rect 11130 9766 11142 9818
rect 11194 9766 11206 9818
rect 11258 9766 20950 9818
rect 21002 9766 21014 9818
rect 21066 9766 21078 9818
rect 21130 9766 21142 9818
rect 21194 9766 21206 9818
rect 21258 9766 30950 9818
rect 31002 9766 31014 9818
rect 31066 9766 31078 9818
rect 31130 9766 31142 9818
rect 31194 9766 31206 9818
rect 31258 9766 33028 9818
rect 1104 9744 33028 9766
rect 15194 9664 15200 9716
rect 15252 9704 15258 9716
rect 17218 9704 17224 9716
rect 15252 9676 17224 9704
rect 15252 9664 15258 9676
rect 17218 9664 17224 9676
rect 17276 9664 17282 9716
rect 21450 9664 21456 9716
rect 21508 9664 21514 9716
rect 19334 9596 19340 9648
rect 19392 9636 19398 9648
rect 19705 9639 19763 9645
rect 19705 9636 19717 9639
rect 19392 9608 19717 9636
rect 19392 9596 19398 9608
rect 19705 9605 19717 9608
rect 19751 9605 19763 9639
rect 19705 9599 19763 9605
rect 19886 9596 19892 9648
rect 19944 9596 19950 9648
rect 21468 9636 21496 9664
rect 20180 9608 21496 9636
rect 3510 9528 3516 9580
rect 3568 9568 3574 9580
rect 3568 9540 4936 9568
rect 3568 9528 3574 9540
rect 1946 9426 1952 9478
rect 2004 9426 2010 9478
rect 3694 9460 3700 9512
rect 3752 9460 3758 9512
rect 4154 9460 4160 9512
rect 4212 9500 4218 9512
rect 4709 9503 4767 9509
rect 4709 9500 4721 9503
rect 4212 9472 4721 9500
rect 4212 9460 4218 9472
rect 4709 9469 4721 9472
rect 4755 9469 4767 9503
rect 4709 9463 4767 9469
rect 4908 9364 4936 9540
rect 6914 9528 6920 9580
rect 6972 9568 6978 9580
rect 6972 9540 7328 9568
rect 6972 9528 6978 9540
rect 7190 9500 7196 9512
rect 6503 9469 6561 9475
rect 6503 9435 6515 9469
rect 6549 9466 6561 9469
rect 6840 9472 7196 9500
rect 6840 9466 6868 9472
rect 6549 9438 6868 9466
rect 7190 9460 7196 9472
rect 7248 9460 7254 9512
rect 7300 9509 7328 9540
rect 9766 9528 9772 9580
rect 9824 9568 9830 9580
rect 10778 9568 10784 9580
rect 9824 9540 10784 9568
rect 9824 9528 9830 9540
rect 10778 9528 10784 9540
rect 10836 9528 10842 9580
rect 15838 9528 15844 9580
rect 15896 9528 15902 9580
rect 16206 9528 16212 9580
rect 16264 9568 16270 9580
rect 17586 9568 17592 9580
rect 16264 9540 17592 9568
rect 16264 9528 16270 9540
rect 17586 9528 17592 9540
rect 17644 9528 17650 9580
rect 7285 9503 7343 9509
rect 7285 9469 7297 9503
rect 7331 9469 7343 9503
rect 10413 9503 10471 9509
rect 10413 9500 10425 9503
rect 7285 9463 7343 9469
rect 9079 9469 9137 9475
rect 6549 9435 6561 9438
rect 6503 9429 6561 9435
rect 9079 9435 9091 9469
rect 9125 9466 9137 9469
rect 9370 9472 10425 9500
rect 9370 9466 9398 9472
rect 9125 9438 9398 9466
rect 10413 9469 10425 9472
rect 10459 9469 10471 9503
rect 10413 9463 10471 9469
rect 9125 9435 9137 9438
rect 9079 9429 9137 9435
rect 12158 9426 12164 9478
rect 12216 9426 12222 9478
rect 13078 9460 13084 9512
rect 13136 9460 13142 9512
rect 15654 9500 15660 9512
rect 14783 9469 14841 9475
rect 14783 9435 14795 9469
rect 14829 9466 14841 9469
rect 15120 9472 15660 9500
rect 15120 9466 15148 9472
rect 14829 9438 15148 9466
rect 15654 9460 15660 9472
rect 15712 9460 15718 9512
rect 17221 9503 17279 9509
rect 17221 9469 17233 9503
rect 17267 9500 17279 9503
rect 17267 9472 17448 9500
rect 17267 9469 17279 9472
rect 17221 9463 17279 9469
rect 14829 9435 14841 9438
rect 14783 9429 14841 9435
rect 16025 9435 16083 9441
rect 16025 9401 16037 9435
rect 16071 9432 16083 9435
rect 17034 9432 17040 9444
rect 16071 9404 17040 9432
rect 16071 9401 16083 9404
rect 16025 9395 16083 9401
rect 17034 9392 17040 9404
rect 17092 9392 17098 9444
rect 5442 9364 5448 9376
rect 4908 9336 5448 9364
rect 5442 9324 5448 9336
rect 5500 9324 5506 9376
rect 15930 9324 15936 9376
rect 15988 9324 15994 9376
rect 16393 9367 16451 9373
rect 16393 9333 16405 9367
rect 16439 9364 16451 9367
rect 16942 9364 16948 9376
rect 16439 9336 16948 9364
rect 16439 9333 16451 9336
rect 16393 9327 16451 9333
rect 16942 9324 16948 9336
rect 17000 9324 17006 9376
rect 17420 9364 17448 9472
rect 18874 9426 18880 9478
rect 18932 9426 18938 9478
rect 19242 9392 19248 9444
rect 19300 9432 19306 9444
rect 20180 9441 20208 9608
rect 20622 9460 20628 9512
rect 20680 9460 20686 9512
rect 20717 9503 20775 9509
rect 20717 9469 20729 9503
rect 20763 9500 20775 9503
rect 21358 9500 21364 9512
rect 20763 9472 21364 9500
rect 20763 9469 20775 9472
rect 20717 9463 20775 9469
rect 21358 9460 21364 9472
rect 21416 9460 21422 9512
rect 21453 9503 21511 9509
rect 21453 9469 21465 9503
rect 21499 9500 21511 9503
rect 24489 9503 24547 9509
rect 21499 9472 21588 9500
rect 21499 9469 21511 9472
rect 21453 9463 21511 9469
rect 20165 9435 20223 9441
rect 20165 9432 20177 9435
rect 19300 9404 20177 9432
rect 19300 9392 19306 9404
rect 20165 9401 20177 9404
rect 20211 9401 20223 9435
rect 20165 9395 20223 9401
rect 17678 9364 17684 9376
rect 17420 9336 17684 9364
rect 17678 9324 17684 9336
rect 17736 9324 17742 9376
rect 21560 9364 21588 9472
rect 23106 9426 23112 9478
rect 23164 9426 23170 9478
rect 24489 9469 24501 9503
rect 24535 9500 24547 9503
rect 26786 9500 26792 9512
rect 24535 9472 24900 9500
rect 24535 9469 24547 9472
rect 24489 9463 24547 9469
rect 22002 9364 22008 9376
rect 21560 9336 22008 9364
rect 22002 9324 22008 9336
rect 22060 9324 22066 9376
rect 24872 9364 24900 9472
rect 26191 9469 26249 9475
rect 26191 9435 26203 9469
rect 26237 9466 26249 9469
rect 26528 9472 26792 9500
rect 26528 9466 26556 9472
rect 26237 9438 26556 9466
rect 26786 9460 26792 9472
rect 26844 9460 26850 9512
rect 26237 9435 26249 9438
rect 26191 9429 26249 9435
rect 27430 9426 27436 9478
rect 27488 9426 27494 9478
rect 29178 9460 29184 9512
rect 29236 9460 29242 9512
rect 29638 9460 29644 9512
rect 29696 9460 29702 9512
rect 31386 9426 31392 9478
rect 31444 9426 31450 9478
rect 25130 9364 25136 9376
rect 24872 9336 25136 9364
rect 25130 9324 25136 9336
rect 25188 9324 25194 9376
rect 1104 9274 33028 9296
rect 1104 9222 11610 9274
rect 11662 9222 11674 9274
rect 11726 9222 11738 9274
rect 11790 9222 11802 9274
rect 11854 9222 11866 9274
rect 11918 9222 21610 9274
rect 21662 9222 21674 9274
rect 21726 9222 21738 9274
rect 21790 9222 21802 9274
rect 21854 9222 21866 9274
rect 21918 9222 31610 9274
rect 31662 9222 31674 9274
rect 31726 9222 31738 9274
rect 31790 9222 31802 9274
rect 31854 9222 31866 9274
rect 31918 9222 33028 9274
rect 1104 9200 33028 9222
rect 5718 9120 5724 9172
rect 5776 9160 5782 9172
rect 5776 9132 6040 9160
rect 5776 9120 5782 9132
rect 1854 9018 1860 9070
rect 1912 9067 1918 9070
rect 1912 9061 1961 9067
rect 1912 9027 1915 9061
rect 1949 9027 1961 9061
rect 1912 9021 1961 9027
rect 3697 9027 3755 9033
rect 1912 9018 1918 9021
rect 3697 8993 3709 9027
rect 3743 9024 3755 9027
rect 3786 9024 3792 9036
rect 3743 8996 3792 9024
rect 3743 8993 3755 8996
rect 3697 8987 3755 8993
rect 3786 8984 3792 8996
rect 3844 8984 3850 9036
rect 4706 9018 4712 9070
rect 4764 9018 4770 9070
rect 6012 8956 6040 9132
rect 6638 9120 6644 9172
rect 6696 9160 6702 9172
rect 7377 9163 7435 9169
rect 7377 9160 7389 9163
rect 6696 9132 7389 9160
rect 6696 9120 6702 9132
rect 7377 9129 7389 9132
rect 7423 9129 7435 9163
rect 7377 9123 7435 9129
rect 8665 9163 8723 9169
rect 8665 9129 8677 9163
rect 8711 9160 8723 9163
rect 9490 9160 9496 9172
rect 8711 9132 9496 9160
rect 8711 9129 8723 9132
rect 8665 9123 8723 9129
rect 9490 9120 9496 9132
rect 9548 9120 9554 9172
rect 11974 9120 11980 9172
rect 12032 9160 12038 9172
rect 12161 9163 12219 9169
rect 12161 9160 12173 9163
rect 12032 9132 12173 9160
rect 12032 9120 12038 9132
rect 12161 9129 12173 9132
rect 12207 9129 12219 9163
rect 22278 9160 22284 9172
rect 12161 9123 12219 9129
rect 21836 9132 22284 9160
rect 9398 9092 9404 9104
rect 6840 9064 9404 9092
rect 6457 9027 6515 9033
rect 6457 8993 6469 9027
rect 6503 9024 6515 9027
rect 6840 9024 6868 9064
rect 9398 9052 9404 9064
rect 9456 9052 9462 9104
rect 6503 8996 6868 9024
rect 6503 8993 6515 8996
rect 6457 8987 6515 8993
rect 6914 8984 6920 9036
rect 6972 9024 6978 9036
rect 7469 9027 7527 9033
rect 7469 9024 7481 9027
rect 6972 8996 7481 9024
rect 6972 8984 6978 8996
rect 7469 8993 7481 8996
rect 7515 8993 7527 9027
rect 7469 8987 7527 8993
rect 9582 8984 9588 9036
rect 9640 8984 9646 9036
rect 11330 9018 11336 9070
rect 11388 9018 11394 9070
rect 11422 9018 11428 9070
rect 11480 9058 11486 9070
rect 11480 9030 11744 9058
rect 11480 9018 11486 9030
rect 11716 9024 11744 9030
rect 12526 9024 12532 9036
rect 11716 8996 12532 9024
rect 12526 8984 12532 8996
rect 12584 8984 12590 9036
rect 13262 8984 13268 9036
rect 13320 8984 13326 9036
rect 15010 9018 15016 9070
rect 15068 9018 15074 9070
rect 16206 9018 16212 9070
rect 16264 9018 16270 9070
rect 17865 9027 17923 9033
rect 17865 8993 17877 9027
rect 17911 9024 17923 9027
rect 18690 9024 18696 9036
rect 17911 8996 18696 9024
rect 17911 8993 17923 8996
rect 17865 8987 17923 8993
rect 18690 8984 18696 8996
rect 18748 8984 18754 9036
rect 18785 9027 18843 9033
rect 18785 8993 18797 9027
rect 18831 8993 18843 9027
rect 20530 9018 20536 9070
rect 20588 9018 20594 9070
rect 21637 9027 21695 9033
rect 18785 8987 18843 8993
rect 21637 8993 21649 9027
rect 21683 9024 21695 9027
rect 21836 9024 21864 9132
rect 22278 9120 22284 9132
rect 22336 9120 22342 9172
rect 27430 9120 27436 9172
rect 27488 9160 27494 9172
rect 29638 9160 29644 9172
rect 27488 9132 29644 9160
rect 27488 9120 27494 9132
rect 29638 9120 29644 9132
rect 29696 9120 29702 9172
rect 30650 9160 30656 9172
rect 30392 9132 30656 9160
rect 24210 9092 24216 9104
rect 21683 8996 21864 9024
rect 23339 9061 23397 9067
rect 23339 9027 23351 9061
rect 23385 9058 23397 9061
rect 23676 9064 24216 9092
rect 23676 9058 23704 9064
rect 23385 9030 23704 9058
rect 24210 9052 24216 9064
rect 24268 9052 24274 9104
rect 26835 9061 26893 9067
rect 23385 9027 23397 9030
rect 23339 9021 23397 9027
rect 21683 8993 21695 8996
rect 21637 8987 21695 8993
rect 7285 8959 7343 8965
rect 6012 8928 6408 8956
rect 6380 8820 6408 8928
rect 7285 8925 7297 8959
rect 7331 8925 7343 8959
rect 8202 8956 8208 8968
rect 7285 8919 7343 8925
rect 7484 8928 8208 8956
rect 7300 8888 7328 8919
rect 7484 8888 7512 8928
rect 8202 8916 8208 8928
rect 8260 8916 8266 8968
rect 8478 8916 8484 8968
rect 8536 8916 8542 8968
rect 8573 8959 8631 8965
rect 8573 8925 8585 8959
rect 8619 8956 8631 8959
rect 10042 8956 10048 8968
rect 8619 8928 8653 8956
rect 8956 8928 10048 8956
rect 8619 8925 8631 8928
rect 8573 8919 8631 8925
rect 7300 8860 7512 8888
rect 7837 8891 7895 8897
rect 7837 8857 7849 8891
rect 7883 8888 7895 8891
rect 8588 8888 8616 8919
rect 8956 8888 8984 8928
rect 10042 8916 10048 8928
rect 10100 8916 10106 8968
rect 17586 8916 17592 8968
rect 17644 8956 17650 8968
rect 18800 8956 18828 8987
rect 24394 8984 24400 9036
rect 24452 8984 24458 9036
rect 24578 8984 24584 9036
rect 24636 9024 24642 9036
rect 25041 9027 25099 9033
rect 25041 9024 25053 9027
rect 24636 8996 25053 9024
rect 24636 8984 24642 8996
rect 25041 8993 25053 8996
rect 25087 8993 25099 9027
rect 26835 9027 26847 9061
rect 26881 9058 26893 9061
rect 26881 9036 27200 9058
rect 27706 9052 27712 9104
rect 27764 9052 27770 9104
rect 28905 9095 28963 9101
rect 28905 9092 28917 9095
rect 27816 9064 28917 9092
rect 26881 9030 27160 9036
rect 26881 9027 26893 9030
rect 26835 9021 26893 9027
rect 25041 8987 25099 8993
rect 27154 8984 27160 9030
rect 27212 8984 27218 9036
rect 27246 8984 27252 9036
rect 27304 9024 27310 9036
rect 27816 9033 27844 9064
rect 28905 9061 28917 9064
rect 28951 9061 28963 9095
rect 28905 9055 28963 9061
rect 27801 9027 27859 9033
rect 27801 9024 27813 9027
rect 27304 8996 27813 9024
rect 27304 8984 27310 8996
rect 27801 8993 27813 8996
rect 27847 8993 27859 9027
rect 27801 8987 27859 8993
rect 28445 9027 28503 9033
rect 28445 8993 28457 9027
rect 28491 8993 28503 9027
rect 28445 8987 28503 8993
rect 30009 9027 30067 9033
rect 30009 8993 30021 9027
rect 30055 9024 30067 9027
rect 30392 9024 30420 9132
rect 30650 9120 30656 9132
rect 30708 9120 30714 9172
rect 30055 8996 30420 9024
rect 31711 9061 31769 9067
rect 31711 9027 31723 9061
rect 31757 9058 31769 9061
rect 31757 9030 32076 9058
rect 31757 9027 31769 9030
rect 31711 9021 31769 9027
rect 32048 9024 32076 9030
rect 32122 9024 32128 9036
rect 32048 8996 32128 9024
rect 30055 8993 30067 8996
rect 30009 8987 30067 8993
rect 19242 8956 19248 8968
rect 17644 8928 18828 8956
rect 18892 8928 19248 8956
rect 17644 8916 17650 8928
rect 7883 8860 8984 8888
rect 9033 8891 9091 8897
rect 7883 8857 7895 8860
rect 7837 8851 7895 8857
rect 9033 8857 9045 8891
rect 9079 8888 9091 8891
rect 9674 8888 9680 8900
rect 9079 8860 9680 8888
rect 9079 8857 9091 8860
rect 9033 8851 9091 8857
rect 9674 8848 9680 8860
rect 9732 8848 9738 8900
rect 17862 8848 17868 8900
rect 17920 8888 17926 8900
rect 18892 8888 18920 8928
rect 19242 8916 19248 8928
rect 19300 8916 19306 8968
rect 21358 8916 21364 8968
rect 21416 8956 21422 8968
rect 22002 8956 22008 8968
rect 21416 8928 22008 8956
rect 21416 8916 21422 8928
rect 22002 8916 22008 8928
rect 22060 8916 22066 8968
rect 24118 8916 24124 8968
rect 24176 8956 24182 8968
rect 24213 8959 24271 8965
rect 24213 8956 24225 8959
rect 24176 8928 24225 8956
rect 24176 8916 24182 8928
rect 24213 8925 24225 8928
rect 24259 8925 24271 8959
rect 24213 8919 24271 8925
rect 27614 8916 27620 8968
rect 27672 8956 27678 8968
rect 28460 8956 28488 8987
rect 32122 8984 32128 8996
rect 32180 8984 32186 9036
rect 28534 8956 28540 8968
rect 27672 8928 28540 8956
rect 27672 8916 27678 8928
rect 28534 8916 28540 8928
rect 28592 8916 28598 8968
rect 17920 8860 18920 8888
rect 17920 8848 17926 8860
rect 27246 8848 27252 8900
rect 27304 8888 27310 8900
rect 29270 8888 29276 8900
rect 27304 8860 29276 8888
rect 27304 8848 27310 8860
rect 29270 8848 29276 8860
rect 29328 8848 29334 8900
rect 9306 8820 9312 8832
rect 6380 8792 9312 8820
rect 9306 8780 9312 8792
rect 9364 8780 9370 8832
rect 11974 8780 11980 8832
rect 12032 8820 12038 8832
rect 12618 8820 12624 8832
rect 12032 8792 12624 8820
rect 12032 8780 12038 8792
rect 12618 8780 12624 8792
rect 12676 8780 12682 8832
rect 23750 8780 23756 8832
rect 23808 8820 23814 8832
rect 24581 8823 24639 8829
rect 24581 8820 24593 8823
rect 23808 8792 24593 8820
rect 23808 8780 23814 8792
rect 24581 8789 24593 8792
rect 24627 8820 24639 8823
rect 24762 8820 24768 8832
rect 24627 8792 24768 8820
rect 24627 8789 24639 8792
rect 24581 8783 24639 8789
rect 24762 8780 24768 8792
rect 24820 8780 24826 8832
rect 28350 8780 28356 8832
rect 28408 8780 28414 8832
rect 1104 8730 33028 8752
rect 1104 8678 10950 8730
rect 11002 8678 11014 8730
rect 11066 8678 11078 8730
rect 11130 8678 11142 8730
rect 11194 8678 11206 8730
rect 11258 8678 20950 8730
rect 21002 8678 21014 8730
rect 21066 8678 21078 8730
rect 21130 8678 21142 8730
rect 21194 8678 21206 8730
rect 21258 8678 30950 8730
rect 31002 8678 31014 8730
rect 31066 8678 31078 8730
rect 31130 8678 31142 8730
rect 31194 8678 31206 8730
rect 31258 8678 33028 8730
rect 1104 8656 33028 8678
rect 5166 8480 5172 8492
rect 3712 8452 5172 8480
rect 3712 8421 3740 8452
rect 5166 8440 5172 8452
rect 5224 8440 5230 8492
rect 14642 8440 14648 8492
rect 14700 8480 14706 8492
rect 14700 8452 15976 8480
rect 14700 8440 14706 8452
rect 3697 8415 3755 8421
rect 1762 8338 1768 8390
rect 1820 8378 1826 8390
rect 1903 8381 1961 8387
rect 1903 8378 1915 8381
rect 1820 8350 1915 8378
rect 1820 8338 1826 8350
rect 1903 8347 1915 8350
rect 1949 8347 1961 8381
rect 3697 8381 3709 8415
rect 3743 8381 3755 8415
rect 3697 8375 3755 8381
rect 4706 8372 4712 8424
rect 4764 8372 4770 8424
rect 7285 8415 7343 8421
rect 7285 8412 7297 8415
rect 6503 8381 6561 8387
rect 1903 8341 1961 8347
rect 6503 8347 6515 8381
rect 6549 8378 6561 8381
rect 6840 8384 7297 8412
rect 6840 8378 6868 8384
rect 6549 8350 6868 8378
rect 7285 8381 7297 8384
rect 7331 8381 7343 8415
rect 9582 8412 9588 8424
rect 7285 8375 7343 8381
rect 9079 8381 9137 8387
rect 6549 8347 6561 8350
rect 6503 8341 6561 8347
rect 9079 8347 9091 8381
rect 9125 8378 9137 8381
rect 9370 8384 9588 8412
rect 9370 8378 9398 8384
rect 9125 8350 9398 8378
rect 9582 8372 9588 8384
rect 9640 8372 9646 8424
rect 10505 8415 10563 8421
rect 10505 8381 10517 8415
rect 10551 8412 10563 8415
rect 10551 8384 10916 8412
rect 10551 8381 10563 8384
rect 10505 8375 10563 8381
rect 9125 8347 9137 8350
rect 9079 8341 9137 8347
rect 10686 8254 10692 8306
rect 10744 8294 10750 8306
rect 10888 8294 10916 8384
rect 12161 8381 12219 8387
rect 12161 8347 12173 8381
rect 12207 8378 12219 8381
rect 12250 8378 12256 8390
rect 12207 8350 12256 8378
rect 12207 8347 12219 8350
rect 12161 8341 12219 8347
rect 12250 8338 12256 8350
rect 12308 8338 12314 8390
rect 13354 8338 13360 8390
rect 13412 8338 13418 8390
rect 15010 8372 15016 8424
rect 15068 8372 15074 8424
rect 15948 8421 15976 8452
rect 15933 8415 15991 8421
rect 15933 8381 15945 8415
rect 15979 8381 15991 8415
rect 18601 8415 18659 8421
rect 15933 8375 15991 8381
rect 17678 8338 17684 8390
rect 17736 8338 17742 8390
rect 18601 8381 18613 8415
rect 18647 8412 18659 8415
rect 18874 8412 18880 8424
rect 18647 8384 18880 8412
rect 18647 8381 18659 8384
rect 18601 8375 18659 8381
rect 18874 8372 18880 8384
rect 18932 8372 18938 8424
rect 21453 8415 21511 8421
rect 20254 8338 20260 8390
rect 20312 8338 20318 8390
rect 21453 8381 21465 8415
rect 21499 8412 21511 8415
rect 23937 8415 23995 8421
rect 23937 8412 23949 8415
rect 21499 8384 21772 8412
rect 21499 8381 21511 8384
rect 21453 8375 21511 8381
rect 10744 8266 10916 8294
rect 21744 8276 21772 8384
rect 23155 8381 23213 8387
rect 23155 8347 23167 8381
rect 23201 8378 23213 8381
rect 23492 8384 23949 8412
rect 23492 8378 23520 8384
rect 23201 8350 23520 8378
rect 23937 8381 23949 8384
rect 23983 8381 23995 8415
rect 23937 8375 23995 8381
rect 25731 8381 25789 8387
rect 23201 8347 23213 8350
rect 23155 8341 23213 8347
rect 25731 8347 25743 8381
rect 25777 8378 25789 8381
rect 25777 8356 26096 8378
rect 27154 8372 27160 8424
rect 27212 8372 27218 8424
rect 25777 8350 26056 8356
rect 25777 8347 25789 8350
rect 25731 8341 25789 8347
rect 26050 8304 26056 8350
rect 26108 8304 26114 8356
rect 28810 8338 28816 8390
rect 28868 8338 28874 8390
rect 29270 8372 29276 8424
rect 29328 8412 29334 8424
rect 29328 8384 30144 8412
rect 29328 8372 29334 8384
rect 30116 8378 30144 8384
rect 30423 8381 30481 8387
rect 30423 8378 30435 8381
rect 30116 8350 30435 8378
rect 30423 8347 30435 8350
rect 30469 8347 30481 8381
rect 32122 8372 32128 8424
rect 32180 8372 32186 8424
rect 30423 8341 30481 8347
rect 22002 8276 22008 8288
rect 10744 8254 10750 8266
rect 21744 8248 22008 8276
rect 22002 8236 22008 8248
rect 22060 8236 22066 8288
rect 1104 8186 33028 8208
rect 1104 8134 11610 8186
rect 11662 8134 11674 8186
rect 11726 8134 11738 8186
rect 11790 8134 11802 8186
rect 11854 8134 11866 8186
rect 11918 8134 21610 8186
rect 21662 8134 21674 8186
rect 21726 8134 21738 8186
rect 21790 8134 21802 8186
rect 21854 8134 21866 8186
rect 21918 8134 31610 8186
rect 31662 8134 31674 8186
rect 31726 8134 31738 8186
rect 31790 8134 31802 8186
rect 31854 8134 31866 8186
rect 31918 8134 33028 8186
rect 1104 8112 33028 8134
rect 11422 8032 11428 8084
rect 11480 8072 11486 8084
rect 13630 8072 13636 8084
rect 11480 8044 13636 8072
rect 11480 8032 11486 8044
rect 13630 8032 13636 8044
rect 13688 8032 13694 8084
rect 14458 8072 14464 8084
rect 14200 8044 14464 8072
rect 6914 8004 6920 8016
rect 2038 7930 2044 7982
rect 2096 7979 2102 7982
rect 2096 7973 2145 7979
rect 2096 7939 2099 7973
rect 2133 7939 2145 7973
rect 6135 7973 6193 7979
rect 2096 7933 2145 7939
rect 2096 7930 2102 7933
rect 3878 7896 3884 7948
rect 3936 7896 3942 7948
rect 4338 7896 4344 7948
rect 4396 7896 4402 7948
rect 6135 7939 6147 7973
rect 6181 7970 6193 7973
rect 6472 7976 6920 8004
rect 6472 7970 6500 7976
rect 6181 7942 6500 7970
rect 6914 7964 6920 7976
rect 6972 7964 6978 8016
rect 7282 7964 7288 8016
rect 7340 8004 7346 8016
rect 8754 8004 8760 8016
rect 7340 7976 8760 8004
rect 7340 7964 7346 7976
rect 8754 7964 8760 7976
rect 8812 7964 8818 8016
rect 11103 7973 11161 7979
rect 6181 7939 6193 7942
rect 6135 7933 6193 7939
rect 6546 7896 6552 7948
rect 6604 7936 6610 7948
rect 7377 7939 7435 7945
rect 7377 7936 7389 7939
rect 6604 7908 7389 7936
rect 6604 7896 6610 7908
rect 7377 7905 7389 7908
rect 7423 7905 7435 7939
rect 7377 7899 7435 7905
rect 7469 7939 7527 7945
rect 7469 7905 7481 7939
rect 7515 7936 7527 7939
rect 9306 7936 9312 7948
rect 7515 7908 9312 7936
rect 7515 7905 7527 7908
rect 7469 7899 7527 7905
rect 7282 7828 7288 7880
rect 7340 7828 7346 7880
rect 7392 7868 7420 7899
rect 9306 7896 9312 7908
rect 9364 7896 9370 7948
rect 9398 7896 9404 7948
rect 9456 7896 9462 7948
rect 11103 7939 11115 7973
rect 11149 7970 11161 7973
rect 11149 7942 11468 7970
rect 11514 7964 11520 8016
rect 11572 8004 11578 8016
rect 11885 8007 11943 8013
rect 11885 8004 11897 8007
rect 11572 7976 11897 8004
rect 11572 7964 11578 7976
rect 11885 7973 11897 7976
rect 11931 8004 11943 8007
rect 13265 8007 13323 8013
rect 13265 8004 13277 8007
rect 11931 7976 13277 8004
rect 11931 7973 11943 7976
rect 11885 7967 11943 7973
rect 13265 7973 13277 7976
rect 13311 7973 13323 8007
rect 13265 7967 13323 7973
rect 11149 7939 11161 7942
rect 11103 7933 11161 7939
rect 11440 7936 11468 7942
rect 11974 7936 11980 7948
rect 11440 7908 11980 7936
rect 11974 7896 11980 7908
rect 12032 7896 12038 7948
rect 12069 7939 12127 7945
rect 12069 7905 12081 7939
rect 12115 7936 12127 7939
rect 13722 7936 13728 7948
rect 12115 7908 13728 7936
rect 12115 7905 12127 7908
rect 12069 7899 12127 7905
rect 13722 7896 13728 7908
rect 13780 7896 13786 7948
rect 13817 7939 13875 7945
rect 13817 7905 13829 7939
rect 13863 7936 13875 7939
rect 14200 7936 14228 8044
rect 14458 8032 14464 8044
rect 14516 8032 14522 8084
rect 15838 8032 15844 8084
rect 15896 8072 15902 8084
rect 17497 8075 17555 8081
rect 17497 8072 17509 8075
rect 15896 8044 17509 8072
rect 15896 8032 15902 8044
rect 17497 8041 17509 8044
rect 17543 8041 17555 8075
rect 17497 8035 17555 8041
rect 17954 8032 17960 8084
rect 18012 8072 18018 8084
rect 18012 8044 19748 8072
rect 18012 8032 18018 8044
rect 16761 8007 16819 8013
rect 13863 7908 14228 7936
rect 15470 7930 15476 7982
rect 15528 7930 15534 7982
rect 16761 7973 16773 8007
rect 16807 8004 16819 8007
rect 19150 8004 19156 8016
rect 16807 7976 19156 8004
rect 16807 7973 16819 7976
rect 16761 7967 16819 7973
rect 19150 7964 19156 7976
rect 19208 7964 19214 8016
rect 16669 7939 16727 7945
rect 13863 7905 13875 7908
rect 13817 7899 13875 7905
rect 16669 7905 16681 7939
rect 16715 7936 16727 7939
rect 16715 7908 16896 7936
rect 16715 7905 16727 7908
rect 16669 7899 16727 7905
rect 7392 7840 8432 7868
rect 6822 7760 6828 7812
rect 6880 7800 6886 7812
rect 8404 7809 8432 7840
rect 8754 7828 8760 7880
rect 8812 7868 8818 7880
rect 9214 7868 9220 7880
rect 8812 7840 9220 7868
rect 8812 7828 8818 7840
rect 9214 7828 9220 7840
rect 9272 7828 9278 7880
rect 9766 7868 9772 7880
rect 9416 7840 9772 7868
rect 8297 7803 8355 7809
rect 8297 7800 8309 7803
rect 6880 7772 8309 7800
rect 6880 7760 6886 7772
rect 8297 7769 8309 7772
rect 8343 7769 8355 7803
rect 8297 7763 8355 7769
rect 8389 7803 8447 7809
rect 8389 7769 8401 7803
rect 8435 7769 8447 7803
rect 8389 7763 8447 7769
rect 7837 7735 7895 7741
rect 7837 7701 7849 7735
rect 7883 7732 7895 7735
rect 9416 7732 9444 7840
rect 9766 7828 9772 7840
rect 9824 7828 9830 7880
rect 12253 7871 12311 7877
rect 12253 7837 12265 7871
rect 12299 7868 12311 7871
rect 12618 7868 12624 7880
rect 12299 7840 12624 7868
rect 12299 7837 12311 7840
rect 12253 7831 12311 7837
rect 12618 7828 12624 7840
rect 12676 7828 12682 7880
rect 12710 7828 12716 7880
rect 12768 7868 12774 7880
rect 14182 7868 14188 7880
rect 12768 7840 14188 7868
rect 12768 7828 12774 7840
rect 14182 7828 14188 7840
rect 14240 7828 14246 7880
rect 11514 7760 11520 7812
rect 11572 7800 11578 7812
rect 11572 7772 12020 7800
rect 11572 7760 11578 7772
rect 7883 7704 9444 7732
rect 11992 7732 12020 7772
rect 12066 7760 12072 7812
rect 12124 7800 12130 7812
rect 12897 7803 12955 7809
rect 12897 7800 12909 7803
rect 12124 7772 12909 7800
rect 12124 7760 12130 7772
rect 12897 7769 12909 7772
rect 12943 7769 12955 7803
rect 16868 7800 16896 7908
rect 17126 7896 17132 7948
rect 17184 7936 17190 7948
rect 19242 7936 19248 7948
rect 17184 7908 19248 7936
rect 17184 7896 17190 7908
rect 19242 7896 19248 7908
rect 19300 7896 19306 7948
rect 16945 7871 17003 7877
rect 16945 7837 16957 7871
rect 16991 7868 17003 7871
rect 16991 7840 17908 7868
rect 16991 7837 17003 7840
rect 16945 7831 17003 7837
rect 17494 7800 17500 7812
rect 16868 7772 17500 7800
rect 12897 7763 12955 7769
rect 17494 7760 17500 7772
rect 17552 7760 17558 7812
rect 17586 7760 17592 7812
rect 17644 7760 17650 7812
rect 17880 7800 17908 7840
rect 17954 7828 17960 7880
rect 18012 7828 18018 7880
rect 18064 7840 18920 7868
rect 18064 7800 18092 7840
rect 17880 7772 18092 7800
rect 18506 7760 18512 7812
rect 18564 7760 18570 7812
rect 18598 7760 18604 7812
rect 18656 7760 18662 7812
rect 18892 7800 18920 7840
rect 18966 7828 18972 7880
rect 19024 7828 19030 7880
rect 19720 7868 19748 8044
rect 22186 8032 22192 8084
rect 22244 8072 22250 8084
rect 24210 8072 24216 8084
rect 22244 8044 24216 8072
rect 22244 8032 22250 8044
rect 24210 8032 24216 8044
rect 24268 8032 24274 8084
rect 25590 8032 25596 8084
rect 25648 8072 25654 8084
rect 25648 8044 25912 8072
rect 25648 8032 25654 8044
rect 22002 8004 22008 8016
rect 21591 7973 21649 7979
rect 19889 7939 19947 7945
rect 19889 7905 19901 7939
rect 19935 7936 19947 7939
rect 20254 7936 20260 7948
rect 19935 7908 20260 7936
rect 19935 7905 19947 7908
rect 19889 7899 19947 7905
rect 20254 7896 20260 7908
rect 20312 7896 20318 7948
rect 21591 7939 21603 7973
rect 21637 7970 21649 7973
rect 21928 7976 22008 8004
rect 21928 7970 21956 7976
rect 21637 7942 21956 7970
rect 22002 7964 22008 7976
rect 22060 7964 22066 8016
rect 22094 7964 22100 8016
rect 22152 8004 22158 8016
rect 22152 7976 23428 8004
rect 22152 7964 22158 7976
rect 21637 7939 21649 7942
rect 21591 7933 21649 7939
rect 22557 7939 22615 7945
rect 22557 7905 22569 7939
rect 22603 7936 22615 7939
rect 23290 7936 23296 7948
rect 22603 7908 23296 7936
rect 22603 7905 22615 7908
rect 22557 7899 22615 7905
rect 23290 7896 23296 7908
rect 23348 7896 23354 7948
rect 23400 7945 23428 7976
rect 23385 7939 23443 7945
rect 23385 7905 23397 7939
rect 23431 7905 23443 7939
rect 24578 7930 24584 7982
rect 24636 7930 24642 7982
rect 23385 7899 23443 7905
rect 20070 7868 20076 7880
rect 19720 7840 20076 7868
rect 20070 7828 20076 7840
rect 20128 7828 20134 7880
rect 22738 7828 22744 7880
rect 22796 7868 22802 7880
rect 23569 7871 23627 7877
rect 23569 7868 23581 7871
rect 22796 7840 23581 7868
rect 22796 7828 22802 7840
rect 23569 7837 23581 7840
rect 23615 7837 23627 7871
rect 25884 7868 25912 8044
rect 26878 8032 26884 8084
rect 26936 8032 26942 8084
rect 28534 8032 28540 8084
rect 28592 8032 28598 8084
rect 29178 7964 29184 8016
rect 29236 8004 29242 8016
rect 29236 7976 30420 8004
rect 29236 7964 29242 7976
rect 30392 7970 30420 7976
rect 30699 7973 30757 7979
rect 30699 7970 30711 7973
rect 26050 7896 26056 7948
rect 26108 7936 26114 7948
rect 26237 7939 26295 7945
rect 26237 7936 26249 7939
rect 26108 7908 26249 7936
rect 26108 7896 26114 7908
rect 26237 7905 26249 7908
rect 26283 7905 26295 7939
rect 26237 7899 26295 7905
rect 26970 7896 26976 7948
rect 27028 7936 27034 7948
rect 27985 7939 28043 7945
rect 30392 7942 30711 7970
rect 27985 7936 27997 7939
rect 27028 7908 27997 7936
rect 27028 7896 27034 7908
rect 27985 7905 27997 7908
rect 28031 7905 28043 7939
rect 30699 7939 30711 7942
rect 30745 7939 30757 7973
rect 30699 7933 30757 7939
rect 27985 7899 28043 7905
rect 32030 7896 32036 7948
rect 32088 7936 32094 7948
rect 32401 7939 32459 7945
rect 32401 7936 32413 7939
rect 32088 7908 32413 7936
rect 32088 7896 32094 7908
rect 32401 7905 32413 7908
rect 32447 7905 32459 7939
rect 32401 7899 32459 7905
rect 27525 7871 27583 7877
rect 27525 7868 27537 7871
rect 25884 7840 27537 7868
rect 23569 7831 23627 7837
rect 27525 7837 27537 7840
rect 27571 7868 27583 7871
rect 29914 7868 29920 7880
rect 27571 7840 29920 7868
rect 27571 7837 27583 7840
rect 27525 7831 27583 7837
rect 29914 7828 29920 7840
rect 29972 7828 29978 7880
rect 19886 7800 19892 7812
rect 18892 7772 19892 7800
rect 19886 7760 19892 7772
rect 19944 7760 19950 7812
rect 22462 7760 22468 7812
rect 22520 7800 22526 7812
rect 24118 7800 24124 7812
rect 22520 7772 24124 7800
rect 22520 7760 22526 7772
rect 24118 7760 24124 7772
rect 24176 7760 24182 7812
rect 26326 7760 26332 7812
rect 26384 7800 26390 7812
rect 29089 7803 29147 7809
rect 29089 7800 29101 7803
rect 26384 7772 29101 7800
rect 26384 7760 26390 7772
rect 29089 7769 29101 7772
rect 29135 7769 29147 7803
rect 29089 7763 29147 7769
rect 12434 7732 12440 7744
rect 11992 7704 12440 7732
rect 7883 7701 7895 7704
rect 7837 7695 7895 7701
rect 12434 7692 12440 7704
rect 12492 7692 12498 7744
rect 12526 7692 12532 7744
rect 12584 7732 12590 7744
rect 12805 7735 12863 7741
rect 12805 7732 12817 7735
rect 12584 7704 12817 7732
rect 12584 7692 12590 7704
rect 12805 7701 12817 7704
rect 12851 7701 12863 7735
rect 12805 7695 12863 7701
rect 13262 7692 13268 7744
rect 13320 7732 13326 7744
rect 13722 7732 13728 7744
rect 13320 7704 13728 7732
rect 13320 7692 13326 7704
rect 13722 7692 13728 7704
rect 13780 7692 13786 7744
rect 15930 7692 15936 7744
rect 15988 7732 15994 7744
rect 16301 7735 16359 7741
rect 16301 7732 16313 7735
rect 15988 7704 16313 7732
rect 15988 7692 15994 7704
rect 16301 7701 16313 7704
rect 16347 7732 16359 7735
rect 19702 7732 19708 7744
rect 16347 7704 19708 7732
rect 16347 7701 16359 7704
rect 16301 7695 16359 7701
rect 19702 7692 19708 7704
rect 19760 7692 19766 7744
rect 22370 7692 22376 7744
rect 22428 7692 22434 7744
rect 23198 7692 23204 7744
rect 23256 7692 23262 7744
rect 26234 7692 26240 7744
rect 26292 7732 26298 7744
rect 28258 7732 28264 7744
rect 26292 7704 28264 7732
rect 26292 7692 26298 7704
rect 28258 7692 28264 7704
rect 28316 7692 28322 7744
rect 1104 7642 33028 7664
rect 1104 7590 10950 7642
rect 11002 7590 11014 7642
rect 11066 7590 11078 7642
rect 11130 7590 11142 7642
rect 11194 7590 11206 7642
rect 11258 7590 20950 7642
rect 21002 7590 21014 7642
rect 21066 7590 21078 7642
rect 21130 7590 21142 7642
rect 21194 7590 21206 7642
rect 21258 7590 30950 7642
rect 31002 7590 31014 7642
rect 31066 7590 31078 7642
rect 31130 7590 31142 7642
rect 31194 7590 31206 7642
rect 31258 7590 33028 7642
rect 1104 7568 33028 7590
rect 1946 7488 1952 7540
rect 2004 7528 2010 7540
rect 4154 7528 4160 7540
rect 2004 7500 4160 7528
rect 2004 7488 2010 7500
rect 4154 7488 4160 7500
rect 4212 7488 4218 7540
rect 10226 7488 10232 7540
rect 10284 7528 10290 7540
rect 11422 7528 11428 7540
rect 10284 7500 11428 7528
rect 10284 7488 10290 7500
rect 11422 7488 11428 7500
rect 11480 7488 11486 7540
rect 11974 7488 11980 7540
rect 12032 7528 12038 7540
rect 12342 7528 12348 7540
rect 12032 7500 12348 7528
rect 12032 7488 12038 7500
rect 12342 7488 12348 7500
rect 12400 7488 12406 7540
rect 14458 7488 14464 7540
rect 14516 7528 14522 7540
rect 17126 7528 17132 7540
rect 14516 7500 17132 7528
rect 14516 7488 14522 7500
rect 17126 7488 17132 7500
rect 17184 7488 17190 7540
rect 19242 7488 19248 7540
rect 19300 7528 19306 7540
rect 22370 7528 22376 7540
rect 19300 7500 22376 7528
rect 19300 7488 19306 7500
rect 22370 7488 22376 7500
rect 22428 7488 22434 7540
rect 25130 7488 25136 7540
rect 25188 7488 25194 7540
rect 27062 7488 27068 7540
rect 27120 7488 27126 7540
rect 28169 7531 28227 7537
rect 28169 7528 28181 7531
rect 27172 7500 28181 7528
rect 1762 7420 1768 7472
rect 1820 7460 1826 7472
rect 4338 7460 4344 7472
rect 1820 7432 4344 7460
rect 1820 7420 1826 7432
rect 4338 7420 4344 7432
rect 4396 7420 4402 7472
rect 9766 7420 9772 7472
rect 9824 7460 9830 7472
rect 10413 7463 10471 7469
rect 10413 7460 10425 7463
rect 9824 7432 10425 7460
rect 9824 7420 9830 7432
rect 2682 7392 2688 7404
rect 1780 7364 2688 7392
rect 1780 7333 1808 7364
rect 2682 7352 2688 7364
rect 2740 7352 2746 7404
rect 3050 7352 3056 7404
rect 3108 7352 3114 7404
rect 6362 7352 6368 7404
rect 6420 7392 6426 7404
rect 6420 7364 7328 7392
rect 6420 7352 6426 7364
rect 1765 7327 1823 7333
rect 1765 7293 1777 7327
rect 1811 7293 1823 7327
rect 1765 7287 1823 7293
rect 1854 7284 1860 7336
rect 1912 7324 1918 7336
rect 2409 7327 2467 7333
rect 2409 7324 2421 7327
rect 1912 7296 2421 7324
rect 1912 7284 1918 7296
rect 2409 7293 2421 7296
rect 2455 7293 2467 7327
rect 2409 7287 2467 7293
rect 1949 7259 2007 7265
rect 1949 7225 1961 7259
rect 1995 7256 2007 7259
rect 2590 7256 2596 7268
rect 1995 7228 2596 7256
rect 1995 7225 2007 7228
rect 1949 7219 2007 7225
rect 2590 7216 2596 7228
rect 2648 7216 2654 7268
rect 5074 7250 5080 7302
rect 5132 7250 5138 7302
rect 6822 7284 6828 7336
rect 6880 7284 6886 7336
rect 7300 7333 7328 7364
rect 7285 7327 7343 7333
rect 7285 7293 7297 7327
rect 7331 7293 7343 7327
rect 9398 7324 9404 7336
rect 7285 7287 7343 7293
rect 9079 7293 9137 7299
rect 9079 7259 9091 7293
rect 9125 7290 9137 7293
rect 9370 7290 9404 7324
rect 9125 7284 9404 7290
rect 9456 7284 9462 7336
rect 10060 7324 10088 7432
rect 10413 7429 10425 7432
rect 10459 7429 10471 7463
rect 11514 7460 11520 7472
rect 10413 7423 10471 7429
rect 10520 7432 11520 7460
rect 10137 7395 10195 7401
rect 10137 7361 10149 7395
rect 10183 7392 10195 7395
rect 10520 7392 10548 7432
rect 10183 7364 10548 7392
rect 10183 7361 10195 7364
rect 10137 7355 10195 7361
rect 10594 7352 10600 7404
rect 10652 7352 10658 7404
rect 11256 7401 11284 7432
rect 11514 7420 11520 7432
rect 11572 7420 11578 7472
rect 14642 7420 14648 7472
rect 14700 7460 14706 7472
rect 17034 7460 17040 7472
rect 14700 7432 17040 7460
rect 14700 7420 14706 7432
rect 17034 7420 17040 7432
rect 17092 7420 17098 7472
rect 19610 7420 19616 7472
rect 19668 7420 19674 7472
rect 19702 7420 19708 7472
rect 19760 7420 19766 7472
rect 21453 7463 21511 7469
rect 21453 7460 21465 7463
rect 19812 7432 21465 7460
rect 11241 7395 11299 7401
rect 10704 7364 11146 7392
rect 10704 7324 10732 7364
rect 10060 7296 10732 7324
rect 11118 7334 11146 7364
rect 11241 7361 11253 7395
rect 11287 7361 11299 7395
rect 12710 7392 12716 7404
rect 11241 7355 11299 7361
rect 11624 7364 12716 7392
rect 11118 7326 11192 7334
rect 11118 7306 11284 7326
rect 11164 7298 11284 7306
rect 9125 7262 9398 7284
rect 9125 7259 9137 7262
rect 9079 7253 9137 7259
rect 11256 7256 11284 7298
rect 11333 7259 11391 7265
rect 11333 7256 11345 7259
rect 11256 7228 11345 7256
rect 11333 7225 11345 7228
rect 11379 7225 11391 7259
rect 11333 7219 11391 7225
rect 11425 7259 11483 7265
rect 11425 7225 11437 7259
rect 11471 7256 11483 7259
rect 11624 7256 11652 7364
rect 12710 7352 12716 7364
rect 12768 7352 12774 7404
rect 14921 7395 14979 7401
rect 14921 7361 14933 7395
rect 14967 7392 14979 7395
rect 14967 7364 17540 7392
rect 14967 7361 14979 7364
rect 14921 7355 14979 7361
rect 12158 7324 12164 7336
rect 11946 7318 12164 7324
rect 11762 7296 12164 7318
rect 11762 7290 11974 7296
rect 11762 7256 11790 7290
rect 12158 7284 12164 7296
rect 12216 7284 12222 7336
rect 12250 7284 12256 7336
rect 12308 7284 12314 7336
rect 11471 7228 11652 7256
rect 11716 7228 11790 7256
rect 13998 7250 14004 7302
rect 14056 7250 14062 7302
rect 14826 7284 14832 7336
rect 14884 7284 14890 7336
rect 15657 7327 15715 7333
rect 15657 7293 15669 7327
rect 15703 7324 15715 7327
rect 15933 7327 15991 7333
rect 15703 7296 15884 7324
rect 15703 7293 15715 7296
rect 15657 7287 15715 7293
rect 11471 7225 11483 7228
rect 11425 7219 11483 7225
rect 1578 7148 1584 7200
rect 1636 7148 1642 7200
rect 3694 7148 3700 7200
rect 3752 7188 3758 7200
rect 4430 7188 4436 7200
rect 3752 7160 4436 7188
rect 3752 7148 3758 7160
rect 4430 7148 4436 7160
rect 4488 7148 4494 7200
rect 9490 7148 9496 7200
rect 9548 7188 9554 7200
rect 11716 7188 11744 7228
rect 14366 7216 14372 7268
rect 14424 7256 14430 7268
rect 15562 7256 15568 7268
rect 14424 7228 15568 7256
rect 14424 7216 14430 7228
rect 15562 7216 15568 7228
rect 15620 7216 15626 7268
rect 15856 7256 15884 7296
rect 15933 7293 15945 7327
rect 15979 7324 15991 7327
rect 16574 7324 16580 7336
rect 15979 7296 16580 7324
rect 15979 7293 15991 7296
rect 15933 7287 15991 7293
rect 16574 7284 16580 7296
rect 16632 7284 16638 7336
rect 17126 7284 17132 7336
rect 17184 7284 17190 7336
rect 16758 7256 16764 7268
rect 15856 7228 16764 7256
rect 16758 7216 16764 7228
rect 16816 7216 16822 7268
rect 9548 7160 11744 7188
rect 11793 7191 11851 7197
rect 9548 7148 9554 7160
rect 11793 7157 11805 7191
rect 11839 7188 11851 7191
rect 11974 7188 11980 7200
rect 11839 7160 11980 7188
rect 11839 7157 11851 7160
rect 11793 7151 11851 7157
rect 11974 7148 11980 7160
rect 12032 7148 12038 7200
rect 17512 7188 17540 7364
rect 18782 7250 18788 7302
rect 18840 7250 18846 7302
rect 19150 7284 19156 7336
rect 19208 7324 19214 7336
rect 19812 7324 19840 7432
rect 21453 7429 21465 7432
rect 21499 7429 21511 7463
rect 22462 7460 22468 7472
rect 21453 7423 21511 7429
rect 21606 7432 22468 7460
rect 20070 7352 20076 7404
rect 20128 7352 20134 7404
rect 20806 7352 20812 7404
rect 20864 7392 20870 7404
rect 21361 7395 21419 7401
rect 21361 7392 21373 7395
rect 20864 7364 21373 7392
rect 20864 7352 20870 7364
rect 21361 7361 21373 7364
rect 21407 7361 21419 7395
rect 21361 7355 21419 7361
rect 19208 7296 19840 7324
rect 19208 7284 19214 7296
rect 20254 7284 20260 7336
rect 20312 7324 20318 7336
rect 20533 7327 20591 7333
rect 20533 7324 20545 7327
rect 20312 7296 20545 7324
rect 20312 7284 20318 7296
rect 20533 7293 20545 7296
rect 20579 7293 20591 7327
rect 20533 7287 20591 7293
rect 19242 7216 19248 7268
rect 19300 7256 19306 7268
rect 20622 7256 20628 7268
rect 19300 7228 20628 7256
rect 19300 7216 19306 7228
rect 20622 7216 20628 7228
rect 20680 7216 20686 7268
rect 21606 7256 21634 7432
rect 22462 7420 22468 7432
rect 22520 7420 22526 7472
rect 21821 7395 21879 7401
rect 21821 7361 21833 7395
rect 21867 7392 21879 7395
rect 22186 7392 22192 7404
rect 21867 7364 22192 7392
rect 21867 7361 21879 7364
rect 21821 7355 21879 7361
rect 22186 7352 22192 7364
rect 22244 7352 22250 7404
rect 24394 7352 24400 7404
rect 24452 7392 24458 7404
rect 26053 7395 26111 7401
rect 26053 7392 26065 7395
rect 24452 7364 26065 7392
rect 24452 7352 24458 7364
rect 26053 7361 26065 7364
rect 26099 7361 26111 7395
rect 27172 7392 27200 7500
rect 28169 7497 28181 7500
rect 28215 7497 28227 7531
rect 28169 7491 28227 7497
rect 28258 7488 28264 7540
rect 28316 7528 28322 7540
rect 30929 7531 30987 7537
rect 30929 7528 30941 7531
rect 28316 7500 30941 7528
rect 28316 7488 28322 7500
rect 30929 7497 30941 7500
rect 30975 7497 30987 7531
rect 30929 7491 30987 7497
rect 26053 7355 26111 7361
rect 26160 7364 27200 7392
rect 21744 7320 22600 7324
rect 20732 7228 21634 7256
rect 21698 7296 22600 7320
rect 21698 7292 21772 7296
rect 17770 7188 17776 7200
rect 17512 7160 17776 7188
rect 17770 7148 17776 7160
rect 17828 7148 17834 7200
rect 19150 7148 19156 7200
rect 19208 7188 19214 7200
rect 20732 7197 20760 7228
rect 20717 7191 20775 7197
rect 20717 7188 20729 7191
rect 19208 7160 20729 7188
rect 19208 7148 19214 7160
rect 20717 7157 20729 7160
rect 20763 7157 20775 7191
rect 20717 7151 20775 7157
rect 20806 7148 20812 7200
rect 20864 7188 20870 7200
rect 21698 7188 21726 7292
rect 22572 7290 22600 7296
rect 22879 7293 22937 7299
rect 22879 7290 22891 7293
rect 22572 7262 22891 7290
rect 22879 7259 22891 7262
rect 22925 7259 22937 7293
rect 24210 7284 24216 7336
rect 24268 7324 24274 7336
rect 24581 7327 24639 7333
rect 24581 7324 24593 7327
rect 24268 7296 24593 7324
rect 24268 7284 24274 7296
rect 24581 7293 24593 7296
rect 24627 7293 24639 7327
rect 24581 7287 24639 7293
rect 25317 7327 25375 7333
rect 25317 7293 25329 7327
rect 25363 7293 25375 7327
rect 25317 7287 25375 7293
rect 22879 7253 22937 7259
rect 25332 7256 25360 7287
rect 25406 7284 25412 7336
rect 25464 7284 25470 7336
rect 25682 7284 25688 7336
rect 25740 7324 25746 7336
rect 26160 7333 26188 7364
rect 27614 7352 27620 7404
rect 27672 7352 27678 7404
rect 26145 7327 26203 7333
rect 26145 7324 26157 7327
rect 25740 7296 26157 7324
rect 25740 7284 25746 7296
rect 26145 7293 26157 7296
rect 26191 7293 26203 7327
rect 26145 7287 26203 7293
rect 26234 7284 26240 7336
rect 26292 7324 26298 7336
rect 29825 7327 29883 7333
rect 29825 7324 29837 7327
rect 26292 7296 29837 7324
rect 26292 7284 26298 7296
rect 29825 7293 29837 7296
rect 29871 7293 29883 7327
rect 29825 7287 29883 7293
rect 28350 7256 28356 7268
rect 25332 7228 28356 7256
rect 28350 7216 28356 7228
rect 28408 7216 28414 7268
rect 30377 7259 30435 7265
rect 30377 7256 30389 7259
rect 28460 7228 30389 7256
rect 20864 7160 21726 7188
rect 20864 7148 20870 7160
rect 24762 7148 24768 7200
rect 24820 7188 24826 7200
rect 28460 7188 28488 7228
rect 30377 7225 30389 7228
rect 30423 7225 30435 7259
rect 30377 7219 30435 7225
rect 24820 7160 28488 7188
rect 24820 7148 24826 7160
rect 28534 7148 28540 7200
rect 28592 7188 28598 7200
rect 28721 7191 28779 7197
rect 28721 7188 28733 7191
rect 28592 7160 28733 7188
rect 28592 7148 28598 7160
rect 28721 7157 28733 7160
rect 28767 7157 28779 7191
rect 28721 7151 28779 7157
rect 28810 7148 28816 7200
rect 28868 7188 28874 7200
rect 29273 7191 29331 7197
rect 29273 7188 29285 7191
rect 28868 7160 29285 7188
rect 28868 7148 28874 7160
rect 29273 7157 29285 7160
rect 29319 7157 29331 7191
rect 29273 7151 29331 7157
rect 1104 7098 33028 7120
rect 1104 7046 11610 7098
rect 11662 7046 11674 7098
rect 11726 7046 11738 7098
rect 11790 7046 11802 7098
rect 11854 7046 11866 7098
rect 11918 7046 21610 7098
rect 21662 7046 21674 7098
rect 21726 7046 21738 7098
rect 21790 7046 21802 7098
rect 21854 7046 21866 7098
rect 21918 7046 31610 7098
rect 31662 7046 31674 7098
rect 31726 7046 31738 7098
rect 31790 7046 31802 7098
rect 31854 7046 31866 7098
rect 31918 7046 33028 7098
rect 1104 7024 33028 7046
rect 2038 6944 2044 6996
rect 2096 6984 2102 6996
rect 2409 6987 2467 6993
rect 2409 6984 2421 6987
rect 2096 6956 2421 6984
rect 2096 6944 2102 6956
rect 2409 6953 2421 6956
rect 2455 6953 2467 6987
rect 2409 6947 2467 6953
rect 3973 6987 4031 6993
rect 3973 6953 3985 6987
rect 4019 6984 4031 6987
rect 4062 6984 4068 6996
rect 4019 6956 4068 6984
rect 4019 6953 4031 6956
rect 3973 6947 4031 6953
rect 4062 6944 4068 6956
rect 4120 6944 4126 6996
rect 9214 6944 9220 6996
rect 9272 6984 9278 6996
rect 10134 6984 10140 6996
rect 9272 6956 10140 6984
rect 9272 6944 9278 6956
rect 10134 6944 10140 6956
rect 10192 6944 10198 6996
rect 11514 6944 11520 6996
rect 11572 6984 11578 6996
rect 11572 6956 11836 6984
rect 11572 6944 11578 6956
rect 3605 6919 3663 6925
rect 3605 6885 3617 6919
rect 3651 6916 3663 6919
rect 4430 6916 4436 6928
rect 3651 6888 4436 6916
rect 3651 6885 3663 6888
rect 3605 6879 3663 6885
rect 4430 6876 4436 6888
rect 4488 6876 4494 6928
rect 2317 6851 2375 6857
rect 2317 6817 2329 6851
rect 2363 6848 2375 6851
rect 4246 6848 4252 6860
rect 2363 6820 4252 6848
rect 2363 6817 2375 6820
rect 2317 6811 2375 6817
rect 4246 6808 4252 6820
rect 4304 6808 4310 6860
rect 4338 6808 4344 6860
rect 4396 6808 4402 6860
rect 4798 6842 4804 6894
rect 4856 6842 4862 6894
rect 6546 6808 6552 6860
rect 6604 6808 6610 6860
rect 7101 6851 7159 6857
rect 7101 6817 7113 6851
rect 7147 6817 7159 6851
rect 8846 6842 8852 6894
rect 8904 6842 8910 6894
rect 10459 6885 10517 6891
rect 10459 6882 10471 6885
rect 7101 6811 7159 6817
rect 2225 6783 2283 6789
rect 2225 6749 2237 6783
rect 2271 6749 2283 6783
rect 2225 6743 2283 6749
rect 2240 6712 2268 6743
rect 3418 6740 3424 6792
rect 3476 6740 3482 6792
rect 3513 6783 3571 6789
rect 3513 6749 3525 6783
rect 3559 6780 3571 6783
rect 4356 6780 4384 6808
rect 3559 6752 4384 6780
rect 3559 6749 3571 6752
rect 3513 6743 3571 6749
rect 6086 6740 6092 6792
rect 6144 6780 6150 6792
rect 7116 6780 7144 6811
rect 9306 6808 9312 6860
rect 9364 6848 9370 6860
rect 10152 6854 10471 6882
rect 10152 6848 10180 6854
rect 9364 6820 10180 6848
rect 10459 6851 10471 6854
rect 10505 6851 10517 6885
rect 10459 6845 10517 6851
rect 9364 6808 9370 6820
rect 6144 6752 7144 6780
rect 11808 6780 11836 6956
rect 17586 6944 17592 6996
rect 17644 6984 17650 6996
rect 19150 6984 19156 6996
rect 17644 6956 17954 6984
rect 17644 6944 17650 6956
rect 12253 6851 12311 6857
rect 12253 6817 12265 6851
rect 12299 6848 12311 6851
rect 12342 6848 12348 6860
rect 12299 6820 12348 6848
rect 12299 6817 12311 6820
rect 12253 6811 12311 6817
rect 12342 6808 12348 6820
rect 12400 6808 12406 6860
rect 12897 6851 12955 6857
rect 12897 6817 12909 6851
rect 12943 6848 12955 6851
rect 12986 6848 12992 6860
rect 12943 6820 12992 6848
rect 12943 6817 12955 6820
rect 12897 6811 12955 6817
rect 12986 6808 12992 6820
rect 13044 6808 13050 6860
rect 14550 6842 14556 6894
rect 14608 6842 14614 6894
rect 15470 6808 15476 6860
rect 15528 6808 15534 6860
rect 17126 6842 17132 6894
rect 17184 6842 17190 6894
rect 13078 6780 13084 6792
rect 11808 6752 13084 6780
rect 6144 6740 6150 6752
rect 13078 6740 13084 6752
rect 13136 6740 13142 6792
rect 17926 6780 17954 6956
rect 18984 6956 19156 6984
rect 18601 6851 18659 6857
rect 18601 6817 18613 6851
rect 18647 6848 18659 6851
rect 18782 6848 18788 6860
rect 18647 6820 18788 6848
rect 18647 6817 18659 6820
rect 18601 6811 18659 6817
rect 18782 6808 18788 6820
rect 18840 6808 18846 6860
rect 18984 6780 19012 6956
rect 19150 6944 19156 6956
rect 19208 6944 19214 6996
rect 23290 6944 23296 6996
rect 23348 6984 23354 6996
rect 25133 6987 25191 6993
rect 25133 6984 25145 6987
rect 23348 6956 25145 6984
rect 23348 6944 23354 6956
rect 25133 6953 25145 6956
rect 25179 6953 25191 6987
rect 28810 6984 28816 6996
rect 25133 6947 25191 6953
rect 27586 6956 28816 6984
rect 20303 6885 20361 6891
rect 20303 6851 20315 6885
rect 20349 6882 20361 6885
rect 20349 6854 20668 6882
rect 20349 6851 20361 6854
rect 20303 6845 20361 6851
rect 20640 6848 20668 6854
rect 21085 6851 21143 6857
rect 21085 6848 21097 6851
rect 20640 6820 21097 6848
rect 21085 6817 21097 6820
rect 21131 6817 21143 6851
rect 22830 6842 22836 6894
rect 22888 6842 22894 6894
rect 24118 6876 24124 6928
rect 24176 6916 24182 6928
rect 24213 6919 24271 6925
rect 24213 6916 24225 6919
rect 24176 6888 24225 6916
rect 24176 6876 24182 6888
rect 24213 6885 24225 6888
rect 24259 6916 24271 6919
rect 27433 6919 27491 6925
rect 27433 6916 27445 6919
rect 24259 6888 27445 6916
rect 24259 6885 24271 6888
rect 24213 6879 24271 6885
rect 27433 6885 27445 6888
rect 27479 6916 27491 6919
rect 27586 6916 27614 6956
rect 28810 6944 28816 6956
rect 28868 6944 28874 6996
rect 29914 6944 29920 6996
rect 29972 6944 29978 6996
rect 27479 6888 27614 6916
rect 27479 6885 27491 6888
rect 27433 6879 27491 6885
rect 24397 6851 24455 6857
rect 21085 6811 21143 6817
rect 24397 6817 24409 6851
rect 24443 6817 24455 6851
rect 24397 6811 24455 6817
rect 17926 6752 19012 6780
rect 23290 6740 23296 6792
rect 23348 6780 23354 6792
rect 24412 6780 24440 6811
rect 25222 6808 25228 6860
rect 25280 6808 25286 6860
rect 25866 6808 25872 6860
rect 25924 6848 25930 6860
rect 28537 6851 28595 6857
rect 28537 6848 28549 6851
rect 25924 6820 28549 6848
rect 25924 6808 25930 6820
rect 28537 6817 28549 6820
rect 28583 6817 28595 6851
rect 28537 6811 28595 6817
rect 23348 6752 24440 6780
rect 24581 6783 24639 6789
rect 23348 6740 23354 6752
rect 24581 6749 24593 6783
rect 24627 6780 24639 6783
rect 24762 6780 24768 6792
rect 24627 6752 24768 6780
rect 24627 6749 24639 6752
rect 24581 6743 24639 6749
rect 24762 6740 24768 6752
rect 24820 6740 24826 6792
rect 25240 6780 25268 6808
rect 27985 6783 28043 6789
rect 27985 6780 27997 6783
rect 25240 6752 27997 6780
rect 27985 6749 27997 6752
rect 28031 6749 28043 6783
rect 27985 6743 28043 6749
rect 4338 6712 4344 6724
rect 2240 6684 4344 6712
rect 4338 6672 4344 6684
rect 4396 6672 4402 6724
rect 26326 6672 26332 6724
rect 26384 6672 26390 6724
rect 29086 6672 29092 6724
rect 29144 6712 29150 6724
rect 32030 6712 32036 6724
rect 29144 6684 32036 6712
rect 29144 6672 29150 6684
rect 32030 6672 32036 6684
rect 32088 6672 32094 6724
rect 2777 6647 2835 6653
rect 2777 6613 2789 6647
rect 2823 6644 2835 6647
rect 3878 6644 3884 6656
rect 2823 6616 3884 6644
rect 2823 6613 2835 6616
rect 2777 6607 2835 6613
rect 3878 6604 3884 6616
rect 3936 6604 3942 6656
rect 24854 6604 24860 6656
rect 24912 6644 24918 6656
rect 25777 6647 25835 6653
rect 25777 6644 25789 6647
rect 24912 6616 25789 6644
rect 24912 6604 24918 6616
rect 25777 6613 25789 6616
rect 25823 6613 25835 6647
rect 25777 6607 25835 6613
rect 26878 6604 26884 6656
rect 26936 6604 26942 6656
rect 1104 6554 33028 6576
rect 1104 6502 10950 6554
rect 11002 6502 11014 6554
rect 11066 6502 11078 6554
rect 11130 6502 11142 6554
rect 11194 6502 11206 6554
rect 11258 6502 20950 6554
rect 21002 6502 21014 6554
rect 21066 6502 21078 6554
rect 21130 6502 21142 6554
rect 21194 6502 21206 6554
rect 21258 6502 30950 6554
rect 31002 6502 31014 6554
rect 31066 6502 31078 6554
rect 31130 6502 31142 6554
rect 31194 6502 31206 6554
rect 31258 6502 33028 6554
rect 1104 6480 33028 6502
rect 4062 6440 4068 6452
rect 2746 6412 4068 6440
rect 2501 6375 2559 6381
rect 2501 6341 2513 6375
rect 2547 6372 2559 6375
rect 2746 6372 2774 6412
rect 4062 6400 4068 6412
rect 4120 6400 4126 6452
rect 16942 6400 16948 6452
rect 17000 6440 17006 6452
rect 17862 6440 17868 6452
rect 17000 6412 17868 6440
rect 17000 6400 17006 6412
rect 17862 6400 17868 6412
rect 17920 6400 17926 6452
rect 20162 6400 20168 6452
rect 20220 6440 20226 6452
rect 20625 6443 20683 6449
rect 20625 6440 20637 6443
rect 20220 6412 20637 6440
rect 20220 6400 20226 6412
rect 20625 6409 20637 6412
rect 20671 6409 20683 6443
rect 20625 6403 20683 6409
rect 30650 6400 30656 6452
rect 30708 6400 30714 6452
rect 4154 6372 4160 6384
rect 2547 6344 2774 6372
rect 3528 6344 4160 6372
rect 2547 6341 2559 6344
rect 2501 6335 2559 6341
rect 1949 6307 2007 6313
rect 1949 6273 1961 6307
rect 1995 6304 2007 6307
rect 3528 6304 3556 6344
rect 4154 6332 4160 6344
rect 4212 6332 4218 6384
rect 15194 6332 15200 6384
rect 15252 6372 15258 6384
rect 15749 6375 15807 6381
rect 15749 6372 15761 6375
rect 15252 6344 15761 6372
rect 15252 6332 15258 6344
rect 15749 6341 15761 6344
rect 15795 6341 15807 6375
rect 15749 6335 15807 6341
rect 16574 6332 16580 6384
rect 16632 6372 16638 6384
rect 16669 6375 16727 6381
rect 16669 6372 16681 6375
rect 16632 6344 16681 6372
rect 16632 6332 16638 6344
rect 16669 6341 16681 6344
rect 16715 6341 16727 6375
rect 16669 6335 16727 6341
rect 16758 6332 16764 6384
rect 16816 6372 16822 6384
rect 18046 6372 18052 6384
rect 16816 6344 18052 6372
rect 16816 6332 16822 6344
rect 18046 6332 18052 6344
rect 18104 6332 18110 6384
rect 1995 6276 3556 6304
rect 3605 6307 3663 6313
rect 1995 6273 2007 6276
rect 1949 6267 2007 6273
rect 3605 6273 3617 6307
rect 3651 6273 3663 6307
rect 3605 6267 3663 6273
rect 2130 6196 2136 6248
rect 2188 6196 2194 6248
rect 3620 6236 3648 6267
rect 12618 6264 12624 6316
rect 12676 6304 12682 6316
rect 13446 6304 13452 6316
rect 12676 6276 13452 6304
rect 12676 6264 12682 6276
rect 13446 6264 13452 6276
rect 13504 6264 13510 6316
rect 15286 6264 15292 6316
rect 15344 6304 15350 6316
rect 15344 6276 16804 6304
rect 15344 6264 15350 6276
rect 4246 6236 4252 6248
rect 3620 6208 4252 6236
rect 4246 6196 4252 6208
rect 4304 6196 4310 6248
rect 6365 6239 6423 6245
rect 2041 6171 2099 6177
rect 2041 6137 2053 6171
rect 2087 6168 2099 6171
rect 3878 6168 3884 6180
rect 2087 6140 3884 6168
rect 2087 6137 2099 6140
rect 2041 6131 2099 6137
rect 3878 6128 3884 6140
rect 3936 6128 3942 6180
rect 4614 6162 4620 6214
rect 4672 6162 4678 6214
rect 6365 6205 6377 6239
rect 6411 6236 6423 6239
rect 6822 6236 6828 6248
rect 6411 6208 6828 6236
rect 6411 6205 6423 6208
rect 6365 6199 6423 6205
rect 6822 6196 6828 6208
rect 6880 6196 6886 6248
rect 6914 6196 6920 6248
rect 6972 6236 6978 6248
rect 7285 6239 7343 6245
rect 7285 6236 7297 6239
rect 6972 6208 7297 6236
rect 6972 6196 6978 6208
rect 7285 6205 7297 6208
rect 7331 6205 7343 6239
rect 10413 6239 10471 6245
rect 10413 6236 10425 6239
rect 7285 6199 7343 6205
rect 9079 6205 9137 6211
rect 9079 6171 9091 6205
rect 9125 6202 9137 6205
rect 9370 6208 10425 6236
rect 9370 6202 9398 6208
rect 9125 6174 9398 6202
rect 10413 6205 10425 6208
rect 10459 6205 10471 6239
rect 13081 6239 13139 6245
rect 10413 6199 10471 6205
rect 12207 6205 12265 6211
rect 9125 6171 9137 6174
rect 9079 6165 9137 6171
rect 12207 6171 12219 6205
rect 12253 6202 12265 6205
rect 13081 6205 13093 6239
rect 13127 6236 13139 6239
rect 13127 6208 13492 6236
rect 13127 6205 13139 6208
rect 12253 6174 12572 6202
rect 13081 6199 13139 6205
rect 12253 6171 12265 6174
rect 12207 6165 12265 6171
rect 12544 6168 12572 6174
rect 12802 6168 12808 6180
rect 12544 6140 12808 6168
rect 12802 6128 12808 6140
rect 12860 6128 12866 6180
rect 2682 6060 2688 6112
rect 2740 6100 2746 6112
rect 2961 6103 3019 6109
rect 2961 6100 2973 6103
rect 2740 6072 2973 6100
rect 2740 6060 2746 6072
rect 2961 6069 2973 6072
rect 3007 6069 3019 6103
rect 2961 6063 3019 6069
rect 3326 6060 3332 6112
rect 3384 6060 3390 6112
rect 3421 6103 3479 6109
rect 3421 6069 3433 6103
rect 3467 6100 3479 6103
rect 3970 6100 3976 6112
rect 3467 6072 3976 6100
rect 3467 6069 3479 6072
rect 3421 6063 3479 6069
rect 3970 6060 3976 6072
rect 4028 6060 4034 6112
rect 9398 6060 9404 6112
rect 9456 6100 9462 6112
rect 10318 6100 10324 6112
rect 9456 6072 10324 6100
rect 9456 6060 9462 6072
rect 10318 6060 10324 6072
rect 10376 6060 10382 6112
rect 13464 6100 13492 6208
rect 14783 6205 14841 6211
rect 14783 6171 14795 6205
rect 14829 6202 14841 6205
rect 14829 6174 15148 6202
rect 15378 6196 15384 6248
rect 15436 6236 15442 6248
rect 16117 6239 16175 6245
rect 16117 6236 16129 6239
rect 15436 6208 16129 6236
rect 15436 6196 15442 6208
rect 16117 6205 16129 6208
rect 16163 6205 16175 6239
rect 16776 6236 16804 6276
rect 27154 6264 27160 6316
rect 27212 6304 27218 6316
rect 28534 6304 28540 6316
rect 27212 6276 28540 6304
rect 27212 6264 27218 6276
rect 28534 6264 28540 6276
rect 28592 6264 28598 6316
rect 17037 6239 17095 6245
rect 17037 6236 17049 6239
rect 16776 6208 17049 6236
rect 16117 6199 16175 6205
rect 17037 6205 17049 6208
rect 17083 6236 17095 6239
rect 17862 6236 17868 6248
rect 17083 6208 17868 6236
rect 17083 6205 17095 6208
rect 17037 6199 17095 6205
rect 17862 6196 17868 6208
rect 17920 6196 17926 6248
rect 17954 6196 17960 6248
rect 18012 6196 18018 6248
rect 14829 6171 14841 6174
rect 14783 6165 14841 6171
rect 15120 6168 15148 6174
rect 15838 6168 15844 6180
rect 15120 6140 15844 6168
rect 15838 6128 15844 6140
rect 15896 6128 15902 6180
rect 19702 6162 19708 6214
rect 19760 6162 19766 6214
rect 20714 6196 20720 6248
rect 20772 6196 20778 6248
rect 21453 6239 21511 6245
rect 21453 6205 21465 6239
rect 21499 6236 21511 6239
rect 24210 6236 24216 6248
rect 21499 6208 21864 6236
rect 21499 6205 21511 6208
rect 21453 6199 21511 6205
rect 13722 6100 13728 6112
rect 13464 6072 13728 6100
rect 13722 6060 13728 6072
rect 13780 6060 13786 6112
rect 15654 6060 15660 6112
rect 15712 6060 15718 6112
rect 16574 6060 16580 6112
rect 16632 6060 16638 6112
rect 21836 6100 21864 6208
rect 23155 6205 23213 6211
rect 23155 6171 23167 6205
rect 23201 6202 23213 6205
rect 23492 6208 24216 6236
rect 23492 6202 23520 6208
rect 23201 6174 23520 6202
rect 24210 6196 24216 6208
rect 24268 6196 24274 6248
rect 24302 6196 24308 6248
rect 24360 6236 24366 6248
rect 24397 6239 24455 6245
rect 24397 6236 24409 6239
rect 24360 6208 24409 6236
rect 24360 6196 24366 6208
rect 24397 6205 24409 6208
rect 24443 6205 24455 6239
rect 24397 6199 24455 6205
rect 26191 6205 26249 6211
rect 23201 6171 23213 6174
rect 23155 6165 23213 6171
rect 26191 6171 26203 6205
rect 26237 6202 26249 6205
rect 26237 6174 26556 6202
rect 27614 6196 27620 6248
rect 27672 6236 27678 6248
rect 28077 6239 28135 6245
rect 28077 6236 28089 6239
rect 27672 6208 28089 6236
rect 27672 6196 27678 6208
rect 28077 6205 28089 6208
rect 28123 6205 28135 6239
rect 28077 6199 28135 6205
rect 26237 6171 26249 6174
rect 26191 6165 26249 6171
rect 26528 6168 26556 6174
rect 26786 6168 26792 6180
rect 26528 6140 26792 6168
rect 26786 6128 26792 6140
rect 26844 6128 26850 6180
rect 29822 6162 29828 6214
rect 29880 6162 29886 6214
rect 22002 6100 22008 6112
rect 21836 6072 22008 6100
rect 22002 6060 22008 6072
rect 22060 6060 22066 6112
rect 1104 6010 33028 6032
rect 1104 5958 11610 6010
rect 11662 5958 11674 6010
rect 11726 5958 11738 6010
rect 11790 5958 11802 6010
rect 11854 5958 11866 6010
rect 11918 5958 21610 6010
rect 21662 5958 21674 6010
rect 21726 5958 21738 6010
rect 21790 5958 21802 6010
rect 21854 5958 21866 6010
rect 21918 5958 31610 6010
rect 31662 5958 31674 6010
rect 31726 5958 31738 6010
rect 31790 5958 31802 6010
rect 31854 5958 31866 6010
rect 31918 5958 33028 6010
rect 1104 5936 33028 5958
rect 3602 5856 3608 5908
rect 3660 5856 3666 5908
rect 3970 5856 3976 5908
rect 4028 5856 4034 5908
rect 2406 5720 2412 5772
rect 2464 5720 2470 5772
rect 4338 5760 4344 5772
rect 2746 5732 4344 5760
rect 2222 5652 2228 5704
rect 2280 5652 2286 5704
rect 2317 5695 2375 5701
rect 2317 5661 2329 5695
rect 2363 5661 2375 5695
rect 2317 5655 2375 5661
rect 2332 5624 2360 5655
rect 2746 5624 2774 5732
rect 4338 5720 4344 5732
rect 4396 5720 4402 5772
rect 4798 5754 4804 5806
rect 4856 5754 4862 5806
rect 9079 5797 9137 5803
rect 6549 5763 6607 5769
rect 6549 5729 6561 5763
rect 6595 5760 6607 5763
rect 7190 5760 7196 5772
rect 6595 5732 7196 5760
rect 6595 5729 6607 5732
rect 6549 5723 6607 5729
rect 7190 5720 7196 5732
rect 7248 5720 7254 5772
rect 7285 5763 7343 5769
rect 7285 5729 7297 5763
rect 7331 5729 7343 5763
rect 9079 5763 9091 5797
rect 9125 5794 9137 5797
rect 11931 5797 11989 5803
rect 9125 5766 9398 5794
rect 9125 5763 9137 5766
rect 9079 5757 9137 5763
rect 9370 5760 9398 5766
rect 9490 5760 9496 5772
rect 9370 5732 9496 5760
rect 7285 5723 7343 5729
rect 3421 5695 3479 5701
rect 3421 5661 3433 5695
rect 3467 5661 3479 5695
rect 3421 5655 3479 5661
rect 3513 5695 3571 5701
rect 3513 5661 3525 5695
rect 3559 5692 3571 5695
rect 4154 5692 4160 5704
rect 3559 5664 4160 5692
rect 3559 5661 3571 5664
rect 3513 5655 3571 5661
rect 2332 5596 2774 5624
rect 3436 5624 3464 5655
rect 4154 5652 4160 5664
rect 4212 5652 4218 5704
rect 6086 5652 6092 5704
rect 6144 5692 6150 5704
rect 7300 5692 7328 5723
rect 9490 5720 9496 5732
rect 9548 5720 9554 5772
rect 10229 5763 10287 5769
rect 10229 5729 10241 5763
rect 10275 5760 10287 5763
rect 10502 5760 10508 5772
rect 10275 5732 10508 5760
rect 10275 5729 10287 5732
rect 10229 5723 10287 5729
rect 10502 5720 10508 5732
rect 10560 5720 10566 5772
rect 11931 5763 11943 5797
rect 11977 5794 11989 5797
rect 11977 5772 12296 5794
rect 11977 5766 12256 5772
rect 11977 5763 11989 5766
rect 11931 5757 11989 5763
rect 12250 5720 12256 5766
rect 12308 5720 12314 5772
rect 12802 5720 12808 5772
rect 12860 5720 12866 5772
rect 14550 5754 14556 5806
rect 14608 5754 14614 5806
rect 17635 5797 17693 5803
rect 15838 5720 15844 5772
rect 15896 5720 15902 5772
rect 17635 5763 17647 5797
rect 17681 5794 17693 5797
rect 17954 5794 17960 5840
rect 17681 5788 17960 5794
rect 18012 5788 18018 5840
rect 21223 5797 21281 5803
rect 17681 5766 18000 5788
rect 17681 5763 17693 5766
rect 17635 5757 17693 5763
rect 18046 5720 18052 5772
rect 18104 5760 18110 5772
rect 18509 5763 18567 5769
rect 18509 5760 18521 5763
rect 18104 5732 18521 5760
rect 18104 5720 18110 5732
rect 18509 5729 18521 5732
rect 18555 5729 18567 5763
rect 18509 5723 18567 5729
rect 19521 5763 19579 5769
rect 19521 5729 19533 5763
rect 19567 5760 19579 5763
rect 19702 5760 19708 5772
rect 19567 5732 19708 5760
rect 19567 5729 19579 5732
rect 19521 5723 19579 5729
rect 19702 5720 19708 5732
rect 19760 5720 19766 5772
rect 21223 5763 21235 5797
rect 21269 5794 21281 5797
rect 21450 5794 21456 5806
rect 21269 5766 21456 5794
rect 21269 5763 21281 5766
rect 21223 5757 21281 5763
rect 21450 5754 21456 5766
rect 21508 5754 21514 5806
rect 22462 5720 22468 5772
rect 22520 5720 22526 5772
rect 23106 5720 23112 5772
rect 23164 5720 23170 5772
rect 23198 5720 23204 5772
rect 23256 5720 23262 5772
rect 23474 5720 23480 5772
rect 23532 5760 23538 5772
rect 24213 5763 24271 5769
rect 24213 5760 24225 5763
rect 23532 5732 24225 5760
rect 23532 5720 23538 5732
rect 24213 5729 24225 5732
rect 24259 5729 24271 5763
rect 25958 5754 25964 5806
rect 26016 5754 26022 5806
rect 28583 5797 28641 5803
rect 24213 5723 24271 5729
rect 26786 5720 26792 5772
rect 26844 5720 26850 5772
rect 28583 5763 28595 5797
rect 28629 5794 28641 5797
rect 31711 5797 31769 5803
rect 28629 5772 28948 5794
rect 28629 5766 28908 5772
rect 28629 5763 28641 5766
rect 28583 5757 28641 5763
rect 28902 5720 28908 5766
rect 28960 5720 28966 5772
rect 29822 5720 29828 5772
rect 29880 5760 29886 5772
rect 29917 5763 29975 5769
rect 29917 5760 29929 5763
rect 29880 5732 29929 5760
rect 29880 5720 29886 5732
rect 29917 5729 29929 5732
rect 29963 5729 29975 5763
rect 31711 5763 31723 5797
rect 31757 5794 31769 5797
rect 32030 5794 32036 5840
rect 31757 5788 32036 5794
rect 32088 5788 32094 5840
rect 31757 5766 32076 5788
rect 31757 5763 31769 5766
rect 31711 5757 31769 5763
rect 29917 5723 29975 5729
rect 6144 5664 7328 5692
rect 6144 5652 6150 5664
rect 18690 5652 18696 5704
rect 18748 5692 18754 5704
rect 19886 5692 19892 5704
rect 18748 5664 19892 5692
rect 18748 5652 18754 5664
rect 19886 5652 19892 5664
rect 19944 5652 19950 5704
rect 22281 5695 22339 5701
rect 22281 5661 22293 5695
rect 22327 5692 22339 5695
rect 22738 5692 22744 5704
rect 22327 5664 22744 5692
rect 22327 5661 22339 5664
rect 22281 5655 22339 5661
rect 22738 5652 22744 5664
rect 22796 5652 22802 5704
rect 3694 5624 3700 5636
rect 3436 5596 3700 5624
rect 3694 5584 3700 5596
rect 3752 5584 3758 5636
rect 4246 5624 4252 5636
rect 3896 5596 4252 5624
rect 2777 5559 2835 5565
rect 2777 5525 2789 5559
rect 2823 5556 2835 5559
rect 3896 5556 3924 5596
rect 4246 5584 4252 5596
rect 4304 5584 4310 5636
rect 22002 5584 22008 5636
rect 22060 5624 22066 5636
rect 22925 5627 22983 5633
rect 22925 5624 22937 5627
rect 22060 5596 22937 5624
rect 22060 5584 22066 5596
rect 22925 5593 22937 5596
rect 22971 5593 22983 5627
rect 22925 5587 22983 5593
rect 2823 5528 3924 5556
rect 2823 5525 2835 5528
rect 2777 5519 2835 5525
rect 6454 5516 6460 5568
rect 6512 5556 6518 5568
rect 7374 5556 7380 5568
rect 6512 5528 7380 5556
rect 6512 5516 6518 5528
rect 7374 5516 7380 5528
rect 7432 5516 7438 5568
rect 18046 5516 18052 5568
rect 18104 5556 18110 5568
rect 19518 5556 19524 5568
rect 18104 5528 19524 5556
rect 18104 5516 18110 5528
rect 19518 5516 19524 5528
rect 19576 5516 19582 5568
rect 1104 5466 33028 5488
rect 1104 5414 10950 5466
rect 11002 5414 11014 5466
rect 11066 5414 11078 5466
rect 11130 5414 11142 5466
rect 11194 5414 11206 5466
rect 11258 5414 20950 5466
rect 21002 5414 21014 5466
rect 21066 5414 21078 5466
rect 21130 5414 21142 5466
rect 21194 5414 21206 5466
rect 21258 5414 30950 5466
rect 31002 5414 31014 5466
rect 31066 5414 31078 5466
rect 31130 5414 31142 5466
rect 31194 5414 31206 5466
rect 31258 5414 33028 5466
rect 1104 5392 33028 5414
rect 4154 5312 4160 5364
rect 4212 5352 4218 5364
rect 5442 5352 5448 5364
rect 4212 5324 5448 5352
rect 4212 5312 4218 5324
rect 5442 5312 5448 5324
rect 5500 5312 5506 5364
rect 15286 5312 15292 5364
rect 15344 5352 15350 5364
rect 16853 5355 16911 5361
rect 16853 5352 16865 5355
rect 15344 5324 16865 5352
rect 15344 5312 15350 5324
rect 16853 5321 16865 5324
rect 16899 5321 16911 5355
rect 17954 5352 17960 5364
rect 16853 5315 16911 5321
rect 17052 5324 17960 5352
rect 3878 5244 3884 5296
rect 3936 5284 3942 5296
rect 5718 5284 5724 5296
rect 3936 5256 5724 5284
rect 3936 5244 3942 5256
rect 5718 5244 5724 5256
rect 5776 5244 5782 5296
rect 9125 5287 9183 5293
rect 9125 5284 9137 5287
rect 7852 5256 9137 5284
rect 1949 5219 2007 5225
rect 1949 5185 1961 5219
rect 1995 5216 2007 5219
rect 1995 5188 4476 5216
rect 1995 5185 2007 5188
rect 1949 5179 2007 5185
rect 1578 5108 1584 5160
rect 1636 5108 1642 5160
rect 1765 5151 1823 5157
rect 1765 5117 1777 5151
rect 1811 5148 1823 5151
rect 2682 5148 2688 5160
rect 1811 5120 2688 5148
rect 1811 5117 1823 5120
rect 1765 5111 1823 5117
rect 2682 5108 2688 5120
rect 2740 5108 2746 5160
rect 3694 5108 3700 5160
rect 3752 5108 3758 5160
rect 4448 5148 4476 5188
rect 4522 5176 4528 5228
rect 4580 5176 4586 5228
rect 4614 5176 4620 5228
rect 4672 5216 4678 5228
rect 4672 5188 4752 5216
rect 4672 5176 4678 5188
rect 4724 5157 4752 5188
rect 7466 5176 7472 5228
rect 7524 5216 7530 5228
rect 7852 5216 7880 5256
rect 9125 5253 9137 5256
rect 9171 5284 9183 5287
rect 9674 5284 9680 5296
rect 9171 5256 9680 5284
rect 9171 5253 9183 5256
rect 9125 5247 9183 5253
rect 9674 5244 9680 5256
rect 9732 5244 9738 5296
rect 15194 5244 15200 5296
rect 15252 5284 15258 5296
rect 16945 5287 17003 5293
rect 16945 5284 16957 5287
rect 15252 5256 16957 5284
rect 15252 5244 15258 5256
rect 16945 5253 16957 5256
rect 16991 5253 17003 5287
rect 16945 5247 17003 5253
rect 7524 5188 7880 5216
rect 8573 5219 8631 5225
rect 7524 5176 7530 5188
rect 8573 5185 8585 5219
rect 8619 5216 8631 5219
rect 10042 5216 10048 5228
rect 8619 5188 10048 5216
rect 8619 5185 8631 5188
rect 8573 5179 8631 5185
rect 10042 5176 10048 5188
rect 10100 5176 10106 5228
rect 16209 5219 16267 5225
rect 16209 5216 16221 5219
rect 15120 5188 16221 5216
rect 15120 5160 15148 5188
rect 16209 5185 16221 5188
rect 16255 5216 16267 5219
rect 17052 5216 17080 5324
rect 17954 5312 17960 5324
rect 18012 5312 18018 5364
rect 20070 5312 20076 5364
rect 20128 5352 20134 5364
rect 20441 5355 20499 5361
rect 20441 5352 20453 5355
rect 20128 5324 20453 5352
rect 20128 5312 20134 5324
rect 20441 5321 20453 5324
rect 20487 5321 20499 5355
rect 20441 5315 20499 5321
rect 18322 5216 18328 5228
rect 16255 5188 17080 5216
rect 17880 5188 18328 5216
rect 16255 5185 16267 5188
rect 16209 5179 16267 5185
rect 4709 5151 4767 5157
rect 4448 5120 4568 5148
rect 1394 5040 1400 5092
rect 1452 5080 1458 5092
rect 2409 5083 2467 5089
rect 2409 5080 2421 5083
rect 1452 5052 2421 5080
rect 1452 5040 1458 5052
rect 2409 5049 2421 5052
rect 2455 5049 2467 5083
rect 2409 5043 2467 5049
rect 2222 4972 2228 5024
rect 2280 5012 2286 5024
rect 4430 5012 4436 5024
rect 2280 4984 4436 5012
rect 2280 4972 2286 4984
rect 4430 4972 4436 4984
rect 4488 4972 4494 5024
rect 4540 5012 4568 5120
rect 4709 5117 4721 5151
rect 4755 5117 4767 5151
rect 4709 5111 4767 5117
rect 5258 5108 5264 5160
rect 5316 5148 5322 5160
rect 5810 5148 5816 5160
rect 5316 5120 5816 5148
rect 5316 5108 5322 5120
rect 5810 5108 5816 5120
rect 5868 5108 5874 5160
rect 6178 5074 6184 5126
rect 6236 5074 6242 5126
rect 7926 5108 7932 5160
rect 7984 5108 7990 5160
rect 8018 5108 8024 5160
rect 8076 5148 8082 5160
rect 9306 5148 9312 5160
rect 8076 5120 9312 5148
rect 8076 5108 8082 5120
rect 9306 5108 9312 5120
rect 9364 5108 9370 5160
rect 9490 5108 9496 5160
rect 9548 5148 9554 5160
rect 9953 5151 10011 5157
rect 9953 5148 9965 5151
rect 9548 5120 9965 5148
rect 9548 5108 9554 5120
rect 9953 5117 9965 5120
rect 9999 5117 10011 5151
rect 9953 5111 10011 5117
rect 11747 5117 11805 5123
rect 8757 5083 8815 5089
rect 8757 5049 8769 5083
rect 8803 5080 8815 5083
rect 9398 5080 9404 5092
rect 8803 5052 9404 5080
rect 8803 5049 8815 5052
rect 8757 5043 8815 5049
rect 9398 5040 9404 5052
rect 9456 5040 9462 5092
rect 11747 5083 11759 5117
rect 11793 5114 11805 5117
rect 12066 5114 12072 5160
rect 11793 5108 12072 5114
rect 12124 5108 12130 5160
rect 12250 5108 12256 5160
rect 12308 5148 12314 5160
rect 12989 5151 13047 5157
rect 12989 5148 13001 5151
rect 12308 5120 13001 5148
rect 12308 5108 12314 5120
rect 12989 5117 13001 5120
rect 13035 5117 13047 5151
rect 12989 5111 13047 5117
rect 11793 5086 12112 5108
rect 11793 5083 11805 5086
rect 11747 5077 11805 5083
rect 14734 5074 14740 5126
rect 14792 5074 14798 5126
rect 15102 5108 15108 5160
rect 15160 5108 15166 5160
rect 16025 5151 16083 5157
rect 16025 5117 16037 5151
rect 16071 5148 16083 5151
rect 17880 5148 17908 5188
rect 18322 5176 18328 5188
rect 18380 5176 18386 5228
rect 20070 5176 20076 5228
rect 20128 5216 20134 5228
rect 20809 5219 20867 5225
rect 20809 5216 20821 5219
rect 20128 5188 20821 5216
rect 20128 5176 20134 5188
rect 20809 5185 20821 5188
rect 20855 5185 20867 5219
rect 20809 5179 20867 5185
rect 28736 5188 30144 5216
rect 16071 5120 17908 5148
rect 17957 5151 18015 5157
rect 16071 5117 16083 5120
rect 16025 5111 16083 5117
rect 17957 5117 17969 5151
rect 18003 5150 18015 5151
rect 18138 5150 18144 5160
rect 18003 5122 18144 5150
rect 18003 5117 18015 5122
rect 17957 5111 18015 5117
rect 18138 5108 18144 5122
rect 18196 5108 18202 5160
rect 15194 5040 15200 5092
rect 15252 5080 15258 5092
rect 16117 5083 16175 5089
rect 16117 5080 16129 5083
rect 15252 5052 16129 5080
rect 15252 5040 15258 5052
rect 16117 5049 16129 5052
rect 16163 5049 16175 5083
rect 16117 5043 16175 5049
rect 16482 5040 16488 5092
rect 16540 5080 16546 5092
rect 17310 5080 17316 5092
rect 16540 5052 17316 5080
rect 16540 5040 16546 5052
rect 17310 5040 17316 5052
rect 17368 5040 17374 5092
rect 19610 5074 19616 5126
rect 19668 5074 19674 5126
rect 19978 5108 19984 5160
rect 20036 5148 20042 5160
rect 20625 5151 20683 5157
rect 20625 5148 20637 5151
rect 20036 5120 20637 5148
rect 20036 5108 20042 5120
rect 20625 5117 20637 5120
rect 20671 5117 20683 5151
rect 20625 5111 20683 5117
rect 21450 5108 21456 5160
rect 21508 5108 21514 5160
rect 23155 5117 23213 5123
rect 23155 5083 23167 5117
rect 23201 5114 23213 5117
rect 23474 5114 23480 5160
rect 23201 5108 23480 5114
rect 23532 5108 23538 5160
rect 23201 5086 23520 5108
rect 23201 5083 23213 5086
rect 23155 5077 23213 5083
rect 24302 5074 24308 5126
rect 24360 5074 24366 5126
rect 25958 5108 25964 5160
rect 26016 5108 26022 5160
rect 27430 5074 27436 5126
rect 27488 5074 27494 5126
rect 4617 5015 4675 5021
rect 4617 5012 4629 5015
rect 4540 4984 4629 5012
rect 4617 4981 4629 4984
rect 4663 5012 4675 5015
rect 4982 5012 4988 5024
rect 4663 4984 4988 5012
rect 4663 4981 4675 4984
rect 4617 4975 4675 4981
rect 4982 4972 4988 4984
rect 5040 4972 5046 5024
rect 5077 5015 5135 5021
rect 5077 4981 5089 5015
rect 5123 5012 5135 5015
rect 5166 5012 5172 5024
rect 5123 4984 5172 5012
rect 5123 4981 5135 4984
rect 5077 4975 5135 4981
rect 5166 4972 5172 4984
rect 5224 5012 5230 5024
rect 5718 5012 5724 5024
rect 5224 4984 5724 5012
rect 5224 4972 5230 4984
rect 5718 4972 5724 4984
rect 5776 4972 5782 5024
rect 8662 4972 8668 5024
rect 8720 4972 8726 5024
rect 15102 4972 15108 5024
rect 15160 5012 15166 5024
rect 15657 5015 15715 5021
rect 15657 5012 15669 5015
rect 15160 4984 15669 5012
rect 15160 4972 15166 4984
rect 15657 4981 15669 4984
rect 15703 4981 15715 5015
rect 15657 4975 15715 4981
rect 28442 4972 28448 5024
rect 28500 5012 28506 5024
rect 28736 5012 28764 5188
rect 28902 5108 28908 5160
rect 28960 5148 28966 5160
rect 29089 5151 29147 5157
rect 29089 5148 29101 5151
rect 28960 5120 29101 5148
rect 28960 5108 28966 5120
rect 29089 5117 29101 5120
rect 29135 5117 29147 5151
rect 29089 5111 29147 5117
rect 30116 5114 30144 5188
rect 32125 5151 32183 5157
rect 32125 5148 32137 5151
rect 30423 5117 30481 5123
rect 30423 5114 30435 5117
rect 30116 5086 30435 5114
rect 30423 5083 30435 5086
rect 30469 5083 30481 5117
rect 30423 5077 30481 5083
rect 31772 5120 32137 5148
rect 28500 4984 28764 5012
rect 28500 4972 28506 4984
rect 31478 4972 31484 5024
rect 31536 5012 31542 5024
rect 31772 5012 31800 5120
rect 32125 5117 32137 5120
rect 32171 5117 32183 5151
rect 32125 5111 32183 5117
rect 31536 4984 31800 5012
rect 31536 4972 31542 4984
rect 1104 4922 33028 4944
rect 1104 4870 11610 4922
rect 11662 4870 11674 4922
rect 11726 4870 11738 4922
rect 11790 4870 11802 4922
rect 11854 4870 11866 4922
rect 11918 4870 21610 4922
rect 21662 4870 21674 4922
rect 21726 4870 21738 4922
rect 21790 4870 21802 4922
rect 21854 4870 21866 4922
rect 21918 4870 31610 4922
rect 31662 4870 31674 4922
rect 31726 4870 31738 4922
rect 31790 4870 31802 4922
rect 31854 4870 31866 4922
rect 31918 4870 33028 4922
rect 1104 4848 33028 4870
rect 4706 4768 4712 4820
rect 4764 4808 4770 4820
rect 5166 4808 5172 4820
rect 4764 4780 5172 4808
rect 4764 4768 4770 4780
rect 5166 4768 5172 4780
rect 5224 4768 5230 4820
rect 8294 4808 8300 4820
rect 8036 4780 8300 4808
rect 2222 4666 2228 4718
rect 2280 4666 2286 4718
rect 3970 4632 3976 4684
rect 4028 4632 4034 4684
rect 4430 4632 4436 4684
rect 4488 4632 4494 4684
rect 6178 4666 6184 4718
rect 6236 4666 6242 4718
rect 7653 4675 7711 4681
rect 7653 4641 7665 4675
rect 7699 4672 7711 4675
rect 8036 4672 8064 4780
rect 8294 4768 8300 4780
rect 8352 4768 8358 4820
rect 13998 4808 14004 4820
rect 13740 4780 14004 4808
rect 7699 4644 8064 4672
rect 9306 4666 9312 4718
rect 9364 4666 9370 4718
rect 11931 4709 11989 4715
rect 10229 4675 10287 4681
rect 7699 4641 7711 4644
rect 7653 4635 7711 4641
rect 10229 4641 10241 4675
rect 10275 4672 10287 4675
rect 10594 4672 10600 4684
rect 10275 4644 10600 4672
rect 10275 4641 10287 4644
rect 10229 4635 10287 4641
rect 10594 4632 10600 4644
rect 10652 4632 10658 4684
rect 11931 4675 11943 4709
rect 11977 4706 11989 4709
rect 11977 4678 12296 4706
rect 11977 4675 11989 4678
rect 11931 4669 11989 4675
rect 12268 4672 12296 4678
rect 13265 4675 13323 4681
rect 13265 4672 13277 4675
rect 12268 4644 13277 4672
rect 13265 4641 13277 4644
rect 13311 4641 13323 4675
rect 13265 4635 13323 4641
rect 6638 4564 6644 4616
rect 6696 4604 6702 4616
rect 8018 4604 8024 4616
rect 6696 4576 8024 4604
rect 6696 4564 6702 4576
rect 8018 4564 8024 4576
rect 8076 4564 8082 4616
rect 12342 4564 12348 4616
rect 12400 4604 12406 4616
rect 13740 4604 13768 4780
rect 13998 4768 14004 4780
rect 14056 4768 14062 4820
rect 23658 4768 23664 4820
rect 23716 4768 23722 4820
rect 18138 4740 18144 4752
rect 15010 4666 15016 4718
rect 15068 4666 15074 4718
rect 17635 4709 17693 4715
rect 15933 4675 15991 4681
rect 15933 4641 15945 4675
rect 15979 4672 15991 4675
rect 16298 4672 16304 4684
rect 15979 4644 16304 4672
rect 15979 4641 15991 4644
rect 15933 4635 15991 4641
rect 16298 4632 16304 4644
rect 16356 4632 16362 4684
rect 17635 4675 17647 4709
rect 17681 4706 17693 4709
rect 17972 4712 18144 4740
rect 17972 4706 18000 4712
rect 17681 4678 18000 4706
rect 18138 4700 18144 4712
rect 18196 4700 18202 4752
rect 21683 4709 21741 4715
rect 17681 4675 17693 4678
rect 17635 4669 17693 4675
rect 18046 4632 18052 4684
rect 18104 4672 18110 4684
rect 19886 4672 19892 4684
rect 18104 4644 19892 4672
rect 18104 4632 18110 4644
rect 19886 4632 19892 4644
rect 19944 4632 19950 4684
rect 19981 4675 20039 4681
rect 19981 4641 19993 4675
rect 20027 4672 20039 4675
rect 20346 4672 20352 4684
rect 20027 4644 20352 4672
rect 20027 4641 20039 4644
rect 19981 4635 20039 4641
rect 20346 4632 20352 4644
rect 20404 4632 20410 4684
rect 21683 4675 21695 4709
rect 21729 4706 21741 4709
rect 21729 4684 22048 4706
rect 21729 4678 22008 4684
rect 21729 4675 21741 4678
rect 21683 4669 21741 4675
rect 22002 4632 22008 4678
rect 22060 4632 22066 4684
rect 22278 4632 22284 4684
rect 22336 4672 22342 4684
rect 22649 4675 22707 4681
rect 22649 4672 22661 4675
rect 22336 4644 22661 4672
rect 22336 4632 22342 4644
rect 22649 4641 22661 4644
rect 22695 4641 22707 4675
rect 22649 4635 22707 4641
rect 22738 4632 22744 4684
rect 22796 4672 22802 4684
rect 23014 4672 23020 4684
rect 22796 4644 23020 4672
rect 22796 4632 22802 4644
rect 23014 4632 23020 4644
rect 23072 4672 23078 4684
rect 23293 4675 23351 4681
rect 23293 4672 23305 4675
rect 23072 4644 23305 4672
rect 23072 4632 23078 4644
rect 23293 4641 23305 4644
rect 23339 4641 23351 4675
rect 23293 4635 23351 4641
rect 23474 4632 23480 4684
rect 23532 4632 23538 4684
rect 23934 4632 23940 4684
rect 23992 4672 23998 4684
rect 24213 4675 24271 4681
rect 24213 4672 24225 4675
rect 23992 4644 24225 4672
rect 23992 4632 23998 4644
rect 24213 4641 24225 4644
rect 24259 4641 24271 4675
rect 25958 4666 25964 4718
rect 26016 4666 26022 4718
rect 24213 4635 24271 4641
rect 26786 4632 26792 4684
rect 26844 4632 26850 4684
rect 28534 4666 28540 4718
rect 28592 4666 28598 4718
rect 31711 4709 31769 4715
rect 29178 4632 29184 4684
rect 29236 4672 29242 4684
rect 29917 4675 29975 4681
rect 29917 4672 29929 4675
rect 29236 4644 29929 4672
rect 29236 4632 29242 4644
rect 29917 4641 29929 4644
rect 29963 4641 29975 4675
rect 31711 4675 31723 4709
rect 31757 4706 31769 4709
rect 31757 4684 32076 4706
rect 31757 4678 32036 4684
rect 31757 4675 31769 4678
rect 31711 4669 31769 4675
rect 29917 4635 29975 4641
rect 32030 4632 32036 4678
rect 32088 4632 32094 4684
rect 12400 4576 13768 4604
rect 12400 4564 12406 4576
rect 18138 4564 18144 4616
rect 18196 4604 18202 4616
rect 18969 4607 19027 4613
rect 18969 4604 18981 4607
rect 18196 4576 18981 4604
rect 18196 4564 18202 4576
rect 18969 4573 18981 4576
rect 19015 4604 19027 4607
rect 19015 4576 20392 4604
rect 19015 4573 19027 4576
rect 18969 4567 19027 4573
rect 20364 4548 20392 4576
rect 18046 4496 18052 4548
rect 18104 4536 18110 4548
rect 18601 4539 18659 4545
rect 18601 4536 18613 4539
rect 18104 4508 18613 4536
rect 18104 4496 18110 4508
rect 18601 4505 18613 4508
rect 18647 4505 18659 4539
rect 18601 4499 18659 4505
rect 20346 4496 20352 4548
rect 20404 4496 20410 4548
rect 18506 4428 18512 4480
rect 18564 4428 18570 4480
rect 22186 4428 22192 4480
rect 22244 4468 22250 4480
rect 22465 4471 22523 4477
rect 22465 4468 22477 4471
rect 22244 4440 22477 4468
rect 22244 4428 22250 4440
rect 22465 4437 22477 4440
rect 22511 4468 22523 4471
rect 23750 4468 23756 4480
rect 22511 4440 23756 4468
rect 22511 4437 22523 4440
rect 22465 4431 22523 4437
rect 23750 4428 23756 4440
rect 23808 4428 23814 4480
rect 1104 4378 33028 4400
rect 1104 4326 10950 4378
rect 11002 4326 11014 4378
rect 11066 4326 11078 4378
rect 11130 4326 11142 4378
rect 11194 4326 11206 4378
rect 11258 4326 20950 4378
rect 21002 4326 21014 4378
rect 21066 4326 21078 4378
rect 21130 4326 21142 4378
rect 21194 4326 21206 4378
rect 21258 4326 30950 4378
rect 31002 4326 31014 4378
rect 31066 4326 31078 4378
rect 31130 4326 31142 4378
rect 31194 4326 31206 4378
rect 31258 4326 33028 4378
rect 1104 4304 33028 4326
rect 3786 4224 3792 4276
rect 3844 4264 3850 4276
rect 4706 4264 4712 4276
rect 3844 4236 4712 4264
rect 3844 4224 3850 4236
rect 4706 4224 4712 4236
rect 4764 4224 4770 4276
rect 4985 4267 5043 4273
rect 4985 4233 4997 4267
rect 5031 4264 5043 4267
rect 5442 4264 5448 4276
rect 5031 4236 5448 4264
rect 5031 4233 5043 4236
rect 4985 4227 5043 4233
rect 5442 4224 5448 4236
rect 5500 4224 5506 4276
rect 6730 4264 6736 4276
rect 5644 4236 6736 4264
rect 5534 4196 5540 4208
rect 4448 4168 5540 4196
rect 4448 4137 4476 4168
rect 5534 4156 5540 4168
rect 5592 4156 5598 4208
rect 4433 4131 4491 4137
rect 4433 4097 4445 4131
rect 4479 4097 4491 4131
rect 4433 4091 4491 4097
rect 4798 4088 4804 4140
rect 4856 4128 4862 4140
rect 5644 4128 5672 4236
rect 6730 4224 6736 4236
rect 6788 4224 6794 4276
rect 5810 4156 5816 4208
rect 5868 4156 5874 4208
rect 4856 4100 5672 4128
rect 5721 4131 5779 4137
rect 4856 4088 4862 4100
rect 5721 4097 5733 4131
rect 5767 4128 5779 4131
rect 5828 4128 5856 4156
rect 6822 4128 6828 4140
rect 5767 4100 5856 4128
rect 6012 4100 6828 4128
rect 5767 4097 5779 4100
rect 5721 4091 5779 4097
rect 3697 4063 3755 4069
rect 1946 3986 1952 4038
rect 2004 3986 2010 4038
rect 3697 4029 3709 4063
rect 3743 4060 3755 4063
rect 3878 4060 3884 4072
rect 3743 4032 3884 4060
rect 3743 4029 3755 4032
rect 3697 4023 3755 4029
rect 3878 4020 3884 4032
rect 3936 4020 3942 4072
rect 4246 4020 4252 4072
rect 4304 4060 4310 4072
rect 4522 4060 4528 4072
rect 4304 4032 4528 4060
rect 4304 4020 4310 4032
rect 4522 4020 4528 4032
rect 4580 4020 4586 4072
rect 5905 3995 5963 4001
rect 5905 3961 5917 3995
rect 5951 3992 5963 3995
rect 6012 3992 6040 4100
rect 6822 4088 6828 4100
rect 6880 4088 6886 4140
rect 8938 4088 8944 4140
rect 8996 4128 9002 4140
rect 10410 4128 10416 4140
rect 8996 4100 10416 4128
rect 8996 4088 9002 4100
rect 10410 4088 10416 4100
rect 10468 4088 10474 4140
rect 14642 4088 14648 4140
rect 14700 4128 14706 4140
rect 14700 4100 16160 4128
rect 14700 4088 14706 4100
rect 6730 4020 6736 4072
rect 6788 4020 6794 4072
rect 5951 3964 6040 3992
rect 8478 3986 8484 4038
rect 8536 3986 8542 4038
rect 9306 4020 9312 4072
rect 9364 4060 9370 4072
rect 9953 4063 10011 4069
rect 9953 4060 9965 4063
rect 9364 4032 9965 4060
rect 9364 4020 9370 4032
rect 9953 4029 9965 4032
rect 9999 4029 10011 4063
rect 9953 4023 10011 4029
rect 11747 4029 11805 4035
rect 11747 3995 11759 4029
rect 11793 4026 11805 4029
rect 12066 4026 12072 4072
rect 11793 4020 12072 4026
rect 12124 4020 12130 4072
rect 11793 3998 12112 4020
rect 11793 3995 11805 3998
rect 11747 3989 11805 3995
rect 13354 3986 13360 4038
rect 13412 3986 13418 4038
rect 15010 4020 15016 4072
rect 15068 4020 15074 4072
rect 16132 4069 16160 4100
rect 16117 4063 16175 4069
rect 16117 4029 16129 4063
rect 16163 4029 16175 4063
rect 18785 4063 18843 4069
rect 16117 4023 16175 4029
rect 17862 3986 17868 4038
rect 17920 3986 17926 4038
rect 18785 4029 18797 4063
rect 18831 4060 18843 4063
rect 19150 4060 19156 4072
rect 18831 4032 19156 4060
rect 18831 4029 18843 4032
rect 18785 4023 18843 4029
rect 19150 4020 19156 4032
rect 19208 4020 19214 4072
rect 21453 4063 21511 4069
rect 20438 3986 20444 4038
rect 20496 3986 20502 4038
rect 21453 4029 21465 4063
rect 21499 4060 21511 4063
rect 23934 4060 23940 4072
rect 21499 4032 21588 4060
rect 21499 4029 21511 4032
rect 21453 4023 21511 4029
rect 5951 3961 5963 3964
rect 5905 3955 5963 3961
rect 4617 3927 4675 3933
rect 4617 3893 4629 3927
rect 4663 3924 4675 3927
rect 5626 3924 5632 3936
rect 4663 3896 5632 3924
rect 4663 3893 4675 3896
rect 4617 3887 4675 3893
rect 5626 3884 5632 3896
rect 5684 3884 5690 3936
rect 5813 3927 5871 3933
rect 5813 3893 5825 3927
rect 5859 3924 5871 3927
rect 6178 3924 6184 3936
rect 5859 3896 6184 3924
rect 5859 3893 5871 3896
rect 5813 3887 5871 3893
rect 6178 3884 6184 3896
rect 6236 3884 6242 3936
rect 6273 3927 6331 3933
rect 6273 3893 6285 3927
rect 6319 3924 6331 3927
rect 6638 3924 6644 3936
rect 6319 3896 6644 3924
rect 6319 3893 6331 3896
rect 6273 3887 6331 3893
rect 6638 3884 6644 3896
rect 6696 3884 6702 3936
rect 9401 3927 9459 3933
rect 9401 3893 9413 3927
rect 9447 3924 9459 3927
rect 9490 3924 9496 3936
rect 9447 3896 9496 3924
rect 9447 3893 9459 3896
rect 9401 3887 9459 3893
rect 9490 3884 9496 3896
rect 9548 3884 9554 3936
rect 21560 3924 21588 4032
rect 23155 4029 23213 4035
rect 23155 3995 23167 4029
rect 23201 4026 23213 4029
rect 23492 4032 23940 4060
rect 23492 4026 23520 4032
rect 23201 3998 23520 4026
rect 23934 4020 23940 4032
rect 23992 4020 23998 4072
rect 23201 3995 23213 3998
rect 23155 3989 23213 3995
rect 24302 3986 24308 4038
rect 24360 3986 24366 4038
rect 25958 4020 25964 4072
rect 26016 4020 26022 4072
rect 27157 4063 27215 4069
rect 27157 4029 27169 4063
rect 27203 4060 27215 4063
rect 27203 4032 27568 4060
rect 27203 4029 27215 4032
rect 27157 4023 27215 4029
rect 22002 3924 22008 3936
rect 21560 3896 22008 3924
rect 22002 3884 22008 3896
rect 22060 3884 22066 3936
rect 27540 3924 27568 4032
rect 28859 4029 28917 4035
rect 28859 3995 28871 4029
rect 28905 4026 28917 4029
rect 29178 4026 29184 4072
rect 28905 4020 29184 4026
rect 29236 4020 29242 4072
rect 31665 4063 31723 4069
rect 28905 3998 29224 4020
rect 28905 3995 28917 3998
rect 28859 3989 28917 3995
rect 30006 3986 30012 4038
rect 30064 3986 30070 4038
rect 31665 4029 31677 4063
rect 31711 4060 31723 4063
rect 32030 4060 32036 4072
rect 31711 4032 32036 4060
rect 31711 4029 31723 4032
rect 31665 4023 31723 4029
rect 32030 4020 32036 4032
rect 32088 4020 32094 4072
rect 27614 3924 27620 3936
rect 27540 3896 27620 3924
rect 27614 3884 27620 3896
rect 27672 3884 27678 3936
rect 1104 3834 33028 3856
rect 1104 3782 11610 3834
rect 11662 3782 11674 3834
rect 11726 3782 11738 3834
rect 11790 3782 11802 3834
rect 11854 3782 11866 3834
rect 11918 3782 21610 3834
rect 21662 3782 21674 3834
rect 21726 3782 21738 3834
rect 21790 3782 21802 3834
rect 21854 3782 21866 3834
rect 21918 3782 31610 3834
rect 31662 3782 31674 3834
rect 31726 3782 31738 3834
rect 31790 3782 31802 3834
rect 31854 3782 31866 3834
rect 31918 3782 33028 3834
rect 1104 3760 33028 3782
rect 1946 3680 1952 3732
rect 2004 3720 2010 3732
rect 4154 3720 4160 3732
rect 2004 3692 4160 3720
rect 2004 3680 2010 3692
rect 4154 3680 4160 3692
rect 4212 3680 4218 3732
rect 6822 3680 6828 3732
rect 6880 3720 6886 3732
rect 8938 3720 8944 3732
rect 6880 3692 8944 3720
rect 6880 3680 6886 3692
rect 8938 3680 8944 3692
rect 8996 3680 9002 3732
rect 11330 3680 11336 3732
rect 11388 3720 11394 3732
rect 12894 3720 12900 3732
rect 11388 3692 12900 3720
rect 11388 3680 11394 3692
rect 12894 3680 12900 3692
rect 12952 3680 12958 3732
rect 13354 3680 13360 3732
rect 13412 3720 13418 3732
rect 14642 3720 14648 3732
rect 13412 3692 14648 3720
rect 13412 3680 13418 3692
rect 14642 3680 14648 3692
rect 14700 3680 14706 3732
rect 19242 3720 19248 3732
rect 18984 3692 19248 3720
rect 1765 3655 1823 3661
rect 1765 3621 1777 3655
rect 1811 3652 1823 3655
rect 4246 3652 4252 3664
rect 1811 3624 4252 3652
rect 1811 3621 1823 3624
rect 1765 3615 1823 3621
rect 4246 3612 4252 3624
rect 4304 3612 4310 3664
rect 2866 3544 2872 3596
rect 2924 3584 2930 3596
rect 3786 3584 3792 3596
rect 2924 3556 3792 3584
rect 2924 3544 2930 3556
rect 3786 3544 3792 3556
rect 3844 3544 3850 3596
rect 3973 3587 4031 3593
rect 3973 3553 3985 3587
rect 4019 3584 4031 3587
rect 4430 3584 4436 3596
rect 4019 3556 4436 3584
rect 4019 3553 4031 3556
rect 3973 3547 4031 3553
rect 4430 3544 4436 3556
rect 4488 3544 4494 3596
rect 4798 3578 4804 3630
rect 4856 3578 4862 3630
rect 6638 3612 6644 3664
rect 6696 3652 6702 3664
rect 8662 3652 8668 3664
rect 6696 3624 8668 3652
rect 6696 3612 6702 3624
rect 8662 3612 8668 3624
rect 8720 3612 8726 3664
rect 12161 3655 12219 3661
rect 12161 3621 12173 3655
rect 12207 3652 12219 3655
rect 14826 3652 14832 3664
rect 12207 3624 14832 3652
rect 12207 3621 12219 3624
rect 6178 3544 6184 3596
rect 6236 3584 6242 3596
rect 6454 3584 6460 3596
rect 6236 3556 6460 3584
rect 6236 3544 6242 3556
rect 6454 3544 6460 3556
rect 6512 3544 6518 3596
rect 6549 3587 6607 3593
rect 6549 3553 6561 3587
rect 6595 3584 6607 3587
rect 6914 3584 6920 3596
rect 6595 3556 6920 3584
rect 6595 3553 6607 3556
rect 6549 3547 6607 3553
rect 6914 3544 6920 3556
rect 6972 3544 6978 3596
rect 7282 3544 7288 3596
rect 7340 3544 7346 3596
rect 8113 3587 8171 3593
rect 8113 3553 8125 3587
rect 8159 3584 8171 3587
rect 9030 3584 9036 3596
rect 8159 3556 9036 3584
rect 8159 3553 8171 3556
rect 8113 3547 8171 3553
rect 9030 3544 9036 3556
rect 9088 3544 9094 3596
rect 9122 3544 9128 3596
rect 9180 3544 9186 3596
rect 10778 3568 10784 3620
rect 10836 3590 10842 3620
rect 12161 3615 12219 3621
rect 14826 3612 14832 3624
rect 14884 3612 14890 3664
rect 10836 3568 11192 3590
rect 10796 3562 11192 3568
rect 2774 3476 2780 3528
rect 2832 3476 2838 3528
rect 6086 3476 6092 3528
rect 6144 3516 6150 3528
rect 8205 3519 8263 3525
rect 8205 3516 8217 3519
rect 6144 3488 8217 3516
rect 6144 3476 6150 3488
rect 2133 3451 2191 3457
rect 2133 3417 2145 3451
rect 2179 3448 2191 3451
rect 4246 3448 4252 3460
rect 2179 3420 4252 3448
rect 2179 3417 2191 3420
rect 2133 3411 2191 3417
rect 4246 3408 4252 3420
rect 4304 3408 4310 3460
rect 7116 3457 7144 3488
rect 8205 3485 8217 3488
rect 8251 3485 8263 3519
rect 8205 3479 8263 3485
rect 8294 3476 8300 3528
rect 8352 3476 8358 3528
rect 11164 3516 11192 3562
rect 11974 3544 11980 3596
rect 12032 3544 12038 3596
rect 14093 3587 14151 3593
rect 14093 3553 14105 3587
rect 14139 3553 14151 3587
rect 14093 3547 14151 3553
rect 11701 3519 11759 3525
rect 11701 3516 11713 3519
rect 11164 3488 11713 3516
rect 11701 3485 11713 3488
rect 11747 3485 11759 3519
rect 11992 3516 12020 3544
rect 11701 3479 11759 3485
rect 11900 3488 12020 3516
rect 7101 3451 7159 3457
rect 7101 3417 7113 3451
rect 7147 3417 7159 3451
rect 7101 3411 7159 3417
rect 7745 3451 7803 3457
rect 7745 3417 7757 3451
rect 7791 3448 7803 3451
rect 8478 3448 8484 3460
rect 7791 3420 8484 3448
rect 7791 3417 7803 3420
rect 7745 3411 7803 3417
rect 2225 3383 2283 3389
rect 2225 3349 2237 3383
rect 2271 3380 2283 3383
rect 3326 3380 3332 3392
rect 2271 3352 3332 3380
rect 2271 3349 2283 3352
rect 2225 3343 2283 3349
rect 3326 3340 3332 3352
rect 3384 3340 3390 3392
rect 6454 3340 6460 3392
rect 6512 3380 6518 3392
rect 7760 3380 7788 3411
rect 8478 3408 8484 3420
rect 8536 3408 8542 3460
rect 10804 3408 10810 3460
rect 10862 3408 10868 3460
rect 11900 3457 11928 3488
rect 13446 3476 13452 3528
rect 13504 3476 13510 3528
rect 14108 3516 14136 3547
rect 14734 3544 14740 3596
rect 14792 3584 14798 3596
rect 14921 3587 14979 3593
rect 14921 3584 14933 3587
rect 14792 3556 14933 3584
rect 14792 3544 14798 3556
rect 14921 3553 14933 3556
rect 14967 3553 14979 3587
rect 16666 3578 16672 3630
rect 16724 3578 16730 3630
rect 14921 3547 14979 3553
rect 17494 3544 17500 3596
rect 17552 3584 17558 3596
rect 17552 3556 18460 3584
rect 17552 3544 17558 3556
rect 15102 3516 15108 3528
rect 14108 3488 15108 3516
rect 15102 3476 15108 3488
rect 15160 3476 15166 3528
rect 17954 3476 17960 3528
rect 18012 3476 18018 3528
rect 18432 3516 18460 3556
rect 18506 3544 18512 3596
rect 18564 3544 18570 3596
rect 18984 3516 19012 3692
rect 19242 3680 19248 3692
rect 19300 3680 19306 3732
rect 20806 3680 20812 3732
rect 20864 3720 20870 3732
rect 21085 3723 21143 3729
rect 21085 3720 21097 3723
rect 20864 3692 21097 3720
rect 20864 3680 20870 3692
rect 21085 3689 21097 3692
rect 21131 3689 21143 3723
rect 21085 3683 21143 3689
rect 22094 3680 22100 3732
rect 22152 3720 22158 3732
rect 22281 3723 22339 3729
rect 22281 3720 22293 3723
rect 22152 3692 22293 3720
rect 22152 3680 22158 3692
rect 22281 3689 22293 3692
rect 22327 3720 22339 3723
rect 22646 3720 22652 3732
rect 22327 3692 22652 3720
rect 22327 3689 22339 3692
rect 22281 3683 22339 3689
rect 22646 3680 22652 3692
rect 22704 3720 22710 3732
rect 23198 3720 23204 3732
rect 22704 3692 23204 3720
rect 22704 3680 22710 3692
rect 23198 3680 23204 3692
rect 23256 3680 23262 3732
rect 27614 3680 27620 3732
rect 27672 3720 27678 3732
rect 28534 3720 28540 3732
rect 27672 3692 28540 3720
rect 27672 3680 27678 3692
rect 28534 3680 28540 3692
rect 28592 3680 28598 3732
rect 30006 3680 30012 3732
rect 30064 3720 30070 3732
rect 31478 3720 31484 3732
rect 30064 3692 31484 3720
rect 30064 3680 30070 3692
rect 31478 3680 31484 3692
rect 31536 3680 31542 3732
rect 26786 3652 26792 3664
rect 20303 3621 20361 3627
rect 20303 3587 20315 3621
rect 20349 3618 20361 3621
rect 26283 3621 26341 3627
rect 20349 3596 20668 3618
rect 20349 3590 20628 3596
rect 20349 3587 20361 3590
rect 20303 3581 20361 3587
rect 20622 3544 20628 3590
rect 20680 3544 20686 3596
rect 21269 3587 21327 3593
rect 21269 3553 21281 3587
rect 21315 3553 21327 3587
rect 21269 3547 21327 3553
rect 18432 3488 19012 3516
rect 11885 3451 11943 3457
rect 11885 3417 11897 3451
rect 11931 3417 11943 3451
rect 11885 3411 11943 3417
rect 11974 3408 11980 3460
rect 12032 3448 12038 3460
rect 14918 3448 14924 3460
rect 12032 3420 14924 3448
rect 12032 3408 12038 3420
rect 14918 3408 14924 3420
rect 14976 3408 14982 3460
rect 17126 3408 17132 3460
rect 17184 3448 17190 3460
rect 17589 3451 17647 3457
rect 17589 3448 17601 3451
rect 17184 3420 17601 3448
rect 17184 3408 17190 3420
rect 17589 3417 17601 3420
rect 17635 3417 17647 3451
rect 17972 3448 18000 3476
rect 18598 3448 18604 3460
rect 17972 3420 18604 3448
rect 17589 3411 17647 3417
rect 18598 3408 18604 3420
rect 18656 3408 18662 3460
rect 21284 3448 21312 3547
rect 22094 3544 22100 3596
rect 22152 3544 22158 3596
rect 22186 3544 22192 3596
rect 22244 3584 22250 3596
rect 22925 3587 22983 3593
rect 22925 3584 22937 3587
rect 22244 3556 22937 3584
rect 22244 3544 22250 3556
rect 22925 3553 22937 3556
rect 22971 3553 22983 3587
rect 22925 3547 22983 3553
rect 23014 3544 23020 3596
rect 23072 3544 23078 3596
rect 24302 3544 24308 3596
rect 24360 3584 24366 3596
rect 24489 3587 24547 3593
rect 24489 3584 24501 3587
rect 24360 3556 24501 3584
rect 24360 3544 24366 3556
rect 24489 3553 24501 3556
rect 24535 3553 24547 3587
rect 26283 3587 26295 3621
rect 26329 3618 26341 3621
rect 26620 3624 26792 3652
rect 26620 3618 26648 3624
rect 26329 3590 26648 3618
rect 26786 3612 26792 3624
rect 26844 3612 26850 3664
rect 27154 3612 27160 3664
rect 27212 3652 27218 3664
rect 29362 3652 29368 3664
rect 27212 3624 29368 3652
rect 27212 3612 27218 3624
rect 29362 3612 29368 3624
rect 29420 3612 29426 3664
rect 26329 3587 26341 3590
rect 26283 3581 26341 3587
rect 24489 3547 24547 3553
rect 26878 3544 26884 3596
rect 26936 3584 26942 3596
rect 28994 3584 29000 3596
rect 26936 3556 29000 3584
rect 26936 3544 26942 3556
rect 28994 3544 29000 3556
rect 29052 3544 29058 3596
rect 21453 3519 21511 3525
rect 21453 3485 21465 3519
rect 21499 3516 21511 3519
rect 21913 3519 21971 3525
rect 21913 3516 21925 3519
rect 21499 3488 21925 3516
rect 21499 3485 21511 3488
rect 21453 3479 21511 3485
rect 21913 3485 21925 3488
rect 21959 3516 21971 3519
rect 23032 3516 23060 3544
rect 24854 3516 24860 3528
rect 21959 3488 23060 3516
rect 23952 3488 24860 3516
rect 21959 3485 21971 3488
rect 21913 3479 21971 3485
rect 23952 3448 23980 3488
rect 24854 3476 24860 3488
rect 24912 3476 24918 3528
rect 21284 3420 23980 3448
rect 6512 3352 7788 3380
rect 6512 3340 6518 3352
rect 8294 3340 8300 3392
rect 8352 3380 8358 3392
rect 9122 3380 9128 3392
rect 8352 3352 9128 3380
rect 8352 3340 8358 3352
rect 9122 3340 9128 3352
rect 9180 3340 9186 3392
rect 11330 3340 11336 3392
rect 11388 3380 11394 3392
rect 15010 3380 15016 3392
rect 11388 3352 15016 3380
rect 11388 3340 11394 3352
rect 15010 3340 15016 3352
rect 15068 3340 15074 3392
rect 17218 3340 17224 3392
rect 17276 3380 17282 3392
rect 17497 3383 17555 3389
rect 17497 3380 17509 3383
rect 17276 3352 17509 3380
rect 17276 3340 17282 3352
rect 17497 3349 17509 3352
rect 17543 3349 17555 3383
rect 17497 3343 17555 3349
rect 20714 3340 20720 3392
rect 20772 3380 20778 3392
rect 22741 3383 22799 3389
rect 22741 3380 22753 3383
rect 20772 3352 22753 3380
rect 20772 3340 20778 3352
rect 22741 3349 22753 3352
rect 22787 3349 22799 3383
rect 22741 3343 22799 3349
rect 23661 3383 23719 3389
rect 23661 3349 23673 3383
rect 23707 3380 23719 3383
rect 23750 3380 23756 3392
rect 23707 3352 23756 3380
rect 23707 3349 23719 3352
rect 23661 3343 23719 3349
rect 23750 3340 23756 3352
rect 23808 3340 23814 3392
rect 27614 3340 27620 3392
rect 27672 3340 27678 3392
rect 1104 3290 33028 3312
rect 1104 3238 10950 3290
rect 11002 3238 11014 3290
rect 11066 3238 11078 3290
rect 11130 3238 11142 3290
rect 11194 3238 11206 3290
rect 11258 3238 20950 3290
rect 21002 3238 21014 3290
rect 21066 3238 21078 3290
rect 21130 3238 21142 3290
rect 21194 3238 21206 3290
rect 21258 3238 30950 3290
rect 31002 3238 31014 3290
rect 31066 3238 31078 3290
rect 31130 3238 31142 3290
rect 31194 3238 31206 3290
rect 31258 3238 33028 3290
rect 1104 3216 33028 3238
rect 3786 3136 3792 3188
rect 3844 3176 3850 3188
rect 4338 3176 4344 3188
rect 3844 3148 4344 3176
rect 3844 3136 3850 3148
rect 4338 3136 4344 3148
rect 4396 3136 4402 3188
rect 15194 3136 15200 3188
rect 15252 3176 15258 3188
rect 16298 3176 16304 3188
rect 15252 3148 16304 3176
rect 15252 3136 15258 3148
rect 16298 3136 16304 3148
rect 16356 3136 16362 3188
rect 16390 3136 16396 3188
rect 16448 3136 16454 3188
rect 16528 3136 16534 3188
rect 16586 3176 16592 3188
rect 17126 3176 17132 3188
rect 16586 3148 17132 3176
rect 16586 3136 16592 3148
rect 17126 3136 17132 3148
rect 17184 3136 17190 3188
rect 22094 3136 22100 3188
rect 22152 3176 22158 3188
rect 23201 3179 23259 3185
rect 23201 3176 23213 3179
rect 22152 3148 23213 3176
rect 22152 3136 22158 3148
rect 23201 3145 23213 3148
rect 23247 3145 23259 3179
rect 23201 3139 23259 3145
rect 23750 3136 23756 3188
rect 23808 3176 23814 3188
rect 27614 3176 27620 3188
rect 23808 3148 27620 3176
rect 23808 3136 23814 3148
rect 27614 3136 27620 3148
rect 27672 3136 27678 3188
rect 15930 3068 15936 3120
rect 15988 3108 15994 3120
rect 17494 3108 17500 3120
rect 15988 3080 17500 3108
rect 15988 3068 15994 3080
rect 17494 3068 17500 3080
rect 17552 3068 17558 3120
rect 19610 3068 19616 3120
rect 19668 3108 19674 3120
rect 20073 3111 20131 3117
rect 20073 3108 20085 3111
rect 19668 3080 20085 3108
rect 19668 3068 19674 3080
rect 20073 3077 20085 3080
rect 20119 3108 20131 3111
rect 23014 3108 23020 3120
rect 20119 3080 23020 3108
rect 20119 3077 20131 3080
rect 20073 3071 20131 3077
rect 23014 3068 23020 3080
rect 23072 3068 23078 3120
rect 27065 3111 27123 3117
rect 27065 3108 27077 3111
rect 23216 3080 27077 3108
rect 23216 3052 23244 3080
rect 27065 3077 27077 3080
rect 27111 3077 27123 3111
rect 27065 3071 27123 3077
rect 15841 3043 15899 3049
rect 15841 3009 15853 3043
rect 15887 3040 15899 3043
rect 17770 3040 17776 3052
rect 15887 3012 17776 3040
rect 15887 3009 15899 3012
rect 15841 3003 15899 3009
rect 17770 3000 17776 3012
rect 17828 3000 17834 3052
rect 20162 3000 20168 3052
rect 20220 3040 20226 3052
rect 20441 3043 20499 3049
rect 20441 3040 20453 3043
rect 20220 3012 20453 3040
rect 20220 3000 20226 3012
rect 20441 3009 20453 3012
rect 20487 3040 20499 3043
rect 20714 3040 20720 3052
rect 20487 3012 20720 3040
rect 20487 3009 20499 3012
rect 20441 3003 20499 3009
rect 20714 3000 20720 3012
rect 20772 3000 20778 3052
rect 22480 3012 22876 3040
rect 1670 2932 1676 2984
rect 1728 2932 1734 2984
rect 3375 2941 3433 2947
rect 3375 2907 3387 2941
rect 3421 2938 3433 2941
rect 3694 2938 3700 2984
rect 3421 2932 3700 2938
rect 3752 2932 3758 2984
rect 3421 2910 3740 2932
rect 3421 2907 3433 2910
rect 3375 2901 3433 2907
rect 5074 2898 5080 2950
rect 5132 2898 5138 2950
rect 6638 2932 6644 2984
rect 6696 2972 6702 2984
rect 6733 2975 6791 2981
rect 6733 2972 6745 2975
rect 6696 2944 6745 2972
rect 6696 2932 6702 2944
rect 6733 2941 6745 2944
rect 6779 2941 6791 2975
rect 6733 2935 6791 2941
rect 7006 2932 7012 2984
rect 7064 2972 7070 2984
rect 7285 2975 7343 2981
rect 7285 2972 7297 2975
rect 7064 2944 7297 2972
rect 7064 2932 7070 2944
rect 7285 2941 7297 2944
rect 7331 2941 7343 2975
rect 7285 2935 7343 2941
rect 9030 2898 9036 2950
rect 9088 2898 9094 2950
rect 9398 2932 9404 2984
rect 9456 2972 9462 2984
rect 9456 2944 10456 2972
rect 9456 2932 9462 2944
rect 10428 2938 10456 2944
rect 10735 2941 10793 2947
rect 10735 2938 10747 2941
rect 10428 2910 10747 2938
rect 10735 2907 10747 2910
rect 10781 2907 10793 2941
rect 12434 2932 12440 2984
rect 12492 2932 12498 2984
rect 13081 2975 13139 2981
rect 13081 2941 13093 2975
rect 13127 2972 13139 2975
rect 13127 2944 13492 2972
rect 13127 2941 13139 2944
rect 13081 2935 13139 2941
rect 10735 2901 10793 2907
rect 13464 2836 13492 2944
rect 14783 2941 14841 2947
rect 14783 2907 14795 2941
rect 14829 2938 14841 2941
rect 14829 2916 15148 2938
rect 15930 2932 15936 2984
rect 15988 2932 15994 2984
rect 16528 2932 16534 2984
rect 16586 2972 16592 2984
rect 17218 2972 17224 2984
rect 16586 2944 17224 2972
rect 16586 2932 16592 2944
rect 17218 2932 17224 2944
rect 17276 2932 17282 2984
rect 17497 2975 17555 2981
rect 17497 2941 17509 2975
rect 17543 2972 17555 2975
rect 17862 2972 17868 2984
rect 17543 2944 17868 2972
rect 17543 2941 17555 2944
rect 17497 2935 17555 2941
rect 17862 2932 17868 2944
rect 17920 2932 17926 2984
rect 14829 2910 15108 2916
rect 14829 2907 14841 2910
rect 14783 2901 14841 2907
rect 15102 2864 15108 2910
rect 15160 2864 15166 2916
rect 15286 2864 15292 2916
rect 15344 2904 15350 2916
rect 16025 2907 16083 2913
rect 16025 2904 16037 2907
rect 15344 2876 16037 2904
rect 15344 2864 15350 2876
rect 16025 2873 16037 2876
rect 16071 2873 16083 2907
rect 16758 2904 16764 2916
rect 16025 2867 16083 2873
rect 16546 2876 16764 2904
rect 13722 2836 13728 2848
rect 13464 2808 13728 2836
rect 13722 2796 13728 2808
rect 13780 2796 13786 2848
rect 15194 2796 15200 2848
rect 15252 2836 15258 2848
rect 16546 2836 16574 2876
rect 16758 2864 16764 2876
rect 16816 2904 16822 2916
rect 16853 2907 16911 2913
rect 16853 2904 16865 2907
rect 16816 2876 16865 2904
rect 16816 2864 16822 2876
rect 16853 2873 16865 2876
rect 16899 2873 16911 2907
rect 19150 2898 19156 2950
rect 19208 2898 19214 2950
rect 21358 2932 21364 2984
rect 21416 2932 21422 2984
rect 22480 2981 22508 3012
rect 22281 2975 22339 2981
rect 22281 2972 22293 2975
rect 21468 2944 22293 2972
rect 16853 2867 16911 2873
rect 19794 2864 19800 2916
rect 19852 2904 19858 2916
rect 21468 2904 21496 2944
rect 22281 2941 22293 2944
rect 22327 2941 22339 2975
rect 22281 2935 22339 2941
rect 22465 2975 22523 2981
rect 22465 2941 22477 2975
rect 22511 2941 22523 2975
rect 22465 2935 22523 2941
rect 22649 2975 22707 2981
rect 22649 2941 22661 2975
rect 22695 2972 22707 2975
rect 22848 2972 22876 3012
rect 23198 3000 23204 3052
rect 23256 3000 23262 3052
rect 25593 3043 25651 3049
rect 25593 3040 25605 3043
rect 23308 3012 25605 3040
rect 23308 2984 23336 3012
rect 25593 3009 25605 3012
rect 25639 3009 25651 3043
rect 25593 3003 25651 3009
rect 22695 2944 22784 2972
rect 22848 2944 23244 2972
rect 22695 2941 22707 2944
rect 22649 2935 22707 2941
rect 19852 2876 21496 2904
rect 21637 2907 21695 2913
rect 19852 2864 19858 2876
rect 21637 2873 21649 2907
rect 21683 2904 21695 2907
rect 22370 2904 22376 2916
rect 21683 2876 22376 2904
rect 21683 2873 21695 2876
rect 21637 2867 21695 2873
rect 15252 2808 16574 2836
rect 15252 2796 15258 2808
rect 19978 2796 19984 2848
rect 20036 2796 20042 2848
rect 20438 2796 20444 2848
rect 20496 2836 20502 2848
rect 21652 2836 21680 2867
rect 22370 2864 22376 2876
rect 22428 2904 22434 2916
rect 22756 2904 22784 2944
rect 22428 2876 22784 2904
rect 23216 2904 23244 2944
rect 23290 2932 23296 2984
rect 23348 2932 23354 2984
rect 23842 2932 23848 2984
rect 23900 2932 23906 2984
rect 23934 2932 23940 2984
rect 23992 2932 23998 2984
rect 24578 2932 24584 2984
rect 24636 2972 24642 2984
rect 26237 2975 26295 2981
rect 26237 2972 26249 2975
rect 24636 2944 26249 2972
rect 24636 2932 24642 2944
rect 26237 2941 26249 2944
rect 26283 2941 26295 2975
rect 26237 2935 26295 2941
rect 24489 2907 24547 2913
rect 24489 2904 24501 2907
rect 23216 2876 24501 2904
rect 22428 2864 22434 2876
rect 24489 2873 24501 2876
rect 24535 2873 24547 2907
rect 24489 2867 24547 2873
rect 20496 2808 21680 2836
rect 20496 2796 20502 2808
rect 23014 2796 23020 2848
rect 23072 2836 23078 2848
rect 25133 2839 25191 2845
rect 25133 2836 25145 2839
rect 23072 2808 25145 2836
rect 23072 2796 23078 2808
rect 25133 2805 25145 2808
rect 25179 2836 25191 2839
rect 26050 2836 26056 2848
rect 25179 2808 26056 2836
rect 25179 2805 25191 2808
rect 25133 2799 25191 2805
rect 26050 2796 26056 2808
rect 26108 2796 26114 2848
rect 27614 2796 27620 2848
rect 27672 2796 27678 2848
rect 1104 2746 33028 2768
rect 1104 2694 11610 2746
rect 11662 2694 11674 2746
rect 11726 2694 11738 2746
rect 11790 2694 11802 2746
rect 11854 2694 11866 2746
rect 11918 2694 21610 2746
rect 21662 2694 21674 2746
rect 21726 2694 21738 2746
rect 21790 2694 21802 2746
rect 21854 2694 21866 2746
rect 21918 2694 31610 2746
rect 31662 2694 31674 2746
rect 31726 2694 31738 2746
rect 31790 2694 31802 2746
rect 31854 2694 31866 2746
rect 31918 2694 33028 2746
rect 1104 2672 33028 2694
rect 5810 2592 5816 2644
rect 5868 2632 5874 2644
rect 8294 2632 8300 2644
rect 5868 2604 6408 2632
rect 5868 2592 5874 2604
rect 1995 2533 2053 2539
rect 1995 2530 2007 2533
rect 1688 2508 2007 2530
rect 1670 2456 1676 2508
rect 1728 2502 2007 2508
rect 1728 2456 1734 2502
rect 1995 2499 2007 2502
rect 2041 2499 2053 2533
rect 1995 2493 2053 2499
rect 3786 2456 3792 2508
rect 3844 2456 3850 2508
rect 4798 2490 4804 2542
rect 4856 2490 4862 2542
rect 6380 2428 6408 2604
rect 8036 2604 8300 2632
rect 6549 2499 6607 2505
rect 6549 2465 6561 2499
rect 6595 2496 6607 2499
rect 6914 2496 6920 2508
rect 6595 2468 6920 2496
rect 6595 2465 6607 2468
rect 6549 2459 6607 2465
rect 6914 2456 6920 2468
rect 6972 2456 6978 2508
rect 7561 2499 7619 2505
rect 7561 2465 7573 2499
rect 7607 2465 7619 2499
rect 7561 2459 7619 2465
rect 7576 2428 7604 2459
rect 8036 2428 8064 2604
rect 8294 2592 8300 2604
rect 8352 2592 8358 2644
rect 20714 2592 20720 2644
rect 20772 2632 20778 2644
rect 20772 2604 23888 2632
rect 20772 2592 20778 2604
rect 12434 2564 12440 2576
rect 9355 2533 9413 2539
rect 9355 2499 9367 2533
rect 9401 2530 9413 2533
rect 11931 2533 11989 2539
rect 9401 2502 9720 2530
rect 9401 2499 9413 2502
rect 9355 2493 9413 2499
rect 9692 2496 9720 2502
rect 10137 2499 10195 2505
rect 10137 2496 10149 2499
rect 9692 2468 10149 2496
rect 10137 2465 10149 2468
rect 10183 2465 10195 2499
rect 11931 2499 11943 2533
rect 11977 2530 11989 2533
rect 12268 2536 12440 2564
rect 12268 2530 12296 2536
rect 11977 2502 12296 2530
rect 12434 2524 12440 2536
rect 12492 2524 12498 2576
rect 18506 2564 18512 2576
rect 11977 2499 11989 2502
rect 11931 2493 11989 2499
rect 10137 2459 10195 2465
rect 12802 2456 12808 2508
rect 12860 2456 12866 2508
rect 14550 2490 14556 2542
rect 14608 2490 14614 2542
rect 17359 2533 17417 2539
rect 15102 2456 15108 2508
rect 15160 2496 15166 2508
rect 15565 2499 15623 2505
rect 15565 2496 15577 2499
rect 15160 2468 15577 2496
rect 15160 2456 15166 2468
rect 15565 2465 15577 2468
rect 15611 2465 15623 2499
rect 17359 2499 17371 2533
rect 17405 2530 17417 2533
rect 17696 2536 18512 2564
rect 17696 2530 17724 2536
rect 17405 2502 17724 2530
rect 18506 2524 18512 2536
rect 18564 2524 18570 2576
rect 22005 2567 22063 2573
rect 22005 2564 22017 2567
rect 17405 2499 17417 2502
rect 17359 2493 17417 2499
rect 18874 2490 18880 2542
rect 18932 2490 18938 2542
rect 20732 2536 22017 2564
rect 15565 2459 15623 2465
rect 20622 2456 20628 2508
rect 20680 2456 20686 2508
rect 6380 2400 7604 2428
rect 7668 2400 8064 2428
rect 7668 2372 7696 2400
rect 20162 2388 20168 2440
rect 20220 2428 20226 2440
rect 20732 2428 20760 2536
rect 22005 2533 22017 2536
rect 22051 2533 22063 2567
rect 23569 2567 23627 2573
rect 23569 2564 23581 2567
rect 22005 2527 22063 2533
rect 22204 2536 23581 2564
rect 22204 2505 22232 2536
rect 23569 2533 23581 2536
rect 23615 2533 23627 2567
rect 23860 2564 23888 2604
rect 23934 2592 23940 2644
rect 23992 2632 23998 2644
rect 24765 2635 24823 2641
rect 24765 2632 24777 2635
rect 23992 2604 24777 2632
rect 23992 2592 23998 2604
rect 24765 2601 24777 2604
rect 24811 2601 24823 2635
rect 24765 2595 24823 2601
rect 25869 2567 25927 2573
rect 25869 2564 25881 2567
rect 23860 2536 25881 2564
rect 23569 2527 23627 2533
rect 25869 2533 25881 2536
rect 25915 2564 25927 2567
rect 26973 2567 27031 2573
rect 26973 2564 26985 2567
rect 25915 2536 26985 2564
rect 25915 2533 25927 2536
rect 25869 2527 25927 2533
rect 26973 2533 26985 2536
rect 27019 2533 27031 2567
rect 26973 2527 27031 2533
rect 22189 2499 22247 2505
rect 22189 2465 22201 2499
rect 22235 2465 22247 2499
rect 22189 2459 22247 2465
rect 22370 2456 22376 2508
rect 22428 2456 22434 2508
rect 22833 2499 22891 2505
rect 22833 2465 22845 2499
rect 22879 2465 22891 2499
rect 22833 2459 22891 2465
rect 20220 2400 20760 2428
rect 20220 2388 20226 2400
rect 20806 2388 20812 2440
rect 20864 2428 20870 2440
rect 21545 2431 21603 2437
rect 21545 2428 21557 2431
rect 20864 2400 21557 2428
rect 20864 2388 20870 2400
rect 21545 2397 21557 2400
rect 21591 2397 21603 2431
rect 21545 2391 21603 2397
rect 7650 2320 7656 2372
rect 7708 2320 7714 2372
rect 20530 2320 20536 2372
rect 20588 2360 20594 2372
rect 21269 2363 21327 2369
rect 21269 2360 21281 2363
rect 20588 2332 21281 2360
rect 20588 2320 20594 2332
rect 21269 2329 21281 2332
rect 21315 2329 21327 2363
rect 21269 2323 21327 2329
rect 20714 2252 20720 2304
rect 20772 2292 20778 2304
rect 21085 2295 21143 2301
rect 21085 2292 21097 2295
rect 20772 2264 21097 2292
rect 20772 2252 20778 2264
rect 21085 2261 21097 2264
rect 21131 2261 21143 2295
rect 21284 2292 21312 2323
rect 22002 2320 22008 2372
rect 22060 2360 22066 2372
rect 22848 2360 22876 2459
rect 23290 2456 23296 2508
rect 23348 2496 23354 2508
rect 23661 2499 23719 2505
rect 23661 2496 23673 2499
rect 23348 2468 23673 2496
rect 23348 2456 23354 2468
rect 23661 2465 23673 2468
rect 23707 2496 23719 2499
rect 25317 2499 25375 2505
rect 25317 2496 25329 2499
rect 23707 2468 25329 2496
rect 23707 2465 23719 2468
rect 23661 2459 23719 2465
rect 25317 2465 25329 2468
rect 25363 2465 25375 2499
rect 25317 2459 25375 2465
rect 22060 2332 22876 2360
rect 22060 2320 22066 2332
rect 23198 2320 23204 2372
rect 23256 2360 23262 2372
rect 26421 2363 26479 2369
rect 26421 2360 26433 2363
rect 23256 2332 26433 2360
rect 23256 2320 23262 2332
rect 26421 2329 26433 2332
rect 26467 2329 26479 2363
rect 26421 2323 26479 2329
rect 22370 2292 22376 2304
rect 21284 2264 22376 2292
rect 21085 2255 21143 2261
rect 22370 2252 22376 2264
rect 22428 2252 22434 2304
rect 22830 2252 22836 2304
rect 22888 2292 22894 2304
rect 22925 2295 22983 2301
rect 22925 2292 22937 2295
rect 22888 2264 22937 2292
rect 22888 2252 22894 2264
rect 22925 2261 22937 2264
rect 22971 2292 22983 2295
rect 23014 2292 23020 2304
rect 22971 2264 23020 2292
rect 22971 2261 22983 2264
rect 22925 2255 22983 2261
rect 23014 2252 23020 2264
rect 23072 2252 23078 2304
rect 24210 2252 24216 2304
rect 24268 2252 24274 2304
rect 1104 2202 33028 2224
rect 1104 2150 10950 2202
rect 11002 2150 11014 2202
rect 11066 2150 11078 2202
rect 11130 2150 11142 2202
rect 11194 2150 11206 2202
rect 11258 2150 20950 2202
rect 21002 2150 21014 2202
rect 21066 2150 21078 2202
rect 21130 2150 21142 2202
rect 21194 2150 21206 2202
rect 21258 2150 30950 2202
rect 31002 2150 31014 2202
rect 31066 2150 31078 2202
rect 31130 2150 31142 2202
rect 31194 2150 31206 2202
rect 31258 2150 33028 2202
rect 1104 2128 33028 2150
rect 15654 2048 15660 2100
rect 15712 2048 15718 2100
rect 22097 2091 22155 2097
rect 22097 2057 22109 2091
rect 22143 2088 22155 2091
rect 22186 2088 22192 2100
rect 22143 2060 22192 2088
rect 22143 2057 22155 2060
rect 22097 2051 22155 2057
rect 22186 2048 22192 2060
rect 22244 2048 22250 2100
rect 22554 2048 22560 2100
rect 22612 2088 22618 2100
rect 22649 2091 22707 2097
rect 22649 2088 22661 2091
rect 22612 2060 22661 2088
rect 22612 2048 22618 2060
rect 22649 2057 22661 2060
rect 22695 2057 22707 2091
rect 22649 2051 22707 2057
rect 23658 2048 23664 2100
rect 23716 2088 23722 2100
rect 25501 2091 25559 2097
rect 25501 2088 25513 2091
rect 23716 2060 25513 2088
rect 23716 2048 23722 2060
rect 25501 2057 25513 2060
rect 25547 2057 25559 2091
rect 25501 2051 25559 2057
rect 26050 2048 26056 2100
rect 26108 2048 26114 2100
rect 15010 1980 15016 2032
rect 15068 2020 15074 2032
rect 15749 2023 15807 2029
rect 15749 2020 15761 2023
rect 15068 1992 15761 2020
rect 15068 1980 15074 1992
rect 15749 1989 15761 1992
rect 15795 1989 15807 2023
rect 15749 1983 15807 1989
rect 16206 1980 16212 2032
rect 16264 2020 16270 2032
rect 16761 2023 16819 2029
rect 16761 2020 16773 2023
rect 16264 1992 16773 2020
rect 16264 1980 16270 1992
rect 16761 1989 16773 1992
rect 16807 2020 16819 2023
rect 17862 2020 17868 2032
rect 16807 1992 17868 2020
rect 16807 1989 16819 1992
rect 16761 1983 16819 1989
rect 17862 1980 17868 1992
rect 17920 1980 17926 2032
rect 20806 1980 20812 2032
rect 20864 1980 20870 2032
rect 21453 2023 21511 2029
rect 21453 1989 21465 2023
rect 21499 2020 21511 2023
rect 22278 2020 22284 2032
rect 21499 1992 22284 2020
rect 21499 1989 21511 1992
rect 21453 1983 21511 1989
rect 22278 1980 22284 1992
rect 22336 1980 22342 2032
rect 22462 1980 22468 2032
rect 22520 2020 22526 2032
rect 23293 2023 23351 2029
rect 23293 2020 23305 2023
rect 22520 1992 23305 2020
rect 22520 1980 22526 1992
rect 23293 1989 23305 1992
rect 23339 2020 23351 2023
rect 24210 2020 24216 2032
rect 23339 1992 24216 2020
rect 23339 1989 23351 1992
rect 23293 1983 23351 1989
rect 24210 1980 24216 1992
rect 24268 1980 24274 2032
rect 14642 1912 14648 1964
rect 14700 1952 14706 1964
rect 16298 1952 16304 1964
rect 14700 1924 16304 1952
rect 14700 1912 14706 1924
rect 16298 1912 16304 1924
rect 16356 1912 16362 1964
rect 17037 1955 17095 1961
rect 17037 1921 17049 1955
rect 17083 1952 17095 1955
rect 17083 1924 18368 1952
rect 17083 1921 17095 1924
rect 17037 1915 17095 1921
rect 1670 1844 1676 1896
rect 1728 1844 1734 1896
rect 3326 1810 3332 1862
rect 3384 1810 3390 1862
rect 5031 1853 5089 1859
rect 5031 1850 5043 1853
rect 4522 1776 4528 1828
rect 4580 1816 4586 1828
rect 4724 1822 5043 1850
rect 4724 1816 4752 1822
rect 4580 1788 4752 1816
rect 5031 1819 5043 1822
rect 5077 1819 5089 1853
rect 6730 1844 6736 1896
rect 6788 1844 6794 1896
rect 5031 1813 5089 1819
rect 7650 1810 7656 1862
rect 7708 1810 7714 1862
rect 9398 1844 9404 1896
rect 9456 1844 9462 1896
rect 9674 1844 9680 1896
rect 9732 1884 9738 1896
rect 10413 1887 10471 1893
rect 10413 1884 10425 1887
rect 9732 1856 10425 1884
rect 9732 1844 9738 1856
rect 10413 1853 10425 1856
rect 10459 1853 10471 1887
rect 12802 1884 12808 1896
rect 10413 1847 10471 1853
rect 12207 1853 12265 1859
rect 12207 1819 12219 1853
rect 12253 1850 12265 1853
rect 12544 1856 12808 1884
rect 12544 1850 12572 1856
rect 12253 1822 12572 1850
rect 12802 1844 12808 1856
rect 12860 1844 12866 1896
rect 12253 1819 12265 1822
rect 12207 1813 12265 1819
rect 13354 1810 13360 1862
rect 13412 1810 13418 1862
rect 15102 1844 15108 1896
rect 15160 1844 15166 1896
rect 17954 1844 17960 1896
rect 18012 1844 18018 1896
rect 4580 1776 4586 1788
rect 16022 1776 16028 1828
rect 16080 1816 16086 1828
rect 16117 1819 16175 1825
rect 16117 1816 16129 1819
rect 16080 1788 16129 1816
rect 16080 1776 16086 1788
rect 16117 1785 16129 1788
rect 16163 1785 16175 1819
rect 16117 1779 16175 1785
rect 15746 1708 15752 1760
rect 15804 1748 15810 1760
rect 16577 1751 16635 1757
rect 16577 1748 16589 1751
rect 15804 1720 16589 1748
rect 15804 1708 15810 1720
rect 16577 1717 16589 1720
rect 16623 1717 16635 1751
rect 16577 1711 16635 1717
rect 16666 1708 16672 1760
rect 16724 1748 16730 1760
rect 17402 1748 17408 1760
rect 16724 1720 17408 1748
rect 16724 1708 16730 1720
rect 17402 1708 17408 1720
rect 17460 1708 17466 1760
rect 18340 1748 18368 1924
rect 20530 1912 20536 1964
rect 20588 1952 20594 1964
rect 24397 1955 24455 1961
rect 24397 1952 24409 1955
rect 20588 1924 24409 1952
rect 20588 1912 20594 1924
rect 19659 1853 19717 1859
rect 19659 1819 19671 1853
rect 19705 1850 19717 1853
rect 19705 1822 20024 1850
rect 20162 1844 20168 1896
rect 20220 1884 20226 1896
rect 20438 1884 20444 1896
rect 20220 1856 20444 1884
rect 20220 1844 20226 1856
rect 20438 1844 20444 1856
rect 20496 1844 20502 1896
rect 21376 1893 21404 1924
rect 24397 1921 24409 1924
rect 24443 1921 24455 1955
rect 24397 1915 24455 1921
rect 20625 1887 20683 1893
rect 20625 1853 20637 1887
rect 20671 1884 20683 1887
rect 21361 1887 21419 1893
rect 20671 1856 21220 1884
rect 20671 1853 20683 1856
rect 20625 1847 20683 1853
rect 19705 1819 19717 1822
rect 19659 1813 19717 1819
rect 19996 1816 20024 1822
rect 20714 1816 20720 1828
rect 19996 1788 20720 1816
rect 20714 1776 20720 1788
rect 20772 1776 20778 1828
rect 21192 1816 21220 1856
rect 21361 1853 21373 1887
rect 21407 1853 21419 1887
rect 21361 1847 21419 1853
rect 22002 1844 22008 1896
rect 22060 1844 22066 1896
rect 22738 1844 22744 1896
rect 22796 1884 22802 1896
rect 22833 1887 22891 1893
rect 22833 1884 22845 1887
rect 22796 1856 22845 1884
rect 22796 1844 22802 1856
rect 22833 1853 22845 1856
rect 22879 1884 22891 1887
rect 24949 1887 25007 1893
rect 24949 1884 24961 1887
rect 22879 1856 24961 1884
rect 22879 1853 22891 1856
rect 22833 1847 22891 1853
rect 24949 1853 24961 1856
rect 24995 1853 25007 1887
rect 24949 1847 25007 1853
rect 21450 1816 21456 1828
rect 21192 1788 21456 1816
rect 21450 1776 21456 1788
rect 21508 1776 21514 1828
rect 23198 1816 23204 1828
rect 22066 1788 23204 1816
rect 18598 1748 18604 1760
rect 18340 1720 18604 1748
rect 18598 1708 18604 1720
rect 18656 1708 18662 1760
rect 19978 1708 19984 1760
rect 20036 1748 20042 1760
rect 22066 1748 22094 1788
rect 23198 1776 23204 1788
rect 23256 1776 23262 1828
rect 20036 1720 22094 1748
rect 20036 1708 20042 1720
rect 22370 1708 22376 1760
rect 22428 1748 22434 1760
rect 23934 1748 23940 1760
rect 22428 1720 23940 1748
rect 22428 1708 22434 1720
rect 23934 1708 23940 1720
rect 23992 1708 23998 1760
rect 1104 1658 33028 1680
rect 1104 1606 11610 1658
rect 11662 1606 11674 1658
rect 11726 1606 11738 1658
rect 11790 1606 11802 1658
rect 11854 1606 11866 1658
rect 11918 1606 21610 1658
rect 21662 1606 21674 1658
rect 21726 1606 21738 1658
rect 21790 1606 21802 1658
rect 21854 1606 21866 1658
rect 21918 1606 31610 1658
rect 31662 1606 31674 1658
rect 31726 1606 31738 1658
rect 31790 1606 31802 1658
rect 31854 1606 31866 1658
rect 31918 1606 33028 1658
rect 1104 1584 33028 1606
rect 6546 1504 6552 1556
rect 6604 1544 6610 1556
rect 16574 1544 16580 1556
rect 6604 1516 6960 1544
rect 6604 1504 6610 1516
rect 3651 1445 3709 1451
rect 1946 1368 1952 1420
rect 2004 1368 2010 1420
rect 3651 1411 3663 1445
rect 3697 1442 3709 1445
rect 6227 1445 6285 1451
rect 3697 1414 4016 1442
rect 3697 1411 3709 1414
rect 3651 1405 3709 1411
rect 3988 1408 4016 1414
rect 4430 1408 4436 1420
rect 3988 1380 4436 1408
rect 4430 1368 4436 1380
rect 4488 1368 4494 1420
rect 4522 1368 4528 1420
rect 4580 1368 4586 1420
rect 6227 1411 6239 1445
rect 6273 1442 6285 1445
rect 6273 1414 6592 1442
rect 6273 1411 6285 1414
rect 6227 1405 6285 1411
rect 6564 1408 6592 1414
rect 6822 1408 6828 1420
rect 6564 1380 6828 1408
rect 6822 1368 6828 1380
rect 6880 1368 6886 1420
rect 6932 1408 6960 1516
rect 16316 1516 16580 1544
rect 9355 1445 9413 1451
rect 7561 1411 7619 1417
rect 7561 1408 7573 1411
rect 6932 1380 7573 1408
rect 7561 1377 7573 1380
rect 7607 1377 7619 1411
rect 9355 1411 9367 1445
rect 9401 1442 9413 1445
rect 9674 1442 9680 1488
rect 9401 1436 9680 1442
rect 9732 1436 9738 1488
rect 9401 1414 9720 1436
rect 9401 1411 9413 1414
rect 9355 1405 9413 1411
rect 10502 1402 10508 1454
rect 10560 1402 10566 1454
rect 14783 1445 14841 1451
rect 7561 1371 7619 1377
rect 12250 1368 12256 1420
rect 12308 1368 12314 1420
rect 12342 1368 12348 1420
rect 12400 1408 12406 1420
rect 12989 1411 13047 1417
rect 12989 1408 13001 1411
rect 12400 1380 13001 1408
rect 12400 1368 12406 1380
rect 12989 1377 13001 1380
rect 13035 1377 13047 1411
rect 14783 1411 14795 1445
rect 14829 1442 14841 1445
rect 15102 1442 15108 1488
rect 14829 1436 15108 1442
rect 15160 1436 15166 1488
rect 14829 1414 15148 1436
rect 14829 1411 14841 1414
rect 14783 1405 14841 1411
rect 15933 1411 15991 1417
rect 12989 1371 13047 1377
rect 15933 1377 15945 1411
rect 15979 1408 15991 1411
rect 16316 1408 16344 1516
rect 16574 1504 16580 1516
rect 16632 1504 16638 1556
rect 21450 1504 21456 1556
rect 21508 1544 21514 1556
rect 21637 1547 21695 1553
rect 21637 1544 21649 1547
rect 21508 1516 21649 1544
rect 21508 1504 21514 1516
rect 21637 1513 21649 1516
rect 21683 1513 21695 1547
rect 21637 1507 21695 1513
rect 22830 1504 22836 1556
rect 22888 1504 22894 1556
rect 15979 1380 16344 1408
rect 17635 1445 17693 1451
rect 17635 1411 17647 1445
rect 17681 1442 17693 1445
rect 17954 1442 17960 1488
rect 17681 1436 17960 1442
rect 18012 1436 18018 1488
rect 19291 1445 19349 1451
rect 19291 1442 19303 1445
rect 17681 1414 18000 1436
rect 18984 1420 19303 1442
rect 17681 1411 17693 1414
rect 17635 1405 17693 1411
rect 15979 1377 15991 1380
rect 15933 1371 15991 1377
rect 18966 1368 18972 1420
rect 19024 1414 19303 1420
rect 19024 1368 19030 1414
rect 19291 1411 19303 1414
rect 19337 1411 19349 1445
rect 22186 1436 22192 1488
rect 22244 1476 22250 1488
rect 23658 1476 23664 1488
rect 22244 1448 23664 1476
rect 22244 1436 22250 1448
rect 23658 1436 23664 1448
rect 23716 1436 23722 1488
rect 19291 1405 19349 1411
rect 20714 1368 20720 1420
rect 20772 1408 20778 1420
rect 20993 1411 21051 1417
rect 20993 1408 21005 1411
rect 20772 1380 21005 1408
rect 20772 1368 20778 1380
rect 20993 1377 21005 1380
rect 21039 1377 21051 1411
rect 20993 1371 21051 1377
rect 21358 1368 21364 1420
rect 21416 1408 21422 1420
rect 21729 1411 21787 1417
rect 21729 1408 21741 1411
rect 21416 1380 21741 1408
rect 21416 1368 21422 1380
rect 21729 1377 21741 1380
rect 21775 1377 21787 1411
rect 21729 1371 21787 1377
rect 12158 1300 12164 1352
rect 12216 1340 12222 1352
rect 13078 1340 13084 1352
rect 12216 1312 13084 1340
rect 12216 1300 12222 1312
rect 13078 1300 13084 1312
rect 13136 1300 13142 1352
rect 22002 1300 22008 1352
rect 22060 1340 22066 1352
rect 24213 1343 24271 1349
rect 24213 1340 24225 1343
rect 22060 1312 24225 1340
rect 22060 1300 22066 1312
rect 24213 1309 24225 1312
rect 24259 1309 24271 1343
rect 24213 1303 24271 1309
rect 24854 1300 24860 1352
rect 24912 1300 24918 1352
rect 22281 1275 22339 1281
rect 22281 1241 22293 1275
rect 22327 1272 22339 1275
rect 22646 1272 22652 1284
rect 22327 1244 22652 1272
rect 22327 1241 22339 1244
rect 22281 1235 22339 1241
rect 22646 1232 22652 1244
rect 22704 1232 22710 1284
rect 23382 1232 23388 1284
rect 23440 1272 23446 1284
rect 26142 1272 26148 1284
rect 23440 1244 26148 1272
rect 23440 1232 23446 1244
rect 26142 1232 26148 1244
rect 26200 1232 26206 1284
rect 1104 1114 33028 1136
rect 1104 1062 10950 1114
rect 11002 1062 11014 1114
rect 11066 1062 11078 1114
rect 11130 1062 11142 1114
rect 11194 1062 11206 1114
rect 11258 1062 20950 1114
rect 21002 1062 21014 1114
rect 21066 1062 21078 1114
rect 21130 1062 21142 1114
rect 21194 1062 21206 1114
rect 21258 1062 30950 1114
rect 31002 1062 31014 1114
rect 31066 1062 31078 1114
rect 31130 1062 31142 1114
rect 31194 1062 31206 1114
rect 31258 1062 33028 1114
rect 1104 1040 33028 1062
rect 12342 960 12348 1012
rect 12400 1000 12406 1012
rect 15286 1000 15292 1012
rect 12400 972 15292 1000
rect 12400 960 12406 972
rect 15286 960 15292 972
rect 15344 960 15350 1012
rect 20162 1000 20168 1012
rect 19352 972 20168 1000
rect 14090 892 14096 944
rect 14148 892 14154 944
rect 19242 932 19248 944
rect 18340 904 19248 932
rect 12989 867 13047 873
rect 12989 833 13001 867
rect 13035 833 13047 867
rect 12989 827 13047 833
rect 1946 722 1952 774
rect 2004 722 2010 774
rect 3326 756 3332 808
rect 3384 796 3390 808
rect 3605 799 3663 805
rect 3605 796 3617 799
rect 3384 768 3617 796
rect 3384 756 3390 768
rect 3605 765 3617 768
rect 3651 765 3663 799
rect 3605 759 3663 765
rect 4430 756 4436 808
rect 4488 756 4494 808
rect 6730 796 6736 808
rect 6227 765 6285 771
rect 6227 731 6239 765
rect 6273 762 6285 765
rect 6564 768 6736 796
rect 6564 762 6592 768
rect 6273 734 6592 762
rect 6730 756 6736 768
rect 6788 756 6794 808
rect 6822 756 6828 808
rect 6880 796 6886 808
rect 7285 799 7343 805
rect 7285 796 7297 799
rect 6880 768 7297 796
rect 6880 756 6886 768
rect 7285 765 7297 768
rect 7331 765 7343 799
rect 10137 799 10195 805
rect 10137 796 10149 799
rect 7285 759 7343 765
rect 9079 765 9137 771
rect 6273 731 6285 734
rect 6227 725 6285 731
rect 9079 731 9091 765
rect 9125 762 9137 765
rect 9416 768 10149 796
rect 9416 762 9444 768
rect 9125 734 9444 762
rect 10137 765 10149 768
rect 10183 765 10195 799
rect 10137 759 10195 765
rect 11931 765 11989 771
rect 9125 731 9137 734
rect 9079 725 9137 731
rect 11931 731 11943 765
rect 11977 762 11989 765
rect 12250 762 12256 808
rect 11977 756 12256 762
rect 12308 756 12314 808
rect 13004 796 13032 827
rect 13078 824 13084 876
rect 13136 824 13142 876
rect 13354 824 13360 876
rect 13412 864 13418 876
rect 13412 836 15700 864
rect 13412 824 13418 836
rect 14826 796 14832 808
rect 13004 768 14832 796
rect 14826 756 14832 768
rect 14884 756 14890 808
rect 14918 756 14924 808
rect 14976 756 14982 808
rect 15010 756 15016 808
rect 15068 756 15074 808
rect 15672 805 15700 836
rect 15657 799 15715 805
rect 15657 765 15669 799
rect 15703 765 15715 799
rect 15657 759 15715 765
rect 11977 734 12296 756
rect 11977 731 11989 734
rect 11931 725 11989 731
rect 14458 688 14464 740
rect 14516 728 14522 740
rect 15028 728 15056 756
rect 14516 700 15056 728
rect 17402 722 17408 774
rect 17460 722 17466 774
rect 14516 688 14522 700
rect 13170 620 13176 672
rect 13228 620 13234 672
rect 13538 620 13544 672
rect 13596 620 13602 672
rect 13998 620 14004 672
rect 14056 620 14062 672
rect 15010 620 15016 672
rect 15068 620 15074 672
rect 17954 620 17960 672
rect 18012 660 18018 672
rect 18340 660 18368 904
rect 19242 892 19248 904
rect 19300 892 19306 944
rect 19352 873 19380 972
rect 20162 960 20168 972
rect 20220 960 20226 1012
rect 20254 960 20260 1012
rect 20312 960 20318 1012
rect 21284 972 21588 1000
rect 21284 932 21312 972
rect 19536 904 21312 932
rect 21453 935 21511 941
rect 18877 867 18935 873
rect 18877 833 18889 867
rect 18923 864 18935 867
rect 19337 867 19395 873
rect 19337 864 19349 867
rect 18923 836 19349 864
rect 18923 833 18935 836
rect 18877 827 18935 833
rect 19337 833 19349 836
rect 19383 833 19395 867
rect 19337 827 19395 833
rect 19536 805 19564 904
rect 21453 901 21465 935
rect 21499 901 21511 935
rect 21560 932 21588 972
rect 23934 960 23940 1012
rect 23992 1000 23998 1012
rect 25317 1003 25375 1009
rect 25317 1000 25329 1003
rect 23992 972 25329 1000
rect 23992 960 23998 972
rect 25317 969 25329 972
rect 25363 969 25375 1003
rect 25317 963 25375 969
rect 23842 932 23848 944
rect 21560 904 23848 932
rect 21453 895 21511 901
rect 21468 864 21496 895
rect 23842 892 23848 904
rect 23900 892 23906 944
rect 20364 836 21496 864
rect 22097 867 22155 873
rect 18693 799 18751 805
rect 18693 765 18705 799
rect 18739 765 18751 799
rect 18693 759 18751 765
rect 19521 799 19579 805
rect 19521 765 19533 799
rect 19567 765 19579 799
rect 19521 759 19579 765
rect 20165 799 20223 805
rect 20165 765 20177 799
rect 20211 796 20223 799
rect 20254 796 20260 808
rect 20211 768 20260 796
rect 20211 765 20223 768
rect 20165 759 20223 765
rect 18414 688 18420 740
rect 18472 728 18478 740
rect 18708 728 18736 759
rect 20254 756 20260 768
rect 20312 756 20318 808
rect 20364 728 20392 836
rect 22097 833 22109 867
rect 22143 864 22155 867
rect 22186 864 22192 876
rect 22143 836 22192 864
rect 22143 833 22155 836
rect 22097 827 22155 833
rect 22186 824 22192 836
rect 22244 824 22250 876
rect 22649 867 22707 873
rect 22649 833 22661 867
rect 22695 864 22707 867
rect 23198 864 23204 876
rect 22695 836 23204 864
rect 22695 833 22707 836
rect 22649 827 22707 833
rect 23198 824 23204 836
rect 23256 824 23262 876
rect 24854 824 24860 876
rect 24912 824 24918 876
rect 21358 756 21364 808
rect 21416 796 21422 808
rect 21521 799 21579 805
rect 21521 796 21533 799
rect 21416 768 21533 796
rect 21416 756 21422 768
rect 21521 765 21533 768
rect 21567 765 21579 799
rect 21521 759 21579 765
rect 24210 756 24216 808
rect 24268 756 24274 808
rect 18472 700 18644 728
rect 18708 700 20392 728
rect 18472 688 18478 700
rect 18509 663 18567 669
rect 18509 660 18521 663
rect 18012 632 18521 660
rect 18012 620 18018 632
rect 18509 629 18521 632
rect 18555 629 18567 663
rect 18616 660 18644 700
rect 22094 688 22100 740
rect 22152 728 22158 740
rect 23109 731 23167 737
rect 23109 728 23121 731
rect 22152 700 23121 728
rect 22152 688 22158 700
rect 23109 697 23121 700
rect 23155 697 23167 731
rect 23109 691 23167 697
rect 19705 663 19763 669
rect 19705 660 19717 663
rect 18616 632 19717 660
rect 18509 623 18567 629
rect 19705 629 19717 632
rect 19751 660 19763 663
rect 23382 660 23388 672
rect 19751 632 23388 660
rect 19751 629 19763 632
rect 19705 623 19763 629
rect 23382 620 23388 632
rect 23440 620 23446 672
rect 1104 570 33028 592
rect 1104 518 11610 570
rect 11662 518 11674 570
rect 11726 518 11738 570
rect 11790 518 11802 570
rect 11854 518 11866 570
rect 11918 518 21610 570
rect 21662 518 21674 570
rect 21726 518 21738 570
rect 21790 518 21802 570
rect 21854 518 21866 570
rect 21918 518 31610 570
rect 31662 518 31674 570
rect 31726 518 31738 570
rect 31790 518 31802 570
rect 31854 518 31866 570
rect 31918 518 33028 570
rect 1104 496 33028 518
rect 9398 416 9404 468
rect 9456 456 9462 468
rect 14642 456 14648 468
rect 9456 428 14648 456
rect 9456 416 9462 428
rect 14642 416 14648 428
rect 14700 416 14706 468
rect 15010 416 15016 468
rect 15068 456 15074 468
rect 23106 456 23112 468
rect 15068 428 23112 456
rect 15068 416 15074 428
rect 23106 416 23112 428
rect 23164 416 23170 468
rect 4246 348 4252 400
rect 4304 388 4310 400
rect 12250 388 12256 400
rect 4304 360 12256 388
rect 4304 348 4310 360
rect 12250 348 12256 360
rect 12308 348 12314 400
rect 12406 360 13124 388
rect 8110 280 8116 332
rect 8168 320 8174 332
rect 11974 320 11980 332
rect 8168 292 11980 320
rect 8168 280 8174 292
rect 11974 280 11980 292
rect 12032 280 12038 332
rect 12406 320 12434 360
rect 12268 292 12434 320
rect 4154 212 4160 264
rect 4212 252 4218 264
rect 12268 252 12296 292
rect 4212 224 12296 252
rect 4212 212 4218 224
rect 12342 212 12348 264
rect 12400 252 12406 264
rect 12986 252 12992 264
rect 12400 224 12992 252
rect 12400 212 12406 224
rect 12986 212 12992 224
rect 13044 212 13050 264
rect 13096 252 13124 360
rect 13170 348 13176 400
rect 13228 388 13234 400
rect 18966 388 18972 400
rect 13228 360 18972 388
rect 13228 348 13234 360
rect 18966 348 18972 360
rect 19024 348 19030 400
rect 13538 280 13544 332
rect 13596 320 13602 332
rect 22002 320 22008 332
rect 13596 292 22008 320
rect 13596 280 13602 292
rect 22002 280 22008 292
rect 22060 280 22066 332
rect 21358 252 21364 264
rect 13096 224 21364 252
rect 21358 212 21364 224
rect 21416 212 21422 264
rect 6638 144 6644 196
rect 6696 184 6702 196
rect 13998 184 14004 196
rect 6696 156 14004 184
rect 6696 144 6702 156
rect 13998 144 14004 156
rect 14056 144 14062 196
rect 14826 144 14832 196
rect 14884 184 14890 196
rect 20806 184 20812 196
rect 14884 156 20812 184
rect 14884 144 14890 156
rect 20806 144 20812 156
rect 20864 144 20870 196
rect 8662 76 8668 128
rect 8720 116 8726 128
rect 14090 116 14096 128
rect 8720 88 14096 116
rect 8720 76 8726 88
rect 14090 76 14096 88
rect 14148 76 14154 128
rect 4982 8 4988 60
rect 5040 48 5046 60
rect 9950 48 9956 60
rect 5040 20 9956 48
rect 5040 8 5046 20
rect 9950 8 9956 20
rect 10008 8 10014 60
rect 10042 8 10048 60
rect 10100 48 10106 60
rect 14458 48 14464 60
rect 10100 20 14464 48
rect 10100 8 10106 20
rect 14458 8 14464 20
rect 14516 8 14522 60
<< via1 >>
rect 4160 11908 4212 11960
rect 22376 11908 22428 11960
rect 30196 11908 30248 11960
rect 3700 11840 3752 11892
rect 12440 11840 12492 11892
rect 12532 11840 12584 11892
rect 20444 11840 20496 11892
rect 1032 11704 1084 11756
rect 3792 11772 3844 11824
rect 3976 11772 4028 11824
rect 20628 11772 20680 11824
rect 2136 11636 2188 11688
rect 12900 11704 12952 11756
rect 12992 11704 13044 11756
rect 14924 11704 14976 11756
rect 3884 11636 3936 11688
rect 21916 11704 21968 11756
rect 30748 11840 30800 11892
rect 15200 11636 15252 11688
rect 22928 11636 22980 11688
rect 29920 11636 29972 11688
rect 940 11568 992 11620
rect 3056 11568 3108 11620
rect 4068 11568 4120 11620
rect 12348 11568 12400 11620
rect 12440 11568 12492 11620
rect 21456 11568 21508 11620
rect 21824 11568 21876 11620
rect 25688 11568 25740 11620
rect 2780 11500 2832 11552
rect 4712 11500 4764 11552
rect 4804 11500 4856 11552
rect 7288 11500 7340 11552
rect 9680 11500 9732 11552
rect 12072 11500 12124 11552
rect 12164 11500 12216 11552
rect 12992 11500 13044 11552
rect 13084 11500 13136 11552
rect 14556 11500 14608 11552
rect 15936 11500 15988 11552
rect 17408 11500 17460 11552
rect 18052 11500 18104 11552
rect 20260 11500 20312 11552
rect 21364 11500 21416 11552
rect 23940 11500 23992 11552
rect 11610 11398 11662 11450
rect 11674 11398 11726 11450
rect 11738 11398 11790 11450
rect 11802 11398 11854 11450
rect 11866 11398 11918 11450
rect 21610 11398 21662 11450
rect 21674 11398 21726 11450
rect 21738 11398 21790 11450
rect 21802 11398 21854 11450
rect 21866 11398 21918 11450
rect 31610 11398 31662 11450
rect 31674 11398 31726 11450
rect 31738 11398 31790 11450
rect 31802 11398 31854 11450
rect 31866 11398 31918 11450
rect 24124 11296 24176 11348
rect 27712 11296 27764 11348
rect 29920 11339 29972 11348
rect 29920 11305 29929 11339
rect 29929 11305 29963 11339
rect 29963 11305 29972 11339
rect 29920 11296 29972 11305
rect 1584 11160 1636 11212
rect 3700 11203 3752 11212
rect 3700 11169 3709 11203
rect 3709 11169 3743 11203
rect 3743 11169 3752 11203
rect 3700 11160 3752 11169
rect 4804 11237 4856 11246
rect 4804 11203 4813 11237
rect 4813 11203 4847 11237
rect 4847 11203 4856 11237
rect 4804 11194 4856 11203
rect 6460 11203 6512 11212
rect 6460 11169 6469 11203
rect 6469 11169 6503 11203
rect 6503 11169 6512 11203
rect 6460 11160 6512 11169
rect 7288 11203 7340 11212
rect 7288 11169 7297 11203
rect 7297 11169 7331 11203
rect 7331 11169 7340 11203
rect 7288 11160 7340 11169
rect 9404 11160 9456 11212
rect 9956 11203 10008 11212
rect 9956 11169 9965 11203
rect 9965 11169 9999 11203
rect 9999 11169 10008 11203
rect 9956 11160 10008 11169
rect 12072 11228 12124 11280
rect 12164 11160 12216 11212
rect 14556 11237 14608 11246
rect 14556 11203 14565 11237
rect 14565 11203 14599 11237
rect 14599 11203 14608 11237
rect 14556 11194 14608 11203
rect 15660 11203 15712 11212
rect 15660 11169 15669 11203
rect 15669 11169 15703 11203
rect 15703 11169 15712 11203
rect 15660 11160 15712 11169
rect 17408 11237 17460 11246
rect 17408 11203 17417 11237
rect 17417 11203 17451 11237
rect 17451 11203 17460 11237
rect 17408 11194 17460 11203
rect 17776 11160 17828 11212
rect 20260 11237 20312 11246
rect 20260 11203 20269 11237
rect 20269 11203 20303 11237
rect 20303 11203 20312 11237
rect 20260 11194 20312 11203
rect 21364 11228 21416 11280
rect 23112 11160 23164 11212
rect 24032 11092 24084 11144
rect 25136 11092 25188 11144
rect 25320 11203 25372 11212
rect 25320 11169 25329 11203
rect 25329 11169 25363 11203
rect 25363 11169 25372 11203
rect 25320 11160 25372 11169
rect 25872 11160 25924 11212
rect 26884 11160 26936 11212
rect 27252 11203 27304 11212
rect 27252 11169 27261 11203
rect 27261 11169 27295 11203
rect 27295 11169 27304 11203
rect 27252 11160 27304 11169
rect 27896 11203 27948 11212
rect 27896 11169 27905 11203
rect 27905 11169 27939 11203
rect 27939 11169 27948 11203
rect 27896 11160 27948 11169
rect 23388 11024 23440 11076
rect 26240 11135 26292 11144
rect 26240 11101 26249 11135
rect 26249 11101 26283 11135
rect 26283 11101 26292 11135
rect 26240 11092 26292 11101
rect 23480 10956 23532 11008
rect 24308 10956 24360 11008
rect 10950 10854 11002 10906
rect 11014 10854 11066 10906
rect 11078 10854 11130 10906
rect 11142 10854 11194 10906
rect 11206 10854 11258 10906
rect 20950 10854 21002 10906
rect 21014 10854 21066 10906
rect 21078 10854 21130 10906
rect 21142 10854 21194 10906
rect 21206 10854 21258 10906
rect 30950 10854 31002 10906
rect 31014 10854 31066 10906
rect 31078 10854 31130 10906
rect 31142 10854 31194 10906
rect 31206 10854 31258 10906
rect 30196 10795 30248 10804
rect 30196 10761 30205 10795
rect 30205 10761 30239 10795
rect 30239 10761 30248 10795
rect 30196 10752 30248 10761
rect 30748 10795 30800 10804
rect 30748 10761 30757 10795
rect 30757 10761 30791 10795
rect 30791 10761 30800 10795
rect 30748 10752 30800 10761
rect 17592 10616 17644 10668
rect 1584 10591 1636 10600
rect 1584 10557 1593 10591
rect 1593 10557 1627 10591
rect 1627 10557 1636 10591
rect 1584 10548 1636 10557
rect 6460 10557 6512 10566
rect 6460 10523 6469 10557
rect 6469 10523 6503 10557
rect 6503 10523 6512 10557
rect 6460 10514 6512 10523
rect 7656 10557 7708 10566
rect 7656 10523 7665 10557
rect 7665 10523 7699 10557
rect 7699 10523 7708 10557
rect 7656 10514 7708 10523
rect 9404 10591 9456 10600
rect 9404 10557 9413 10591
rect 9413 10557 9447 10591
rect 9447 10557 9456 10591
rect 9404 10548 9456 10557
rect 10784 10548 10836 10600
rect 12532 10480 12584 10532
rect 13360 10557 13412 10566
rect 13360 10523 13369 10557
rect 13369 10523 13403 10557
rect 13403 10523 13412 10557
rect 13360 10514 13412 10523
rect 15016 10591 15068 10600
rect 15016 10557 15025 10591
rect 15025 10557 15059 10591
rect 15059 10557 15068 10591
rect 15016 10548 15068 10557
rect 16304 10557 16356 10566
rect 16304 10523 16313 10557
rect 16313 10523 16347 10557
rect 16347 10523 16356 10557
rect 16304 10514 16356 10523
rect 18052 10591 18104 10600
rect 18052 10557 18061 10591
rect 18061 10557 18095 10591
rect 18095 10557 18104 10591
rect 18052 10548 18104 10557
rect 20720 10616 20772 10668
rect 23112 10557 23164 10566
rect 23112 10523 23121 10557
rect 23121 10523 23155 10557
rect 23155 10523 23164 10557
rect 23112 10514 23164 10523
rect 23940 10591 23992 10600
rect 23940 10557 23949 10591
rect 23949 10557 23983 10591
rect 23983 10557 23992 10591
rect 23940 10548 23992 10557
rect 25688 10557 25740 10566
rect 25688 10523 25697 10557
rect 25697 10523 25731 10557
rect 25731 10523 25740 10557
rect 25688 10514 25740 10523
rect 22008 10412 22060 10464
rect 26056 10412 26108 10464
rect 29920 10480 29972 10532
rect 28356 10412 28408 10464
rect 11610 10310 11662 10362
rect 11674 10310 11726 10362
rect 11738 10310 11790 10362
rect 11802 10310 11854 10362
rect 11866 10310 11918 10362
rect 21610 10310 21662 10362
rect 21674 10310 21726 10362
rect 21738 10310 21790 10362
rect 21802 10310 21854 10362
rect 21866 10310 21918 10362
rect 31610 10310 31662 10362
rect 31674 10310 31726 10362
rect 31738 10310 31790 10362
rect 31802 10310 31854 10362
rect 31866 10310 31918 10362
rect 17960 10208 18012 10260
rect 19064 10208 19116 10260
rect 2228 10149 2280 10158
rect 2228 10115 2237 10149
rect 2237 10115 2271 10149
rect 2271 10115 2280 10149
rect 2228 10106 2280 10115
rect 4160 10072 4212 10124
rect 3516 10004 3568 10056
rect 6828 10072 6880 10124
rect 7196 10072 7248 10124
rect 9956 10140 10008 10192
rect 9772 10072 9824 10124
rect 11980 10106 12032 10158
rect 12532 10072 12584 10124
rect 15016 10149 15068 10158
rect 15016 10115 15025 10149
rect 15025 10115 15059 10149
rect 15059 10115 15068 10149
rect 15016 10106 15068 10115
rect 15936 10115 15988 10124
rect 15936 10081 15945 10115
rect 15945 10081 15979 10115
rect 15979 10081 15988 10115
rect 15936 10072 15988 10081
rect 18052 10140 18104 10192
rect 19800 10072 19852 10124
rect 20536 10208 20588 10260
rect 22008 10208 22060 10260
rect 22100 10140 22152 10192
rect 23388 10140 23440 10192
rect 22008 10072 22060 10124
rect 24124 10072 24176 10124
rect 24216 10115 24268 10124
rect 24216 10081 24225 10115
rect 24225 10081 24259 10115
rect 24259 10081 24268 10115
rect 24216 10072 24268 10081
rect 25964 10149 26016 10158
rect 25964 10115 25973 10149
rect 25973 10115 26007 10149
rect 26007 10115 26016 10149
rect 25964 10106 26016 10115
rect 26792 10115 26844 10124
rect 26792 10081 26801 10115
rect 26801 10081 26835 10115
rect 26835 10081 26844 10115
rect 26792 10072 26844 10081
rect 28540 10149 28592 10158
rect 28540 10115 28549 10149
rect 28549 10115 28583 10149
rect 28583 10115 28592 10149
rect 28540 10106 28592 10115
rect 29920 10115 29972 10124
rect 29920 10081 29929 10115
rect 29929 10081 29963 10115
rect 29963 10081 29972 10115
rect 29920 10072 29972 10081
rect 32036 10072 32088 10124
rect 20260 10004 20312 10056
rect 22376 10047 22428 10056
rect 22376 10013 22385 10047
rect 22385 10013 22419 10047
rect 22419 10013 22428 10047
rect 22376 10004 22428 10013
rect 22100 9936 22152 9988
rect 24124 9936 24176 9988
rect 18052 9868 18104 9920
rect 18972 9868 19024 9920
rect 19156 9868 19208 9920
rect 10950 9766 11002 9818
rect 11014 9766 11066 9818
rect 11078 9766 11130 9818
rect 11142 9766 11194 9818
rect 11206 9766 11258 9818
rect 20950 9766 21002 9818
rect 21014 9766 21066 9818
rect 21078 9766 21130 9818
rect 21142 9766 21194 9818
rect 21206 9766 21258 9818
rect 30950 9766 31002 9818
rect 31014 9766 31066 9818
rect 31078 9766 31130 9818
rect 31142 9766 31194 9818
rect 31206 9766 31258 9818
rect 15200 9664 15252 9716
rect 17224 9664 17276 9716
rect 21456 9664 21508 9716
rect 19340 9596 19392 9648
rect 19892 9639 19944 9648
rect 19892 9605 19901 9639
rect 19901 9605 19935 9639
rect 19935 9605 19944 9639
rect 19892 9596 19944 9605
rect 3516 9528 3568 9580
rect 1952 9469 2004 9478
rect 1952 9435 1961 9469
rect 1961 9435 1995 9469
rect 1995 9435 2004 9469
rect 1952 9426 2004 9435
rect 3700 9503 3752 9512
rect 3700 9469 3709 9503
rect 3709 9469 3743 9503
rect 3743 9469 3752 9503
rect 3700 9460 3752 9469
rect 4160 9460 4212 9512
rect 6920 9528 6972 9580
rect 7196 9460 7248 9512
rect 9772 9528 9824 9580
rect 10784 9528 10836 9580
rect 15844 9571 15896 9580
rect 15844 9537 15853 9571
rect 15853 9537 15887 9571
rect 15887 9537 15896 9571
rect 15844 9528 15896 9537
rect 16212 9528 16264 9580
rect 17592 9528 17644 9580
rect 12164 9469 12216 9478
rect 12164 9435 12173 9469
rect 12173 9435 12207 9469
rect 12207 9435 12216 9469
rect 12164 9426 12216 9435
rect 13084 9503 13136 9512
rect 13084 9469 13093 9503
rect 13093 9469 13127 9503
rect 13127 9469 13136 9503
rect 13084 9460 13136 9469
rect 15660 9460 15712 9512
rect 17040 9392 17092 9444
rect 5448 9324 5500 9376
rect 15936 9367 15988 9376
rect 15936 9333 15945 9367
rect 15945 9333 15979 9367
rect 15979 9333 15988 9367
rect 15936 9324 15988 9333
rect 16948 9324 17000 9376
rect 18880 9469 18932 9478
rect 18880 9435 18889 9469
rect 18889 9435 18923 9469
rect 18923 9435 18932 9469
rect 18880 9426 18932 9435
rect 19248 9392 19300 9444
rect 20628 9503 20680 9512
rect 20628 9469 20637 9503
rect 20637 9469 20671 9503
rect 20671 9469 20680 9503
rect 20628 9460 20680 9469
rect 21364 9460 21416 9512
rect 17684 9324 17736 9376
rect 23112 9469 23164 9478
rect 23112 9435 23121 9469
rect 23121 9435 23155 9469
rect 23155 9435 23164 9469
rect 23112 9426 23164 9435
rect 22008 9324 22060 9376
rect 26792 9460 26844 9512
rect 27436 9469 27488 9478
rect 27436 9435 27445 9469
rect 27445 9435 27479 9469
rect 27479 9435 27488 9469
rect 27436 9426 27488 9435
rect 29184 9503 29236 9512
rect 29184 9469 29193 9503
rect 29193 9469 29227 9503
rect 29227 9469 29236 9503
rect 29184 9460 29236 9469
rect 29644 9503 29696 9512
rect 29644 9469 29653 9503
rect 29653 9469 29687 9503
rect 29687 9469 29696 9503
rect 29644 9460 29696 9469
rect 31392 9469 31444 9478
rect 31392 9435 31401 9469
rect 31401 9435 31435 9469
rect 31435 9435 31444 9469
rect 31392 9426 31444 9435
rect 25136 9324 25188 9376
rect 11610 9222 11662 9274
rect 11674 9222 11726 9274
rect 11738 9222 11790 9274
rect 11802 9222 11854 9274
rect 11866 9222 11918 9274
rect 21610 9222 21662 9274
rect 21674 9222 21726 9274
rect 21738 9222 21790 9274
rect 21802 9222 21854 9274
rect 21866 9222 21918 9274
rect 31610 9222 31662 9274
rect 31674 9222 31726 9274
rect 31738 9222 31790 9274
rect 31802 9222 31854 9274
rect 31866 9222 31918 9274
rect 5724 9120 5776 9172
rect 1860 9018 1912 9070
rect 3792 8984 3844 9036
rect 4712 9061 4764 9070
rect 4712 9027 4721 9061
rect 4721 9027 4755 9061
rect 4755 9027 4764 9061
rect 4712 9018 4764 9027
rect 6644 9120 6696 9172
rect 9496 9120 9548 9172
rect 11980 9120 12032 9172
rect 9404 9052 9456 9104
rect 6920 8984 6972 9036
rect 9588 9027 9640 9036
rect 9588 8993 9597 9027
rect 9597 8993 9631 9027
rect 9631 8993 9640 9027
rect 9588 8984 9640 8993
rect 11336 9061 11388 9070
rect 11336 9027 11345 9061
rect 11345 9027 11379 9061
rect 11379 9027 11388 9061
rect 11336 9018 11388 9027
rect 11428 9018 11480 9070
rect 12532 8984 12584 9036
rect 13268 9027 13320 9036
rect 13268 8993 13277 9027
rect 13277 8993 13311 9027
rect 13311 8993 13320 9027
rect 13268 8984 13320 8993
rect 15016 9061 15068 9070
rect 15016 9027 15025 9061
rect 15025 9027 15059 9061
rect 15059 9027 15068 9061
rect 15016 9018 15068 9027
rect 16212 9061 16264 9070
rect 16212 9027 16221 9061
rect 16221 9027 16255 9061
rect 16255 9027 16264 9061
rect 16212 9018 16264 9027
rect 18696 8984 18748 9036
rect 20536 9061 20588 9070
rect 20536 9027 20545 9061
rect 20545 9027 20579 9061
rect 20579 9027 20588 9061
rect 20536 9018 20588 9027
rect 22284 9120 22336 9172
rect 27436 9120 27488 9172
rect 29644 9120 29696 9172
rect 24216 9052 24268 9104
rect 8208 8916 8260 8968
rect 8484 8959 8536 8968
rect 8484 8925 8493 8959
rect 8493 8925 8527 8959
rect 8527 8925 8536 8959
rect 8484 8916 8536 8925
rect 10048 8916 10100 8968
rect 17592 8916 17644 8968
rect 24400 9027 24452 9036
rect 24400 8993 24409 9027
rect 24409 8993 24443 9027
rect 24443 8993 24452 9027
rect 24400 8984 24452 8993
rect 24584 8984 24636 9036
rect 27712 9095 27764 9104
rect 27712 9061 27721 9095
rect 27721 9061 27755 9095
rect 27755 9061 27764 9095
rect 27712 9052 27764 9061
rect 27160 8984 27212 9036
rect 27252 8984 27304 9036
rect 30656 9120 30708 9172
rect 9680 8848 9732 8900
rect 17868 8848 17920 8900
rect 19248 8916 19300 8968
rect 21364 8916 21416 8968
rect 22008 8916 22060 8968
rect 24124 8916 24176 8968
rect 27620 8916 27672 8968
rect 32128 8984 32180 9036
rect 28540 8916 28592 8968
rect 27252 8848 27304 8900
rect 29276 8848 29328 8900
rect 9312 8780 9364 8832
rect 11980 8780 12032 8832
rect 12624 8780 12676 8832
rect 23756 8780 23808 8832
rect 24768 8780 24820 8832
rect 28356 8823 28408 8832
rect 28356 8789 28365 8823
rect 28365 8789 28399 8823
rect 28399 8789 28408 8823
rect 28356 8780 28408 8789
rect 10950 8678 11002 8730
rect 11014 8678 11066 8730
rect 11078 8678 11130 8730
rect 11142 8678 11194 8730
rect 11206 8678 11258 8730
rect 20950 8678 21002 8730
rect 21014 8678 21066 8730
rect 21078 8678 21130 8730
rect 21142 8678 21194 8730
rect 21206 8678 21258 8730
rect 30950 8678 31002 8730
rect 31014 8678 31066 8730
rect 31078 8678 31130 8730
rect 31142 8678 31194 8730
rect 31206 8678 31258 8730
rect 5172 8440 5224 8492
rect 14648 8440 14700 8492
rect 1768 8338 1820 8390
rect 4712 8415 4764 8424
rect 4712 8381 4721 8415
rect 4721 8381 4755 8415
rect 4755 8381 4764 8415
rect 4712 8372 4764 8381
rect 9588 8372 9640 8424
rect 10692 8254 10744 8306
rect 12256 8338 12308 8390
rect 13360 8381 13412 8390
rect 13360 8347 13369 8381
rect 13369 8347 13403 8381
rect 13403 8347 13412 8381
rect 13360 8338 13412 8347
rect 15016 8415 15068 8424
rect 15016 8381 15025 8415
rect 15025 8381 15059 8415
rect 15059 8381 15068 8415
rect 15016 8372 15068 8381
rect 17684 8381 17736 8390
rect 17684 8347 17693 8381
rect 17693 8347 17727 8381
rect 17727 8347 17736 8381
rect 17684 8338 17736 8347
rect 18880 8372 18932 8424
rect 20260 8381 20312 8390
rect 20260 8347 20269 8381
rect 20269 8347 20303 8381
rect 20303 8347 20312 8381
rect 20260 8338 20312 8347
rect 27160 8415 27212 8424
rect 27160 8381 27169 8415
rect 27169 8381 27203 8415
rect 27203 8381 27212 8415
rect 27160 8372 27212 8381
rect 26056 8304 26108 8356
rect 28816 8381 28868 8390
rect 28816 8347 28825 8381
rect 28825 8347 28859 8381
rect 28859 8347 28868 8381
rect 28816 8338 28868 8347
rect 29276 8372 29328 8424
rect 32128 8415 32180 8424
rect 32128 8381 32137 8415
rect 32137 8381 32171 8415
rect 32171 8381 32180 8415
rect 32128 8372 32180 8381
rect 22008 8236 22060 8288
rect 11610 8134 11662 8186
rect 11674 8134 11726 8186
rect 11738 8134 11790 8186
rect 11802 8134 11854 8186
rect 11866 8134 11918 8186
rect 21610 8134 21662 8186
rect 21674 8134 21726 8186
rect 21738 8134 21790 8186
rect 21802 8134 21854 8186
rect 21866 8134 21918 8186
rect 31610 8134 31662 8186
rect 31674 8134 31726 8186
rect 31738 8134 31790 8186
rect 31802 8134 31854 8186
rect 31866 8134 31918 8186
rect 11428 8032 11480 8084
rect 13636 8032 13688 8084
rect 2044 7930 2096 7982
rect 3884 7939 3936 7948
rect 3884 7905 3893 7939
rect 3893 7905 3927 7939
rect 3927 7905 3936 7939
rect 3884 7896 3936 7905
rect 4344 7939 4396 7948
rect 4344 7905 4353 7939
rect 4353 7905 4387 7939
rect 4387 7905 4396 7939
rect 4344 7896 4396 7905
rect 6920 7964 6972 8016
rect 7288 7964 7340 8016
rect 8760 7964 8812 8016
rect 6552 7896 6604 7948
rect 7288 7871 7340 7880
rect 7288 7837 7297 7871
rect 7297 7837 7331 7871
rect 7331 7837 7340 7871
rect 7288 7828 7340 7837
rect 9312 7896 9364 7948
rect 9404 7939 9456 7948
rect 9404 7905 9413 7939
rect 9413 7905 9447 7939
rect 9447 7905 9456 7939
rect 9404 7896 9456 7905
rect 11520 7964 11572 8016
rect 11980 7896 12032 7948
rect 13728 7896 13780 7948
rect 14464 8032 14516 8084
rect 15844 8032 15896 8084
rect 17960 8032 18012 8084
rect 15476 7973 15528 7982
rect 15476 7939 15485 7973
rect 15485 7939 15519 7973
rect 15519 7939 15528 7973
rect 15476 7930 15528 7939
rect 19156 7964 19208 8016
rect 6828 7760 6880 7812
rect 8760 7871 8812 7880
rect 8760 7837 8769 7871
rect 8769 7837 8803 7871
rect 8803 7837 8812 7871
rect 8760 7828 8812 7837
rect 9220 7828 9272 7880
rect 9772 7828 9824 7880
rect 12624 7828 12676 7880
rect 12716 7828 12768 7880
rect 14188 7828 14240 7880
rect 11520 7760 11572 7812
rect 12072 7760 12124 7812
rect 17132 7896 17184 7948
rect 19248 7896 19300 7948
rect 17500 7760 17552 7812
rect 17592 7803 17644 7812
rect 17592 7769 17601 7803
rect 17601 7769 17635 7803
rect 17635 7769 17644 7803
rect 17592 7760 17644 7769
rect 17960 7871 18012 7880
rect 17960 7837 17969 7871
rect 17969 7837 18003 7871
rect 18003 7837 18012 7871
rect 17960 7828 18012 7837
rect 18512 7803 18564 7812
rect 18512 7769 18521 7803
rect 18521 7769 18555 7803
rect 18555 7769 18564 7803
rect 18512 7760 18564 7769
rect 18604 7803 18656 7812
rect 18604 7769 18613 7803
rect 18613 7769 18647 7803
rect 18647 7769 18656 7803
rect 18604 7760 18656 7769
rect 18972 7871 19024 7880
rect 18972 7837 18981 7871
rect 18981 7837 19015 7871
rect 19015 7837 19024 7871
rect 18972 7828 19024 7837
rect 22192 8032 22244 8084
rect 24216 8032 24268 8084
rect 25596 8032 25648 8084
rect 20260 7896 20312 7948
rect 22008 7964 22060 8016
rect 22100 7964 22152 8016
rect 23296 7896 23348 7948
rect 24584 7973 24636 7982
rect 24584 7939 24593 7973
rect 24593 7939 24627 7973
rect 24627 7939 24636 7973
rect 24584 7930 24636 7939
rect 20076 7828 20128 7880
rect 22744 7871 22796 7880
rect 22744 7837 22753 7871
rect 22753 7837 22787 7871
rect 22787 7837 22796 7871
rect 22744 7828 22796 7837
rect 26884 8075 26936 8084
rect 26884 8041 26893 8075
rect 26893 8041 26927 8075
rect 26927 8041 26936 8075
rect 26884 8032 26936 8041
rect 28540 8075 28592 8084
rect 28540 8041 28549 8075
rect 28549 8041 28583 8075
rect 28583 8041 28592 8075
rect 28540 8032 28592 8041
rect 29184 7964 29236 8016
rect 26056 7896 26108 7948
rect 26976 7939 27028 7948
rect 26976 7905 26985 7939
rect 26985 7905 27019 7939
rect 27019 7905 27028 7939
rect 26976 7896 27028 7905
rect 32036 7896 32088 7948
rect 29920 7828 29972 7880
rect 19892 7760 19944 7812
rect 22468 7760 22520 7812
rect 24124 7760 24176 7812
rect 26332 7760 26384 7812
rect 12440 7692 12492 7744
rect 12532 7692 12584 7744
rect 13268 7692 13320 7744
rect 13728 7692 13780 7744
rect 15936 7692 15988 7744
rect 19708 7692 19760 7744
rect 22376 7735 22428 7744
rect 22376 7701 22385 7735
rect 22385 7701 22419 7735
rect 22419 7701 22428 7735
rect 22376 7692 22428 7701
rect 23204 7735 23256 7744
rect 23204 7701 23213 7735
rect 23213 7701 23247 7735
rect 23247 7701 23256 7735
rect 23204 7692 23256 7701
rect 26240 7692 26292 7744
rect 28264 7692 28316 7744
rect 10950 7590 11002 7642
rect 11014 7590 11066 7642
rect 11078 7590 11130 7642
rect 11142 7590 11194 7642
rect 11206 7590 11258 7642
rect 20950 7590 21002 7642
rect 21014 7590 21066 7642
rect 21078 7590 21130 7642
rect 21142 7590 21194 7642
rect 21206 7590 21258 7642
rect 30950 7590 31002 7642
rect 31014 7590 31066 7642
rect 31078 7590 31130 7642
rect 31142 7590 31194 7642
rect 31206 7590 31258 7642
rect 1952 7488 2004 7540
rect 4160 7488 4212 7540
rect 10232 7488 10284 7540
rect 11428 7488 11480 7540
rect 11980 7488 12032 7540
rect 12348 7488 12400 7540
rect 14464 7488 14516 7540
rect 17132 7488 17184 7540
rect 19248 7488 19300 7540
rect 22376 7488 22428 7540
rect 25136 7531 25188 7540
rect 25136 7497 25145 7531
rect 25145 7497 25179 7531
rect 25179 7497 25188 7531
rect 25136 7488 25188 7497
rect 27068 7531 27120 7540
rect 27068 7497 27077 7531
rect 27077 7497 27111 7531
rect 27111 7497 27120 7531
rect 27068 7488 27120 7497
rect 1768 7420 1820 7472
rect 4344 7420 4396 7472
rect 9772 7420 9824 7472
rect 2688 7352 2740 7404
rect 3056 7395 3108 7404
rect 3056 7361 3065 7395
rect 3065 7361 3099 7395
rect 3099 7361 3108 7395
rect 3056 7352 3108 7361
rect 6368 7352 6420 7404
rect 1860 7284 1912 7336
rect 2596 7216 2648 7268
rect 5080 7293 5132 7302
rect 5080 7259 5089 7293
rect 5089 7259 5123 7293
rect 5123 7259 5132 7293
rect 5080 7250 5132 7259
rect 6828 7327 6880 7336
rect 6828 7293 6837 7327
rect 6837 7293 6871 7327
rect 6871 7293 6880 7327
rect 6828 7284 6880 7293
rect 9404 7284 9456 7336
rect 10600 7395 10652 7404
rect 10600 7361 10609 7395
rect 10609 7361 10643 7395
rect 10643 7361 10652 7395
rect 10600 7352 10652 7361
rect 11520 7420 11572 7472
rect 14648 7420 14700 7472
rect 17040 7420 17092 7472
rect 19616 7463 19668 7472
rect 19616 7429 19625 7463
rect 19625 7429 19659 7463
rect 19659 7429 19668 7463
rect 19616 7420 19668 7429
rect 19708 7463 19760 7472
rect 19708 7429 19717 7463
rect 19717 7429 19751 7463
rect 19751 7429 19760 7463
rect 19708 7420 19760 7429
rect 12716 7352 12768 7404
rect 12164 7284 12216 7336
rect 12256 7327 12308 7336
rect 12256 7293 12265 7327
rect 12265 7293 12299 7327
rect 12299 7293 12308 7327
rect 12256 7284 12308 7293
rect 14004 7293 14056 7302
rect 14004 7259 14013 7293
rect 14013 7259 14047 7293
rect 14047 7259 14056 7293
rect 14004 7250 14056 7259
rect 14832 7327 14884 7336
rect 14832 7293 14841 7327
rect 14841 7293 14875 7327
rect 14875 7293 14884 7327
rect 14832 7284 14884 7293
rect 1584 7191 1636 7200
rect 1584 7157 1593 7191
rect 1593 7157 1627 7191
rect 1627 7157 1636 7191
rect 1584 7148 1636 7157
rect 3700 7148 3752 7200
rect 4436 7148 4488 7200
rect 9496 7148 9548 7200
rect 14372 7216 14424 7268
rect 15568 7216 15620 7268
rect 16580 7284 16632 7336
rect 17132 7327 17184 7336
rect 17132 7293 17141 7327
rect 17141 7293 17175 7327
rect 17175 7293 17184 7327
rect 17132 7284 17184 7293
rect 16764 7216 16816 7268
rect 11980 7148 12032 7200
rect 18788 7293 18840 7302
rect 18788 7259 18797 7293
rect 18797 7259 18831 7293
rect 18831 7259 18840 7293
rect 18788 7250 18840 7259
rect 19156 7284 19208 7336
rect 20076 7395 20128 7404
rect 20076 7361 20085 7395
rect 20085 7361 20119 7395
rect 20119 7361 20128 7395
rect 20076 7352 20128 7361
rect 20812 7352 20864 7404
rect 20260 7284 20312 7336
rect 19248 7216 19300 7268
rect 20628 7216 20680 7268
rect 22468 7420 22520 7472
rect 22192 7352 22244 7404
rect 24400 7352 24452 7404
rect 28264 7488 28316 7540
rect 17776 7148 17828 7200
rect 19156 7148 19208 7200
rect 20812 7148 20864 7200
rect 24216 7284 24268 7336
rect 25412 7327 25464 7336
rect 25412 7293 25421 7327
rect 25421 7293 25455 7327
rect 25455 7293 25464 7327
rect 25412 7284 25464 7293
rect 25688 7284 25740 7336
rect 27620 7395 27672 7404
rect 27620 7361 27629 7395
rect 27629 7361 27663 7395
rect 27663 7361 27672 7395
rect 27620 7352 27672 7361
rect 26240 7284 26292 7336
rect 28356 7216 28408 7268
rect 24768 7148 24820 7200
rect 28540 7148 28592 7200
rect 28816 7148 28868 7200
rect 11610 7046 11662 7098
rect 11674 7046 11726 7098
rect 11738 7046 11790 7098
rect 11802 7046 11854 7098
rect 11866 7046 11918 7098
rect 21610 7046 21662 7098
rect 21674 7046 21726 7098
rect 21738 7046 21790 7098
rect 21802 7046 21854 7098
rect 21866 7046 21918 7098
rect 31610 7046 31662 7098
rect 31674 7046 31726 7098
rect 31738 7046 31790 7098
rect 31802 7046 31854 7098
rect 31866 7046 31918 7098
rect 2044 6944 2096 6996
rect 4068 6944 4120 6996
rect 9220 6944 9272 6996
rect 10140 6944 10192 6996
rect 11520 6944 11572 6996
rect 4436 6876 4488 6928
rect 4252 6808 4304 6860
rect 4344 6808 4396 6860
rect 4804 6885 4856 6894
rect 4804 6851 4813 6885
rect 4813 6851 4847 6885
rect 4847 6851 4856 6885
rect 4804 6842 4856 6851
rect 6552 6851 6604 6860
rect 6552 6817 6561 6851
rect 6561 6817 6595 6851
rect 6595 6817 6604 6851
rect 6552 6808 6604 6817
rect 8852 6885 8904 6894
rect 8852 6851 8861 6885
rect 8861 6851 8895 6885
rect 8895 6851 8904 6885
rect 8852 6842 8904 6851
rect 3424 6783 3476 6792
rect 3424 6749 3433 6783
rect 3433 6749 3467 6783
rect 3467 6749 3476 6783
rect 3424 6740 3476 6749
rect 6092 6740 6144 6792
rect 9312 6808 9364 6860
rect 17592 6944 17644 6996
rect 12348 6808 12400 6860
rect 12992 6808 13044 6860
rect 14556 6885 14608 6894
rect 14556 6851 14565 6885
rect 14565 6851 14599 6885
rect 14599 6851 14608 6885
rect 14556 6842 14608 6851
rect 15476 6851 15528 6860
rect 15476 6817 15485 6851
rect 15485 6817 15519 6851
rect 15519 6817 15528 6851
rect 15476 6808 15528 6817
rect 17132 6885 17184 6894
rect 17132 6851 17141 6885
rect 17141 6851 17175 6885
rect 17175 6851 17184 6885
rect 17132 6842 17184 6851
rect 13084 6740 13136 6792
rect 18788 6808 18840 6860
rect 19156 6944 19208 6996
rect 23296 6944 23348 6996
rect 22836 6885 22888 6894
rect 22836 6851 22845 6885
rect 22845 6851 22879 6885
rect 22879 6851 22888 6885
rect 22836 6842 22888 6851
rect 24124 6876 24176 6928
rect 28816 6944 28868 6996
rect 29920 6987 29972 6996
rect 29920 6953 29929 6987
rect 29929 6953 29963 6987
rect 29963 6953 29972 6987
rect 29920 6944 29972 6953
rect 23296 6740 23348 6792
rect 25228 6851 25280 6860
rect 25228 6817 25237 6851
rect 25237 6817 25271 6851
rect 25271 6817 25280 6851
rect 25228 6808 25280 6817
rect 25872 6851 25924 6860
rect 25872 6817 25881 6851
rect 25881 6817 25915 6851
rect 25915 6817 25924 6851
rect 25872 6808 25924 6817
rect 24768 6740 24820 6792
rect 4344 6672 4396 6724
rect 26332 6715 26384 6724
rect 26332 6681 26341 6715
rect 26341 6681 26375 6715
rect 26375 6681 26384 6715
rect 26332 6672 26384 6681
rect 29092 6715 29144 6724
rect 29092 6681 29101 6715
rect 29101 6681 29135 6715
rect 29135 6681 29144 6715
rect 29092 6672 29144 6681
rect 32036 6672 32088 6724
rect 3884 6604 3936 6656
rect 24860 6604 24912 6656
rect 26884 6647 26936 6656
rect 26884 6613 26893 6647
rect 26893 6613 26927 6647
rect 26927 6613 26936 6647
rect 26884 6604 26936 6613
rect 10950 6502 11002 6554
rect 11014 6502 11066 6554
rect 11078 6502 11130 6554
rect 11142 6502 11194 6554
rect 11206 6502 11258 6554
rect 20950 6502 21002 6554
rect 21014 6502 21066 6554
rect 21078 6502 21130 6554
rect 21142 6502 21194 6554
rect 21206 6502 21258 6554
rect 30950 6502 31002 6554
rect 31014 6502 31066 6554
rect 31078 6502 31130 6554
rect 31142 6502 31194 6554
rect 31206 6502 31258 6554
rect 4068 6400 4120 6452
rect 16948 6400 17000 6452
rect 17868 6400 17920 6452
rect 20168 6400 20220 6452
rect 30656 6443 30708 6452
rect 30656 6409 30665 6443
rect 30665 6409 30699 6443
rect 30699 6409 30708 6443
rect 30656 6400 30708 6409
rect 4160 6332 4212 6384
rect 15200 6332 15252 6384
rect 16580 6332 16632 6384
rect 16764 6332 16816 6384
rect 18052 6332 18104 6384
rect 2136 6239 2188 6248
rect 2136 6205 2145 6239
rect 2145 6205 2179 6239
rect 2179 6205 2188 6239
rect 2136 6196 2188 6205
rect 12624 6264 12676 6316
rect 13452 6264 13504 6316
rect 15292 6264 15344 6316
rect 4252 6196 4304 6248
rect 3884 6128 3936 6180
rect 4620 6205 4672 6214
rect 4620 6171 4629 6205
rect 4629 6171 4663 6205
rect 4663 6171 4672 6205
rect 4620 6162 4672 6171
rect 6828 6196 6880 6248
rect 6920 6196 6972 6248
rect 12808 6128 12860 6180
rect 2688 6060 2740 6112
rect 3332 6103 3384 6112
rect 3332 6069 3341 6103
rect 3341 6069 3375 6103
rect 3375 6069 3384 6103
rect 3332 6060 3384 6069
rect 3976 6060 4028 6112
rect 9404 6060 9456 6112
rect 10324 6060 10376 6112
rect 15384 6196 15436 6248
rect 27160 6307 27212 6316
rect 27160 6273 27169 6307
rect 27169 6273 27203 6307
rect 27203 6273 27212 6307
rect 27160 6264 27212 6273
rect 28540 6264 28592 6316
rect 17868 6196 17920 6248
rect 17960 6239 18012 6248
rect 17960 6205 17969 6239
rect 17969 6205 18003 6239
rect 18003 6205 18012 6239
rect 17960 6196 18012 6205
rect 15844 6128 15896 6180
rect 19708 6205 19760 6214
rect 19708 6171 19717 6205
rect 19717 6171 19751 6205
rect 19751 6171 19760 6205
rect 19708 6162 19760 6171
rect 20720 6239 20772 6248
rect 20720 6205 20729 6239
rect 20729 6205 20763 6239
rect 20763 6205 20772 6239
rect 20720 6196 20772 6205
rect 13728 6060 13780 6112
rect 15660 6103 15712 6112
rect 15660 6069 15669 6103
rect 15669 6069 15703 6103
rect 15703 6069 15712 6103
rect 15660 6060 15712 6069
rect 16580 6103 16632 6112
rect 16580 6069 16589 6103
rect 16589 6069 16623 6103
rect 16623 6069 16632 6103
rect 16580 6060 16632 6069
rect 24216 6196 24268 6248
rect 24308 6196 24360 6248
rect 27620 6196 27672 6248
rect 26792 6128 26844 6180
rect 29828 6205 29880 6214
rect 29828 6171 29837 6205
rect 29837 6171 29871 6205
rect 29871 6171 29880 6205
rect 29828 6162 29880 6171
rect 22008 6060 22060 6112
rect 11610 5958 11662 6010
rect 11674 5958 11726 6010
rect 11738 5958 11790 6010
rect 11802 5958 11854 6010
rect 11866 5958 11918 6010
rect 21610 5958 21662 6010
rect 21674 5958 21726 6010
rect 21738 5958 21790 6010
rect 21802 5958 21854 6010
rect 21866 5958 21918 6010
rect 31610 5958 31662 6010
rect 31674 5958 31726 6010
rect 31738 5958 31790 6010
rect 31802 5958 31854 6010
rect 31866 5958 31918 6010
rect 3608 5899 3660 5908
rect 3608 5865 3617 5899
rect 3617 5865 3651 5899
rect 3651 5865 3660 5899
rect 3608 5856 3660 5865
rect 3976 5899 4028 5908
rect 3976 5865 3985 5899
rect 3985 5865 4019 5899
rect 4019 5865 4028 5899
rect 3976 5856 4028 5865
rect 2412 5763 2464 5772
rect 2412 5729 2421 5763
rect 2421 5729 2455 5763
rect 2455 5729 2464 5763
rect 2412 5720 2464 5729
rect 2228 5695 2280 5704
rect 2228 5661 2237 5695
rect 2237 5661 2271 5695
rect 2271 5661 2280 5695
rect 2228 5652 2280 5661
rect 4344 5720 4396 5772
rect 4804 5797 4856 5806
rect 4804 5763 4813 5797
rect 4813 5763 4847 5797
rect 4847 5763 4856 5797
rect 4804 5754 4856 5763
rect 7196 5720 7248 5772
rect 4160 5652 4212 5704
rect 6092 5652 6144 5704
rect 9496 5720 9548 5772
rect 10508 5720 10560 5772
rect 12256 5720 12308 5772
rect 12808 5763 12860 5772
rect 12808 5729 12817 5763
rect 12817 5729 12851 5763
rect 12851 5729 12860 5763
rect 12808 5720 12860 5729
rect 14556 5797 14608 5806
rect 14556 5763 14565 5797
rect 14565 5763 14599 5797
rect 14599 5763 14608 5797
rect 14556 5754 14608 5763
rect 15844 5763 15896 5772
rect 15844 5729 15853 5763
rect 15853 5729 15887 5763
rect 15887 5729 15896 5763
rect 15844 5720 15896 5729
rect 17960 5788 18012 5840
rect 18052 5720 18104 5772
rect 19708 5720 19760 5772
rect 21456 5754 21508 5806
rect 22468 5763 22520 5772
rect 22468 5729 22477 5763
rect 22477 5729 22511 5763
rect 22511 5729 22520 5763
rect 22468 5720 22520 5729
rect 23112 5763 23164 5772
rect 23112 5729 23121 5763
rect 23121 5729 23155 5763
rect 23155 5729 23164 5763
rect 23112 5720 23164 5729
rect 23204 5763 23256 5772
rect 23204 5729 23213 5763
rect 23213 5729 23247 5763
rect 23247 5729 23256 5763
rect 23204 5720 23256 5729
rect 23480 5720 23532 5772
rect 25964 5797 26016 5806
rect 25964 5763 25973 5797
rect 25973 5763 26007 5797
rect 26007 5763 26016 5797
rect 25964 5754 26016 5763
rect 26792 5763 26844 5772
rect 26792 5729 26801 5763
rect 26801 5729 26835 5763
rect 26835 5729 26844 5763
rect 26792 5720 26844 5729
rect 28908 5720 28960 5772
rect 29828 5720 29880 5772
rect 32036 5788 32088 5840
rect 18696 5695 18748 5704
rect 18696 5661 18705 5695
rect 18705 5661 18739 5695
rect 18739 5661 18748 5695
rect 18696 5652 18748 5661
rect 19892 5652 19944 5704
rect 22744 5652 22796 5704
rect 3700 5584 3752 5636
rect 4252 5584 4304 5636
rect 22008 5584 22060 5636
rect 6460 5516 6512 5568
rect 7380 5516 7432 5568
rect 18052 5516 18104 5568
rect 19524 5516 19576 5568
rect 10950 5414 11002 5466
rect 11014 5414 11066 5466
rect 11078 5414 11130 5466
rect 11142 5414 11194 5466
rect 11206 5414 11258 5466
rect 20950 5414 21002 5466
rect 21014 5414 21066 5466
rect 21078 5414 21130 5466
rect 21142 5414 21194 5466
rect 21206 5414 21258 5466
rect 30950 5414 31002 5466
rect 31014 5414 31066 5466
rect 31078 5414 31130 5466
rect 31142 5414 31194 5466
rect 31206 5414 31258 5466
rect 4160 5312 4212 5364
rect 5448 5312 5500 5364
rect 15292 5312 15344 5364
rect 3884 5244 3936 5296
rect 5724 5244 5776 5296
rect 1584 5151 1636 5160
rect 1584 5117 1593 5151
rect 1593 5117 1627 5151
rect 1627 5117 1636 5151
rect 1584 5108 1636 5117
rect 2688 5108 2740 5160
rect 3700 5151 3752 5160
rect 3700 5117 3709 5151
rect 3709 5117 3743 5151
rect 3743 5117 3752 5151
rect 3700 5108 3752 5117
rect 4528 5219 4580 5228
rect 4528 5185 4537 5219
rect 4537 5185 4571 5219
rect 4571 5185 4580 5219
rect 4528 5176 4580 5185
rect 4620 5176 4672 5228
rect 7472 5176 7524 5228
rect 9680 5244 9732 5296
rect 15200 5244 15252 5296
rect 10048 5176 10100 5228
rect 17960 5312 18012 5364
rect 20076 5312 20128 5364
rect 1400 5040 1452 5092
rect 2228 4972 2280 5024
rect 4436 4972 4488 5024
rect 5264 5108 5316 5160
rect 5816 5108 5868 5160
rect 6184 5117 6236 5126
rect 6184 5083 6193 5117
rect 6193 5083 6227 5117
rect 6227 5083 6236 5117
rect 6184 5074 6236 5083
rect 7932 5151 7984 5160
rect 7932 5117 7941 5151
rect 7941 5117 7975 5151
rect 7975 5117 7984 5151
rect 7932 5108 7984 5117
rect 8024 5108 8076 5160
rect 9312 5108 9364 5160
rect 9496 5108 9548 5160
rect 9404 5040 9456 5092
rect 12072 5108 12124 5160
rect 12256 5108 12308 5160
rect 14740 5117 14792 5126
rect 14740 5083 14749 5117
rect 14749 5083 14783 5117
rect 14783 5083 14792 5117
rect 14740 5074 14792 5083
rect 15108 5108 15160 5160
rect 18328 5176 18380 5228
rect 20076 5176 20128 5228
rect 18144 5108 18196 5160
rect 15200 5040 15252 5092
rect 16488 5040 16540 5092
rect 17316 5083 17368 5092
rect 17316 5049 17325 5083
rect 17325 5049 17359 5083
rect 17359 5049 17368 5083
rect 17316 5040 17368 5049
rect 19616 5117 19668 5126
rect 19616 5083 19625 5117
rect 19625 5083 19659 5117
rect 19659 5083 19668 5117
rect 19616 5074 19668 5083
rect 19984 5108 20036 5160
rect 21456 5151 21508 5160
rect 21456 5117 21465 5151
rect 21465 5117 21499 5151
rect 21499 5117 21508 5151
rect 21456 5108 21508 5117
rect 23480 5108 23532 5160
rect 24308 5117 24360 5126
rect 24308 5083 24317 5117
rect 24317 5083 24351 5117
rect 24351 5083 24360 5117
rect 24308 5074 24360 5083
rect 25964 5151 26016 5160
rect 25964 5117 25973 5151
rect 25973 5117 26007 5151
rect 26007 5117 26016 5151
rect 25964 5108 26016 5117
rect 27436 5117 27488 5126
rect 27436 5083 27445 5117
rect 27445 5083 27479 5117
rect 27479 5083 27488 5117
rect 27436 5074 27488 5083
rect 4988 4972 5040 5024
rect 5172 4972 5224 5024
rect 5724 4972 5776 5024
rect 8668 5015 8720 5024
rect 8668 4981 8677 5015
rect 8677 4981 8711 5015
rect 8711 4981 8720 5015
rect 8668 4972 8720 4981
rect 15108 4972 15160 5024
rect 28448 4972 28500 5024
rect 28908 5108 28960 5160
rect 31484 4972 31536 5024
rect 11610 4870 11662 4922
rect 11674 4870 11726 4922
rect 11738 4870 11790 4922
rect 11802 4870 11854 4922
rect 11866 4870 11918 4922
rect 21610 4870 21662 4922
rect 21674 4870 21726 4922
rect 21738 4870 21790 4922
rect 21802 4870 21854 4922
rect 21866 4870 21918 4922
rect 31610 4870 31662 4922
rect 31674 4870 31726 4922
rect 31738 4870 31790 4922
rect 31802 4870 31854 4922
rect 31866 4870 31918 4922
rect 4712 4768 4764 4820
rect 5172 4768 5224 4820
rect 2228 4709 2280 4718
rect 2228 4675 2237 4709
rect 2237 4675 2271 4709
rect 2271 4675 2280 4709
rect 2228 4666 2280 4675
rect 3976 4675 4028 4684
rect 3976 4641 3985 4675
rect 3985 4641 4019 4675
rect 4019 4641 4028 4675
rect 3976 4632 4028 4641
rect 4436 4675 4488 4684
rect 4436 4641 4445 4675
rect 4445 4641 4479 4675
rect 4479 4641 4488 4675
rect 4436 4632 4488 4641
rect 6184 4709 6236 4718
rect 6184 4675 6193 4709
rect 6193 4675 6227 4709
rect 6227 4675 6236 4709
rect 6184 4666 6236 4675
rect 8300 4768 8352 4820
rect 9312 4709 9364 4718
rect 9312 4675 9321 4709
rect 9321 4675 9355 4709
rect 9355 4675 9364 4709
rect 9312 4666 9364 4675
rect 10600 4632 10652 4684
rect 6644 4564 6696 4616
rect 8024 4564 8076 4616
rect 12348 4564 12400 4616
rect 14004 4768 14056 4820
rect 23664 4811 23716 4820
rect 23664 4777 23673 4811
rect 23673 4777 23707 4811
rect 23707 4777 23716 4811
rect 23664 4768 23716 4777
rect 15016 4709 15068 4718
rect 15016 4675 15025 4709
rect 15025 4675 15059 4709
rect 15059 4675 15068 4709
rect 15016 4666 15068 4675
rect 16304 4632 16356 4684
rect 18144 4700 18196 4752
rect 18052 4632 18104 4684
rect 19892 4632 19944 4684
rect 20352 4632 20404 4684
rect 22008 4632 22060 4684
rect 22284 4632 22336 4684
rect 22744 4675 22796 4684
rect 22744 4641 22753 4675
rect 22753 4641 22787 4675
rect 22787 4641 22796 4675
rect 22744 4632 22796 4641
rect 23020 4632 23072 4684
rect 23480 4675 23532 4684
rect 23480 4641 23489 4675
rect 23489 4641 23523 4675
rect 23523 4641 23532 4675
rect 23480 4632 23532 4641
rect 23940 4632 23992 4684
rect 25964 4709 26016 4718
rect 25964 4675 25973 4709
rect 25973 4675 26007 4709
rect 26007 4675 26016 4709
rect 25964 4666 26016 4675
rect 26792 4675 26844 4684
rect 26792 4641 26801 4675
rect 26801 4641 26835 4675
rect 26835 4641 26844 4675
rect 26792 4632 26844 4641
rect 28540 4709 28592 4718
rect 28540 4675 28549 4709
rect 28549 4675 28583 4709
rect 28583 4675 28592 4709
rect 28540 4666 28592 4675
rect 29184 4632 29236 4684
rect 32036 4632 32088 4684
rect 18144 4564 18196 4616
rect 18052 4496 18104 4548
rect 20352 4496 20404 4548
rect 18512 4471 18564 4480
rect 18512 4437 18521 4471
rect 18521 4437 18555 4471
rect 18555 4437 18564 4471
rect 18512 4428 18564 4437
rect 22192 4428 22244 4480
rect 23756 4428 23808 4480
rect 10950 4326 11002 4378
rect 11014 4326 11066 4378
rect 11078 4326 11130 4378
rect 11142 4326 11194 4378
rect 11206 4326 11258 4378
rect 20950 4326 21002 4378
rect 21014 4326 21066 4378
rect 21078 4326 21130 4378
rect 21142 4326 21194 4378
rect 21206 4326 21258 4378
rect 30950 4326 31002 4378
rect 31014 4326 31066 4378
rect 31078 4326 31130 4378
rect 31142 4326 31194 4378
rect 31206 4326 31258 4378
rect 3792 4224 3844 4276
rect 4712 4224 4764 4276
rect 5448 4224 5500 4276
rect 5540 4156 5592 4208
rect 4804 4088 4856 4140
rect 6736 4224 6788 4276
rect 5816 4156 5868 4208
rect 1952 4029 2004 4038
rect 1952 3995 1961 4029
rect 1961 3995 1995 4029
rect 1995 3995 2004 4029
rect 1952 3986 2004 3995
rect 3884 4020 3936 4072
rect 4252 4020 4304 4072
rect 4528 4063 4580 4072
rect 4528 4029 4537 4063
rect 4537 4029 4571 4063
rect 4571 4029 4580 4063
rect 4528 4020 4580 4029
rect 6828 4088 6880 4140
rect 8944 4088 8996 4140
rect 10416 4088 10468 4140
rect 14648 4088 14700 4140
rect 6736 4063 6788 4072
rect 6736 4029 6745 4063
rect 6745 4029 6779 4063
rect 6779 4029 6788 4063
rect 6736 4020 6788 4029
rect 8484 4029 8536 4038
rect 8484 3995 8493 4029
rect 8493 3995 8527 4029
rect 8527 3995 8536 4029
rect 8484 3986 8536 3995
rect 9312 4020 9364 4072
rect 12072 4020 12124 4072
rect 13360 4029 13412 4038
rect 13360 3995 13369 4029
rect 13369 3995 13403 4029
rect 13403 3995 13412 4029
rect 13360 3986 13412 3995
rect 15016 4063 15068 4072
rect 15016 4029 15025 4063
rect 15025 4029 15059 4063
rect 15059 4029 15068 4063
rect 15016 4020 15068 4029
rect 17868 4029 17920 4038
rect 17868 3995 17877 4029
rect 17877 3995 17911 4029
rect 17911 3995 17920 4029
rect 17868 3986 17920 3995
rect 19156 4020 19208 4072
rect 20444 4029 20496 4038
rect 20444 3995 20453 4029
rect 20453 3995 20487 4029
rect 20487 3995 20496 4029
rect 20444 3986 20496 3995
rect 5632 3884 5684 3936
rect 6184 3884 6236 3936
rect 6644 3884 6696 3936
rect 9496 3884 9548 3936
rect 23940 4020 23992 4072
rect 24308 4029 24360 4038
rect 24308 3995 24317 4029
rect 24317 3995 24351 4029
rect 24351 3995 24360 4029
rect 24308 3986 24360 3995
rect 25964 4063 26016 4072
rect 25964 4029 25973 4063
rect 25973 4029 26007 4063
rect 26007 4029 26016 4063
rect 25964 4020 26016 4029
rect 22008 3884 22060 3936
rect 29184 4020 29236 4072
rect 30012 4029 30064 4038
rect 30012 3995 30021 4029
rect 30021 3995 30055 4029
rect 30055 3995 30064 4029
rect 30012 3986 30064 3995
rect 32036 4020 32088 4072
rect 27620 3884 27672 3936
rect 11610 3782 11662 3834
rect 11674 3782 11726 3834
rect 11738 3782 11790 3834
rect 11802 3782 11854 3834
rect 11866 3782 11918 3834
rect 21610 3782 21662 3834
rect 21674 3782 21726 3834
rect 21738 3782 21790 3834
rect 21802 3782 21854 3834
rect 21866 3782 21918 3834
rect 31610 3782 31662 3834
rect 31674 3782 31726 3834
rect 31738 3782 31790 3834
rect 31802 3782 31854 3834
rect 31866 3782 31918 3834
rect 1952 3680 2004 3732
rect 4160 3680 4212 3732
rect 6828 3680 6880 3732
rect 8944 3680 8996 3732
rect 11336 3680 11388 3732
rect 12900 3680 12952 3732
rect 13360 3680 13412 3732
rect 14648 3680 14700 3732
rect 4252 3612 4304 3664
rect 2872 3544 2924 3596
rect 3792 3544 3844 3596
rect 4436 3544 4488 3596
rect 4804 3621 4856 3630
rect 4804 3587 4813 3621
rect 4813 3587 4847 3621
rect 4847 3587 4856 3621
rect 4804 3578 4856 3587
rect 6644 3612 6696 3664
rect 8668 3612 8720 3664
rect 6184 3544 6236 3596
rect 6460 3544 6512 3596
rect 6920 3544 6972 3596
rect 7288 3587 7340 3596
rect 7288 3553 7297 3587
rect 7297 3553 7331 3587
rect 7331 3553 7340 3587
rect 7288 3544 7340 3553
rect 9036 3544 9088 3596
rect 9128 3587 9180 3596
rect 9128 3553 9137 3587
rect 9137 3553 9171 3587
rect 9171 3553 9180 3587
rect 9128 3544 9180 3553
rect 10784 3568 10836 3620
rect 14832 3612 14884 3664
rect 2780 3519 2832 3528
rect 2780 3485 2789 3519
rect 2789 3485 2823 3519
rect 2823 3485 2832 3519
rect 2780 3476 2832 3485
rect 6092 3476 6144 3528
rect 4252 3408 4304 3460
rect 8300 3519 8352 3528
rect 8300 3485 8309 3519
rect 8309 3485 8343 3519
rect 8343 3485 8352 3519
rect 8300 3476 8352 3485
rect 11980 3544 12032 3596
rect 3332 3340 3384 3392
rect 6460 3340 6512 3392
rect 8484 3408 8536 3460
rect 10810 3451 10862 3460
rect 10810 3417 10819 3451
rect 10819 3417 10853 3451
rect 10853 3417 10862 3451
rect 10810 3408 10862 3417
rect 13452 3519 13504 3528
rect 13452 3485 13461 3519
rect 13461 3485 13495 3519
rect 13495 3485 13504 3519
rect 13452 3476 13504 3485
rect 14740 3544 14792 3596
rect 16672 3621 16724 3630
rect 16672 3587 16681 3621
rect 16681 3587 16715 3621
rect 16715 3587 16724 3621
rect 16672 3578 16724 3587
rect 17500 3544 17552 3596
rect 15108 3476 15160 3528
rect 17960 3519 18012 3528
rect 17960 3485 17969 3519
rect 17969 3485 18003 3519
rect 18003 3485 18012 3519
rect 17960 3476 18012 3485
rect 18512 3587 18564 3596
rect 18512 3553 18521 3587
rect 18521 3553 18555 3587
rect 18555 3553 18564 3587
rect 18512 3544 18564 3553
rect 19248 3680 19300 3732
rect 20812 3680 20864 3732
rect 22100 3680 22152 3732
rect 22652 3680 22704 3732
rect 23204 3680 23256 3732
rect 27620 3680 27672 3732
rect 28540 3680 28592 3732
rect 30012 3680 30064 3732
rect 31484 3680 31536 3732
rect 20628 3544 20680 3596
rect 11980 3408 12032 3460
rect 14924 3408 14976 3460
rect 17132 3408 17184 3460
rect 18604 3408 18656 3460
rect 22100 3587 22152 3596
rect 22100 3553 22109 3587
rect 22109 3553 22143 3587
rect 22143 3553 22152 3587
rect 22100 3544 22152 3553
rect 22192 3544 22244 3596
rect 23020 3587 23072 3596
rect 23020 3553 23029 3587
rect 23029 3553 23063 3587
rect 23063 3553 23072 3587
rect 23020 3544 23072 3553
rect 24308 3544 24360 3596
rect 26792 3612 26844 3664
rect 27160 3655 27212 3664
rect 27160 3621 27169 3655
rect 27169 3621 27203 3655
rect 27203 3621 27212 3655
rect 27160 3612 27212 3621
rect 29368 3612 29420 3664
rect 26884 3544 26936 3596
rect 29000 3544 29052 3596
rect 24860 3476 24912 3528
rect 8300 3340 8352 3392
rect 9128 3340 9180 3392
rect 11336 3340 11388 3392
rect 15016 3340 15068 3392
rect 17224 3340 17276 3392
rect 20720 3340 20772 3392
rect 23756 3340 23808 3392
rect 27620 3383 27672 3392
rect 27620 3349 27629 3383
rect 27629 3349 27663 3383
rect 27663 3349 27672 3383
rect 27620 3340 27672 3349
rect 10950 3238 11002 3290
rect 11014 3238 11066 3290
rect 11078 3238 11130 3290
rect 11142 3238 11194 3290
rect 11206 3238 11258 3290
rect 20950 3238 21002 3290
rect 21014 3238 21066 3290
rect 21078 3238 21130 3290
rect 21142 3238 21194 3290
rect 21206 3238 21258 3290
rect 30950 3238 31002 3290
rect 31014 3238 31066 3290
rect 31078 3238 31130 3290
rect 31142 3238 31194 3290
rect 31206 3238 31258 3290
rect 3792 3136 3844 3188
rect 4344 3136 4396 3188
rect 15200 3136 15252 3188
rect 16304 3136 16356 3188
rect 16396 3179 16448 3188
rect 16396 3145 16405 3179
rect 16405 3145 16439 3179
rect 16439 3145 16448 3179
rect 16396 3136 16448 3145
rect 16534 3136 16586 3188
rect 17132 3136 17184 3188
rect 22100 3136 22152 3188
rect 23756 3136 23808 3188
rect 27620 3136 27672 3188
rect 15936 3068 15988 3120
rect 17500 3068 17552 3120
rect 19616 3068 19668 3120
rect 23020 3068 23072 3120
rect 17776 3000 17828 3052
rect 20168 3000 20220 3052
rect 20720 3000 20772 3052
rect 1676 2975 1728 2984
rect 1676 2941 1685 2975
rect 1685 2941 1719 2975
rect 1719 2941 1728 2975
rect 1676 2932 1728 2941
rect 3700 2932 3752 2984
rect 5080 2941 5132 2950
rect 5080 2907 5089 2941
rect 5089 2907 5123 2941
rect 5123 2907 5132 2941
rect 5080 2898 5132 2907
rect 6644 2932 6696 2984
rect 7012 2932 7064 2984
rect 9036 2941 9088 2950
rect 9036 2907 9045 2941
rect 9045 2907 9079 2941
rect 9079 2907 9088 2941
rect 9036 2898 9088 2907
rect 9404 2932 9456 2984
rect 12440 2975 12492 2984
rect 12440 2941 12449 2975
rect 12449 2941 12483 2975
rect 12483 2941 12492 2975
rect 12440 2932 12492 2941
rect 15936 2975 15988 2984
rect 15936 2941 15945 2975
rect 15945 2941 15979 2975
rect 15979 2941 15988 2975
rect 15936 2932 15988 2941
rect 16534 2932 16586 2984
rect 17224 2932 17276 2984
rect 17868 2932 17920 2984
rect 15108 2864 15160 2916
rect 15292 2864 15344 2916
rect 13728 2796 13780 2848
rect 15200 2796 15252 2848
rect 16764 2864 16816 2916
rect 19156 2941 19208 2950
rect 19156 2907 19165 2941
rect 19165 2907 19199 2941
rect 19199 2907 19208 2941
rect 19156 2898 19208 2907
rect 21364 2975 21416 2984
rect 21364 2941 21373 2975
rect 21373 2941 21407 2975
rect 21407 2941 21416 2975
rect 21364 2932 21416 2941
rect 19800 2864 19852 2916
rect 23204 3000 23256 3052
rect 19984 2839 20036 2848
rect 19984 2805 19993 2839
rect 19993 2805 20027 2839
rect 20027 2805 20036 2839
rect 19984 2796 20036 2805
rect 20444 2796 20496 2848
rect 22376 2864 22428 2916
rect 23296 2975 23348 2984
rect 23296 2941 23305 2975
rect 23305 2941 23339 2975
rect 23339 2941 23348 2975
rect 23296 2932 23348 2941
rect 23848 2975 23900 2984
rect 23848 2941 23857 2975
rect 23857 2941 23891 2975
rect 23891 2941 23900 2975
rect 23848 2932 23900 2941
rect 23940 2975 23992 2984
rect 23940 2941 23949 2975
rect 23949 2941 23983 2975
rect 23983 2941 23992 2975
rect 23940 2932 23992 2941
rect 24584 2975 24636 2984
rect 24584 2941 24593 2975
rect 24593 2941 24627 2975
rect 24627 2941 24636 2975
rect 24584 2932 24636 2941
rect 23020 2796 23072 2848
rect 26056 2796 26108 2848
rect 27620 2839 27672 2848
rect 27620 2805 27629 2839
rect 27629 2805 27663 2839
rect 27663 2805 27672 2839
rect 27620 2796 27672 2805
rect 11610 2694 11662 2746
rect 11674 2694 11726 2746
rect 11738 2694 11790 2746
rect 11802 2694 11854 2746
rect 11866 2694 11918 2746
rect 21610 2694 21662 2746
rect 21674 2694 21726 2746
rect 21738 2694 21790 2746
rect 21802 2694 21854 2746
rect 21866 2694 21918 2746
rect 31610 2694 31662 2746
rect 31674 2694 31726 2746
rect 31738 2694 31790 2746
rect 31802 2694 31854 2746
rect 31866 2694 31918 2746
rect 5816 2592 5868 2644
rect 1676 2456 1728 2508
rect 3792 2499 3844 2508
rect 3792 2465 3801 2499
rect 3801 2465 3835 2499
rect 3835 2465 3844 2499
rect 3792 2456 3844 2465
rect 4804 2533 4856 2542
rect 4804 2499 4813 2533
rect 4813 2499 4847 2533
rect 4847 2499 4856 2533
rect 4804 2490 4856 2499
rect 6920 2456 6972 2508
rect 8300 2592 8352 2644
rect 20720 2592 20772 2644
rect 12440 2524 12492 2576
rect 12808 2499 12860 2508
rect 12808 2465 12817 2499
rect 12817 2465 12851 2499
rect 12851 2465 12860 2499
rect 12808 2456 12860 2465
rect 14556 2533 14608 2542
rect 14556 2499 14565 2533
rect 14565 2499 14599 2533
rect 14599 2499 14608 2533
rect 14556 2490 14608 2499
rect 15108 2456 15160 2508
rect 18512 2524 18564 2576
rect 18880 2533 18932 2542
rect 18880 2499 18889 2533
rect 18889 2499 18923 2533
rect 18923 2499 18932 2533
rect 18880 2490 18932 2499
rect 20628 2499 20680 2508
rect 20628 2465 20637 2499
rect 20637 2465 20671 2499
rect 20671 2465 20680 2499
rect 20628 2456 20680 2465
rect 20168 2388 20220 2440
rect 23940 2592 23992 2644
rect 22376 2499 22428 2508
rect 22376 2465 22385 2499
rect 22385 2465 22419 2499
rect 22419 2465 22428 2499
rect 22376 2456 22428 2465
rect 20812 2388 20864 2440
rect 7656 2320 7708 2372
rect 20536 2320 20588 2372
rect 20720 2252 20772 2304
rect 22008 2320 22060 2372
rect 23296 2456 23348 2508
rect 23204 2320 23256 2372
rect 22376 2252 22428 2304
rect 22836 2252 22888 2304
rect 23020 2252 23072 2304
rect 24216 2295 24268 2304
rect 24216 2261 24225 2295
rect 24225 2261 24259 2295
rect 24259 2261 24268 2295
rect 24216 2252 24268 2261
rect 10950 2150 11002 2202
rect 11014 2150 11066 2202
rect 11078 2150 11130 2202
rect 11142 2150 11194 2202
rect 11206 2150 11258 2202
rect 20950 2150 21002 2202
rect 21014 2150 21066 2202
rect 21078 2150 21130 2202
rect 21142 2150 21194 2202
rect 21206 2150 21258 2202
rect 30950 2150 31002 2202
rect 31014 2150 31066 2202
rect 31078 2150 31130 2202
rect 31142 2150 31194 2202
rect 31206 2150 31258 2202
rect 15660 2091 15712 2100
rect 15660 2057 15669 2091
rect 15669 2057 15703 2091
rect 15703 2057 15712 2091
rect 15660 2048 15712 2057
rect 22192 2048 22244 2100
rect 22560 2048 22612 2100
rect 23664 2048 23716 2100
rect 26056 2091 26108 2100
rect 26056 2057 26065 2091
rect 26065 2057 26099 2091
rect 26099 2057 26108 2091
rect 26056 2048 26108 2057
rect 15016 1980 15068 2032
rect 16212 1980 16264 2032
rect 17868 1980 17920 2032
rect 20812 2023 20864 2032
rect 20812 1989 20821 2023
rect 20821 1989 20855 2023
rect 20855 1989 20864 2023
rect 20812 1980 20864 1989
rect 22284 1980 22336 2032
rect 22468 1980 22520 2032
rect 24216 1980 24268 2032
rect 14648 1912 14700 1964
rect 16304 1912 16356 1964
rect 1676 1887 1728 1896
rect 1676 1853 1685 1887
rect 1685 1853 1719 1887
rect 1719 1853 1728 1887
rect 1676 1844 1728 1853
rect 3332 1853 3384 1862
rect 3332 1819 3341 1853
rect 3341 1819 3375 1853
rect 3375 1819 3384 1853
rect 3332 1810 3384 1819
rect 4528 1776 4580 1828
rect 6736 1887 6788 1896
rect 6736 1853 6745 1887
rect 6745 1853 6779 1887
rect 6779 1853 6788 1887
rect 6736 1844 6788 1853
rect 7656 1853 7708 1862
rect 7656 1819 7665 1853
rect 7665 1819 7699 1853
rect 7699 1819 7708 1853
rect 7656 1810 7708 1819
rect 9404 1887 9456 1896
rect 9404 1853 9413 1887
rect 9413 1853 9447 1887
rect 9447 1853 9456 1887
rect 9404 1844 9456 1853
rect 9680 1844 9732 1896
rect 12808 1844 12860 1896
rect 13360 1853 13412 1862
rect 13360 1819 13369 1853
rect 13369 1819 13403 1853
rect 13403 1819 13412 1853
rect 13360 1810 13412 1819
rect 15108 1887 15160 1896
rect 15108 1853 15117 1887
rect 15117 1853 15151 1887
rect 15151 1853 15160 1887
rect 15108 1844 15160 1853
rect 17960 1887 18012 1896
rect 17960 1853 17969 1887
rect 17969 1853 18003 1887
rect 18003 1853 18012 1887
rect 17960 1844 18012 1853
rect 16028 1776 16080 1828
rect 15752 1708 15804 1760
rect 16672 1708 16724 1760
rect 17408 1708 17460 1760
rect 20536 1912 20588 1964
rect 20168 1844 20220 1896
rect 20444 1887 20496 1896
rect 20444 1853 20453 1887
rect 20453 1853 20487 1887
rect 20487 1853 20496 1887
rect 20444 1844 20496 1853
rect 20720 1776 20772 1828
rect 22008 1887 22060 1896
rect 22008 1853 22017 1887
rect 22017 1853 22051 1887
rect 22051 1853 22060 1887
rect 22008 1844 22060 1853
rect 22744 1844 22796 1896
rect 21456 1776 21508 1828
rect 18604 1708 18656 1760
rect 19984 1708 20036 1760
rect 23204 1776 23256 1828
rect 22376 1708 22428 1760
rect 23940 1751 23992 1760
rect 23940 1717 23949 1751
rect 23949 1717 23983 1751
rect 23983 1717 23992 1751
rect 23940 1708 23992 1717
rect 11610 1606 11662 1658
rect 11674 1606 11726 1658
rect 11738 1606 11790 1658
rect 11802 1606 11854 1658
rect 11866 1606 11918 1658
rect 21610 1606 21662 1658
rect 21674 1606 21726 1658
rect 21738 1606 21790 1658
rect 21802 1606 21854 1658
rect 21866 1606 21918 1658
rect 31610 1606 31662 1658
rect 31674 1606 31726 1658
rect 31738 1606 31790 1658
rect 31802 1606 31854 1658
rect 31866 1606 31918 1658
rect 6552 1504 6604 1556
rect 1952 1411 2004 1420
rect 1952 1377 1961 1411
rect 1961 1377 1995 1411
rect 1995 1377 2004 1411
rect 1952 1368 2004 1377
rect 4436 1368 4488 1420
rect 4528 1411 4580 1420
rect 4528 1377 4537 1411
rect 4537 1377 4571 1411
rect 4571 1377 4580 1411
rect 4528 1368 4580 1377
rect 6828 1368 6880 1420
rect 9680 1436 9732 1488
rect 10508 1445 10560 1454
rect 10508 1411 10517 1445
rect 10517 1411 10551 1445
rect 10551 1411 10560 1445
rect 10508 1402 10560 1411
rect 12256 1411 12308 1420
rect 12256 1377 12265 1411
rect 12265 1377 12299 1411
rect 12299 1377 12308 1411
rect 12256 1368 12308 1377
rect 12348 1368 12400 1420
rect 15108 1436 15160 1488
rect 16580 1504 16632 1556
rect 21456 1504 21508 1556
rect 22836 1547 22888 1556
rect 22836 1513 22845 1547
rect 22845 1513 22879 1547
rect 22879 1513 22888 1547
rect 22836 1504 22888 1513
rect 17960 1436 18012 1488
rect 18972 1368 19024 1420
rect 22192 1436 22244 1488
rect 23664 1436 23716 1488
rect 20720 1368 20772 1420
rect 21364 1368 21416 1420
rect 12164 1300 12216 1352
rect 13084 1300 13136 1352
rect 22008 1300 22060 1352
rect 24860 1343 24912 1352
rect 24860 1309 24869 1343
rect 24869 1309 24903 1343
rect 24903 1309 24912 1343
rect 24860 1300 24912 1309
rect 22652 1232 22704 1284
rect 23388 1275 23440 1284
rect 23388 1241 23397 1275
rect 23397 1241 23431 1275
rect 23431 1241 23440 1275
rect 23388 1232 23440 1241
rect 26148 1232 26200 1284
rect 10950 1062 11002 1114
rect 11014 1062 11066 1114
rect 11078 1062 11130 1114
rect 11142 1062 11194 1114
rect 11206 1062 11258 1114
rect 20950 1062 21002 1114
rect 21014 1062 21066 1114
rect 21078 1062 21130 1114
rect 21142 1062 21194 1114
rect 21206 1062 21258 1114
rect 30950 1062 31002 1114
rect 31014 1062 31066 1114
rect 31078 1062 31130 1114
rect 31142 1062 31194 1114
rect 31206 1062 31258 1114
rect 12348 960 12400 1012
rect 15292 960 15344 1012
rect 14096 935 14148 944
rect 14096 901 14105 935
rect 14105 901 14139 935
rect 14139 901 14148 935
rect 14096 892 14148 901
rect 1952 765 2004 774
rect 1952 731 1961 765
rect 1961 731 1995 765
rect 1995 731 2004 765
rect 1952 722 2004 731
rect 3332 756 3384 808
rect 4436 799 4488 808
rect 4436 765 4445 799
rect 4445 765 4479 799
rect 4479 765 4488 799
rect 4436 756 4488 765
rect 6736 756 6788 808
rect 6828 756 6880 808
rect 12256 756 12308 808
rect 13084 867 13136 876
rect 13084 833 13093 867
rect 13093 833 13127 867
rect 13127 833 13136 867
rect 13084 824 13136 833
rect 13360 824 13412 876
rect 14832 756 14884 808
rect 14924 799 14976 808
rect 14924 765 14933 799
rect 14933 765 14967 799
rect 14967 765 14976 799
rect 14924 756 14976 765
rect 15016 756 15068 808
rect 14464 731 14516 740
rect 14464 697 14473 731
rect 14473 697 14507 731
rect 14507 697 14516 731
rect 17408 765 17460 774
rect 17408 731 17417 765
rect 17417 731 17451 765
rect 17451 731 17460 765
rect 17408 722 17460 731
rect 14464 688 14516 697
rect 13176 663 13228 672
rect 13176 629 13185 663
rect 13185 629 13219 663
rect 13219 629 13228 663
rect 13176 620 13228 629
rect 13544 663 13596 672
rect 13544 629 13553 663
rect 13553 629 13587 663
rect 13587 629 13596 663
rect 13544 620 13596 629
rect 14004 663 14056 672
rect 14004 629 14013 663
rect 14013 629 14047 663
rect 14047 629 14056 663
rect 14004 620 14056 629
rect 15016 663 15068 672
rect 15016 629 15025 663
rect 15025 629 15059 663
rect 15059 629 15068 663
rect 15016 620 15068 629
rect 17960 620 18012 672
rect 19248 892 19300 944
rect 20168 960 20220 1012
rect 20260 1003 20312 1012
rect 20260 969 20269 1003
rect 20269 969 20303 1003
rect 20303 969 20312 1003
rect 20260 960 20312 969
rect 23940 960 23992 1012
rect 23848 892 23900 944
rect 18420 688 18472 740
rect 20260 756 20312 808
rect 22192 824 22244 876
rect 23204 824 23256 876
rect 24860 867 24912 876
rect 24860 833 24869 867
rect 24869 833 24903 867
rect 24903 833 24912 867
rect 24860 824 24912 833
rect 21364 756 21416 808
rect 24216 799 24268 808
rect 24216 765 24225 799
rect 24225 765 24259 799
rect 24259 765 24268 799
rect 24216 756 24268 765
rect 22100 688 22152 740
rect 23388 620 23440 672
rect 11610 518 11662 570
rect 11674 518 11726 570
rect 11738 518 11790 570
rect 11802 518 11854 570
rect 11866 518 11918 570
rect 21610 518 21662 570
rect 21674 518 21726 570
rect 21738 518 21790 570
rect 21802 518 21854 570
rect 21866 518 21918 570
rect 31610 518 31662 570
rect 31674 518 31726 570
rect 31738 518 31790 570
rect 31802 518 31854 570
rect 31866 518 31918 570
rect 9404 416 9456 468
rect 14648 416 14700 468
rect 15016 416 15068 468
rect 23112 416 23164 468
rect 4252 348 4304 400
rect 12256 348 12308 400
rect 8116 280 8168 332
rect 11980 280 12032 332
rect 4160 212 4212 264
rect 12348 212 12400 264
rect 12992 212 13044 264
rect 13176 348 13228 400
rect 18972 348 19024 400
rect 13544 280 13596 332
rect 22008 280 22060 332
rect 21364 212 21416 264
rect 6644 144 6696 196
rect 14004 144 14056 196
rect 14832 144 14884 196
rect 20812 144 20864 196
rect 8668 76 8720 128
rect 14096 76 14148 128
rect 4988 8 5040 60
rect 9956 8 10008 60
rect 10048 8 10100 60
rect 14464 8 14516 60
<< metal2 >>
rect 4160 11960 4212 11966
rect 22376 11960 22428 11966
rect 4160 11902 4212 11908
rect 12438 11928 12494 11937
rect 3700 11892 3752 11898
rect 3700 11834 3752 11840
rect 1032 11756 1084 11762
rect 1032 11698 1084 11704
rect 938 11656 994 11665
rect 938 11591 940 11600
rect 992 11591 994 11600
rect 940 11562 992 11568
rect 1044 11257 1072 11698
rect 2136 11688 2188 11694
rect 2136 11630 2188 11636
rect 1030 11248 1086 11257
rect 1030 11183 1086 11192
rect 1584 11212 1636 11218
rect 1584 11154 1636 11160
rect 1596 10606 1624 11154
rect 1584 10600 1636 10606
rect 1584 10542 1636 10548
rect 938 9752 994 9761
rect 938 9687 994 9696
rect 952 8809 980 9687
rect 1952 9478 2004 9484
rect 1952 9420 2004 9426
rect 1860 9070 1912 9076
rect 1860 9012 1912 9018
rect 938 8800 994 8809
rect 938 8735 994 8744
rect 1768 8390 1820 8396
rect 1768 8332 1820 8338
rect 1780 7478 1808 8332
rect 1768 7472 1820 7478
rect 1768 7414 1820 7420
rect 1872 7342 1900 9012
rect 1964 7546 1992 9420
rect 2044 7982 2096 7988
rect 2044 7924 2096 7930
rect 1952 7540 2004 7546
rect 1952 7482 2004 7488
rect 1860 7336 1912 7342
rect 1860 7278 1912 7284
rect 1584 7200 1636 7206
rect 1584 7142 1636 7148
rect 1596 5166 1624 7142
rect 2056 7002 2084 7924
rect 2044 6996 2096 7002
rect 2044 6938 2096 6944
rect 2148 6254 2176 11630
rect 3056 11620 3108 11626
rect 3056 11562 3108 11568
rect 2780 11552 2832 11558
rect 2780 11494 2832 11500
rect 2226 10160 2282 10169
rect 2226 10095 2282 10104
rect 2226 9888 2282 9897
rect 2226 9823 2282 9832
rect 2136 6248 2188 6254
rect 2136 6190 2188 6196
rect 2240 5710 2268 9823
rect 2792 9761 2820 11494
rect 2778 9752 2834 9761
rect 2778 9687 2834 9696
rect 2870 8256 2926 8265
rect 2870 8191 2926 8200
rect 2594 8120 2650 8129
rect 2594 8055 2650 8064
rect 2608 7274 2636 8055
rect 2686 7440 2742 7449
rect 2686 7375 2688 7384
rect 2740 7375 2742 7384
rect 2688 7346 2740 7352
rect 2596 7268 2648 7274
rect 2596 7210 2648 7216
rect 2688 6112 2740 6118
rect 2688 6054 2740 6060
rect 2412 5772 2464 5778
rect 2412 5714 2464 5720
rect 2228 5704 2280 5710
rect 2424 5681 2452 5714
rect 2228 5646 2280 5652
rect 2410 5672 2466 5681
rect 2410 5607 2466 5616
rect 2700 5166 2728 6054
rect 1584 5160 1636 5166
rect 1584 5102 1636 5108
rect 2688 5160 2740 5166
rect 2688 5102 2740 5108
rect 1400 5092 1452 5098
rect 1400 5034 1452 5040
rect 938 4992 994 5001
rect 938 4927 994 4936
rect 952 4185 980 4927
rect 938 4176 994 4185
rect 938 4111 994 4120
rect 1412 649 1440 5034
rect 2228 5024 2280 5030
rect 2228 4966 2280 4972
rect 2240 4724 2268 4966
rect 2228 4718 2280 4724
rect 2228 4660 2280 4666
rect 1952 4038 2004 4044
rect 1952 3980 2004 3986
rect 1964 3738 1992 3980
rect 1952 3732 2004 3738
rect 1952 3674 2004 3680
rect 2884 3602 2912 8191
rect 3068 7410 3096 11562
rect 3606 11520 3662 11529
rect 3606 11455 3662 11464
rect 3514 10160 3570 10169
rect 3514 10095 3570 10104
rect 3528 10062 3556 10095
rect 3516 10056 3568 10062
rect 3516 9998 3568 10004
rect 3516 9580 3568 9586
rect 3516 9522 3568 9528
rect 3528 8945 3556 9522
rect 3514 8936 3570 8945
rect 3514 8871 3570 8880
rect 3620 7585 3648 11455
rect 3712 11218 3740 11834
rect 3792 11824 3844 11830
rect 3792 11766 3844 11772
rect 3976 11824 4028 11830
rect 3976 11766 4028 11772
rect 3804 11665 3832 11766
rect 3884 11688 3936 11694
rect 3790 11656 3846 11665
rect 3884 11630 3936 11636
rect 3790 11591 3846 11600
rect 3700 11212 3752 11218
rect 3700 11154 3752 11160
rect 3700 9512 3752 9518
rect 3700 9454 3752 9460
rect 3712 8945 3740 9454
rect 3804 9042 3832 11591
rect 3896 10033 3924 11630
rect 3988 10441 4016 11766
rect 4068 11620 4120 11626
rect 4068 11562 4120 11568
rect 4080 10849 4108 11562
rect 4066 10840 4122 10849
rect 4066 10775 4122 10784
rect 3974 10432 4030 10441
rect 3974 10367 4030 10376
rect 4172 10130 4200 11902
rect 20810 11928 20866 11937
rect 12438 11863 12440 11872
rect 12492 11863 12494 11872
rect 12532 11892 12584 11898
rect 12440 11834 12492 11840
rect 12532 11834 12584 11840
rect 20444 11892 20496 11898
rect 22376 11902 22428 11908
rect 30196 11960 30248 11966
rect 30196 11902 30248 11908
rect 20810 11863 20866 11872
rect 20444 11834 20496 11840
rect 12544 11801 12572 11834
rect 9310 11792 9366 11801
rect 9310 11727 9366 11736
rect 12530 11792 12586 11801
rect 14936 11762 15240 11778
rect 12530 11727 12586 11736
rect 12900 11756 12952 11762
rect 4712 11552 4764 11558
rect 4712 11494 4764 11500
rect 4804 11552 4856 11558
rect 4804 11494 4856 11500
rect 7288 11552 7340 11558
rect 7288 11494 7340 11500
rect 4724 11393 4752 11494
rect 4710 11384 4766 11393
rect 4710 11319 4766 11328
rect 4816 11252 4844 11494
rect 4804 11246 4856 11252
rect 7300 11218 7328 11494
rect 4804 11188 4856 11194
rect 6460 11212 6512 11218
rect 6460 11154 6512 11160
rect 7288 11212 7340 11218
rect 7288 11154 7340 11160
rect 4434 10704 4490 10713
rect 4434 10639 4490 10648
rect 4160 10124 4212 10130
rect 4160 10066 4212 10072
rect 3882 10024 3938 10033
rect 3882 9959 3938 9968
rect 4250 9752 4306 9761
rect 4250 9687 4306 9696
rect 4160 9512 4212 9518
rect 4160 9454 4212 9460
rect 3792 9036 3844 9042
rect 3792 8978 3844 8984
rect 3698 8936 3754 8945
rect 3698 8871 3754 8880
rect 3882 7984 3938 7993
rect 3882 7919 3884 7928
rect 3936 7919 3938 7928
rect 3884 7890 3936 7896
rect 4066 7848 4122 7857
rect 4066 7783 4122 7792
rect 3606 7576 3662 7585
rect 3606 7511 3662 7520
rect 3882 7576 3938 7585
rect 3882 7511 3938 7520
rect 3056 7404 3108 7410
rect 3056 7346 3108 7352
rect 3700 7200 3752 7206
rect 3700 7142 3752 7148
rect 3424 6792 3476 6798
rect 3424 6734 3476 6740
rect 3332 6112 3384 6118
rect 3436 6089 3464 6734
rect 3332 6054 3384 6060
rect 3422 6080 3478 6089
rect 2962 5944 3018 5953
rect 2962 5879 3018 5888
rect 2872 3596 2924 3602
rect 2872 3538 2924 3544
rect 2780 3528 2832 3534
rect 2780 3470 2832 3476
rect 1676 2984 1728 2990
rect 1676 2926 1728 2932
rect 1688 2825 1716 2926
rect 1674 2816 1730 2825
rect 1596 2774 1674 2802
rect 1398 640 1454 649
rect 1398 575 1454 584
rect 1596 241 1624 2774
rect 1674 2751 1730 2760
rect 1676 2508 1728 2514
rect 1676 2450 1728 2456
rect 1688 1902 1716 2450
rect 1676 1896 1728 1902
rect 2792 1873 2820 3470
rect 2976 1873 3004 5879
rect 3344 5545 3372 6054
rect 3422 6015 3478 6024
rect 3606 5944 3662 5953
rect 3606 5879 3608 5888
rect 3660 5879 3662 5888
rect 3608 5850 3660 5856
rect 3712 5642 3740 7142
rect 3896 6905 3924 7511
rect 3974 7032 4030 7041
rect 4080 7002 4108 7783
rect 4172 7546 4200 9454
rect 4160 7540 4212 7546
rect 4160 7482 4212 7488
rect 3974 6967 4030 6976
rect 4068 6996 4120 7002
rect 3882 6896 3938 6905
rect 3882 6831 3938 6840
rect 3884 6656 3936 6662
rect 3884 6598 3936 6604
rect 3896 6497 3924 6598
rect 3882 6488 3938 6497
rect 3882 6423 3938 6432
rect 3884 6180 3936 6186
rect 3884 6122 3936 6128
rect 3700 5636 3752 5642
rect 3700 5578 3752 5584
rect 3146 5536 3202 5545
rect 3146 5471 3202 5480
rect 3330 5536 3386 5545
rect 3330 5471 3386 5480
rect 3160 5386 3188 5471
rect 3160 5358 3556 5386
rect 3054 4176 3110 4185
rect 3054 4111 3110 4120
rect 1676 1838 1728 1844
rect 2778 1864 2834 1873
rect 2778 1799 2834 1808
rect 2962 1864 3018 1873
rect 2962 1799 3018 1808
rect 1952 1420 2004 1426
rect 1952 1362 2004 1368
rect 1964 780 1992 1362
rect 1952 774 2004 780
rect 1952 716 2004 722
rect 3068 649 3096 4111
rect 3332 3392 3384 3398
rect 3332 3334 3384 3340
rect 3344 2417 3372 3334
rect 3422 3088 3478 3097
rect 3422 3023 3478 3032
rect 3330 2408 3386 2417
rect 3330 2343 3386 2352
rect 3332 1862 3384 1868
rect 3332 1804 3384 1810
rect 3344 814 3372 1804
rect 3332 808 3384 814
rect 3332 750 3384 756
rect 3054 640 3110 649
rect 3054 575 3110 584
rect 3436 513 3464 3023
rect 3528 2774 3556 5358
rect 3896 5302 3924 6122
rect 3988 6118 4016 6967
rect 4068 6938 4120 6944
rect 4264 6866 4292 9687
rect 4344 7948 4396 7954
rect 4344 7890 4396 7896
rect 4356 7478 4384 7890
rect 4344 7472 4396 7478
rect 4344 7414 4396 7420
rect 4448 7206 4476 10639
rect 6472 10572 6500 11154
rect 6642 11112 6698 11121
rect 6642 11047 6698 11056
rect 6460 10566 6512 10572
rect 6460 10508 6512 10514
rect 5448 9376 5500 9382
rect 5448 9318 5500 9324
rect 5460 9194 5488 9318
rect 5460 9178 5764 9194
rect 6656 9178 6684 11047
rect 7654 10568 7710 10577
rect 7654 10503 7710 10512
rect 6828 10124 6880 10130
rect 6828 10066 6880 10072
rect 7196 10124 7248 10130
rect 7196 10066 7248 10072
rect 6840 9602 6868 10066
rect 6840 9586 6960 9602
rect 6840 9580 6972 9586
rect 6840 9574 6920 9580
rect 6920 9522 6972 9528
rect 7208 9518 7236 10066
rect 8206 10024 8262 10033
rect 8206 9959 8262 9968
rect 7196 9512 7248 9518
rect 7196 9454 7248 9460
rect 5460 9172 5776 9178
rect 5460 9166 5724 9172
rect 5724 9114 5776 9120
rect 6644 9172 6696 9178
rect 6644 9114 6696 9120
rect 4712 9070 4764 9076
rect 4712 9012 4764 9018
rect 4724 8430 4752 9012
rect 5172 8492 5224 8498
rect 5172 8434 5224 8440
rect 4712 8424 4764 8430
rect 4712 8366 4764 8372
rect 5184 8265 5212 8434
rect 5170 8256 5226 8265
rect 5170 8191 5226 8200
rect 6552 7948 6604 7954
rect 6552 7890 6604 7896
rect 6564 7857 6592 7890
rect 6550 7848 6606 7857
rect 6550 7783 6606 7792
rect 6274 7712 6330 7721
rect 6274 7647 6330 7656
rect 6550 7712 6606 7721
rect 6550 7647 6606 7656
rect 5078 7304 5134 7313
rect 5078 7239 5134 7248
rect 4436 7200 4488 7206
rect 4436 7142 4488 7148
rect 4356 6990 4568 7018
rect 4356 6866 4384 6990
rect 4436 6928 4488 6934
rect 4436 6870 4488 6876
rect 4252 6860 4304 6866
rect 4252 6802 4304 6808
rect 4344 6860 4396 6866
rect 4344 6802 4396 6808
rect 4448 6769 4476 6870
rect 4434 6760 4490 6769
rect 4344 6724 4396 6730
rect 4540 6746 4568 6990
rect 6288 6905 6316 7647
rect 6368 7404 6420 7410
rect 6368 7346 6420 7352
rect 6380 7313 6408 7346
rect 6366 7304 6422 7313
rect 6366 7239 6422 7248
rect 4802 6896 4858 6905
rect 4802 6831 4858 6840
rect 6090 6896 6146 6905
rect 6090 6831 6146 6840
rect 6274 6896 6330 6905
rect 6564 6866 6592 7647
rect 6274 6831 6330 6840
rect 6552 6860 6604 6866
rect 6104 6798 6132 6831
rect 6552 6802 6604 6808
rect 6092 6792 6144 6798
rect 4540 6718 5212 6746
rect 6092 6734 6144 6740
rect 4434 6695 4490 6704
rect 4344 6666 4396 6672
rect 4356 6633 4384 6666
rect 4342 6624 4398 6633
rect 4342 6559 4398 6568
rect 4080 6458 4936 6474
rect 4068 6452 4936 6458
rect 4120 6446 4936 6452
rect 4068 6394 4120 6400
rect 4160 6384 4212 6390
rect 4212 6332 4752 6338
rect 4160 6326 4752 6332
rect 4172 6310 4752 6326
rect 4252 6248 4304 6254
rect 4250 6216 4252 6225
rect 4304 6216 4306 6225
rect 4250 6151 4306 6160
rect 4620 6214 4672 6220
rect 4620 6156 4672 6162
rect 3976 6112 4028 6118
rect 3976 6054 4028 6060
rect 3988 5914 4016 6054
rect 3976 5908 4028 5914
rect 3976 5850 4028 5856
rect 4344 5772 4396 5778
rect 4344 5714 4396 5720
rect 4160 5704 4212 5710
rect 4160 5646 4212 5652
rect 4172 5370 4200 5646
rect 4252 5636 4304 5642
rect 4252 5578 4304 5584
rect 4160 5364 4212 5370
rect 4160 5306 4212 5312
rect 3884 5296 3936 5302
rect 3884 5238 3936 5244
rect 3700 5160 3752 5166
rect 3700 5102 3752 5108
rect 3712 2990 3740 5102
rect 3790 4856 3846 4865
rect 3790 4791 3846 4800
rect 3804 4282 3832 4791
rect 3976 4684 4028 4690
rect 3976 4626 4028 4632
rect 3792 4276 3844 4282
rect 3792 4218 3844 4224
rect 3884 4072 3936 4078
rect 3884 4014 3936 4020
rect 3792 3596 3844 3602
rect 3792 3538 3844 3544
rect 3804 3194 3832 3538
rect 3792 3188 3844 3194
rect 3792 3130 3844 3136
rect 3700 2984 3752 2990
rect 3700 2926 3752 2932
rect 3528 2746 3648 2774
rect 3620 785 3648 2746
rect 3792 2508 3844 2514
rect 3792 2450 3844 2456
rect 3606 776 3662 785
rect 3606 711 3662 720
rect 3422 504 3478 513
rect 3422 439 3478 448
rect 3804 377 3832 2450
rect 3896 1329 3924 4014
rect 3882 1320 3938 1329
rect 3882 1255 3938 1264
rect 3988 1193 4016 4626
rect 4264 4078 4292 5578
rect 4356 4570 4384 5714
rect 4632 5234 4660 6156
rect 4528 5228 4580 5234
rect 4528 5170 4580 5176
rect 4620 5228 4672 5234
rect 4620 5170 4672 5176
rect 4436 5024 4488 5030
rect 4436 4966 4488 4972
rect 4448 4690 4476 4966
rect 4540 4865 4568 5170
rect 4526 4856 4582 4865
rect 4724 4826 4752 6310
rect 4802 5808 4858 5817
rect 4802 5743 4858 5752
rect 4526 4791 4582 4800
rect 4712 4820 4764 4826
rect 4712 4762 4764 4768
rect 4436 4684 4488 4690
rect 4436 4626 4488 4632
rect 4356 4542 4660 4570
rect 4252 4072 4304 4078
rect 4252 4014 4304 4020
rect 4528 4072 4580 4078
rect 4528 4014 4580 4020
rect 4160 3732 4212 3738
rect 4160 3674 4212 3680
rect 4172 2774 4200 3674
rect 4252 3664 4304 3670
rect 4250 3632 4252 3641
rect 4304 3632 4306 3641
rect 4250 3567 4306 3576
rect 4436 3596 4488 3602
rect 4436 3538 4488 3544
rect 4250 3496 4306 3505
rect 4250 3431 4252 3440
rect 4304 3431 4306 3440
rect 4252 3402 4304 3408
rect 4344 3188 4396 3194
rect 4344 3130 4396 3136
rect 4172 2746 4292 2774
rect 4066 2680 4122 2689
rect 4122 2638 4200 2666
rect 4066 2615 4122 2624
rect 3974 1184 4030 1193
rect 3974 1119 4030 1128
rect 3790 368 3846 377
rect 3790 303 3846 312
rect 4172 270 4200 2638
rect 4264 406 4292 2746
rect 4356 921 4384 3130
rect 4448 2961 4476 3538
rect 4434 2952 4490 2961
rect 4434 2887 4490 2896
rect 4540 2145 4568 4014
rect 4632 3233 4660 4542
rect 4712 4276 4764 4282
rect 4712 4218 4764 4224
rect 4618 3224 4674 3233
rect 4618 3159 4674 3168
rect 4526 2136 4582 2145
rect 4526 2071 4582 2080
rect 4724 2009 4752 4218
rect 4804 4140 4856 4146
rect 4804 4082 4856 4088
rect 4816 3636 4844 4082
rect 4804 3630 4856 3636
rect 4804 3572 4856 3578
rect 4802 2544 4858 2553
rect 4802 2479 4858 2488
rect 4710 2000 4766 2009
rect 4710 1935 4766 1944
rect 4528 1828 4580 1834
rect 4528 1770 4580 1776
rect 4540 1426 4568 1770
rect 4908 1737 4936 6446
rect 5184 5030 5212 6718
rect 6656 6497 6684 9114
rect 6920 9036 6972 9042
rect 6920 8978 6972 8984
rect 6932 8022 6960 8978
rect 8220 8974 8248 9959
rect 8208 8968 8260 8974
rect 8208 8910 8260 8916
rect 8484 8968 8536 8974
rect 8484 8910 8536 8916
rect 6920 8016 6972 8022
rect 6920 7958 6972 7964
rect 7288 8016 7340 8022
rect 7288 7958 7340 7964
rect 7300 7886 7328 7958
rect 7288 7880 7340 7886
rect 8496 7857 8524 8910
rect 9324 8838 9352 11727
rect 12900 11698 12952 11704
rect 12992 11756 13044 11762
rect 12992 11698 13044 11704
rect 14924 11756 15240 11762
rect 14976 11750 15240 11756
rect 14924 11698 14976 11704
rect 12162 11656 12218 11665
rect 12162 11591 12218 11600
rect 12348 11620 12400 11626
rect 12176 11558 12204 11591
rect 12348 11562 12400 11568
rect 12440 11620 12492 11626
rect 12440 11562 12492 11568
rect 9680 11552 9732 11558
rect 9680 11494 9732 11500
rect 12072 11552 12124 11558
rect 12072 11494 12124 11500
rect 12164 11552 12216 11558
rect 12164 11494 12216 11500
rect 9404 11212 9456 11218
rect 9404 11154 9456 11160
rect 9416 10606 9444 11154
rect 9404 10600 9456 10606
rect 9404 10542 9456 10548
rect 9402 10296 9458 10305
rect 9402 10231 9458 10240
rect 9416 9110 9444 10231
rect 9692 9194 9720 11494
rect 9956 11212 10008 11218
rect 9956 11154 10008 11160
rect 9770 10568 9826 10577
rect 9770 10503 9826 10512
rect 9784 10130 9812 10503
rect 9968 10198 9996 11154
rect 10598 10976 10654 10985
rect 10598 10911 10654 10920
rect 10322 10840 10378 10849
rect 10322 10775 10378 10784
rect 9956 10192 10008 10198
rect 9956 10134 10008 10140
rect 9772 10124 9824 10130
rect 9772 10066 9824 10072
rect 9772 9580 9824 9586
rect 9772 9522 9824 9528
rect 9508 9178 9720 9194
rect 9496 9172 9720 9178
rect 9548 9166 9720 9172
rect 9496 9114 9548 9120
rect 9404 9104 9456 9110
rect 9404 9046 9456 9052
rect 9588 9036 9640 9042
rect 9588 8978 9640 8984
rect 9312 8832 9364 8838
rect 9312 8774 9364 8780
rect 9600 8430 9628 8978
rect 9784 8922 9812 9522
rect 9692 8906 9812 8922
rect 10048 8968 10100 8974
rect 10048 8910 10100 8916
rect 9680 8900 9812 8906
rect 9732 8894 9812 8900
rect 9680 8842 9732 8848
rect 9588 8424 9640 8430
rect 9588 8366 9640 8372
rect 10060 8265 10088 8910
rect 9862 8256 9918 8265
rect 9862 8191 9918 8200
rect 10046 8256 10102 8265
rect 10046 8191 10102 8200
rect 8760 8016 8812 8022
rect 8760 7958 8812 7964
rect 8772 7886 8800 7958
rect 9312 7948 9364 7954
rect 9312 7890 9364 7896
rect 9404 7948 9456 7954
rect 9404 7890 9456 7896
rect 8760 7880 8812 7886
rect 7288 7822 7340 7828
rect 8482 7848 8538 7857
rect 6828 7812 6880 7818
rect 8760 7822 8812 7828
rect 9220 7880 9272 7886
rect 9220 7822 9272 7828
rect 8482 7783 8538 7792
rect 6828 7754 6880 7760
rect 6840 7342 6868 7754
rect 6828 7336 6880 7342
rect 6828 7278 6880 7284
rect 9232 7002 9260 7822
rect 9220 6996 9272 7002
rect 9220 6938 9272 6944
rect 8852 6894 8904 6900
rect 9324 6866 9352 7890
rect 9416 7342 9444 7890
rect 9772 7880 9824 7886
rect 9772 7822 9824 7828
rect 9494 7576 9550 7585
rect 9550 7534 9720 7562
rect 9494 7511 9550 7520
rect 9494 7440 9550 7449
rect 9494 7375 9550 7384
rect 9404 7336 9456 7342
rect 9404 7278 9456 7284
rect 9508 7206 9536 7375
rect 9692 7290 9720 7534
rect 9784 7478 9812 7822
rect 9772 7472 9824 7478
rect 9876 7449 9904 8191
rect 10232 7540 10284 7546
rect 10232 7482 10284 7488
rect 9772 7414 9824 7420
rect 9862 7440 9918 7449
rect 9862 7375 9918 7384
rect 9770 7304 9826 7313
rect 9692 7262 9770 7290
rect 9770 7239 9826 7248
rect 9496 7200 9548 7206
rect 9496 7142 9548 7148
rect 9954 7168 10010 7177
rect 9954 7103 10010 7112
rect 9968 6905 9996 7103
rect 10140 6996 10192 7002
rect 10140 6938 10192 6944
rect 10152 6905 10180 6938
rect 9954 6896 10010 6905
rect 8852 6836 8904 6842
rect 9312 6860 9364 6866
rect 8864 6769 8892 6836
rect 9954 6831 10010 6840
rect 10138 6896 10194 6905
rect 10138 6831 10194 6840
rect 9312 6802 9364 6808
rect 8850 6760 8906 6769
rect 8850 6695 8906 6704
rect 9586 6624 9642 6633
rect 9586 6559 9642 6568
rect 6642 6488 6698 6497
rect 6642 6423 6698 6432
rect 6826 6488 6882 6497
rect 6826 6423 6882 6432
rect 6840 6254 6868 6423
rect 6828 6248 6880 6254
rect 6828 6190 6880 6196
rect 6920 6248 6972 6254
rect 6920 6190 6972 6196
rect 6090 5808 6146 5817
rect 6090 5743 6146 5752
rect 6104 5710 6132 5743
rect 6092 5704 6144 5710
rect 5262 5672 5318 5681
rect 5262 5607 5318 5616
rect 5446 5672 5502 5681
rect 6092 5646 6144 5652
rect 5446 5607 5502 5616
rect 5276 5166 5304 5607
rect 5460 5370 5488 5607
rect 6460 5568 6512 5574
rect 6380 5516 6460 5522
rect 6380 5510 6512 5516
rect 6380 5494 6500 5510
rect 6380 5386 6408 5494
rect 5448 5364 5500 5370
rect 5448 5306 5500 5312
rect 5736 5358 6408 5386
rect 5264 5160 5316 5166
rect 5264 5102 5316 5108
rect 4988 5024 5040 5030
rect 4988 4966 5040 4972
rect 5172 5024 5224 5030
rect 5172 4966 5224 4972
rect 5000 3913 5028 4966
rect 5172 4820 5224 4826
rect 5172 4762 5224 4768
rect 4986 3904 5042 3913
rect 4986 3839 5042 3848
rect 5184 3346 5212 4762
rect 5460 4282 5488 5306
rect 5736 5302 5764 5358
rect 5724 5296 5776 5302
rect 5724 5238 5776 5244
rect 5816 5160 5868 5166
rect 5868 5120 6132 5148
rect 5816 5102 5868 5108
rect 5724 5024 5776 5030
rect 6104 5012 6132 5120
rect 6184 5126 6236 5132
rect 6932 5114 6960 6190
rect 9404 6112 9456 6118
rect 7010 6080 7066 6089
rect 7010 6015 7066 6024
rect 7194 6080 7250 6089
rect 9404 6054 9456 6060
rect 7194 6015 7250 6024
rect 7024 5817 7052 6015
rect 7010 5808 7066 5817
rect 7208 5778 7236 6015
rect 7010 5743 7066 5752
rect 7196 5772 7248 5778
rect 7196 5714 7248 5720
rect 7380 5568 7432 5574
rect 7380 5510 7432 5516
rect 7392 5386 7420 5510
rect 7392 5358 7512 5386
rect 7484 5234 7512 5358
rect 9416 5250 9444 6054
rect 9496 5772 9548 5778
rect 9496 5714 9548 5720
rect 7472 5228 7524 5234
rect 7472 5170 7524 5176
rect 9324 5222 9444 5250
rect 9324 5166 9352 5222
rect 9508 5166 9536 5714
rect 9600 5545 9628 6559
rect 10244 5817 10272 7482
rect 10336 6118 10364 10775
rect 10612 7410 10640 10911
rect 10944 10906 11264 11472
rect 10944 10854 10950 10906
rect 11002 10854 11014 10906
rect 11066 10854 11078 10906
rect 11130 10854 11142 10906
rect 11194 10854 11206 10906
rect 11258 10854 11264 10906
rect 10784 10600 10836 10606
rect 10690 10568 10746 10577
rect 10784 10542 10836 10548
rect 10690 10503 10746 10512
rect 10704 8312 10732 10503
rect 10796 10441 10824 10542
rect 10782 10432 10838 10441
rect 10782 10367 10838 10376
rect 10782 10160 10838 10169
rect 10782 10095 10838 10104
rect 10796 9586 10824 10095
rect 10944 9818 11264 10854
rect 11604 11450 11924 11472
rect 11604 11398 11610 11450
rect 11662 11398 11674 11450
rect 11726 11398 11738 11450
rect 11790 11398 11802 11450
rect 11854 11398 11866 11450
rect 11918 11398 11924 11450
rect 11334 10568 11390 10577
rect 11334 10503 11390 10512
rect 10944 9766 10950 9818
rect 11002 9766 11014 9818
rect 11066 9766 11078 9818
rect 11130 9766 11142 9818
rect 11194 9766 11206 9818
rect 11258 9766 11264 9818
rect 10784 9580 10836 9586
rect 10784 9522 10836 9528
rect 10944 8730 11264 9766
rect 11348 9076 11376 10503
rect 11604 10362 11924 11398
rect 12084 11286 12112 11494
rect 12072 11280 12124 11286
rect 12360 11257 12388 11562
rect 12452 11393 12480 11562
rect 12438 11384 12494 11393
rect 12438 11319 12494 11328
rect 12072 11222 12124 11228
rect 12346 11248 12402 11257
rect 12164 11212 12216 11218
rect 12346 11183 12402 11192
rect 12164 11154 12216 11160
rect 12070 10840 12126 10849
rect 12070 10775 12126 10784
rect 11978 10432 12034 10441
rect 11978 10367 12034 10376
rect 11604 10310 11610 10362
rect 11662 10310 11674 10362
rect 11726 10310 11738 10362
rect 11790 10310 11802 10362
rect 11854 10310 11866 10362
rect 11918 10310 11924 10362
rect 11604 9352 11924 10310
rect 11992 10164 12020 10367
rect 11980 10158 12032 10164
rect 11980 10100 12032 10106
rect 11978 9752 12034 9761
rect 11978 9687 12034 9696
rect 11604 9274 11616 9352
rect 11912 9274 11924 9352
rect 11604 9222 11610 9274
rect 11918 9222 11924 9274
rect 11336 9070 11388 9076
rect 11336 9012 11388 9018
rect 11428 9070 11480 9076
rect 11428 9012 11480 9018
rect 11604 9056 11616 9222
rect 11912 9056 11924 9222
rect 11992 9178 12020 9687
rect 11980 9172 12032 9178
rect 11980 9114 12032 9120
rect 10944 8678 10950 8730
rect 11002 8692 11014 8730
rect 11066 8692 11078 8730
rect 11130 8692 11142 8730
rect 11194 8692 11206 8730
rect 11258 8678 11264 8730
rect 10944 8396 10956 8678
rect 11252 8396 11264 8678
rect 10692 8306 10744 8312
rect 10692 8248 10744 8254
rect 10944 7642 11264 8396
rect 11440 8242 11468 9012
rect 11348 8214 11468 8242
rect 11348 7721 11376 8214
rect 11604 8186 11924 9056
rect 11980 8832 12032 8838
rect 11980 8774 12032 8780
rect 11992 8265 12020 8774
rect 11978 8256 12034 8265
rect 11978 8191 12034 8200
rect 11604 8134 11610 8186
rect 11662 8134 11674 8186
rect 11726 8134 11738 8186
rect 11790 8134 11802 8186
rect 11854 8134 11866 8186
rect 11918 8134 11924 8186
rect 11426 8120 11482 8129
rect 11426 8055 11428 8064
rect 11480 8055 11482 8064
rect 11428 8026 11480 8032
rect 11520 8016 11572 8022
rect 11440 7964 11520 7970
rect 11440 7958 11572 7964
rect 11440 7942 11560 7958
rect 11334 7712 11390 7721
rect 11334 7647 11390 7656
rect 10944 7590 10950 7642
rect 11002 7590 11014 7642
rect 11066 7590 11078 7642
rect 11130 7590 11142 7642
rect 11194 7590 11206 7642
rect 11258 7590 11264 7642
rect 10600 7404 10652 7410
rect 10600 7346 10652 7352
rect 10944 6554 11264 7590
rect 11440 7546 11468 7942
rect 11520 7812 11572 7818
rect 11520 7754 11572 7760
rect 11428 7540 11480 7546
rect 11428 7482 11480 7488
rect 11532 7478 11560 7754
rect 11520 7472 11572 7478
rect 11520 7414 11572 7420
rect 11604 7098 11924 8134
rect 11980 7948 12032 7954
rect 11980 7890 12032 7896
rect 11992 7546 12020 7890
rect 12084 7818 12112 10775
rect 12176 9484 12204 11154
rect 12912 10985 12940 11698
rect 13004 11558 13032 11698
rect 15212 11694 15240 11750
rect 15200 11688 15252 11694
rect 15200 11630 15252 11636
rect 17498 11656 17554 11665
rect 17498 11591 17554 11600
rect 12992 11552 13044 11558
rect 12992 11494 13044 11500
rect 13084 11552 13136 11558
rect 13084 11494 13136 11500
rect 14556 11552 14608 11558
rect 14556 11494 14608 11500
rect 15936 11552 15988 11558
rect 15936 11494 15988 11500
rect 17408 11552 17460 11558
rect 17408 11494 17460 11500
rect 12898 10976 12954 10985
rect 12898 10911 12954 10920
rect 12990 10840 13046 10849
rect 12990 10775 13046 10784
rect 12532 10532 12584 10538
rect 12532 10474 12584 10480
rect 12438 10432 12494 10441
rect 12438 10367 12494 10376
rect 12346 10296 12402 10305
rect 12346 10231 12402 10240
rect 12360 9761 12388 10231
rect 12346 9752 12402 9761
rect 12346 9687 12402 9696
rect 12164 9478 12216 9484
rect 12164 9420 12216 9426
rect 12256 8390 12308 8396
rect 12256 8332 12308 8338
rect 12072 7812 12124 7818
rect 12072 7754 12124 7760
rect 11980 7540 12032 7546
rect 11980 7482 12032 7488
rect 12268 7342 12296 8332
rect 12452 8265 12480 10367
rect 12544 10130 12572 10474
rect 12532 10124 12584 10130
rect 12532 10066 12584 10072
rect 12622 9752 12678 9761
rect 12622 9687 12678 9696
rect 12532 9036 12584 9042
rect 12532 8978 12584 8984
rect 12438 8256 12494 8265
rect 12438 8191 12494 8200
rect 12438 8120 12494 8129
rect 12438 8055 12494 8064
rect 12452 7857 12480 8055
rect 12438 7848 12494 7857
rect 12438 7783 12494 7792
rect 12544 7750 12572 8978
rect 12636 8838 12664 9687
rect 12624 8832 12676 8838
rect 12624 8774 12676 8780
rect 12636 7942 12940 7970
rect 12636 7886 12664 7942
rect 12624 7880 12676 7886
rect 12624 7822 12676 7828
rect 12716 7880 12768 7886
rect 12716 7822 12768 7828
rect 12806 7848 12862 7857
rect 12440 7744 12492 7750
rect 12440 7686 12492 7692
rect 12532 7744 12584 7750
rect 12532 7686 12584 7692
rect 12452 7562 12480 7686
rect 12728 7562 12756 7822
rect 12806 7783 12862 7792
rect 12348 7540 12400 7546
rect 12452 7534 12756 7562
rect 12348 7482 12400 7488
rect 12164 7336 12216 7342
rect 12164 7278 12216 7284
rect 12256 7336 12308 7342
rect 12256 7278 12308 7284
rect 11980 7200 12032 7206
rect 11980 7142 12032 7148
rect 11604 7046 11610 7098
rect 11662 7046 11674 7098
rect 11726 7046 11738 7098
rect 11790 7046 11802 7098
rect 11854 7046 11866 7098
rect 11918 7046 11924 7098
rect 11334 7032 11390 7041
rect 11390 7002 11560 7018
rect 11390 6996 11572 7002
rect 11390 6990 11520 6996
rect 11334 6967 11390 6976
rect 11520 6938 11572 6944
rect 11334 6896 11390 6905
rect 11334 6831 11390 6840
rect 10944 6502 10950 6554
rect 11002 6502 11014 6554
rect 11066 6502 11078 6554
rect 11130 6502 11142 6554
rect 11194 6502 11206 6554
rect 11258 6502 11264 6554
rect 10324 6112 10376 6118
rect 10324 6054 10376 6060
rect 10230 5808 10286 5817
rect 10230 5743 10286 5752
rect 10506 5808 10562 5817
rect 10506 5743 10508 5752
rect 10560 5743 10562 5752
rect 10508 5714 10560 5720
rect 9586 5536 9642 5545
rect 9586 5471 9642 5480
rect 10944 5466 11264 6502
rect 10944 5414 10950 5466
rect 11002 5414 11014 5466
rect 11066 5414 11078 5466
rect 11130 5414 11142 5466
rect 11194 5414 11206 5466
rect 11258 5414 11264 5466
rect 9680 5296 9732 5302
rect 9680 5238 9732 5244
rect 6236 5086 6960 5114
rect 7932 5160 7984 5166
rect 7932 5102 7984 5108
rect 8024 5160 8076 5166
rect 8024 5102 8076 5108
rect 9312 5160 9364 5166
rect 9312 5102 9364 5108
rect 9496 5160 9548 5166
rect 9496 5102 9548 5108
rect 6184 5068 6236 5074
rect 6104 4984 6224 5012
rect 5724 4966 5776 4972
rect 5736 4570 5764 4966
rect 6196 4724 6224 4984
rect 7944 4865 7972 5102
rect 7746 4856 7802 4865
rect 7746 4791 7802 4800
rect 7930 4856 7986 4865
rect 7930 4791 7986 4800
rect 6184 4718 6236 4724
rect 6184 4660 6236 4666
rect 6644 4616 6696 4622
rect 5736 4564 6644 4570
rect 5736 4558 6696 4564
rect 5736 4542 6684 4558
rect 5722 4312 5778 4321
rect 5448 4276 5500 4282
rect 5722 4247 5778 4256
rect 6736 4276 6788 4282
rect 5448 4218 5500 4224
rect 5540 4208 5592 4214
rect 5538 4176 5540 4185
rect 5592 4176 5594 4185
rect 5538 4111 5594 4120
rect 5630 4040 5686 4049
rect 5630 3975 5686 3984
rect 5644 3942 5672 3975
rect 5632 3936 5684 3942
rect 5632 3878 5684 3884
rect 5446 3632 5502 3641
rect 5446 3567 5502 3576
rect 5460 3369 5488 3567
rect 5736 3482 5764 4247
rect 6736 4218 6788 4224
rect 5816 4208 5868 4214
rect 5816 4150 5868 4156
rect 5828 3641 5856 4150
rect 6748 4078 6776 4218
rect 6828 4140 6880 4146
rect 6828 4082 6880 4088
rect 6736 4072 6788 4078
rect 6736 4014 6788 4020
rect 6184 3936 6236 3942
rect 6184 3878 6236 3884
rect 6644 3936 6696 3942
rect 6644 3878 6696 3884
rect 5814 3632 5870 3641
rect 6196 3602 6224 3878
rect 6656 3670 6684 3878
rect 6840 3738 6868 4082
rect 6918 4040 6974 4049
rect 6918 3975 6974 3984
rect 6828 3732 6880 3738
rect 6828 3674 6880 3680
rect 6644 3664 6696 3670
rect 6644 3606 6696 3612
rect 6932 3602 6960 3975
rect 7760 3777 7788 4791
rect 8036 4622 8064 5102
rect 9404 5092 9456 5098
rect 9404 5034 9456 5040
rect 8668 5024 8720 5030
rect 8668 4966 8720 4972
rect 8300 4820 8352 4826
rect 8300 4762 8352 4768
rect 8024 4616 8076 4622
rect 8024 4558 8076 4564
rect 8312 4026 8340 4762
rect 8484 4038 8536 4044
rect 8312 3998 8484 4026
rect 8484 3980 8536 3986
rect 7562 3768 7618 3777
rect 7562 3703 7618 3712
rect 7746 3768 7802 3777
rect 7746 3703 7802 3712
rect 5814 3567 5870 3576
rect 6184 3596 6236 3602
rect 6184 3538 6236 3544
rect 6460 3596 6512 3602
rect 6460 3538 6512 3544
rect 6920 3596 6972 3602
rect 6920 3538 6972 3544
rect 7288 3596 7340 3602
rect 7288 3538 7340 3544
rect 6092 3528 6144 3534
rect 6090 3496 6092 3505
rect 6144 3496 6146 3505
rect 5736 3454 5948 3482
rect 5000 3318 5212 3346
rect 5446 3360 5502 3369
rect 4894 1728 4950 1737
rect 4894 1663 4950 1672
rect 4436 1420 4488 1426
rect 4436 1362 4488 1368
rect 4528 1420 4580 1426
rect 4528 1362 4580 1368
rect 4342 912 4398 921
rect 4342 847 4398 856
rect 4448 814 4476 1362
rect 4436 808 4488 814
rect 4436 750 4488 756
rect 4252 400 4304 406
rect 4252 342 4304 348
rect 4160 264 4212 270
rect 1582 232 1638 241
rect 4160 206 4212 212
rect 1582 167 1638 176
rect 5000 66 5028 3318
rect 5446 3295 5502 3304
rect 5080 2950 5132 2956
rect 5132 2910 5580 2938
rect 5080 2892 5132 2898
rect 5552 2774 5580 2910
rect 5552 2746 5856 2774
rect 5828 2650 5856 2746
rect 5816 2644 5868 2650
rect 5816 2586 5868 2592
rect 5920 2281 5948 3454
rect 6090 3431 6146 3440
rect 6472 3398 6500 3538
rect 7300 3505 7328 3538
rect 7286 3496 7342 3505
rect 7286 3431 7342 3440
rect 6460 3392 6512 3398
rect 6460 3334 6512 3340
rect 6644 2984 6696 2990
rect 6644 2926 6696 2932
rect 7012 2984 7064 2990
rect 7576 2961 7604 3703
rect 8680 3670 8708 4966
rect 9312 4718 9364 4724
rect 9312 4660 9364 4666
rect 8944 4140 8996 4146
rect 8944 4082 8996 4088
rect 8956 3738 8984 4082
rect 9324 4078 9352 4660
rect 9312 4072 9364 4078
rect 9312 4014 9364 4020
rect 8944 3732 8996 3738
rect 8944 3674 8996 3680
rect 8668 3664 8720 3670
rect 8668 3606 8720 3612
rect 8300 3528 8352 3534
rect 8220 3476 8300 3482
rect 8220 3470 8352 3476
rect 8220 3454 8340 3470
rect 8484 3460 8536 3466
rect 8220 3369 8248 3454
rect 8484 3402 8536 3408
rect 8300 3392 8352 3398
rect 8206 3360 8262 3369
rect 8496 3369 8524 3402
rect 8300 3334 8352 3340
rect 8482 3360 8538 3369
rect 8206 3295 8262 3304
rect 7012 2926 7064 2932
rect 7378 2952 7434 2961
rect 6550 2544 6606 2553
rect 6550 2479 6606 2488
rect 5906 2272 5962 2281
rect 5906 2207 5962 2216
rect 6564 1562 6592 2479
rect 6552 1556 6604 1562
rect 6552 1498 6604 1504
rect 6656 202 6684 2926
rect 6918 2544 6974 2553
rect 6918 2479 6920 2488
rect 6972 2479 6974 2488
rect 6920 2450 6972 2456
rect 7024 2417 7052 2926
rect 7378 2887 7434 2896
rect 7562 2952 7618 2961
rect 7562 2887 7618 2896
rect 7392 2417 7420 2887
rect 8220 2774 8248 3295
rect 8128 2746 8248 2774
rect 7010 2408 7066 2417
rect 7010 2343 7066 2352
rect 7378 2408 7434 2417
rect 7378 2343 7434 2352
rect 7656 2372 7708 2378
rect 7656 2314 7708 2320
rect 6736 1896 6788 1902
rect 7668 1868 7696 2314
rect 6736 1838 6788 1844
rect 7656 1862 7708 1868
rect 6748 814 6776 1838
rect 7656 1804 7708 1810
rect 6828 1420 6880 1426
rect 6828 1362 6880 1368
rect 6840 814 6868 1362
rect 6736 808 6788 814
rect 6736 750 6788 756
rect 6828 808 6880 814
rect 6828 750 6880 756
rect 8128 338 8156 2746
rect 8312 2650 8340 3334
rect 8482 3295 8538 3304
rect 8300 2644 8352 2650
rect 8300 2586 8352 2592
rect 8116 332 8168 338
rect 8116 274 8168 280
rect 6644 196 6696 202
rect 6644 138 6696 144
rect 8680 134 8708 3606
rect 9036 3596 9088 3602
rect 9036 3538 9088 3544
rect 9128 3596 9180 3602
rect 9128 3538 9180 3544
rect 9048 2956 9076 3538
rect 9140 3398 9168 3538
rect 9128 3392 9180 3398
rect 9128 3334 9180 3340
rect 9416 2990 9444 5034
rect 9496 3936 9548 3942
rect 9496 3878 9548 3884
rect 9404 2984 9456 2990
rect 9036 2950 9088 2956
rect 9404 2926 9456 2932
rect 9036 2892 9088 2898
rect 9508 2689 9536 3878
rect 9692 2689 9720 5238
rect 10048 5228 10100 5234
rect 10048 5170 10100 5176
rect 9494 2680 9550 2689
rect 9494 2615 9550 2624
rect 9678 2680 9734 2689
rect 9678 2615 9734 2624
rect 9404 1896 9456 1902
rect 9404 1838 9456 1844
rect 9416 474 9444 1838
rect 9404 468 9456 474
rect 9404 410 9456 416
rect 8668 128 8720 134
rect 9508 105 9536 2615
rect 9680 1896 9732 1902
rect 9680 1838 9732 1844
rect 9692 1494 9720 1838
rect 9680 1488 9732 1494
rect 9680 1430 9732 1436
rect 9954 232 10010 241
rect 9954 167 10010 176
rect 8668 70 8720 76
rect 9494 96 9550 105
rect 4988 60 5040 66
rect 9968 66 9996 167
rect 10060 66 10088 5170
rect 10944 4692 11264 5414
rect 10600 4684 10652 4690
rect 10600 4626 10652 4632
rect 10416 4140 10468 4146
rect 10416 4082 10468 4088
rect 10428 3448 10456 4082
rect 10612 3618 10640 4626
rect 10944 4396 10956 4692
rect 11252 4396 11264 4692
rect 10944 4378 11264 4396
rect 10944 4326 10950 4378
rect 11002 4326 11014 4378
rect 11066 4326 11078 4378
rect 11130 4326 11142 4378
rect 11194 4326 11206 4378
rect 11258 4326 11264 4378
rect 10784 3620 10836 3626
rect 10612 3590 10784 3618
rect 10784 3562 10836 3568
rect 10810 3460 10862 3466
rect 10428 3420 10810 3448
rect 10810 3402 10862 3408
rect 10944 3290 11264 4326
rect 11348 3738 11376 6831
rect 11604 6010 11924 7046
rect 11604 5958 11610 6010
rect 11662 5958 11674 6010
rect 11726 5958 11738 6010
rect 11790 5958 11802 6010
rect 11854 5958 11866 6010
rect 11918 5958 11924 6010
rect 11604 5352 11924 5958
rect 11604 5056 11616 5352
rect 11912 5056 11924 5352
rect 11604 4922 11924 5056
rect 11604 4870 11610 4922
rect 11662 4870 11674 4922
rect 11726 4870 11738 4922
rect 11790 4870 11802 4922
rect 11854 4870 11866 4922
rect 11918 4870 11924 4922
rect 11604 3834 11924 4870
rect 11604 3782 11610 3834
rect 11662 3782 11674 3834
rect 11726 3782 11738 3834
rect 11790 3782 11802 3834
rect 11854 3782 11866 3834
rect 11918 3782 11924 3834
rect 11336 3732 11388 3738
rect 11336 3674 11388 3680
rect 11336 3392 11388 3398
rect 11334 3360 11336 3369
rect 11388 3360 11390 3369
rect 11334 3295 11390 3304
rect 10944 3238 10950 3290
rect 11002 3238 11014 3290
rect 11066 3238 11078 3290
rect 11130 3238 11142 3290
rect 11194 3238 11206 3290
rect 11258 3238 11264 3290
rect 10944 2202 11264 3238
rect 10944 2150 10950 2202
rect 11002 2150 11014 2202
rect 11066 2150 11078 2202
rect 11130 2150 11142 2202
rect 11194 2150 11206 2202
rect 11258 2150 11264 2202
rect 10506 1456 10562 1465
rect 10506 1391 10562 1400
rect 10944 1114 11264 2150
rect 10944 1062 10950 1114
rect 11002 1062 11014 1114
rect 11066 1062 11078 1114
rect 11130 1062 11142 1114
rect 11194 1062 11206 1114
rect 11258 1062 11264 1114
rect 10944 496 11264 1062
rect 11604 2746 11924 3782
rect 11992 4706 12020 7142
rect 12176 7041 12204 7278
rect 12162 7032 12218 7041
rect 12162 6967 12218 6976
rect 12360 6866 12388 7482
rect 12716 7404 12768 7410
rect 12716 7346 12768 7352
rect 12728 7313 12756 7346
rect 12714 7304 12770 7313
rect 12714 7239 12770 7248
rect 12820 7177 12848 7783
rect 12806 7168 12862 7177
rect 12806 7103 12862 7112
rect 12348 6860 12400 6866
rect 12348 6802 12400 6808
rect 12530 6760 12586 6769
rect 12912 6746 12940 7942
rect 13004 6866 13032 10775
rect 13096 9518 13124 11494
rect 14568 11252 14596 11494
rect 14556 11246 14608 11252
rect 14556 11188 14608 11194
rect 15660 11212 15712 11218
rect 15660 11154 15712 11160
rect 13174 11112 13230 11121
rect 13174 11047 13230 11056
rect 13358 11112 13414 11121
rect 13358 11047 13414 11056
rect 13084 9512 13136 9518
rect 13084 9454 13136 9460
rect 13188 7177 13216 11047
rect 13372 10572 13400 11047
rect 15016 10600 15068 10606
rect 13360 10566 13412 10572
rect 15016 10542 15068 10548
rect 13360 10508 13412 10514
rect 15028 10164 15056 10542
rect 15016 10158 15068 10164
rect 15016 10100 15068 10106
rect 15198 9752 15254 9761
rect 15198 9687 15200 9696
rect 15252 9687 15254 9696
rect 15200 9658 15252 9664
rect 15672 9518 15700 11154
rect 15842 10432 15898 10441
rect 15842 10367 15898 10376
rect 15856 9586 15884 10367
rect 15948 10130 15976 11494
rect 17420 11252 17448 11494
rect 17408 11246 17460 11252
rect 17408 11188 17460 11194
rect 16486 10704 16542 10713
rect 16486 10639 16542 10648
rect 17222 10704 17278 10713
rect 17222 10639 17278 10648
rect 16302 10568 16358 10577
rect 16302 10503 16358 10512
rect 15936 10124 15988 10130
rect 15936 10066 15988 10072
rect 15844 9580 15896 9586
rect 15844 9522 15896 9528
rect 16212 9580 16264 9586
rect 16212 9522 16264 9528
rect 15660 9512 15712 9518
rect 15660 9454 15712 9460
rect 15936 9376 15988 9382
rect 15936 9318 15988 9324
rect 15016 9070 15068 9076
rect 13268 9036 13320 9042
rect 15016 9012 15068 9018
rect 13268 8978 13320 8984
rect 13280 7750 13308 8978
rect 14648 8492 14700 8498
rect 14648 8434 14700 8440
rect 13360 8390 13412 8396
rect 14660 8378 14688 8434
rect 15028 8430 15056 9012
rect 13412 8350 14688 8378
rect 15016 8424 15068 8430
rect 15016 8366 15068 8372
rect 13360 8332 13412 8338
rect 13636 8084 13688 8090
rect 13636 8026 13688 8032
rect 14464 8084 14516 8090
rect 15844 8084 15896 8090
rect 14516 8044 14596 8072
rect 14464 8026 14516 8032
rect 13268 7744 13320 7750
rect 13648 7721 13676 8026
rect 13728 7948 13780 7954
rect 13780 7908 14136 7936
rect 13728 7890 13780 7896
rect 13728 7744 13780 7750
rect 13268 7686 13320 7692
rect 13634 7712 13690 7721
rect 13728 7686 13780 7692
rect 13634 7647 13690 7656
rect 13740 7290 13768 7686
rect 14108 7460 14136 7908
rect 14188 7880 14240 7886
rect 14188 7822 14240 7828
rect 14200 7528 14228 7822
rect 14464 7540 14516 7546
rect 14200 7500 14464 7528
rect 14464 7482 14516 7488
rect 14108 7432 14412 7460
rect 14004 7302 14056 7308
rect 13740 7262 14004 7290
rect 14384 7274 14412 7432
rect 14004 7244 14056 7250
rect 14372 7268 14424 7274
rect 14372 7210 14424 7216
rect 13174 7168 13230 7177
rect 13174 7103 13230 7112
rect 14568 6900 14596 8044
rect 15844 8026 15896 8032
rect 15856 7993 15884 8026
rect 15476 7982 15528 7988
rect 15476 7924 15528 7930
rect 15842 7984 15898 7993
rect 14830 7848 14886 7857
rect 14830 7783 14886 7792
rect 14844 7585 14872 7783
rect 14646 7576 14702 7585
rect 14646 7511 14702 7520
rect 14830 7576 14886 7585
rect 14830 7511 14886 7520
rect 14660 7478 14688 7511
rect 14648 7472 14700 7478
rect 14648 7414 14700 7420
rect 14844 7342 14872 7511
rect 14832 7336 14884 7342
rect 14832 7278 14884 7284
rect 14556 6894 14608 6900
rect 12992 6860 13044 6866
rect 15488 6866 15516 7924
rect 15842 7919 15898 7928
rect 15566 7848 15622 7857
rect 15566 7783 15622 7792
rect 15580 7274 15608 7783
rect 15948 7750 15976 9318
rect 16224 9076 16252 9522
rect 16212 9070 16264 9076
rect 16212 9012 16264 9018
rect 15936 7744 15988 7750
rect 15936 7686 15988 7692
rect 15568 7268 15620 7274
rect 15568 7210 15620 7216
rect 14556 6836 14608 6842
rect 15476 6860 15528 6866
rect 12992 6802 13044 6808
rect 15476 6802 15528 6808
rect 13084 6792 13136 6798
rect 12912 6718 13032 6746
rect 13084 6734 13136 6740
rect 12530 6695 12586 6704
rect 12254 6624 12310 6633
rect 12310 6582 12388 6610
rect 12254 6559 12310 6568
rect 12254 6488 12310 6497
rect 12360 6474 12388 6582
rect 12544 6474 12572 6695
rect 12714 6624 12770 6633
rect 12714 6559 12770 6568
rect 12360 6446 12572 6474
rect 12254 6423 12310 6432
rect 12268 6100 12296 6423
rect 12624 6316 12676 6322
rect 12624 6258 12676 6264
rect 12530 6216 12586 6225
rect 12636 6202 12664 6258
rect 12728 6225 12756 6559
rect 12898 6488 12954 6497
rect 12898 6423 12954 6432
rect 12586 6174 12664 6202
rect 12714 6216 12770 6225
rect 12530 6151 12586 6160
rect 12714 6151 12770 6160
rect 12808 6180 12860 6186
rect 12808 6122 12860 6128
rect 12268 6089 12572 6100
rect 12268 6080 12586 6089
rect 12268 6072 12530 6080
rect 12530 6015 12586 6024
rect 12070 5808 12126 5817
rect 12820 5778 12848 6122
rect 12070 5743 12126 5752
rect 12256 5772 12308 5778
rect 12084 5166 12112 5743
rect 12256 5714 12308 5720
rect 12808 5772 12860 5778
rect 12808 5714 12860 5720
rect 12268 5166 12296 5714
rect 12072 5160 12124 5166
rect 12072 5102 12124 5108
rect 12256 5160 12308 5166
rect 12256 5102 12308 5108
rect 11992 4678 12388 4706
rect 11992 3602 12020 4678
rect 12360 4622 12388 4678
rect 12348 4616 12400 4622
rect 12348 4558 12400 4564
rect 12070 4176 12126 4185
rect 12254 4176 12310 4185
rect 12070 4111 12126 4120
rect 12176 4134 12254 4162
rect 12084 4078 12112 4111
rect 12072 4072 12124 4078
rect 12072 4014 12124 4020
rect 12070 3904 12126 3913
rect 12176 3890 12204 4134
rect 12254 4111 12310 4120
rect 12126 3862 12204 3890
rect 12070 3839 12126 3848
rect 12912 3738 12940 6423
rect 13004 5681 13032 6718
rect 13096 6633 13124 6734
rect 13082 6624 13138 6633
rect 13082 6559 13138 6568
rect 14568 6446 15332 6474
rect 14568 6338 14596 6446
rect 15200 6384 15252 6390
rect 13464 6322 14596 6338
rect 13452 6316 14596 6322
rect 13504 6310 14596 6316
rect 14660 6332 15200 6338
rect 14660 6326 15252 6332
rect 14660 6310 15240 6326
rect 15304 6322 15332 6446
rect 15292 6316 15344 6322
rect 13452 6258 13504 6264
rect 13728 6112 13780 6118
rect 13780 6060 14596 6066
rect 13728 6054 14596 6060
rect 13740 6038 14596 6054
rect 14568 5812 14596 6038
rect 14556 5806 14608 5812
rect 14556 5748 14608 5754
rect 12990 5672 13046 5681
rect 12990 5607 13046 5616
rect 13818 4856 13874 4865
rect 13818 4791 13874 4800
rect 14002 4856 14058 4865
rect 14002 4791 14004 4800
rect 13832 4185 13860 4791
rect 14056 4791 14058 4800
rect 14004 4762 14056 4768
rect 14660 4298 14688 6310
rect 15292 6258 15344 6264
rect 15384 6248 15436 6254
rect 15384 6190 15436 6196
rect 15290 5944 15346 5953
rect 15290 5879 15346 5888
rect 15198 5536 15254 5545
rect 15198 5471 15254 5480
rect 15212 5302 15240 5471
rect 15304 5370 15332 5879
rect 15396 5545 15424 6190
rect 15844 6180 15896 6186
rect 15844 6122 15896 6128
rect 15660 6112 15712 6118
rect 15658 6080 15660 6089
rect 15712 6080 15714 6089
rect 15658 6015 15714 6024
rect 15856 5778 15884 6122
rect 15844 5772 15896 5778
rect 15844 5714 15896 5720
rect 15382 5536 15438 5545
rect 15382 5471 15438 5480
rect 15292 5364 15344 5370
rect 15292 5306 15344 5312
rect 15200 5296 15252 5302
rect 15200 5238 15252 5244
rect 15108 5160 15160 5166
rect 14740 5126 14792 5132
rect 14740 5068 14792 5074
rect 14936 5120 15108 5148
rect 13924 4270 14688 4298
rect 13634 4176 13690 4185
rect 13634 4111 13690 4120
rect 13818 4176 13874 4185
rect 13818 4111 13874 4120
rect 13360 4038 13412 4044
rect 13648 4026 13676 4111
rect 13924 4026 13952 4270
rect 14648 4140 14700 4146
rect 14648 4082 14700 4088
rect 13648 3998 13952 4026
rect 13360 3980 13412 3986
rect 13372 3738 13400 3980
rect 14554 3768 14610 3777
rect 12900 3732 12952 3738
rect 12900 3674 12952 3680
rect 13360 3732 13412 3738
rect 14660 3738 14688 4082
rect 14554 3703 14610 3712
rect 14648 3732 14700 3738
rect 13360 3674 13412 3680
rect 13450 3632 13506 3641
rect 11980 3596 12032 3602
rect 13450 3567 13506 3576
rect 11980 3538 12032 3544
rect 13464 3534 13492 3567
rect 13452 3528 13504 3534
rect 11978 3496 12034 3505
rect 13452 3470 13504 3476
rect 11978 3431 11980 3440
rect 12032 3431 12034 3440
rect 11980 3402 12032 3408
rect 14568 3369 14596 3703
rect 14648 3674 14700 3680
rect 14752 3602 14780 5068
rect 14832 3664 14884 3670
rect 14936 3652 14964 5120
rect 15108 5102 15160 5108
rect 15200 5092 15252 5098
rect 15200 5034 15252 5040
rect 15108 5024 15160 5030
rect 15108 4966 15160 4972
rect 15016 4718 15068 4724
rect 15016 4660 15068 4666
rect 15028 4078 15056 4660
rect 15016 4072 15068 4078
rect 15016 4014 15068 4020
rect 14884 3624 14964 3652
rect 14832 3606 14884 3612
rect 14740 3596 14792 3602
rect 14740 3538 14792 3544
rect 15120 3534 15148 4966
rect 15212 4865 15240 5034
rect 15198 4856 15254 4865
rect 15198 4791 15254 4800
rect 15396 3913 15424 5471
rect 16500 5098 16528 10639
rect 16854 9752 16910 9761
rect 17236 9722 17264 10639
rect 17406 10296 17462 10305
rect 17406 10231 17462 10240
rect 16854 9687 16910 9696
rect 17224 9716 17276 9722
rect 16868 8945 16896 9687
rect 17224 9658 17276 9664
rect 17040 9444 17092 9450
rect 17040 9386 17092 9392
rect 16948 9376 17000 9382
rect 16948 9318 17000 9324
rect 16854 8936 16910 8945
rect 16854 8871 16910 8880
rect 16578 7984 16634 7993
rect 16578 7919 16634 7928
rect 16592 7342 16620 7919
rect 16580 7336 16632 7342
rect 16580 7278 16632 7284
rect 16764 7268 16816 7274
rect 16764 7210 16816 7216
rect 16578 6624 16634 6633
rect 16578 6559 16634 6568
rect 16592 6390 16620 6559
rect 16776 6390 16804 7210
rect 16960 6458 16988 9318
rect 17052 8945 17080 9386
rect 17038 8936 17094 8945
rect 17038 8871 17094 8880
rect 17132 7948 17184 7954
rect 17132 7890 17184 7896
rect 17144 7546 17172 7890
rect 17420 7698 17448 10231
rect 17512 7818 17540 11591
rect 18052 11552 18104 11558
rect 18052 11494 18104 11500
rect 20260 11552 20312 11558
rect 20260 11494 20312 11500
rect 17776 11212 17828 11218
rect 17776 11154 17828 11160
rect 17788 11121 17816 11154
rect 17774 11112 17830 11121
rect 17774 11047 17830 11056
rect 17958 10976 18014 10985
rect 17958 10911 18014 10920
rect 17592 10668 17644 10674
rect 17592 10610 17644 10616
rect 17604 10577 17632 10610
rect 17590 10568 17646 10577
rect 17590 10503 17646 10512
rect 17866 10432 17922 10441
rect 17866 10367 17922 10376
rect 17880 9738 17908 10367
rect 17972 10266 18000 10911
rect 18064 10606 18092 11494
rect 20272 11252 20300 11494
rect 20260 11246 20312 11252
rect 20260 11188 20312 11194
rect 20456 11121 20484 11834
rect 20628 11824 20680 11830
rect 20628 11766 20680 11772
rect 20442 11112 20498 11121
rect 20442 11047 20498 11056
rect 20640 10985 20668 11766
rect 20718 11520 20774 11529
rect 20718 11455 20774 11464
rect 20626 10976 20682 10985
rect 20626 10911 20682 10920
rect 19890 10704 19946 10713
rect 20732 10674 20760 11455
rect 20824 10713 20852 11863
rect 21916 11756 21968 11762
rect 21968 11716 22048 11744
rect 21916 11698 21968 11704
rect 21638 11656 21694 11665
rect 21456 11620 21508 11626
rect 21694 11626 21864 11642
rect 21694 11620 21876 11626
rect 21694 11614 21824 11620
rect 21638 11591 21694 11600
rect 21456 11562 21508 11568
rect 21824 11562 21876 11568
rect 21364 11552 21416 11558
rect 21364 11494 21416 11500
rect 20944 10906 21264 11472
rect 21376 11286 21404 11494
rect 21468 11393 21496 11562
rect 21604 11450 21924 11472
rect 21604 11398 21610 11450
rect 21662 11398 21674 11450
rect 21726 11398 21738 11450
rect 21790 11398 21802 11450
rect 21854 11398 21866 11450
rect 21918 11398 21924 11450
rect 21454 11384 21510 11393
rect 21454 11319 21510 11328
rect 21364 11280 21416 11286
rect 21364 11222 21416 11228
rect 20944 10854 20950 10906
rect 21002 10854 21014 10906
rect 21066 10854 21078 10906
rect 21130 10854 21142 10906
rect 21194 10854 21206 10906
rect 21258 10854 21264 10906
rect 20810 10704 20866 10713
rect 19890 10639 19946 10648
rect 20720 10668 20772 10674
rect 18052 10600 18104 10606
rect 18052 10542 18104 10548
rect 18970 10296 19026 10305
rect 17960 10260 18012 10266
rect 18970 10231 19026 10240
rect 19064 10260 19116 10266
rect 17960 10202 18012 10208
rect 18052 10192 18104 10198
rect 18050 10160 18052 10169
rect 18104 10160 18106 10169
rect 18050 10095 18106 10104
rect 18050 10024 18106 10033
rect 18050 9959 18106 9968
rect 18064 9926 18092 9959
rect 18984 9926 19012 10231
rect 19064 10202 19116 10208
rect 18052 9920 18104 9926
rect 18052 9862 18104 9868
rect 18972 9920 19024 9926
rect 18972 9862 19024 9868
rect 17880 9710 18000 9738
rect 17592 9580 17644 9586
rect 17592 9522 17644 9528
rect 17604 8974 17632 9522
rect 17684 9376 17736 9382
rect 17684 9318 17736 9324
rect 17592 8968 17644 8974
rect 17592 8910 17644 8916
rect 17696 8396 17724 9318
rect 17868 8900 17920 8906
rect 17868 8842 17920 8848
rect 17684 8390 17736 8396
rect 17684 8332 17736 8338
rect 17880 8129 17908 8842
rect 17866 8120 17922 8129
rect 17972 8090 18000 9710
rect 18880 9478 18932 9484
rect 18880 9420 18932 9426
rect 18696 9036 18748 9042
rect 18696 8978 18748 8984
rect 18708 8265 18736 8978
rect 18892 8430 18920 9420
rect 18880 8424 18932 8430
rect 18880 8366 18932 8372
rect 18694 8256 18750 8265
rect 18694 8191 18750 8200
rect 17866 8055 17922 8064
rect 17960 8084 18012 8090
rect 17960 8026 18012 8032
rect 18984 7886 19012 9862
rect 17960 7880 18012 7886
rect 17960 7822 18012 7828
rect 18972 7880 19024 7886
rect 18972 7822 19024 7828
rect 17500 7812 17552 7818
rect 17500 7754 17552 7760
rect 17592 7812 17644 7818
rect 17592 7754 17644 7760
rect 17604 7698 17632 7754
rect 17420 7670 17632 7698
rect 17132 7540 17184 7546
rect 17132 7482 17184 7488
rect 17040 7472 17092 7478
rect 17092 7420 17448 7426
rect 17040 7414 17448 7420
rect 17052 7398 17448 7414
rect 17132 7336 17184 7342
rect 17132 7278 17184 7284
rect 17144 6900 17172 7278
rect 17420 6905 17448 7398
rect 17604 7002 17632 7670
rect 17776 7200 17828 7206
rect 17776 7142 17828 7148
rect 17592 6996 17644 7002
rect 17592 6938 17644 6944
rect 17132 6894 17184 6900
rect 17132 6836 17184 6842
rect 17222 6896 17278 6905
rect 17222 6831 17278 6840
rect 17406 6896 17462 6905
rect 17406 6831 17462 6840
rect 17038 6624 17094 6633
rect 17038 6559 17094 6568
rect 16948 6452 17000 6458
rect 16948 6394 17000 6400
rect 16580 6384 16632 6390
rect 16580 6326 16632 6332
rect 16764 6384 16816 6390
rect 16764 6326 16816 6332
rect 16580 6112 16632 6118
rect 16580 6054 16632 6060
rect 16488 5092 16540 5098
rect 16488 5034 16540 5040
rect 16304 4684 16356 4690
rect 16356 4644 16528 4672
rect 16304 4626 16356 4632
rect 15382 3904 15438 3913
rect 15382 3839 15438 3848
rect 16210 3768 16266 3777
rect 16210 3703 16266 3712
rect 15108 3528 15160 3534
rect 15108 3470 15160 3476
rect 14924 3460 14976 3466
rect 14924 3402 14976 3408
rect 14936 3369 14964 3402
rect 15016 3392 15068 3398
rect 14554 3360 14610 3369
rect 14554 3295 14610 3304
rect 14922 3360 14978 3369
rect 15068 3352 15240 3380
rect 15016 3334 15068 3340
rect 14922 3295 14978 3304
rect 12254 3224 12310 3233
rect 15212 3194 15240 3352
rect 15934 3224 15990 3233
rect 12254 3159 12310 3168
rect 15200 3188 15252 3194
rect 11604 2694 11610 2746
rect 11662 2694 11674 2746
rect 11726 2694 11738 2746
rect 11790 2694 11802 2746
rect 11854 2694 11866 2746
rect 11918 2694 11924 2746
rect 11604 1658 11924 2694
rect 12268 2417 12296 3159
rect 15934 3159 15990 3168
rect 15200 3130 15252 3136
rect 15948 3126 15976 3159
rect 15936 3120 15988 3126
rect 15936 3062 15988 3068
rect 16224 3074 16252 3703
rect 16500 3618 16528 4644
rect 16592 4185 16620 6054
rect 16578 4176 16634 4185
rect 16578 4111 16634 4120
rect 16776 3777 16804 6326
rect 17052 6225 17080 6559
rect 17038 6216 17094 6225
rect 17038 6151 17094 6160
rect 17236 5953 17264 6831
rect 17222 5944 17278 5953
rect 17222 5879 17278 5888
rect 17788 5250 17816 7142
rect 17972 6633 18000 7822
rect 18512 7812 18564 7818
rect 18512 7754 18564 7760
rect 18604 7812 18656 7818
rect 18604 7754 18656 7760
rect 18524 7449 18552 7754
rect 18510 7440 18566 7449
rect 18510 7375 18566 7384
rect 18616 7177 18644 7754
rect 18788 7302 18840 7308
rect 18788 7244 18840 7250
rect 18602 7168 18658 7177
rect 18602 7103 18658 7112
rect 18800 6866 18828 7244
rect 18788 6860 18840 6866
rect 18788 6802 18840 6808
rect 17958 6624 18014 6633
rect 17958 6559 18014 6568
rect 17866 6488 17922 6497
rect 17866 6423 17868 6432
rect 17920 6423 17922 6432
rect 19076 6474 19104 10202
rect 19800 10124 19852 10130
rect 19800 10066 19852 10072
rect 19812 10033 19840 10066
rect 19798 10024 19854 10033
rect 19798 9959 19854 9968
rect 19156 9920 19208 9926
rect 19156 9862 19208 9868
rect 19168 8022 19196 9862
rect 19338 9752 19394 9761
rect 19338 9687 19394 9696
rect 19352 9654 19380 9687
rect 19904 9654 19932 10639
rect 20810 10639 20866 10648
rect 20720 10610 20772 10616
rect 20732 10418 20760 10610
rect 20640 10390 20760 10418
rect 20536 10260 20588 10266
rect 20536 10202 20588 10208
rect 20258 10160 20314 10169
rect 20258 10095 20314 10104
rect 20272 10062 20300 10095
rect 20260 10056 20312 10062
rect 20260 9998 20312 10004
rect 19340 9648 19392 9654
rect 19340 9590 19392 9596
rect 19892 9648 19944 9654
rect 19892 9590 19944 9596
rect 19248 9444 19300 9450
rect 19248 9386 19300 9392
rect 19260 8974 19288 9386
rect 20548 9076 20576 10202
rect 20640 9518 20668 10390
rect 20628 9512 20680 9518
rect 20628 9454 20680 9460
rect 20536 9070 20588 9076
rect 20536 9012 20588 9018
rect 19248 8968 19300 8974
rect 19248 8910 19300 8916
rect 20260 8390 20312 8396
rect 20260 8332 20312 8338
rect 19614 8120 19670 8129
rect 19614 8055 19670 8064
rect 19890 8120 19946 8129
rect 19890 8055 19946 8064
rect 19156 8016 19208 8022
rect 19156 7958 19208 7964
rect 19168 7342 19196 7958
rect 19248 7948 19300 7954
rect 19248 7890 19300 7896
rect 19260 7546 19288 7890
rect 19248 7540 19300 7546
rect 19248 7482 19300 7488
rect 19628 7478 19656 8055
rect 19904 7818 19932 8055
rect 20272 7954 20300 8332
rect 20260 7948 20312 7954
rect 20260 7890 20312 7896
rect 20076 7880 20128 7886
rect 19982 7848 20038 7857
rect 19892 7812 19944 7818
rect 20076 7822 20128 7828
rect 20258 7848 20314 7857
rect 19982 7783 20038 7792
rect 19892 7754 19944 7760
rect 19708 7744 19760 7750
rect 19708 7686 19760 7692
rect 19720 7478 19748 7686
rect 19616 7472 19668 7478
rect 19616 7414 19668 7420
rect 19708 7472 19760 7478
rect 19708 7414 19760 7420
rect 19156 7336 19208 7342
rect 19156 7278 19208 7284
rect 19248 7268 19300 7274
rect 19248 7210 19300 7216
rect 19156 7200 19208 7206
rect 19260 7177 19288 7210
rect 19156 7142 19208 7148
rect 19246 7168 19302 7177
rect 19168 7002 19196 7142
rect 19246 7103 19302 7112
rect 19430 7168 19486 7177
rect 19430 7103 19486 7112
rect 19444 7018 19472 7103
rect 19156 6996 19208 7002
rect 19156 6938 19208 6944
rect 19260 6990 19472 7018
rect 19260 6633 19288 6990
rect 19246 6624 19302 6633
rect 19246 6559 19302 6568
rect 19430 6624 19486 6633
rect 19430 6559 19486 6568
rect 19444 6474 19472 6559
rect 19076 6446 19472 6474
rect 17868 6394 17920 6400
rect 18052 6384 18104 6390
rect 17866 6352 17922 6361
rect 18052 6326 18104 6332
rect 17866 6287 17922 6296
rect 17880 6254 17908 6287
rect 17868 6248 17920 6254
rect 17868 6190 17920 6196
rect 17960 6248 18012 6254
rect 17960 6190 18012 6196
rect 17972 5846 18000 6190
rect 17960 5840 18012 5846
rect 17960 5782 18012 5788
rect 18064 5778 18092 6326
rect 18052 5772 18104 5778
rect 18052 5714 18104 5720
rect 18696 5704 18748 5710
rect 18694 5672 18696 5681
rect 18748 5672 18750 5681
rect 18694 5607 18750 5616
rect 18052 5568 18104 5574
rect 18052 5510 18104 5516
rect 18064 5386 18092 5510
rect 17972 5370 18092 5386
rect 17960 5364 18092 5370
rect 18012 5358 18092 5364
rect 17960 5306 18012 5312
rect 17788 5222 18092 5250
rect 17316 5092 17368 5098
rect 17316 5034 17368 5040
rect 17328 4185 17356 5034
rect 18064 4690 18092 5222
rect 18328 5228 18380 5234
rect 18328 5170 18380 5176
rect 18144 5160 18196 5166
rect 18144 5102 18196 5108
rect 18156 4758 18184 5102
rect 18340 4865 18368 5170
rect 18326 4856 18382 4865
rect 18326 4791 18382 4800
rect 18144 4752 18196 4758
rect 18144 4694 18196 4700
rect 18052 4684 18104 4690
rect 18052 4626 18104 4632
rect 18144 4616 18196 4622
rect 18144 4558 18196 4564
rect 18052 4548 18104 4554
rect 18052 4490 18104 4496
rect 17314 4176 17370 4185
rect 17314 4111 17370 4120
rect 17868 4038 17920 4044
rect 17868 3980 17920 3986
rect 16762 3768 16818 3777
rect 16762 3703 16818 3712
rect 16672 3630 16724 3636
rect 16500 3590 16672 3618
rect 16672 3572 16724 3578
rect 16316 3318 16574 3346
rect 16316 3194 16344 3318
rect 16546 3194 16574 3318
rect 16304 3188 16356 3194
rect 16304 3130 16356 3136
rect 16396 3188 16448 3194
rect 16396 3130 16448 3136
rect 16534 3188 16586 3194
rect 16534 3130 16586 3136
rect 16408 3074 16436 3130
rect 15948 2990 15976 3062
rect 16224 3046 16436 3074
rect 12440 2984 12492 2990
rect 12440 2926 12492 2932
rect 15936 2984 15988 2990
rect 15936 2926 15988 2932
rect 12452 2582 12480 2926
rect 15108 2916 15160 2922
rect 15108 2858 15160 2864
rect 15292 2916 15344 2922
rect 15292 2858 15344 2864
rect 13728 2848 13780 2854
rect 13728 2790 13780 2796
rect 12440 2576 12492 2582
rect 12440 2518 12492 2524
rect 13740 2530 13768 2790
rect 15014 2680 15070 2689
rect 15014 2615 15070 2624
rect 14556 2542 14608 2548
rect 12808 2508 12860 2514
rect 13740 2502 14556 2530
rect 14556 2484 14608 2490
rect 12808 2450 12860 2456
rect 12254 2408 12310 2417
rect 12254 2343 12310 2352
rect 12392 2408 12448 2417
rect 12392 2343 12448 2352
rect 12406 2258 12434 2343
rect 12268 2230 12434 2258
rect 12268 1873 12296 2230
rect 12820 1902 12848 2450
rect 15028 2038 15056 2615
rect 15120 2514 15148 2858
rect 15200 2848 15252 2854
rect 15200 2790 15252 2796
rect 15108 2508 15160 2514
rect 15108 2450 15160 2456
rect 15016 2032 15068 2038
rect 15016 1974 15068 1980
rect 14648 1964 14700 1970
rect 14648 1906 14700 1912
rect 12808 1896 12860 1902
rect 12254 1864 12310 1873
rect 12808 1838 12860 1844
rect 13082 1864 13138 1873
rect 12254 1799 12310 1808
rect 13082 1799 13138 1808
rect 13360 1862 13412 1868
rect 13360 1804 13412 1810
rect 12162 1728 12218 1737
rect 12162 1663 12218 1672
rect 12990 1728 13046 1737
rect 12990 1663 13046 1672
rect 11604 1606 11610 1658
rect 11662 1606 11674 1658
rect 11726 1606 11738 1658
rect 11790 1606 11802 1658
rect 11854 1606 11866 1658
rect 11918 1606 11924 1658
rect 11604 570 11924 1606
rect 12176 1358 12204 1663
rect 12346 1456 12402 1465
rect 12256 1420 12308 1426
rect 12346 1391 12348 1400
rect 12256 1362 12308 1368
rect 12400 1391 12402 1400
rect 12348 1362 12400 1368
rect 12164 1352 12216 1358
rect 12164 1294 12216 1300
rect 12268 814 12296 1362
rect 12348 1012 12400 1018
rect 12348 954 12400 960
rect 12256 808 12308 814
rect 12256 750 12308 756
rect 12360 626 12388 954
rect 11604 518 11610 570
rect 11662 518 11674 570
rect 11726 518 11738 570
rect 11790 518 11802 570
rect 11854 518 11866 570
rect 11918 518 11924 570
rect 11604 496 11924 518
rect 12268 598 12388 626
rect 12268 406 12296 598
rect 12256 400 12308 406
rect 12256 342 12308 348
rect 11980 332 12032 338
rect 11980 274 12032 280
rect 11992 82 12020 274
rect 13004 270 13032 1663
rect 13096 1358 13124 1799
rect 13084 1352 13136 1358
rect 13084 1294 13136 1300
rect 13096 882 13124 1294
rect 13372 882 13400 1804
rect 14096 944 14148 950
rect 14096 886 14148 892
rect 13084 876 13136 882
rect 13084 818 13136 824
rect 13360 876 13412 882
rect 13360 818 13412 824
rect 13176 672 13228 678
rect 13176 614 13228 620
rect 13544 672 13596 678
rect 13544 614 13596 620
rect 14004 672 14056 678
rect 14004 614 14056 620
rect 13188 406 13216 614
rect 13176 400 13228 406
rect 13176 342 13228 348
rect 13556 338 13584 614
rect 13544 332 13596 338
rect 13544 274 13596 280
rect 12348 264 12400 270
rect 12070 232 12126 241
rect 12126 212 12348 218
rect 12126 206 12400 212
rect 12992 264 13044 270
rect 12992 206 13044 212
rect 12126 190 12388 206
rect 14016 202 14044 614
rect 14004 196 14056 202
rect 12070 167 12126 176
rect 14004 138 14056 144
rect 14108 134 14136 886
rect 14464 740 14516 746
rect 14464 682 14516 688
rect 14096 128 14148 134
rect 12346 96 12402 105
rect 9494 31 9550 40
rect 9956 60 10008 66
rect 4988 2 5040 8
rect 9956 2 10008 8
rect 10048 60 10100 66
rect 11992 54 12346 82
rect 14096 70 14148 76
rect 14476 66 14504 682
rect 14660 474 14688 1906
rect 15108 1896 15160 1902
rect 15108 1838 15160 1844
rect 15120 1494 15148 1838
rect 15108 1488 15160 1494
rect 15014 1456 15070 1465
rect 15108 1430 15160 1436
rect 15014 1391 15070 1400
rect 14922 912 14978 921
rect 14922 847 14978 856
rect 14936 814 14964 847
rect 15028 814 15056 1391
rect 14832 808 14884 814
rect 14832 750 14884 756
rect 14924 808 14976 814
rect 14924 750 14976 756
rect 15016 808 15068 814
rect 15016 750 15068 756
rect 14648 468 14700 474
rect 14648 410 14700 416
rect 14844 202 14872 750
rect 15016 672 15068 678
rect 15016 614 15068 620
rect 15028 474 15056 614
rect 15016 468 15068 474
rect 15016 410 15068 416
rect 15212 241 15240 2790
rect 15304 1018 15332 2858
rect 15658 2544 15714 2553
rect 15658 2479 15714 2488
rect 15842 2544 15898 2553
rect 15842 2479 15898 2488
rect 15672 2106 15700 2479
rect 15660 2100 15712 2106
rect 15660 2042 15712 2048
rect 15856 1873 15884 2479
rect 16224 2038 16252 3046
rect 16534 2984 16586 2990
rect 16316 2944 16534 2972
rect 16212 2032 16264 2038
rect 16212 1974 16264 1980
rect 16316 1970 16344 2944
rect 16534 2926 16586 2932
rect 16776 2922 16804 3703
rect 17500 3596 17552 3602
rect 17500 3538 17552 3544
rect 17132 3460 17184 3466
rect 17132 3402 17184 3408
rect 17144 3194 17172 3402
rect 17224 3392 17276 3398
rect 17224 3334 17276 3340
rect 17132 3188 17184 3194
rect 17132 3130 17184 3136
rect 17236 2990 17264 3334
rect 17314 3224 17370 3233
rect 17314 3159 17370 3168
rect 17224 2984 17276 2990
rect 17328 2961 17356 3159
rect 17512 3126 17540 3538
rect 17500 3120 17552 3126
rect 17500 3062 17552 3068
rect 17776 3052 17828 3058
rect 17776 2994 17828 3000
rect 17788 2961 17816 2994
rect 17880 2990 17908 3980
rect 17960 3528 18012 3534
rect 17958 3496 17960 3505
rect 18012 3496 18014 3505
rect 17958 3431 18014 3440
rect 17868 2984 17920 2990
rect 17224 2926 17276 2932
rect 17314 2952 17370 2961
rect 16764 2916 16816 2922
rect 17314 2887 17370 2896
rect 17774 2952 17830 2961
rect 17868 2926 17920 2932
rect 17774 2887 17830 2896
rect 16764 2858 16816 2864
rect 18064 2145 18092 4490
rect 18156 4321 18184 4558
rect 18512 4480 18564 4486
rect 18512 4422 18564 4428
rect 18142 4312 18198 4321
rect 18142 4247 18198 4256
rect 18524 4049 18552 4422
rect 18510 4040 18566 4049
rect 18510 3975 18566 3984
rect 18512 3596 18564 3602
rect 18512 3538 18564 3544
rect 18524 2582 18552 3538
rect 18604 3460 18656 3466
rect 18604 3402 18656 3408
rect 18512 2576 18564 2582
rect 18512 2518 18564 2524
rect 18616 2417 18644 3402
rect 19076 2774 19104 6446
rect 19996 6440 20024 7783
rect 20088 7721 20116 7822
rect 20258 7783 20314 7792
rect 20074 7712 20130 7721
rect 20074 7647 20130 7656
rect 20088 7410 20116 7647
rect 20076 7404 20128 7410
rect 20076 7346 20128 7352
rect 20272 7342 20300 7783
rect 20824 7410 20852 10639
rect 20944 9818 21264 10854
rect 20944 9766 20950 9818
rect 21002 9766 21014 9818
rect 21066 9766 21078 9818
rect 21130 9766 21142 9818
rect 21194 9766 21206 9818
rect 21258 9766 21264 9818
rect 20944 8730 21264 9766
rect 21604 10362 21924 11398
rect 22020 11257 22048 11716
rect 22006 11248 22062 11257
rect 22006 11183 22062 11192
rect 22008 10464 22060 10470
rect 22006 10432 22008 10441
rect 22060 10432 22062 10441
rect 22006 10367 22062 10376
rect 21604 10310 21610 10362
rect 21662 10310 21674 10362
rect 21726 10310 21738 10362
rect 21790 10310 21802 10362
rect 21854 10310 21866 10362
rect 21918 10310 21924 10362
rect 21454 9752 21510 9761
rect 21454 9687 21456 9696
rect 21508 9687 21510 9696
rect 21456 9658 21508 9664
rect 21364 9512 21416 9518
rect 21364 9454 21416 9460
rect 21376 8974 21404 9454
rect 21604 9352 21924 10310
rect 22006 10296 22062 10305
rect 22006 10231 22008 10240
rect 22060 10231 22062 10240
rect 22008 10202 22060 10208
rect 22100 10192 22152 10198
rect 22098 10160 22100 10169
rect 22152 10160 22154 10169
rect 22008 10124 22060 10130
rect 22098 10095 22154 10104
rect 22008 10066 22060 10072
rect 22020 9382 22048 10066
rect 22388 10062 22416 11902
rect 22928 11688 22980 11694
rect 22928 11630 22980 11636
rect 29920 11688 29972 11694
rect 29920 11630 29972 11636
rect 22940 10713 22968 11630
rect 25688 11620 25740 11626
rect 25688 11562 25740 11568
rect 23940 11552 23992 11558
rect 23940 11494 23992 11500
rect 23112 11212 23164 11218
rect 23112 11154 23164 11160
rect 22926 10704 22982 10713
rect 22926 10639 22982 10648
rect 23124 10572 23152 11154
rect 23388 11076 23440 11082
rect 23388 11018 23440 11024
rect 23112 10566 23164 10572
rect 23112 10508 23164 10514
rect 23400 10198 23428 11018
rect 23480 11008 23532 11014
rect 23480 10950 23532 10956
rect 23388 10192 23440 10198
rect 23388 10134 23440 10140
rect 22376 10056 22428 10062
rect 22098 10024 22154 10033
rect 22376 9998 22428 10004
rect 22098 9959 22100 9968
rect 22152 9959 22154 9968
rect 22100 9930 22152 9936
rect 23492 9761 23520 10950
rect 23952 10606 23980 11494
rect 25042 11384 25098 11393
rect 24124 11348 24176 11354
rect 25042 11319 25098 11328
rect 24124 11290 24176 11296
rect 24032 11144 24084 11150
rect 24032 11086 24084 11092
rect 23940 10600 23992 10606
rect 23940 10542 23992 10548
rect 23662 10160 23718 10169
rect 23662 10095 23718 10104
rect 23478 9752 23534 9761
rect 23478 9687 23534 9696
rect 23112 9478 23164 9484
rect 23032 9438 23112 9466
rect 21604 9274 21616 9352
rect 21912 9274 21924 9352
rect 22008 9376 22060 9382
rect 22008 9318 22060 9324
rect 21604 9222 21610 9274
rect 21918 9222 21924 9274
rect 21604 9056 21616 9222
rect 21912 9056 21924 9222
rect 23032 9194 23060 9438
rect 23112 9420 23164 9426
rect 22296 9178 23060 9194
rect 22284 9172 23060 9178
rect 22336 9166 23060 9172
rect 22284 9114 22336 9120
rect 21364 8968 21416 8974
rect 21364 8910 21416 8916
rect 20944 8678 20950 8730
rect 21002 8692 21014 8730
rect 21066 8692 21078 8730
rect 21130 8692 21142 8730
rect 21194 8692 21206 8730
rect 21258 8678 21264 8730
rect 20944 8396 20956 8678
rect 21252 8396 21264 8678
rect 20944 7642 21264 8396
rect 20944 7590 20950 7642
rect 21002 7590 21014 7642
rect 21066 7590 21078 7642
rect 21130 7590 21142 7642
rect 21194 7590 21206 7642
rect 21258 7590 21264 7642
rect 20812 7404 20864 7410
rect 20812 7346 20864 7352
rect 20260 7336 20312 7342
rect 20260 7278 20312 7284
rect 20810 7304 20866 7313
rect 20168 6452 20220 6458
rect 19996 6412 20168 6440
rect 20168 6394 20220 6400
rect 19708 6214 19760 6220
rect 19708 6156 19760 6162
rect 19614 5808 19670 5817
rect 19720 5778 19748 6156
rect 19890 5808 19946 5817
rect 19614 5743 19670 5752
rect 19708 5772 19760 5778
rect 19522 5672 19578 5681
rect 19522 5607 19578 5616
rect 19536 5574 19564 5607
rect 19524 5568 19576 5574
rect 19524 5510 19576 5516
rect 19628 5132 19656 5743
rect 19890 5743 19946 5752
rect 19708 5714 19760 5720
rect 19904 5710 19932 5743
rect 19892 5704 19944 5710
rect 19892 5646 19944 5652
rect 19904 5250 19932 5646
rect 20074 5536 20130 5545
rect 20074 5471 20130 5480
rect 20088 5370 20116 5471
rect 20076 5364 20128 5370
rect 20076 5306 20128 5312
rect 19904 5234 20116 5250
rect 19904 5228 20128 5234
rect 19904 5222 20076 5228
rect 20076 5170 20128 5176
rect 19984 5160 20036 5166
rect 19616 5126 19668 5132
rect 19616 5068 19668 5074
rect 19904 5120 19984 5148
rect 19904 4690 19932 5120
rect 19984 5102 20036 5108
rect 19892 4684 19944 4690
rect 19892 4626 19944 4632
rect 19156 4072 19208 4078
rect 19156 4014 19208 4020
rect 19168 2956 19196 4014
rect 19248 3732 19300 3738
rect 19300 3692 19656 3720
rect 19248 3674 19300 3680
rect 19628 3126 19656 3692
rect 19616 3120 19668 3126
rect 19616 3062 19668 3068
rect 20168 3052 20220 3058
rect 20168 2994 20220 3000
rect 20180 2961 20208 2994
rect 19156 2950 19208 2956
rect 20166 2952 20222 2961
rect 19156 2892 19208 2898
rect 19800 2916 19852 2922
rect 20166 2887 20222 2896
rect 19800 2858 19852 2864
rect 18892 2746 19104 2774
rect 18892 2548 18920 2746
rect 19246 2680 19302 2689
rect 19246 2615 19302 2624
rect 18880 2542 18932 2548
rect 18880 2484 18932 2490
rect 18602 2408 18658 2417
rect 18602 2343 18658 2352
rect 18050 2136 18106 2145
rect 18050 2071 18106 2080
rect 17868 2032 17920 2038
rect 17868 1974 17920 1980
rect 16304 1964 16356 1970
rect 16304 1906 16356 1912
rect 17880 1873 17908 1974
rect 17960 1896 18012 1902
rect 15842 1864 15898 1873
rect 17866 1864 17922 1873
rect 15842 1799 15898 1808
rect 16028 1828 16080 1834
rect 17960 1838 18012 1844
rect 17866 1799 17922 1808
rect 16028 1770 16080 1776
rect 15752 1760 15804 1766
rect 16040 1737 16068 1770
rect 16672 1760 16724 1766
rect 15752 1702 15804 1708
rect 16026 1728 16082 1737
rect 15764 1193 15792 1702
rect 16026 1663 16082 1672
rect 16592 1720 16672 1748
rect 16592 1562 16620 1720
rect 16672 1702 16724 1708
rect 17408 1760 17460 1766
rect 17408 1702 17460 1708
rect 16580 1556 16632 1562
rect 16580 1498 16632 1504
rect 15750 1184 15806 1193
rect 15750 1119 15806 1128
rect 15292 1012 15344 1018
rect 15292 954 15344 960
rect 17420 780 17448 1702
rect 17972 1494 18000 1838
rect 18604 1760 18656 1766
rect 18418 1728 18474 1737
rect 18418 1663 18474 1672
rect 18602 1728 18604 1737
rect 18656 1728 18658 1737
rect 18602 1663 18658 1672
rect 17960 1488 18012 1494
rect 17960 1430 18012 1436
rect 17408 774 17460 780
rect 18432 746 18460 1663
rect 18972 1420 19024 1426
rect 18972 1362 19024 1368
rect 17408 716 17460 722
rect 18420 740 18472 746
rect 18420 682 18472 688
rect 17960 672 18012 678
rect 17960 614 18012 620
rect 15198 232 15254 241
rect 14832 196 14884 202
rect 15198 167 15254 176
rect 14832 138 14884 144
rect 17972 105 18000 614
rect 18984 406 19012 1362
rect 19260 950 19288 2615
rect 19812 1465 19840 2858
rect 19984 2848 20036 2854
rect 19984 2790 20036 2796
rect 19996 1986 20024 2790
rect 20168 2440 20220 2446
rect 20166 2408 20168 2417
rect 20220 2408 20222 2417
rect 20166 2343 20222 2352
rect 19904 1958 20024 1986
rect 19798 1456 19854 1465
rect 19798 1391 19854 1400
rect 19904 1329 19932 1958
rect 20168 1896 20220 1902
rect 19982 1864 20038 1873
rect 20168 1838 20220 1844
rect 19982 1799 20038 1808
rect 19996 1766 20024 1799
rect 19984 1760 20036 1766
rect 19984 1702 20036 1708
rect 19890 1320 19946 1329
rect 19890 1255 19946 1264
rect 20180 1018 20208 1838
rect 20272 1601 20300 7278
rect 20628 7268 20680 7274
rect 20810 7239 20866 7248
rect 20628 7210 20680 7216
rect 20534 6352 20590 6361
rect 20534 6287 20590 6296
rect 20548 5545 20576 6287
rect 20534 5536 20590 5545
rect 20534 5471 20590 5480
rect 20352 4684 20404 4690
rect 20404 4644 20484 4672
rect 20352 4626 20404 4632
rect 20352 4548 20404 4554
rect 20352 4490 20404 4496
rect 20364 4321 20392 4490
rect 20350 4312 20406 4321
rect 20350 4247 20406 4256
rect 20456 4044 20484 4644
rect 20640 4049 20668 7210
rect 20824 7206 20852 7239
rect 20812 7200 20864 7206
rect 20812 7142 20864 7148
rect 20718 6896 20774 6905
rect 20718 6831 20774 6840
rect 20732 6361 20760 6831
rect 20944 6554 21264 7590
rect 21604 8186 21924 9056
rect 22008 8968 22060 8974
rect 22008 8910 22060 8916
rect 22020 8378 22048 8910
rect 22020 8350 22140 8378
rect 22008 8288 22060 8294
rect 22008 8230 22060 8236
rect 21604 8134 21610 8186
rect 21662 8134 21674 8186
rect 21726 8134 21738 8186
rect 21790 8134 21802 8186
rect 21854 8134 21866 8186
rect 21918 8134 21924 8186
rect 21362 7576 21418 7585
rect 21362 7511 21418 7520
rect 21376 7177 21404 7511
rect 21362 7168 21418 7177
rect 21362 7103 21418 7112
rect 21604 7098 21924 8134
rect 22020 8022 22048 8230
rect 22112 8022 22140 8350
rect 22190 8120 22246 8129
rect 22190 8055 22192 8064
rect 22244 8055 22246 8064
rect 22192 8026 22244 8032
rect 22008 8016 22060 8022
rect 22008 7958 22060 7964
rect 22100 8016 22152 8022
rect 22100 7958 22152 7964
rect 22204 7410 22232 8026
rect 23296 7948 23348 7954
rect 23296 7890 23348 7896
rect 22744 7880 22796 7886
rect 22744 7822 22796 7828
rect 22468 7812 22520 7818
rect 22468 7754 22520 7760
rect 22376 7744 22428 7750
rect 22376 7686 22428 7692
rect 22388 7546 22416 7686
rect 22376 7540 22428 7546
rect 22376 7482 22428 7488
rect 22480 7478 22508 7754
rect 22650 7576 22706 7585
rect 22650 7511 22706 7520
rect 22468 7472 22520 7478
rect 22468 7414 22520 7420
rect 22192 7404 22244 7410
rect 22192 7346 22244 7352
rect 22664 7290 22692 7511
rect 22388 7262 22692 7290
rect 22388 7177 22416 7262
rect 22374 7168 22430 7177
rect 22374 7103 22430 7112
rect 21604 7046 21610 7098
rect 21662 7046 21674 7098
rect 21726 7046 21738 7098
rect 21790 7046 21802 7098
rect 21854 7046 21866 7098
rect 21918 7046 21924 7098
rect 21362 6896 21418 6905
rect 21362 6831 21418 6840
rect 21376 6633 21404 6831
rect 21362 6624 21418 6633
rect 21362 6559 21418 6568
rect 20944 6502 20950 6554
rect 21002 6502 21014 6554
rect 21066 6502 21078 6554
rect 21130 6502 21142 6554
rect 21194 6502 21206 6554
rect 21258 6502 21264 6554
rect 20718 6352 20774 6361
rect 20718 6287 20774 6296
rect 20732 6254 20760 6287
rect 20720 6248 20772 6254
rect 20720 6190 20772 6196
rect 20810 5536 20866 5545
rect 20810 5471 20866 5480
rect 20444 4038 20496 4044
rect 20444 3980 20496 3986
rect 20626 4040 20682 4049
rect 20626 3975 20682 3984
rect 20824 3738 20852 5471
rect 20944 5466 21264 6502
rect 21604 6010 21924 7046
rect 22006 6624 22062 6633
rect 22006 6559 22062 6568
rect 22020 6118 22048 6559
rect 22008 6112 22060 6118
rect 22008 6054 22060 6060
rect 21604 5958 21610 6010
rect 21662 5958 21674 6010
rect 21726 5958 21738 6010
rect 21790 5958 21802 6010
rect 21854 5958 21866 6010
rect 21918 5958 21924 6010
rect 21456 5806 21508 5812
rect 21456 5748 21508 5754
rect 20944 5414 20950 5466
rect 21002 5414 21014 5466
rect 21066 5414 21078 5466
rect 21130 5414 21142 5466
rect 21194 5414 21206 5466
rect 21258 5414 21264 5466
rect 20944 4692 21264 5414
rect 21468 5166 21496 5748
rect 21604 5352 21924 5958
rect 22468 5772 22520 5778
rect 22468 5714 22520 5720
rect 22006 5672 22062 5681
rect 22006 5607 22008 5616
rect 22060 5607 22062 5616
rect 22008 5578 22060 5584
rect 21456 5160 21508 5166
rect 21456 5102 21508 5108
rect 20944 4396 20956 4692
rect 21252 4396 21264 4692
rect 20944 4378 21264 4396
rect 20944 4326 20950 4378
rect 21002 4326 21014 4378
rect 21066 4326 21078 4378
rect 21130 4326 21142 4378
rect 21194 4326 21206 4378
rect 21258 4326 21264 4378
rect 20812 3732 20864 3738
rect 20812 3674 20864 3680
rect 20628 3596 20680 3602
rect 20628 3538 20680 3544
rect 20350 2952 20406 2961
rect 20350 2887 20406 2896
rect 20258 1592 20314 1601
rect 20258 1527 20314 1536
rect 20258 1184 20314 1193
rect 20258 1119 20314 1128
rect 20272 1018 20300 1119
rect 20168 1012 20220 1018
rect 20168 954 20220 960
rect 20260 1012 20312 1018
rect 20260 954 20312 960
rect 19248 944 19300 950
rect 19248 886 19300 892
rect 20260 808 20312 814
rect 20364 785 20392 2887
rect 20444 2848 20496 2854
rect 20444 2790 20496 2796
rect 20456 1902 20484 2790
rect 20534 2544 20590 2553
rect 20640 2514 20668 3538
rect 20720 3392 20772 3398
rect 20720 3334 20772 3340
rect 20732 3058 20760 3334
rect 20944 3290 21264 4326
rect 21604 5056 21616 5352
rect 21912 5056 21924 5352
rect 21604 4922 21924 5056
rect 21604 4870 21610 4922
rect 21662 4870 21674 4922
rect 21726 4870 21738 4922
rect 21790 4870 21802 4922
rect 21854 4870 21866 4922
rect 21918 4870 21924 4922
rect 21604 3834 21924 4870
rect 22008 4684 22060 4690
rect 22008 4626 22060 4632
rect 22284 4684 22336 4690
rect 22284 4626 22336 4632
rect 22020 3942 22048 4626
rect 22192 4480 22244 4486
rect 22192 4422 22244 4428
rect 22098 4312 22154 4321
rect 22098 4247 22154 4256
rect 22008 3936 22060 3942
rect 22008 3878 22060 3884
rect 21604 3782 21610 3834
rect 21662 3782 21674 3834
rect 21726 3782 21738 3834
rect 21790 3782 21802 3834
rect 21854 3782 21866 3834
rect 21918 3782 21924 3834
rect 21362 3768 21418 3777
rect 21362 3703 21418 3712
rect 20944 3238 20950 3290
rect 21002 3238 21014 3290
rect 21066 3238 21078 3290
rect 21130 3238 21142 3290
rect 21194 3238 21206 3290
rect 21258 3238 21264 3290
rect 20720 3052 20772 3058
rect 20720 2994 20772 3000
rect 20718 2680 20774 2689
rect 20718 2615 20720 2624
rect 20772 2615 20774 2624
rect 20720 2586 20772 2592
rect 20534 2479 20590 2488
rect 20628 2508 20680 2514
rect 20548 2378 20576 2479
rect 20628 2450 20680 2456
rect 20812 2440 20864 2446
rect 20812 2382 20864 2388
rect 20536 2372 20588 2378
rect 20536 2314 20588 2320
rect 20720 2304 20772 2310
rect 20534 2272 20590 2281
rect 20720 2246 20772 2252
rect 20534 2207 20590 2216
rect 20548 1970 20576 2207
rect 20732 1986 20760 2246
rect 20824 2038 20852 2382
rect 20944 2202 21264 3238
rect 21376 2990 21404 3703
rect 21364 2984 21416 2990
rect 21364 2926 21416 2932
rect 20944 2150 20950 2202
rect 21002 2150 21014 2202
rect 21066 2150 21078 2202
rect 21130 2150 21142 2202
rect 21194 2150 21206 2202
rect 21258 2150 21264 2202
rect 20536 1964 20588 1970
rect 20536 1906 20588 1912
rect 20640 1958 20760 1986
rect 20812 2032 20864 2038
rect 20812 1974 20864 1980
rect 20444 1896 20496 1902
rect 20444 1838 20496 1844
rect 20640 1306 20668 1958
rect 20720 1828 20772 1834
rect 20720 1770 20772 1776
rect 20732 1426 20760 1770
rect 20720 1420 20772 1426
rect 20720 1362 20772 1368
rect 20640 1278 20760 1306
rect 20260 750 20312 756
rect 20350 776 20406 785
rect 20272 649 20300 750
rect 20350 711 20406 720
rect 20258 640 20314 649
rect 20258 575 20314 584
rect 18972 400 19024 406
rect 20732 377 20760 1278
rect 18972 342 19024 348
rect 20718 368 20774 377
rect 20718 303 20774 312
rect 20824 202 20852 1974
rect 20944 1114 21264 2150
rect 21604 2746 21924 3782
rect 22112 3738 22140 4247
rect 22204 4185 22232 4422
rect 22190 4176 22246 4185
rect 22190 4111 22246 4120
rect 22100 3732 22152 3738
rect 22100 3674 22152 3680
rect 22100 3596 22152 3602
rect 22100 3538 22152 3544
rect 22192 3596 22244 3602
rect 22192 3538 22244 3544
rect 22112 3194 22140 3538
rect 22100 3188 22152 3194
rect 22100 3130 22152 3136
rect 21604 2694 21610 2746
rect 21662 2694 21674 2746
rect 21726 2694 21738 2746
rect 21790 2694 21802 2746
rect 21854 2694 21866 2746
rect 21918 2694 21924 2746
rect 21362 2136 21418 2145
rect 21362 2071 21418 2080
rect 21376 1465 21404 2071
rect 21456 1828 21508 1834
rect 21456 1770 21508 1776
rect 21468 1562 21496 1770
rect 21604 1658 21924 2694
rect 22008 2372 22060 2378
rect 22008 2314 22060 2320
rect 22020 2122 22048 2314
rect 22020 2094 22140 2122
rect 22204 2106 22232 3538
rect 22006 2000 22062 2009
rect 22006 1935 22062 1944
rect 22020 1902 22048 1935
rect 22008 1896 22060 1902
rect 22008 1838 22060 1844
rect 21604 1606 21610 1658
rect 21662 1606 21674 1658
rect 21726 1606 21738 1658
rect 21790 1606 21802 1658
rect 21854 1606 21866 1658
rect 21918 1606 21924 1658
rect 21456 1556 21508 1562
rect 21456 1498 21508 1504
rect 21362 1456 21418 1465
rect 21362 1391 21364 1400
rect 21416 1391 21418 1400
rect 21364 1362 21416 1368
rect 20944 1062 20950 1114
rect 21002 1062 21014 1114
rect 21066 1062 21078 1114
rect 21130 1062 21142 1114
rect 21194 1062 21206 1114
rect 21258 1062 21264 1114
rect 20944 496 21264 1062
rect 21364 808 21416 814
rect 21362 776 21364 785
rect 21416 776 21418 785
rect 21362 711 21418 720
rect 21376 270 21404 711
rect 21604 570 21924 1606
rect 22020 1358 22048 1838
rect 22008 1352 22060 1358
rect 22008 1294 22060 1300
rect 22112 1170 22140 2094
rect 22192 2100 22244 2106
rect 22192 2042 22244 2048
rect 22296 2038 22324 4626
rect 22480 3777 22508 5714
rect 22664 5658 22692 7262
rect 22756 5817 22784 7822
rect 23204 7744 23256 7750
rect 23204 7686 23256 7692
rect 22836 6894 22888 6900
rect 22836 6836 22888 6842
rect 22848 6633 22876 6836
rect 22834 6624 22890 6633
rect 22834 6559 22890 6568
rect 23216 6225 23244 7686
rect 23308 7002 23336 7890
rect 23296 6996 23348 7002
rect 23296 6938 23348 6944
rect 23296 6792 23348 6798
rect 23296 6734 23348 6740
rect 23308 6497 23336 6734
rect 23294 6488 23350 6497
rect 23294 6423 23350 6432
rect 23202 6216 23258 6225
rect 23202 6151 23258 6160
rect 22742 5808 22798 5817
rect 23202 5808 23258 5817
rect 22742 5743 22798 5752
rect 23112 5772 23164 5778
rect 23202 5743 23204 5752
rect 23112 5714 23164 5720
rect 23256 5743 23258 5752
rect 23480 5772 23532 5778
rect 23204 5714 23256 5720
rect 23480 5714 23532 5720
rect 22572 5630 22692 5658
rect 22744 5704 22796 5710
rect 22744 5646 22796 5652
rect 22466 3768 22522 3777
rect 22466 3703 22522 3712
rect 22376 2916 22428 2922
rect 22376 2858 22428 2864
rect 22388 2514 22416 2858
rect 22376 2508 22428 2514
rect 22376 2450 22428 2456
rect 22376 2304 22428 2310
rect 22376 2246 22428 2252
rect 22284 2032 22336 2038
rect 22284 1974 22336 1980
rect 22388 1766 22416 2246
rect 22480 2038 22508 3703
rect 22572 2106 22600 5630
rect 22756 4690 22784 5646
rect 22744 4684 22796 4690
rect 22744 4626 22796 4632
rect 23020 4684 23072 4690
rect 23020 4626 23072 4632
rect 22652 3732 22704 3738
rect 22652 3674 22704 3680
rect 22560 2100 22612 2106
rect 22560 2042 22612 2048
rect 22468 2032 22520 2038
rect 22468 1974 22520 1980
rect 22376 1760 22428 1766
rect 22190 1728 22246 1737
rect 22376 1702 22428 1708
rect 22190 1663 22246 1672
rect 22204 1494 22232 1663
rect 22192 1488 22244 1494
rect 22192 1430 22244 1436
rect 21604 518 21610 570
rect 21662 518 21674 570
rect 21726 518 21738 570
rect 21790 518 21802 570
rect 21854 518 21866 570
rect 21918 518 21924 570
rect 21604 496 21924 518
rect 22020 1142 22140 1170
rect 22020 338 22048 1142
rect 22204 882 22232 1430
rect 22664 1290 22692 3674
rect 23032 3602 23060 4626
rect 23020 3596 23072 3602
rect 23020 3538 23072 3544
rect 23020 3120 23072 3126
rect 23020 3062 23072 3068
rect 23032 2854 23060 3062
rect 23020 2848 23072 2854
rect 23020 2790 23072 2796
rect 23032 2310 23060 2790
rect 22836 2304 22888 2310
rect 22836 2246 22888 2252
rect 23020 2304 23072 2310
rect 23020 2246 23072 2252
rect 22744 1896 22796 1902
rect 22744 1838 22796 1844
rect 22652 1284 22704 1290
rect 22652 1226 22704 1232
rect 22756 1057 22784 1838
rect 22848 1562 22876 2246
rect 22836 1556 22888 1562
rect 22836 1498 22888 1504
rect 22742 1048 22798 1057
rect 22742 983 22798 992
rect 22192 876 22244 882
rect 22192 818 22244 824
rect 22100 740 22152 746
rect 22100 682 22152 688
rect 22112 649 22140 682
rect 22098 640 22154 649
rect 22098 575 22154 584
rect 23124 474 23152 5714
rect 23492 5166 23520 5714
rect 23480 5160 23532 5166
rect 23480 5102 23532 5108
rect 23676 4826 23704 10095
rect 24044 10010 24072 11086
rect 24136 10130 24164 11290
rect 24308 11008 24360 11014
rect 24308 10950 24360 10956
rect 24124 10124 24176 10130
rect 24124 10066 24176 10072
rect 24216 10124 24268 10130
rect 24216 10066 24268 10072
rect 24044 9994 24164 10010
rect 24044 9988 24176 9994
rect 24044 9982 24124 9988
rect 24124 9930 24176 9936
rect 24136 8974 24164 9930
rect 24228 9110 24256 10066
rect 24216 9104 24268 9110
rect 24216 9046 24268 9052
rect 24124 8968 24176 8974
rect 24124 8910 24176 8916
rect 23756 8832 23808 8838
rect 23756 8774 23808 8780
rect 23768 7313 23796 8774
rect 24136 7993 24164 8910
rect 24216 8084 24268 8090
rect 24320 8072 24348 10950
rect 24400 9036 24452 9042
rect 24400 8978 24452 8984
rect 24584 9036 24636 9042
rect 24584 8978 24636 8984
rect 24268 8044 24348 8072
rect 24216 8026 24268 8032
rect 24122 7984 24178 7993
rect 24122 7919 24178 7928
rect 24124 7812 24176 7818
rect 24124 7754 24176 7760
rect 23754 7304 23810 7313
rect 23754 7239 23810 7248
rect 24136 6934 24164 7754
rect 24412 7410 24440 8978
rect 24596 7988 24624 8978
rect 24768 8832 24820 8838
rect 24768 8774 24820 8780
rect 24780 8106 24808 8774
rect 25056 8242 25084 11319
rect 25320 11212 25372 11218
rect 25320 11154 25372 11160
rect 25136 11144 25188 11150
rect 25332 11098 25360 11154
rect 25188 11092 25360 11098
rect 25136 11086 25360 11092
rect 25148 11070 25360 11086
rect 25700 10572 25728 11562
rect 29932 11354 29960 11630
rect 27712 11348 27764 11354
rect 27712 11290 27764 11296
rect 29920 11348 29972 11354
rect 29920 11290 29972 11296
rect 27250 11248 27306 11257
rect 25872 11212 25924 11218
rect 25872 11154 25924 11160
rect 26884 11212 26936 11218
rect 27250 11183 27252 11192
rect 26884 11154 26936 11160
rect 27304 11183 27306 11192
rect 27252 11154 27304 11160
rect 25884 11098 25912 11154
rect 26240 11144 26292 11150
rect 25884 11092 26240 11098
rect 25884 11086 26292 11092
rect 25884 11070 26280 11086
rect 25688 10566 25740 10572
rect 25688 10508 25740 10514
rect 26056 10464 26108 10470
rect 26054 10432 26056 10441
rect 26108 10432 26110 10441
rect 26054 10367 26110 10376
rect 25964 10158 26016 10164
rect 25148 10118 25964 10146
rect 25148 9382 25176 10118
rect 25964 10100 26016 10106
rect 26792 10124 26844 10130
rect 26792 10066 26844 10072
rect 26804 9518 26832 10066
rect 26792 9512 26844 9518
rect 26792 9454 26844 9460
rect 25136 9376 25188 9382
rect 25136 9318 25188 9324
rect 26056 8356 26108 8362
rect 26056 8298 26108 8304
rect 25056 8214 25728 8242
rect 24780 8090 25636 8106
rect 24780 8084 25648 8090
rect 24780 8078 25596 8084
rect 25596 8026 25648 8032
rect 24584 7982 24636 7988
rect 24584 7924 24636 7930
rect 25410 7984 25466 7993
rect 25410 7919 25466 7928
rect 25134 7712 25190 7721
rect 25134 7647 25190 7656
rect 25148 7546 25176 7647
rect 25136 7540 25188 7546
rect 25136 7482 25188 7488
rect 24400 7404 24452 7410
rect 24400 7346 24452 7352
rect 25424 7342 25452 7919
rect 25700 7342 25728 8214
rect 26068 7954 26096 8298
rect 26896 8090 26924 11154
rect 27250 11112 27306 11121
rect 27250 11047 27306 11056
rect 26974 9616 27030 9625
rect 26974 9551 27030 9560
rect 26884 8084 26936 8090
rect 26884 8026 26936 8032
rect 26988 7954 27016 9551
rect 27264 9042 27292 11047
rect 27618 10840 27674 10849
rect 27618 10775 27674 10784
rect 27436 9478 27488 9484
rect 27436 9420 27488 9426
rect 27448 9178 27476 9420
rect 27436 9172 27488 9178
rect 27436 9114 27488 9120
rect 27160 9036 27212 9042
rect 27160 8978 27212 8984
rect 27252 9036 27304 9042
rect 27252 8978 27304 8984
rect 27172 8430 27200 8978
rect 27632 8974 27660 10775
rect 27724 9110 27752 11290
rect 27896 11212 27948 11218
rect 27896 11154 27948 11160
rect 27908 10985 27936 11154
rect 27894 10976 27950 10985
rect 27894 10911 27950 10920
rect 30208 10810 30236 11902
rect 30748 11892 30800 11898
rect 30748 11834 30800 11840
rect 30760 10810 30788 11834
rect 30944 10906 31264 11472
rect 30944 10854 30950 10906
rect 31002 10854 31014 10906
rect 31066 10854 31078 10906
rect 31130 10854 31142 10906
rect 31194 10854 31206 10906
rect 31258 10854 31264 10906
rect 30196 10804 30248 10810
rect 30196 10746 30248 10752
rect 30748 10804 30800 10810
rect 30748 10746 30800 10752
rect 29920 10532 29972 10538
rect 29920 10474 29972 10480
rect 28356 10464 28408 10470
rect 28408 10424 28580 10452
rect 28356 10406 28408 10412
rect 28552 10164 28580 10424
rect 28540 10158 28592 10164
rect 29932 10130 29960 10474
rect 28540 10100 28592 10106
rect 29920 10124 29972 10130
rect 29920 10066 29972 10072
rect 30944 9818 31264 10854
rect 30944 9766 30950 9818
rect 31002 9766 31014 9818
rect 31066 9766 31078 9818
rect 31130 9766 31142 9818
rect 31194 9766 31206 9818
rect 31258 9766 31264 9818
rect 30654 9616 30710 9625
rect 30654 9551 30710 9560
rect 29184 9512 29236 9518
rect 29184 9454 29236 9460
rect 29644 9512 29696 9518
rect 29644 9454 29696 9460
rect 27712 9104 27764 9110
rect 27712 9046 27764 9052
rect 27620 8968 27672 8974
rect 27250 8936 27306 8945
rect 27620 8910 27672 8916
rect 28540 8968 28592 8974
rect 28540 8910 28592 8916
rect 27250 8871 27252 8880
rect 27304 8871 27306 8880
rect 27252 8842 27304 8848
rect 28356 8832 28408 8838
rect 28356 8774 28408 8780
rect 27160 8424 27212 8430
rect 27160 8366 27212 8372
rect 26056 7948 26108 7954
rect 26056 7890 26108 7896
rect 26976 7948 27028 7954
rect 26976 7890 27028 7896
rect 27066 7848 27122 7857
rect 26332 7812 26384 7818
rect 27066 7783 27122 7792
rect 26332 7754 26384 7760
rect 26240 7744 26292 7750
rect 26240 7686 26292 7692
rect 26252 7585 26280 7686
rect 26238 7576 26294 7585
rect 26238 7511 26294 7520
rect 24216 7336 24268 7342
rect 24216 7278 24268 7284
rect 25412 7336 25464 7342
rect 25412 7278 25464 7284
rect 25688 7336 25740 7342
rect 26240 7336 26292 7342
rect 25688 7278 25740 7284
rect 26160 7284 26240 7290
rect 26160 7278 26292 7284
rect 24124 6928 24176 6934
rect 24124 6870 24176 6876
rect 24228 6254 24256 7278
rect 26160 7262 26280 7278
rect 24768 7200 24820 7206
rect 24768 7142 24820 7148
rect 24780 7041 24808 7142
rect 24766 7032 24822 7041
rect 24766 6967 24822 6976
rect 24780 6798 24808 6967
rect 25228 6860 25280 6866
rect 25228 6802 25280 6808
rect 25872 6860 25924 6866
rect 25872 6802 25924 6808
rect 24768 6792 24820 6798
rect 24768 6734 24820 6740
rect 24860 6656 24912 6662
rect 24860 6598 24912 6604
rect 24216 6248 24268 6254
rect 24216 6190 24268 6196
rect 24308 6248 24360 6254
rect 24308 6190 24360 6196
rect 24320 5132 24348 6190
rect 24308 5126 24360 5132
rect 24308 5068 24360 5074
rect 23664 4820 23716 4826
rect 23664 4762 23716 4768
rect 23480 4684 23532 4690
rect 23480 4626 23532 4632
rect 23204 3732 23256 3738
rect 23204 3674 23256 3680
rect 23216 3058 23244 3674
rect 23204 3052 23256 3058
rect 23204 2994 23256 3000
rect 23296 2984 23348 2990
rect 23294 2952 23296 2961
rect 23348 2952 23350 2961
rect 23294 2887 23350 2896
rect 23296 2508 23348 2514
rect 23296 2450 23348 2456
rect 23204 2372 23256 2378
rect 23204 2314 23256 2320
rect 23216 1834 23244 2314
rect 23204 1828 23256 1834
rect 23204 1770 23256 1776
rect 23216 882 23244 1770
rect 23204 876 23256 882
rect 23204 818 23256 824
rect 23308 513 23336 2450
rect 23388 1284 23440 1290
rect 23388 1226 23440 1232
rect 23400 678 23428 1226
rect 23492 1193 23520 4626
rect 23676 2106 23704 4762
rect 23940 4684 23992 4690
rect 23940 4626 23992 4632
rect 23756 4480 23808 4486
rect 23756 4422 23808 4428
rect 23768 3398 23796 4422
rect 23952 4078 23980 4626
rect 23940 4072 23992 4078
rect 23940 4014 23992 4020
rect 24308 4038 24360 4044
rect 24308 3980 24360 3986
rect 24320 3602 24348 3980
rect 24308 3596 24360 3602
rect 24308 3538 24360 3544
rect 24872 3534 24900 6598
rect 25240 5953 25268 6802
rect 25884 6089 25912 6802
rect 25870 6080 25926 6089
rect 25870 6015 25926 6024
rect 25226 5944 25282 5953
rect 25226 5879 25282 5888
rect 25964 5806 26016 5812
rect 25964 5748 26016 5754
rect 25976 5166 26004 5748
rect 25964 5160 26016 5166
rect 25964 5102 26016 5108
rect 25964 4718 26016 4724
rect 25964 4660 26016 4666
rect 25976 4078 26004 4660
rect 25964 4072 26016 4078
rect 25964 4014 26016 4020
rect 24860 3528 24912 3534
rect 24860 3470 24912 3476
rect 23756 3392 23808 3398
rect 23756 3334 23808 3340
rect 23768 3194 23796 3334
rect 23938 3224 23994 3233
rect 23756 3188 23808 3194
rect 23938 3159 23994 3168
rect 23756 3130 23808 3136
rect 23952 2990 23980 3159
rect 24582 3088 24638 3097
rect 24582 3023 24638 3032
rect 24596 2990 24624 3023
rect 23848 2984 23900 2990
rect 23848 2926 23900 2932
rect 23940 2984 23992 2990
rect 23940 2926 23992 2932
rect 24584 2984 24636 2990
rect 24584 2926 24636 2932
rect 23664 2100 23716 2106
rect 23664 2042 23716 2048
rect 23676 1494 23704 2042
rect 23664 1488 23716 1494
rect 23664 1430 23716 1436
rect 23478 1184 23534 1193
rect 23478 1119 23534 1128
rect 23860 950 23888 2926
rect 23952 2650 23980 2926
rect 26056 2848 26108 2854
rect 26056 2790 26108 2796
rect 23940 2644 23992 2650
rect 23940 2586 23992 2592
rect 24216 2304 24268 2310
rect 24216 2246 24268 2252
rect 24228 2038 24256 2246
rect 26068 2106 26096 2790
rect 26056 2100 26108 2106
rect 26056 2042 26108 2048
rect 24216 2032 24268 2038
rect 24216 1974 24268 1980
rect 23940 1760 23992 1766
rect 23940 1702 23992 1708
rect 23952 1018 23980 1702
rect 24858 1456 24914 1465
rect 24858 1391 24914 1400
rect 24872 1358 24900 1391
rect 24860 1352 24912 1358
rect 24860 1294 24912 1300
rect 26160 1290 26188 7262
rect 26344 6730 26372 7754
rect 27080 7546 27108 7783
rect 28264 7744 28316 7750
rect 28264 7686 28316 7692
rect 28276 7546 28304 7686
rect 27068 7540 27120 7546
rect 27068 7482 27120 7488
rect 28264 7540 28316 7546
rect 28264 7482 28316 7488
rect 27618 7440 27674 7449
rect 27618 7375 27620 7384
rect 27672 7375 27674 7384
rect 27620 7346 27672 7352
rect 28368 7274 28396 8774
rect 28552 8090 28580 8910
rect 28816 8390 28868 8396
rect 28816 8332 28868 8338
rect 28828 8265 28856 8332
rect 28814 8256 28870 8265
rect 28814 8191 28870 8200
rect 28540 8084 28592 8090
rect 28540 8026 28592 8032
rect 29196 8022 29224 9454
rect 29656 9178 29684 9454
rect 30668 9178 30696 9551
rect 29644 9172 29696 9178
rect 29644 9114 29696 9120
rect 30656 9172 30708 9178
rect 30656 9114 30708 9120
rect 29366 8936 29422 8945
rect 29276 8900 29328 8906
rect 29366 8871 29422 8880
rect 29276 8842 29328 8848
rect 29288 8430 29316 8842
rect 29276 8424 29328 8430
rect 29276 8366 29328 8372
rect 29184 8016 29236 8022
rect 29184 7958 29236 7964
rect 28356 7268 28408 7274
rect 28356 7210 28408 7216
rect 28540 7200 28592 7206
rect 28540 7142 28592 7148
rect 28816 7200 28868 7206
rect 28816 7142 28868 7148
rect 26332 6724 26384 6730
rect 26332 6666 26384 6672
rect 26344 4049 26372 6666
rect 26884 6656 26936 6662
rect 26884 6598 26936 6604
rect 26896 6361 26924 6598
rect 26882 6352 26938 6361
rect 28552 6322 28580 7142
rect 28828 7002 28856 7142
rect 28816 6996 28868 7002
rect 28816 6938 28868 6944
rect 29090 6760 29146 6769
rect 29090 6695 29092 6704
rect 29144 6695 29146 6704
rect 29092 6666 29144 6672
rect 26882 6287 26938 6296
rect 27160 6316 27212 6322
rect 27160 6258 27212 6264
rect 28540 6316 28592 6322
rect 28540 6258 28592 6264
rect 26792 6180 26844 6186
rect 26792 6122 26844 6128
rect 26804 5778 26832 6122
rect 26792 5772 26844 5778
rect 26792 5714 26844 5720
rect 27172 5545 27200 6258
rect 27620 6248 27672 6254
rect 27620 6190 27672 6196
rect 27158 5536 27214 5545
rect 27158 5471 27214 5480
rect 27436 5126 27488 5132
rect 27632 5114 27660 6190
rect 28908 5772 28960 5778
rect 28908 5714 28960 5720
rect 28920 5166 28948 5714
rect 27488 5086 27660 5114
rect 28908 5160 28960 5166
rect 28908 5102 28960 5108
rect 27436 5068 27488 5074
rect 28448 5024 28500 5030
rect 28448 4966 28500 4972
rect 28460 4865 28488 4966
rect 28446 4856 28502 4865
rect 28446 4791 28502 4800
rect 28540 4718 28592 4724
rect 26792 4684 26844 4690
rect 28540 4660 28592 4666
rect 29184 4684 29236 4690
rect 26792 4626 26844 4632
rect 26330 4040 26386 4049
rect 26330 3975 26386 3984
rect 26804 3670 26832 4626
rect 27620 3936 27672 3942
rect 27620 3878 27672 3884
rect 27632 3738 27660 3878
rect 28552 3738 28580 4660
rect 29184 4626 29236 4632
rect 29196 4078 29224 4626
rect 29184 4072 29236 4078
rect 29184 4014 29236 4020
rect 27620 3732 27672 3738
rect 27620 3674 27672 3680
rect 28540 3732 28592 3738
rect 28540 3674 28592 3680
rect 29380 3670 29408 8871
rect 30944 8730 31264 9766
rect 31604 11450 31924 11472
rect 31604 11398 31610 11450
rect 31662 11398 31674 11450
rect 31726 11398 31738 11450
rect 31790 11398 31802 11450
rect 31854 11398 31866 11450
rect 31918 11398 31924 11450
rect 31604 10362 31924 11398
rect 31604 10310 31610 10362
rect 31662 10310 31674 10362
rect 31726 10310 31738 10362
rect 31790 10310 31802 10362
rect 31854 10310 31866 10362
rect 31918 10310 31924 10362
rect 31390 9616 31446 9625
rect 31390 9551 31446 9560
rect 31404 9484 31432 9551
rect 31392 9478 31444 9484
rect 31392 9420 31444 9426
rect 30944 8678 30950 8730
rect 31002 8692 31014 8730
rect 31066 8692 31078 8730
rect 31130 8692 31142 8730
rect 31194 8692 31206 8730
rect 31258 8678 31264 8730
rect 30944 8396 30956 8678
rect 31252 8396 31264 8678
rect 29920 7880 29972 7886
rect 29920 7822 29972 7828
rect 29932 7002 29960 7822
rect 30944 7642 31264 8396
rect 30944 7590 30950 7642
rect 31002 7590 31014 7642
rect 31066 7590 31078 7642
rect 31130 7590 31142 7642
rect 31194 7590 31206 7642
rect 31258 7590 31264 7642
rect 29920 6996 29972 7002
rect 29920 6938 29972 6944
rect 30654 6896 30710 6905
rect 30654 6831 30710 6840
rect 30668 6458 30696 6831
rect 30944 6554 31264 7590
rect 30944 6502 30950 6554
rect 31002 6502 31014 6554
rect 31066 6502 31078 6554
rect 31130 6502 31142 6554
rect 31194 6502 31206 6554
rect 31258 6502 31264 6554
rect 30656 6452 30708 6458
rect 30656 6394 30708 6400
rect 29828 6214 29880 6220
rect 29828 6156 29880 6162
rect 29840 5778 29868 6156
rect 29828 5772 29880 5778
rect 29828 5714 29880 5720
rect 30944 5466 31264 6502
rect 30944 5414 30950 5466
rect 31002 5414 31014 5466
rect 31066 5414 31078 5466
rect 31130 5414 31142 5466
rect 31194 5414 31206 5466
rect 31258 5414 31264 5466
rect 30944 4692 31264 5414
rect 31604 9352 31924 10310
rect 32036 10124 32088 10130
rect 32036 10066 32088 10072
rect 31604 9274 31616 9352
rect 31912 9274 31924 9352
rect 31604 9222 31610 9274
rect 31918 9222 31924 9274
rect 31604 9056 31616 9222
rect 31912 9056 31924 9222
rect 31604 8186 31924 9056
rect 31604 8134 31610 8186
rect 31662 8134 31674 8186
rect 31726 8134 31738 8186
rect 31790 8134 31802 8186
rect 31854 8134 31866 8186
rect 31918 8134 31924 8186
rect 31604 7098 31924 8134
rect 32048 7954 32076 10066
rect 32128 9036 32180 9042
rect 32128 8978 32180 8984
rect 32140 8430 32168 8978
rect 32128 8424 32180 8430
rect 32128 8366 32180 8372
rect 32036 7948 32088 7954
rect 32036 7890 32088 7896
rect 31604 7046 31610 7098
rect 31662 7046 31674 7098
rect 31726 7046 31738 7098
rect 31790 7046 31802 7098
rect 31854 7046 31866 7098
rect 31918 7046 31924 7098
rect 31604 6010 31924 7046
rect 32036 6724 32088 6730
rect 32036 6666 32088 6672
rect 31604 5958 31610 6010
rect 31662 5958 31674 6010
rect 31726 5958 31738 6010
rect 31790 5958 31802 6010
rect 31854 5958 31866 6010
rect 31918 5958 31924 6010
rect 31604 5352 31924 5958
rect 32048 5846 32076 6666
rect 32036 5840 32088 5846
rect 32036 5782 32088 5788
rect 31604 5056 31616 5352
rect 31912 5056 31924 5352
rect 31484 5024 31536 5030
rect 31484 4966 31536 4972
rect 30944 4396 30956 4692
rect 31252 4396 31264 4692
rect 30944 4378 31264 4396
rect 30944 4326 30950 4378
rect 31002 4326 31014 4378
rect 31066 4326 31078 4378
rect 31130 4326 31142 4378
rect 31194 4326 31206 4378
rect 31258 4326 31264 4378
rect 30012 4038 30064 4044
rect 30012 3980 30064 3986
rect 30024 3738 30052 3980
rect 30012 3732 30064 3738
rect 30012 3674 30064 3680
rect 26792 3664 26844 3670
rect 27160 3664 27212 3670
rect 26792 3606 26844 3612
rect 26882 3632 26938 3641
rect 27160 3606 27212 3612
rect 29368 3664 29420 3670
rect 29368 3606 29420 3612
rect 26882 3567 26884 3576
rect 26936 3567 26938 3576
rect 26884 3538 26936 3544
rect 27172 3369 27200 3606
rect 29000 3596 29052 3602
rect 29000 3538 29052 3544
rect 27620 3392 27672 3398
rect 27158 3360 27214 3369
rect 27620 3334 27672 3340
rect 27158 3295 27214 3304
rect 27632 3194 27660 3334
rect 27620 3188 27672 3194
rect 27620 3130 27672 3136
rect 29012 2961 29040 3538
rect 30944 3290 31264 4326
rect 31496 3738 31524 4966
rect 31604 4922 31924 5056
rect 31604 4870 31610 4922
rect 31662 4870 31674 4922
rect 31726 4870 31738 4922
rect 31790 4870 31802 4922
rect 31854 4870 31866 4922
rect 31918 4870 31924 4922
rect 31604 3834 31924 4870
rect 32036 4684 32088 4690
rect 32036 4626 32088 4632
rect 32048 4078 32076 4626
rect 32036 4072 32088 4078
rect 32036 4014 32088 4020
rect 31604 3782 31610 3834
rect 31662 3782 31674 3834
rect 31726 3782 31738 3834
rect 31790 3782 31802 3834
rect 31854 3782 31866 3834
rect 31918 3782 31924 3834
rect 31484 3732 31536 3738
rect 31484 3674 31536 3680
rect 30944 3238 30950 3290
rect 31002 3238 31014 3290
rect 31066 3238 31078 3290
rect 31130 3238 31142 3290
rect 31194 3238 31206 3290
rect 31258 3238 31264 3290
rect 28998 2952 29054 2961
rect 28998 2887 29054 2896
rect 27620 2848 27672 2854
rect 27618 2816 27620 2825
rect 27672 2816 27674 2825
rect 27618 2751 27674 2760
rect 30944 2202 31264 3238
rect 30944 2150 30950 2202
rect 31002 2150 31014 2202
rect 31066 2150 31078 2202
rect 31130 2150 31142 2202
rect 31194 2150 31206 2202
rect 31258 2150 31264 2202
rect 26148 1284 26200 1290
rect 26148 1226 26200 1232
rect 30944 1114 31264 2150
rect 30944 1062 30950 1114
rect 31002 1062 31014 1114
rect 31066 1062 31078 1114
rect 31130 1062 31142 1114
rect 31194 1062 31206 1114
rect 31258 1062 31264 1114
rect 23940 1012 23992 1018
rect 23940 954 23992 960
rect 23848 944 23900 950
rect 23848 886 23900 892
rect 24858 912 24914 921
rect 24858 847 24860 856
rect 24912 847 24914 856
rect 24860 818 24912 824
rect 24216 808 24268 814
rect 24214 776 24216 785
rect 24268 776 24270 785
rect 24214 711 24270 720
rect 23388 672 23440 678
rect 23388 614 23440 620
rect 23294 504 23350 513
rect 23112 468 23164 474
rect 30944 496 31264 1062
rect 31604 2746 31924 3782
rect 31604 2694 31610 2746
rect 31662 2694 31674 2746
rect 31726 2694 31738 2746
rect 31790 2694 31802 2746
rect 31854 2694 31866 2746
rect 31918 2694 31924 2746
rect 31604 1658 31924 2694
rect 31604 1606 31610 1658
rect 31662 1606 31674 1658
rect 31726 1606 31738 1658
rect 31790 1606 31802 1658
rect 31854 1606 31866 1658
rect 31918 1606 31924 1658
rect 31604 570 31924 1606
rect 31604 518 31610 570
rect 31662 518 31674 570
rect 31726 518 31738 570
rect 31790 518 31802 570
rect 31854 518 31866 570
rect 31918 518 31924 570
rect 31604 496 31924 518
rect 23294 439 23350 448
rect 23112 410 23164 416
rect 22008 332 22060 338
rect 22008 274 22060 280
rect 21364 264 21416 270
rect 21364 206 21416 212
rect 20812 196 20864 202
rect 20812 138 20864 144
rect 17958 96 18014 105
rect 12346 31 12402 40
rect 14464 60 14516 66
rect 10048 2 10100 8
rect 17958 31 18014 40
rect 14464 2 14516 8
<< via2 >>
rect 938 11620 994 11656
rect 938 11600 940 11620
rect 940 11600 992 11620
rect 992 11600 994 11620
rect 1030 11192 1086 11248
rect 938 9696 994 9752
rect 938 8744 994 8800
rect 2226 10158 2282 10160
rect 2226 10106 2228 10158
rect 2228 10106 2280 10158
rect 2280 10106 2282 10158
rect 2226 10104 2282 10106
rect 2226 9832 2282 9888
rect 2778 9696 2834 9752
rect 2870 8200 2926 8256
rect 2594 8064 2650 8120
rect 2686 7404 2742 7440
rect 2686 7384 2688 7404
rect 2688 7384 2740 7404
rect 2740 7384 2742 7404
rect 2410 5616 2466 5672
rect 938 4936 994 4992
rect 938 4120 994 4176
rect 3606 11464 3662 11520
rect 3514 10104 3570 10160
rect 3514 8880 3570 8936
rect 3790 11600 3846 11656
rect 4066 10784 4122 10840
rect 3974 10376 4030 10432
rect 12438 11892 12494 11928
rect 12438 11872 12440 11892
rect 12440 11872 12492 11892
rect 12492 11872 12494 11892
rect 20810 11872 20866 11928
rect 9310 11736 9366 11792
rect 12530 11736 12586 11792
rect 4710 11328 4766 11384
rect 4434 10648 4490 10704
rect 3882 9968 3938 10024
rect 4250 9696 4306 9752
rect 3698 8880 3754 8936
rect 3882 7948 3938 7984
rect 3882 7928 3884 7948
rect 3884 7928 3936 7948
rect 3936 7928 3938 7948
rect 4066 7792 4122 7848
rect 3606 7520 3662 7576
rect 3882 7520 3938 7576
rect 2962 5888 3018 5944
rect 1398 584 1454 640
rect 1674 2760 1730 2816
rect 3422 6024 3478 6080
rect 3606 5908 3662 5944
rect 3606 5888 3608 5908
rect 3608 5888 3660 5908
rect 3660 5888 3662 5908
rect 3974 6976 4030 7032
rect 3882 6840 3938 6896
rect 3882 6432 3938 6488
rect 3146 5480 3202 5536
rect 3330 5480 3386 5536
rect 3054 4120 3110 4176
rect 2778 1808 2834 1864
rect 2962 1808 3018 1864
rect 3422 3032 3478 3088
rect 3330 2352 3386 2408
rect 3054 584 3110 640
rect 6642 11056 6698 11112
rect 7654 10566 7710 10568
rect 7654 10514 7656 10566
rect 7656 10514 7708 10566
rect 7708 10514 7710 10566
rect 7654 10512 7710 10514
rect 8206 9968 8262 10024
rect 5170 8200 5226 8256
rect 6550 7792 6606 7848
rect 6274 7656 6330 7712
rect 6550 7656 6606 7712
rect 5078 7302 5134 7304
rect 5078 7250 5080 7302
rect 5080 7250 5132 7302
rect 5132 7250 5134 7302
rect 5078 7248 5134 7250
rect 4434 6704 4490 6760
rect 6366 7248 6422 7304
rect 4802 6894 4858 6896
rect 4802 6842 4804 6894
rect 4804 6842 4856 6894
rect 4856 6842 4858 6894
rect 4802 6840 4858 6842
rect 6090 6840 6146 6896
rect 6274 6840 6330 6896
rect 4342 6568 4398 6624
rect 4250 6196 4252 6216
rect 4252 6196 4304 6216
rect 4304 6196 4306 6216
rect 4250 6160 4306 6196
rect 3790 4800 3846 4856
rect 3606 720 3662 776
rect 3422 448 3478 504
rect 3882 1264 3938 1320
rect 4526 4800 4582 4856
rect 4802 5806 4858 5808
rect 4802 5754 4804 5806
rect 4804 5754 4856 5806
rect 4856 5754 4858 5806
rect 4802 5752 4858 5754
rect 4250 3612 4252 3632
rect 4252 3612 4304 3632
rect 4304 3612 4306 3632
rect 4250 3576 4306 3612
rect 4250 3460 4306 3496
rect 4250 3440 4252 3460
rect 4252 3440 4304 3460
rect 4304 3440 4306 3460
rect 4066 2624 4122 2680
rect 3974 1128 4030 1184
rect 3790 312 3846 368
rect 4434 2896 4490 2952
rect 4618 3168 4674 3224
rect 4526 2080 4582 2136
rect 4802 2542 4858 2544
rect 4802 2490 4804 2542
rect 4804 2490 4856 2542
rect 4856 2490 4858 2542
rect 4802 2488 4858 2490
rect 4710 1944 4766 2000
rect 12162 11600 12218 11656
rect 9402 10240 9458 10296
rect 9770 10512 9826 10568
rect 10598 10920 10654 10976
rect 10322 10784 10378 10840
rect 9862 8200 9918 8256
rect 10046 8200 10102 8256
rect 8482 7792 8538 7848
rect 9494 7520 9550 7576
rect 9494 7384 9550 7440
rect 9862 7384 9918 7440
rect 9770 7248 9826 7304
rect 9954 7112 10010 7168
rect 9954 6840 10010 6896
rect 10138 6840 10194 6896
rect 8850 6704 8906 6760
rect 9586 6568 9642 6624
rect 6642 6432 6698 6488
rect 6826 6432 6882 6488
rect 6090 5752 6146 5808
rect 5262 5616 5318 5672
rect 5446 5616 5502 5672
rect 4986 3848 5042 3904
rect 7010 6024 7066 6080
rect 7194 6024 7250 6080
rect 7010 5752 7066 5808
rect 10690 10512 10746 10568
rect 10782 10376 10838 10432
rect 10782 10104 10838 10160
rect 11334 10512 11390 10568
rect 12438 11328 12494 11384
rect 12346 11192 12402 11248
rect 12070 10784 12126 10840
rect 11978 10376 12034 10432
rect 11978 9696 12034 9752
rect 11616 9274 11912 9352
rect 11616 9222 11662 9274
rect 11662 9222 11674 9274
rect 11674 9222 11726 9274
rect 11726 9222 11738 9274
rect 11738 9222 11790 9274
rect 11790 9222 11802 9274
rect 11802 9222 11854 9274
rect 11854 9222 11866 9274
rect 11866 9222 11912 9274
rect 11616 9056 11912 9222
rect 10956 8678 11002 8692
rect 11002 8678 11014 8692
rect 11014 8678 11066 8692
rect 11066 8678 11078 8692
rect 11078 8678 11130 8692
rect 11130 8678 11142 8692
rect 11142 8678 11194 8692
rect 11194 8678 11206 8692
rect 11206 8678 11252 8692
rect 10956 8396 11252 8678
rect 11978 8200 12034 8256
rect 11426 8084 11482 8120
rect 11426 8064 11428 8084
rect 11428 8064 11480 8084
rect 11480 8064 11482 8084
rect 11334 7656 11390 7712
rect 17498 11600 17554 11656
rect 12898 10920 12954 10976
rect 12990 10784 13046 10840
rect 12438 10376 12494 10432
rect 12346 10240 12402 10296
rect 12346 9696 12402 9752
rect 12622 9696 12678 9752
rect 12438 8200 12494 8256
rect 12438 8064 12494 8120
rect 12438 7792 12494 7848
rect 12806 7792 12862 7848
rect 11334 6976 11390 7032
rect 11334 6840 11390 6896
rect 10230 5752 10286 5808
rect 10506 5772 10562 5808
rect 10506 5752 10508 5772
rect 10508 5752 10560 5772
rect 10560 5752 10562 5772
rect 9586 5480 9642 5536
rect 7746 4800 7802 4856
rect 7930 4800 7986 4856
rect 5722 4256 5778 4312
rect 5538 4156 5540 4176
rect 5540 4156 5592 4176
rect 5592 4156 5594 4176
rect 5538 4120 5594 4156
rect 5630 3984 5686 4040
rect 5446 3576 5502 3632
rect 5814 3576 5870 3632
rect 6918 3984 6974 4040
rect 7562 3712 7618 3768
rect 7746 3712 7802 3768
rect 4894 1672 4950 1728
rect 4342 856 4398 912
rect 1582 176 1638 232
rect 5446 3304 5502 3360
rect 6090 3476 6092 3496
rect 6092 3476 6144 3496
rect 6144 3476 6146 3496
rect 6090 3440 6146 3476
rect 7286 3440 7342 3496
rect 8206 3304 8262 3360
rect 6550 2488 6606 2544
rect 5906 2216 5962 2272
rect 6918 2508 6974 2544
rect 6918 2488 6920 2508
rect 6920 2488 6972 2508
rect 6972 2488 6974 2508
rect 7378 2896 7434 2952
rect 7562 2896 7618 2952
rect 7010 2352 7066 2408
rect 7378 2352 7434 2408
rect 8482 3304 8538 3360
rect 9494 2624 9550 2680
rect 9678 2624 9734 2680
rect 9954 176 10010 232
rect 9494 40 9550 96
rect 10956 4396 11252 4692
rect 11616 5056 11912 5352
rect 11334 3340 11336 3360
rect 11336 3340 11388 3360
rect 11388 3340 11390 3360
rect 11334 3304 11390 3340
rect 10506 1454 10562 1456
rect 10506 1402 10508 1454
rect 10508 1402 10560 1454
rect 10560 1402 10562 1454
rect 10506 1400 10562 1402
rect 12162 6976 12218 7032
rect 12714 7248 12770 7304
rect 12806 7112 12862 7168
rect 12530 6704 12586 6760
rect 13174 11056 13230 11112
rect 13358 11056 13414 11112
rect 15198 9716 15254 9752
rect 15198 9696 15200 9716
rect 15200 9696 15252 9716
rect 15252 9696 15254 9716
rect 15842 10376 15898 10432
rect 16486 10648 16542 10704
rect 17222 10648 17278 10704
rect 16302 10566 16358 10568
rect 16302 10514 16304 10566
rect 16304 10514 16356 10566
rect 16356 10514 16358 10566
rect 16302 10512 16358 10514
rect 13634 7656 13690 7712
rect 13174 7112 13230 7168
rect 15842 7928 15898 7984
rect 14830 7792 14886 7848
rect 14646 7520 14702 7576
rect 14830 7520 14886 7576
rect 15566 7792 15622 7848
rect 12254 6568 12310 6624
rect 12254 6432 12310 6488
rect 12714 6568 12770 6624
rect 12530 6160 12586 6216
rect 12898 6432 12954 6488
rect 12714 6160 12770 6216
rect 12530 6024 12586 6080
rect 12070 5752 12126 5808
rect 12070 4120 12126 4176
rect 12070 3848 12126 3904
rect 12254 4120 12310 4176
rect 13082 6568 13138 6624
rect 12990 5616 13046 5672
rect 13818 4800 13874 4856
rect 14002 4820 14058 4856
rect 14002 4800 14004 4820
rect 14004 4800 14056 4820
rect 14056 4800 14058 4820
rect 15290 5888 15346 5944
rect 15198 5480 15254 5536
rect 15658 6060 15660 6080
rect 15660 6060 15712 6080
rect 15712 6060 15714 6080
rect 15658 6024 15714 6060
rect 15382 5480 15438 5536
rect 13634 4120 13690 4176
rect 13818 4120 13874 4176
rect 14554 3712 14610 3768
rect 13450 3576 13506 3632
rect 11978 3460 12034 3496
rect 11978 3440 11980 3460
rect 11980 3440 12032 3460
rect 12032 3440 12034 3460
rect 15198 4800 15254 4856
rect 16854 9696 16910 9752
rect 17406 10240 17462 10296
rect 16854 8880 16910 8936
rect 16578 7928 16634 7984
rect 16578 6568 16634 6624
rect 17038 8880 17094 8936
rect 17774 11056 17830 11112
rect 17958 10920 18014 10976
rect 17590 10512 17646 10568
rect 17866 10376 17922 10432
rect 20442 11056 20498 11112
rect 20718 11464 20774 11520
rect 20626 10920 20682 10976
rect 19890 10648 19946 10704
rect 21638 11600 21694 11656
rect 21454 11328 21510 11384
rect 18970 10240 19026 10296
rect 18050 10140 18052 10160
rect 18052 10140 18104 10160
rect 18104 10140 18106 10160
rect 18050 10104 18106 10140
rect 18050 9968 18106 10024
rect 17866 8064 17922 8120
rect 18694 8200 18750 8256
rect 17222 6840 17278 6896
rect 17406 6840 17462 6896
rect 17038 6568 17094 6624
rect 15382 3848 15438 3904
rect 16210 3712 16266 3768
rect 14554 3304 14610 3360
rect 14922 3304 14978 3360
rect 12254 3168 12310 3224
rect 15934 3168 15990 3224
rect 16578 4120 16634 4176
rect 17038 6160 17094 6216
rect 17222 5888 17278 5944
rect 18510 7384 18566 7440
rect 18602 7112 18658 7168
rect 17958 6568 18014 6624
rect 17866 6452 17922 6488
rect 17866 6432 17868 6452
rect 17868 6432 17920 6452
rect 17920 6432 17922 6452
rect 19798 9968 19854 10024
rect 19338 9696 19394 9752
rect 20810 10648 20866 10704
rect 20258 10104 20314 10160
rect 19614 8064 19670 8120
rect 19890 8064 19946 8120
rect 19982 7792 20038 7848
rect 19246 7112 19302 7168
rect 19430 7112 19486 7168
rect 19246 6568 19302 6624
rect 19430 6568 19486 6624
rect 17866 6296 17922 6352
rect 18694 5652 18696 5672
rect 18696 5652 18748 5672
rect 18748 5652 18750 5672
rect 18694 5616 18750 5652
rect 18326 4800 18382 4856
rect 17314 4120 17370 4176
rect 16762 3712 16818 3768
rect 15014 2624 15070 2680
rect 12254 2352 12310 2408
rect 12392 2352 12448 2408
rect 12254 1808 12310 1864
rect 13082 1808 13138 1864
rect 12162 1672 12218 1728
rect 12990 1672 13046 1728
rect 12346 1420 12402 1456
rect 12346 1400 12348 1420
rect 12348 1400 12400 1420
rect 12400 1400 12402 1420
rect 12070 176 12126 232
rect 12346 40 12402 96
rect 15014 1400 15070 1456
rect 14922 856 14978 912
rect 15658 2488 15714 2544
rect 15842 2488 15898 2544
rect 17314 3168 17370 3224
rect 17958 3476 17960 3496
rect 17960 3476 18012 3496
rect 18012 3476 18014 3496
rect 17958 3440 18014 3476
rect 17314 2896 17370 2952
rect 17774 2896 17830 2952
rect 18142 4256 18198 4312
rect 18510 3984 18566 4040
rect 20258 7792 20314 7848
rect 20074 7656 20130 7712
rect 22006 11192 22062 11248
rect 22006 10412 22008 10432
rect 22008 10412 22060 10432
rect 22060 10412 22062 10432
rect 22006 10376 22062 10412
rect 21454 9716 21510 9752
rect 21454 9696 21456 9716
rect 21456 9696 21508 9716
rect 21508 9696 21510 9716
rect 22006 10260 22062 10296
rect 22006 10240 22008 10260
rect 22008 10240 22060 10260
rect 22060 10240 22062 10260
rect 22098 10140 22100 10160
rect 22100 10140 22152 10160
rect 22152 10140 22154 10160
rect 22098 10104 22154 10140
rect 22926 10648 22982 10704
rect 22098 9988 22154 10024
rect 22098 9968 22100 9988
rect 22100 9968 22152 9988
rect 22152 9968 22154 9988
rect 25042 11328 25098 11384
rect 23662 10104 23718 10160
rect 23478 9696 23534 9752
rect 21616 9274 21912 9352
rect 21616 9222 21662 9274
rect 21662 9222 21674 9274
rect 21674 9222 21726 9274
rect 21726 9222 21738 9274
rect 21738 9222 21790 9274
rect 21790 9222 21802 9274
rect 21802 9222 21854 9274
rect 21854 9222 21866 9274
rect 21866 9222 21912 9274
rect 21616 9056 21912 9222
rect 20956 8678 21002 8692
rect 21002 8678 21014 8692
rect 21014 8678 21066 8692
rect 21066 8678 21078 8692
rect 21078 8678 21130 8692
rect 21130 8678 21142 8692
rect 21142 8678 21194 8692
rect 21194 8678 21206 8692
rect 21206 8678 21252 8692
rect 20956 8396 21252 8678
rect 19614 5752 19670 5808
rect 19522 5616 19578 5672
rect 19890 5752 19946 5808
rect 20074 5480 20130 5536
rect 20166 2896 20222 2952
rect 19246 2624 19302 2680
rect 18602 2352 18658 2408
rect 18050 2080 18106 2136
rect 15842 1808 15898 1864
rect 17866 1808 17922 1864
rect 16026 1672 16082 1728
rect 15750 1128 15806 1184
rect 18418 1672 18474 1728
rect 18602 1708 18604 1728
rect 18604 1708 18656 1728
rect 18656 1708 18658 1728
rect 18602 1672 18658 1708
rect 15198 176 15254 232
rect 20166 2388 20168 2408
rect 20168 2388 20220 2408
rect 20220 2388 20222 2408
rect 20166 2352 20222 2388
rect 19798 1400 19854 1456
rect 19982 1808 20038 1864
rect 19890 1264 19946 1320
rect 20810 7248 20866 7304
rect 20534 6296 20590 6352
rect 20534 5480 20590 5536
rect 20350 4256 20406 4312
rect 20718 6840 20774 6896
rect 21362 7520 21418 7576
rect 21362 7112 21418 7168
rect 22190 8084 22246 8120
rect 22190 8064 22192 8084
rect 22192 8064 22244 8084
rect 22244 8064 22246 8084
rect 22650 7520 22706 7576
rect 22374 7112 22430 7168
rect 21362 6840 21418 6896
rect 21362 6568 21418 6624
rect 20718 6296 20774 6352
rect 20810 5480 20866 5536
rect 20626 3984 20682 4040
rect 22006 6568 22062 6624
rect 22006 5636 22062 5672
rect 22006 5616 22008 5636
rect 22008 5616 22060 5636
rect 22060 5616 22062 5636
rect 20956 4396 21252 4692
rect 20350 2896 20406 2952
rect 20258 1536 20314 1592
rect 20258 1128 20314 1184
rect 20534 2488 20590 2544
rect 21616 5056 21912 5352
rect 22098 4256 22154 4312
rect 21362 3712 21418 3768
rect 20718 2644 20774 2680
rect 20718 2624 20720 2644
rect 20720 2624 20772 2644
rect 20772 2624 20774 2644
rect 20534 2216 20590 2272
rect 20350 720 20406 776
rect 20258 584 20314 640
rect 20718 312 20774 368
rect 22190 4120 22246 4176
rect 21362 2080 21418 2136
rect 22006 1944 22062 2000
rect 21362 1420 21418 1456
rect 21362 1400 21364 1420
rect 21364 1400 21416 1420
rect 21416 1400 21418 1420
rect 21362 756 21364 776
rect 21364 756 21416 776
rect 21416 756 21418 776
rect 21362 720 21418 756
rect 22834 6568 22890 6624
rect 23294 6432 23350 6488
rect 23202 6160 23258 6216
rect 22742 5752 22798 5808
rect 23202 5772 23258 5808
rect 23202 5752 23204 5772
rect 23204 5752 23256 5772
rect 23256 5752 23258 5772
rect 22466 3712 22522 3768
rect 22190 1672 22246 1728
rect 22742 992 22798 1048
rect 22098 584 22154 640
rect 24122 7928 24178 7984
rect 23754 7248 23810 7304
rect 27250 11212 27306 11248
rect 27250 11192 27252 11212
rect 27252 11192 27304 11212
rect 27304 11192 27306 11212
rect 26054 10412 26056 10432
rect 26056 10412 26108 10432
rect 26108 10412 26110 10432
rect 26054 10376 26110 10412
rect 25410 7928 25466 7984
rect 25134 7656 25190 7712
rect 27250 11056 27306 11112
rect 26974 9560 27030 9616
rect 27618 10784 27674 10840
rect 27894 10920 27950 10976
rect 30654 9560 30710 9616
rect 27250 8900 27306 8936
rect 27250 8880 27252 8900
rect 27252 8880 27304 8900
rect 27304 8880 27306 8900
rect 27066 7792 27122 7848
rect 26238 7520 26294 7576
rect 24766 6976 24822 7032
rect 23294 2932 23296 2952
rect 23296 2932 23348 2952
rect 23348 2932 23350 2952
rect 23294 2896 23350 2932
rect 25870 6024 25926 6080
rect 25226 5888 25282 5944
rect 23938 3168 23994 3224
rect 24582 3032 24638 3088
rect 23478 1128 23534 1184
rect 24858 1400 24914 1456
rect 27618 7404 27674 7440
rect 27618 7384 27620 7404
rect 27620 7384 27672 7404
rect 27672 7384 27674 7404
rect 28814 8200 28870 8256
rect 29366 8880 29422 8936
rect 26882 6296 26938 6352
rect 29090 6724 29146 6760
rect 29090 6704 29092 6724
rect 29092 6704 29144 6724
rect 29144 6704 29146 6724
rect 27158 5480 27214 5536
rect 28446 4800 28502 4856
rect 26330 3984 26386 4040
rect 31390 9560 31446 9616
rect 30956 8678 31002 8692
rect 31002 8678 31014 8692
rect 31014 8678 31066 8692
rect 31066 8678 31078 8692
rect 31078 8678 31130 8692
rect 31130 8678 31142 8692
rect 31142 8678 31194 8692
rect 31194 8678 31206 8692
rect 31206 8678 31252 8692
rect 30956 8396 31252 8678
rect 30654 6840 30710 6896
rect 31616 9274 31912 9352
rect 31616 9222 31662 9274
rect 31662 9222 31674 9274
rect 31674 9222 31726 9274
rect 31726 9222 31738 9274
rect 31738 9222 31790 9274
rect 31790 9222 31802 9274
rect 31802 9222 31854 9274
rect 31854 9222 31866 9274
rect 31866 9222 31912 9274
rect 31616 9056 31912 9222
rect 31616 5056 31912 5352
rect 30956 4396 31252 4692
rect 26882 3596 26938 3632
rect 26882 3576 26884 3596
rect 26884 3576 26936 3596
rect 26936 3576 26938 3596
rect 27158 3304 27214 3360
rect 28998 2896 29054 2952
rect 27618 2796 27620 2816
rect 27620 2796 27672 2816
rect 27672 2796 27674 2816
rect 27618 2760 27674 2796
rect 24858 876 24914 912
rect 24858 856 24860 876
rect 24860 856 24912 876
rect 24912 856 24914 876
rect 24214 756 24216 776
rect 24216 756 24268 776
rect 24268 756 24270 776
rect 24214 720 24270 756
rect 23294 448 23350 504
rect 17958 40 18014 96
<< metal3 >>
rect 12433 11930 12499 11933
rect 20805 11930 20871 11933
rect 12433 11928 20871 11930
rect 12433 11872 12438 11928
rect 12494 11872 20810 11928
rect 20866 11872 20871 11928
rect 12433 11870 20871 11872
rect 12433 11867 12499 11870
rect 20805 11867 20871 11870
rect 9305 11794 9371 11797
rect 12525 11794 12591 11797
rect 9305 11792 12591 11794
rect 9305 11736 9310 11792
rect 9366 11736 12530 11792
rect 12586 11736 12591 11792
rect 9305 11734 12591 11736
rect 9305 11731 9371 11734
rect 12525 11731 12591 11734
rect 0 11658 800 11688
rect 933 11658 999 11661
rect 0 11656 999 11658
rect 0 11600 938 11656
rect 994 11600 999 11656
rect 0 11598 999 11600
rect 0 11568 800 11598
rect 933 11595 999 11598
rect 3785 11658 3851 11661
rect 12157 11658 12223 11661
rect 3785 11656 12223 11658
rect 3785 11600 3790 11656
rect 3846 11600 12162 11656
rect 12218 11600 12223 11656
rect 3785 11598 12223 11600
rect 3785 11595 3851 11598
rect 12157 11595 12223 11598
rect 17493 11658 17559 11661
rect 21633 11658 21699 11661
rect 17493 11656 21699 11658
rect 17493 11600 17498 11656
rect 17554 11600 21638 11656
rect 21694 11600 21699 11656
rect 17493 11598 21699 11600
rect 17493 11595 17559 11598
rect 21633 11595 21699 11598
rect 3601 11522 3667 11525
rect 20713 11522 20779 11525
rect 3601 11520 20779 11522
rect 3601 11464 3606 11520
rect 3662 11464 20718 11520
rect 20774 11464 20779 11520
rect 3601 11462 20779 11464
rect 3601 11459 3667 11462
rect 20713 11459 20779 11462
rect 4705 11386 4771 11389
rect 12433 11386 12499 11389
rect 4705 11384 12499 11386
rect 4705 11328 4710 11384
rect 4766 11328 12438 11384
rect 12494 11328 12499 11384
rect 4705 11326 12499 11328
rect 4705 11323 4771 11326
rect 12433 11323 12499 11326
rect 21449 11386 21515 11389
rect 25037 11386 25103 11389
rect 21449 11384 25103 11386
rect 21449 11328 21454 11384
rect 21510 11328 25042 11384
rect 25098 11328 25103 11384
rect 21449 11326 25103 11328
rect 21449 11323 21515 11326
rect 25037 11323 25103 11326
rect 0 11250 800 11280
rect 1025 11250 1091 11253
rect 0 11248 1091 11250
rect 0 11192 1030 11248
rect 1086 11192 1091 11248
rect 0 11190 1091 11192
rect 0 11160 800 11190
rect 1025 11187 1091 11190
rect 12341 11250 12407 11253
rect 22001 11250 22067 11253
rect 27245 11250 27311 11253
rect 12341 11248 19350 11250
rect 12341 11192 12346 11248
rect 12402 11192 19350 11248
rect 12341 11190 19350 11192
rect 12341 11187 12407 11190
rect 6637 11114 6703 11117
rect 13169 11114 13235 11117
rect 6637 11112 13235 11114
rect 6637 11056 6642 11112
rect 6698 11056 13174 11112
rect 13230 11056 13235 11112
rect 6637 11054 13235 11056
rect 6637 11051 6703 11054
rect 13169 11051 13235 11054
rect 13353 11114 13419 11117
rect 17769 11114 17835 11117
rect 13353 11112 17835 11114
rect 13353 11056 13358 11112
rect 13414 11056 17774 11112
rect 17830 11056 17835 11112
rect 13353 11054 17835 11056
rect 13353 11051 13419 11054
rect 17769 11051 17835 11054
rect 10593 10978 10659 10981
rect 12893 10978 12959 10981
rect 17953 10978 18019 10981
rect 10593 10976 12818 10978
rect 10593 10920 10598 10976
rect 10654 10920 12818 10976
rect 10593 10918 12818 10920
rect 10593 10915 10659 10918
rect 0 10842 800 10872
rect 4061 10842 4127 10845
rect 0 10840 4127 10842
rect 0 10784 4066 10840
rect 4122 10784 4127 10840
rect 0 10782 4127 10784
rect 0 10752 800 10782
rect 4061 10779 4127 10782
rect 10317 10842 10383 10845
rect 12065 10842 12131 10845
rect 10317 10840 12131 10842
rect 10317 10784 10322 10840
rect 10378 10784 12070 10840
rect 12126 10784 12131 10840
rect 10317 10782 12131 10784
rect 12758 10842 12818 10918
rect 12893 10976 18019 10978
rect 12893 10920 12898 10976
rect 12954 10920 17958 10976
rect 18014 10920 18019 10976
rect 12893 10918 18019 10920
rect 12893 10915 12959 10918
rect 17953 10915 18019 10918
rect 12985 10842 13051 10845
rect 12758 10840 13051 10842
rect 12758 10784 12990 10840
rect 13046 10784 13051 10840
rect 12758 10782 13051 10784
rect 19290 10842 19350 11190
rect 22001 11248 27311 11250
rect 22001 11192 22006 11248
rect 22062 11192 27250 11248
rect 27306 11192 27311 11248
rect 22001 11190 27311 11192
rect 22001 11187 22067 11190
rect 27245 11187 27311 11190
rect 20437 11114 20503 11117
rect 27245 11114 27311 11117
rect 20437 11112 27311 11114
rect 20437 11056 20442 11112
rect 20498 11056 27250 11112
rect 27306 11056 27311 11112
rect 20437 11054 27311 11056
rect 20437 11051 20503 11054
rect 27245 11051 27311 11054
rect 20621 10978 20687 10981
rect 27889 10978 27955 10981
rect 20621 10976 27955 10978
rect 20621 10920 20626 10976
rect 20682 10920 27894 10976
rect 27950 10920 27955 10976
rect 20621 10918 27955 10920
rect 20621 10915 20687 10918
rect 27889 10915 27955 10918
rect 27613 10842 27679 10845
rect 19290 10840 27679 10842
rect 19290 10784 27618 10840
rect 27674 10784 27679 10840
rect 19290 10782 27679 10784
rect 10317 10779 10383 10782
rect 12065 10779 12131 10782
rect 12985 10779 13051 10782
rect 27613 10779 27679 10782
rect 4429 10706 4495 10709
rect 16481 10706 16547 10709
rect 4429 10704 16547 10706
rect 4429 10648 4434 10704
rect 4490 10648 16486 10704
rect 16542 10648 16547 10704
rect 4429 10646 16547 10648
rect 4429 10643 4495 10646
rect 16481 10643 16547 10646
rect 17217 10706 17283 10709
rect 19885 10706 19951 10709
rect 17217 10704 19951 10706
rect 17217 10648 17222 10704
rect 17278 10648 19890 10704
rect 19946 10648 19951 10704
rect 17217 10646 19951 10648
rect 17217 10643 17283 10646
rect 19885 10643 19951 10646
rect 20805 10706 20871 10709
rect 22921 10706 22987 10709
rect 20805 10704 22987 10706
rect 20805 10648 20810 10704
rect 20866 10648 22926 10704
rect 22982 10648 22987 10704
rect 20805 10646 22987 10648
rect 20805 10643 20871 10646
rect 22921 10643 22987 10646
rect 7649 10570 7715 10573
rect 9765 10570 9831 10573
rect 7649 10568 9831 10570
rect 7649 10512 7654 10568
rect 7710 10512 9770 10568
rect 9826 10512 9831 10568
rect 7649 10510 9831 10512
rect 7649 10507 7715 10510
rect 9765 10507 9831 10510
rect 10685 10570 10751 10573
rect 11329 10570 11395 10573
rect 10685 10568 11395 10570
rect 10685 10512 10690 10568
rect 10746 10512 11334 10568
rect 11390 10512 11395 10568
rect 10685 10510 11395 10512
rect 10685 10507 10751 10510
rect 11329 10507 11395 10510
rect 16297 10570 16363 10573
rect 17585 10570 17651 10573
rect 16297 10568 17651 10570
rect 16297 10512 16302 10568
rect 16358 10512 17590 10568
rect 17646 10512 17651 10568
rect 16297 10510 17651 10512
rect 16297 10507 16363 10510
rect 17585 10507 17651 10510
rect 0 10434 800 10464
rect 3969 10434 4035 10437
rect 0 10432 4035 10434
rect 0 10376 3974 10432
rect 4030 10376 4035 10432
rect 0 10374 4035 10376
rect 0 10344 800 10374
rect 3969 10371 4035 10374
rect 10777 10434 10843 10437
rect 11973 10434 12039 10437
rect 12433 10434 12499 10437
rect 10777 10432 12039 10434
rect 10777 10376 10782 10432
rect 10838 10376 11978 10432
rect 12034 10376 12039 10432
rect 10777 10374 12039 10376
rect 10777 10371 10843 10374
rect 11973 10371 12039 10374
rect 12206 10432 12499 10434
rect 12206 10376 12438 10432
rect 12494 10376 12499 10432
rect 12206 10374 12499 10376
rect 9397 10298 9463 10301
rect 12206 10298 12266 10374
rect 12433 10371 12499 10374
rect 15837 10434 15903 10437
rect 17861 10434 17927 10437
rect 15837 10432 17927 10434
rect 15837 10376 15842 10432
rect 15898 10376 17866 10432
rect 17922 10376 17927 10432
rect 15837 10374 17927 10376
rect 15837 10371 15903 10374
rect 17861 10371 17927 10374
rect 22001 10434 22067 10437
rect 26049 10434 26115 10437
rect 22001 10432 26115 10434
rect 22001 10376 22006 10432
rect 22062 10376 26054 10432
rect 26110 10376 26115 10432
rect 22001 10374 26115 10376
rect 22001 10371 22067 10374
rect 26049 10371 26115 10374
rect 9397 10296 12266 10298
rect 9397 10240 9402 10296
rect 9458 10240 12266 10296
rect 9397 10238 12266 10240
rect 12341 10298 12407 10301
rect 17401 10298 17467 10301
rect 12341 10296 17467 10298
rect 12341 10240 12346 10296
rect 12402 10240 17406 10296
rect 17462 10240 17467 10296
rect 12341 10238 17467 10240
rect 9397 10235 9463 10238
rect 12341 10235 12407 10238
rect 17401 10235 17467 10238
rect 18965 10298 19031 10301
rect 22001 10298 22067 10301
rect 18965 10296 22067 10298
rect 18965 10240 18970 10296
rect 19026 10240 22006 10296
rect 22062 10240 22067 10296
rect 18965 10238 22067 10240
rect 18965 10235 19031 10238
rect 22001 10235 22067 10238
rect 2221 10162 2287 10165
rect 3509 10162 3575 10165
rect 2221 10160 3575 10162
rect 2221 10104 2226 10160
rect 2282 10104 3514 10160
rect 3570 10104 3575 10160
rect 2221 10102 3575 10104
rect 2221 10099 2287 10102
rect 3509 10099 3575 10102
rect 10777 10162 10843 10165
rect 18045 10162 18111 10165
rect 10777 10160 18111 10162
rect 10777 10104 10782 10160
rect 10838 10104 18050 10160
rect 18106 10104 18111 10160
rect 10777 10102 18111 10104
rect 10777 10099 10843 10102
rect 18045 10099 18111 10102
rect 20253 10162 20319 10165
rect 22093 10162 22159 10165
rect 23657 10162 23723 10165
rect 20253 10160 22159 10162
rect 20253 10104 20258 10160
rect 20314 10104 22098 10160
rect 22154 10104 22159 10160
rect 20253 10102 22159 10104
rect 20253 10099 20319 10102
rect 22093 10099 22159 10102
rect 23062 10160 23723 10162
rect 23062 10104 23662 10160
rect 23718 10104 23723 10160
rect 23062 10102 23723 10104
rect 0 10026 800 10056
rect 3877 10026 3943 10029
rect 0 10024 3943 10026
rect 0 9968 3882 10024
rect 3938 9968 3943 10024
rect 0 9966 3943 9968
rect 0 9936 800 9966
rect 3877 9963 3943 9966
rect 8201 10026 8267 10029
rect 18045 10026 18111 10029
rect 8201 10024 18111 10026
rect 8201 9968 8206 10024
rect 8262 9968 18050 10024
rect 18106 9968 18111 10024
rect 8201 9966 18111 9968
rect 8201 9963 8267 9966
rect 18045 9963 18111 9966
rect 19793 10026 19859 10029
rect 22093 10026 22159 10029
rect 19793 10024 22159 10026
rect 19793 9968 19798 10024
rect 19854 9968 22098 10024
rect 22154 9968 22159 10024
rect 19793 9966 22159 9968
rect 19793 9963 19859 9966
rect 22093 9963 22159 9966
rect 2221 9890 2287 9893
rect 23062 9890 23122 10102
rect 23657 10099 23723 10102
rect 2221 9888 23122 9890
rect 2221 9832 2226 9888
rect 2282 9832 23122 9888
rect 2221 9830 23122 9832
rect 2221 9827 2287 9830
rect 933 9754 999 9757
rect 2773 9754 2839 9757
rect 933 9752 2839 9754
rect 933 9696 938 9752
rect 994 9696 2778 9752
rect 2834 9696 2839 9752
rect 933 9694 2839 9696
rect 933 9691 999 9694
rect 2773 9691 2839 9694
rect 4245 9754 4311 9757
rect 11973 9754 12039 9757
rect 12341 9754 12407 9757
rect 4245 9752 12407 9754
rect 4245 9696 4250 9752
rect 4306 9696 11978 9752
rect 12034 9696 12346 9752
rect 12402 9696 12407 9752
rect 4245 9694 12407 9696
rect 4245 9691 4311 9694
rect 11973 9691 12039 9694
rect 12341 9691 12407 9694
rect 12617 9754 12683 9757
rect 15193 9754 15259 9757
rect 12617 9752 15259 9754
rect 12617 9696 12622 9752
rect 12678 9696 15198 9752
rect 15254 9696 15259 9752
rect 12617 9694 15259 9696
rect 12617 9691 12683 9694
rect 15193 9691 15259 9694
rect 16849 9754 16915 9757
rect 19333 9754 19399 9757
rect 16849 9752 19399 9754
rect 16849 9696 16854 9752
rect 16910 9696 19338 9752
rect 19394 9696 19399 9752
rect 16849 9694 19399 9696
rect 16849 9691 16915 9694
rect 19333 9691 19399 9694
rect 21449 9754 21515 9757
rect 23473 9754 23539 9757
rect 21449 9752 23539 9754
rect 21449 9696 21454 9752
rect 21510 9696 23478 9752
rect 23534 9696 23539 9752
rect 21449 9694 23539 9696
rect 21449 9691 21515 9694
rect 23473 9691 23539 9694
rect 0 9618 800 9648
rect 26969 9618 27035 9621
rect 0 9616 27035 9618
rect 0 9560 26974 9616
rect 27030 9560 27035 9616
rect 0 9558 27035 9560
rect 0 9528 800 9558
rect 26969 9555 27035 9558
rect 30649 9618 30715 9621
rect 31385 9618 31451 9621
rect 30649 9616 31451 9618
rect 30649 9560 30654 9616
rect 30710 9560 31390 9616
rect 31446 9560 31451 9616
rect 30649 9558 31451 9560
rect 30649 9555 30715 9558
rect 31385 9555 31451 9558
rect 1056 9352 33076 9364
rect 0 9210 800 9240
rect 0 9120 858 9210
rect 798 8972 858 9120
rect 1056 9056 11616 9352
rect 11912 9056 21616 9352
rect 21912 9056 31616 9352
rect 31912 9056 33076 9352
rect 1056 9044 33076 9056
rect 798 8938 1042 8972
rect 3509 8938 3575 8941
rect 798 8936 3575 8938
rect 798 8912 3514 8936
rect 982 8880 3514 8912
rect 3570 8880 3575 8936
rect 982 8878 3575 8880
rect 3509 8875 3575 8878
rect 3693 8938 3759 8941
rect 16849 8938 16915 8941
rect 3693 8936 16915 8938
rect 3693 8880 3698 8936
rect 3754 8880 16854 8936
rect 16910 8880 16915 8936
rect 3693 8878 16915 8880
rect 3693 8875 3759 8878
rect 16849 8875 16915 8878
rect 17033 8938 17099 8941
rect 27245 8938 27311 8941
rect 17033 8936 27311 8938
rect 17033 8880 17038 8936
rect 17094 8880 27250 8936
rect 27306 8880 27311 8936
rect 17033 8878 27311 8880
rect 17033 8875 17099 8878
rect 27245 8875 27311 8878
rect 29361 8938 29427 8941
rect 33400 8938 34200 8968
rect 29361 8936 34200 8938
rect 29361 8880 29366 8936
rect 29422 8880 34200 8936
rect 29361 8878 34200 8880
rect 29361 8875 29427 8878
rect 33400 8848 34200 8878
rect 0 8802 800 8832
rect 933 8802 999 8805
rect 0 8800 999 8802
rect 0 8744 938 8800
rect 994 8744 999 8800
rect 0 8742 999 8744
rect 0 8712 800 8742
rect 933 8739 999 8742
rect 1056 8692 33076 8704
rect 0 8394 800 8424
rect 1056 8396 10956 8692
rect 11252 8396 20956 8692
rect 21252 8396 30956 8692
rect 31252 8396 33076 8692
rect 0 8304 858 8394
rect 1056 8384 33076 8396
rect 798 8258 858 8304
rect 2865 8258 2931 8261
rect 798 8256 2931 8258
rect 798 8200 2870 8256
rect 2926 8200 2931 8256
rect 798 8198 2931 8200
rect 2865 8195 2931 8198
rect 5165 8258 5231 8261
rect 9857 8258 9923 8261
rect 5165 8256 9923 8258
rect 5165 8200 5170 8256
rect 5226 8200 9862 8256
rect 9918 8200 9923 8256
rect 5165 8198 9923 8200
rect 5165 8195 5231 8198
rect 9857 8195 9923 8198
rect 10041 8258 10107 8261
rect 11973 8258 12039 8261
rect 10041 8256 12039 8258
rect 10041 8200 10046 8256
rect 10102 8200 11978 8256
rect 12034 8200 12039 8256
rect 10041 8198 12039 8200
rect 10041 8195 10107 8198
rect 11973 8195 12039 8198
rect 12433 8258 12499 8261
rect 18689 8258 18755 8261
rect 28809 8258 28875 8261
rect 12433 8256 18522 8258
rect 12433 8200 12438 8256
rect 12494 8200 18522 8256
rect 12433 8198 18522 8200
rect 12433 8195 12499 8198
rect 2589 8122 2655 8125
rect 11421 8122 11487 8125
rect 2589 8120 11487 8122
rect 2589 8064 2594 8120
rect 2650 8064 11426 8120
rect 11482 8064 11487 8120
rect 12433 8122 12499 8125
rect 17861 8122 17927 8125
rect 12433 8120 17927 8122
rect 2589 8062 11487 8064
rect 2589 8059 2655 8062
rect 11421 8059 11487 8062
rect 11654 8028 12220 8088
rect 12433 8064 12438 8120
rect 12494 8064 17866 8120
rect 17922 8064 17927 8120
rect 12433 8062 17927 8064
rect 18462 8122 18522 8198
rect 18689 8256 28875 8258
rect 18689 8200 18694 8256
rect 18750 8200 28814 8256
rect 28870 8200 28875 8256
rect 18689 8198 28875 8200
rect 18689 8195 18755 8198
rect 28809 8195 28875 8198
rect 19609 8122 19675 8125
rect 18462 8120 19675 8122
rect 18462 8064 19614 8120
rect 19670 8064 19675 8120
rect 18462 8062 19675 8064
rect 12433 8059 12499 8062
rect 17861 8059 17927 8062
rect 19609 8059 19675 8062
rect 19885 8122 19951 8125
rect 22185 8122 22251 8125
rect 19885 8120 22251 8122
rect 19885 8064 19890 8120
rect 19946 8064 22190 8120
rect 22246 8064 22251 8120
rect 19885 8062 22251 8064
rect 19885 8059 19951 8062
rect 22185 8059 22251 8062
rect 0 7986 800 8016
rect 3877 7986 3943 7989
rect 11654 7986 11714 8028
rect 0 7926 2790 7986
rect 0 7896 800 7926
rect 2730 7714 2790 7926
rect 3877 7984 11714 7986
rect 3877 7928 3882 7984
rect 3938 7928 11714 7984
rect 3877 7926 11714 7928
rect 12160 7986 12220 8028
rect 15837 7986 15903 7989
rect 12160 7984 15903 7986
rect 12160 7928 15842 7984
rect 15898 7928 15903 7984
rect 12160 7926 15903 7928
rect 3877 7923 3943 7926
rect 15837 7923 15903 7926
rect 16573 7986 16639 7989
rect 24117 7986 24183 7989
rect 25405 7986 25471 7989
rect 16573 7984 25471 7986
rect 16573 7928 16578 7984
rect 16634 7928 24122 7984
rect 24178 7928 25410 7984
rect 25466 7928 25471 7984
rect 16573 7926 25471 7928
rect 16573 7923 16639 7926
rect 24117 7923 24183 7926
rect 25405 7923 25471 7926
rect 4061 7850 4127 7853
rect 6545 7850 6611 7853
rect 4061 7848 6611 7850
rect 4061 7792 4066 7848
rect 4122 7792 6550 7848
rect 6606 7792 6611 7848
rect 4061 7790 6611 7792
rect 4061 7787 4127 7790
rect 6545 7787 6611 7790
rect 8477 7850 8543 7853
rect 12433 7850 12499 7853
rect 8477 7848 11530 7850
rect 8477 7792 8482 7848
rect 8538 7792 11530 7848
rect 12206 7848 12499 7850
rect 12206 7816 12438 7848
rect 8477 7790 11530 7792
rect 8477 7787 8543 7790
rect 6269 7714 6335 7717
rect 2730 7712 6335 7714
rect 2730 7656 6274 7712
rect 6330 7656 6335 7712
rect 2730 7654 6335 7656
rect 6269 7651 6335 7654
rect 6545 7714 6611 7717
rect 11329 7714 11395 7717
rect 6545 7712 11395 7714
rect 6545 7656 6550 7712
rect 6606 7656 11334 7712
rect 11390 7656 11395 7712
rect 6545 7654 11395 7656
rect 11470 7714 11530 7790
rect 11838 7792 12438 7816
rect 12494 7792 12499 7848
rect 11838 7790 12499 7792
rect 11838 7756 12266 7790
rect 12433 7787 12499 7790
rect 12801 7850 12867 7853
rect 14825 7850 14891 7853
rect 12801 7848 14891 7850
rect 12801 7792 12806 7848
rect 12862 7792 14830 7848
rect 14886 7792 14891 7848
rect 12801 7790 14891 7792
rect 12801 7787 12867 7790
rect 14825 7787 14891 7790
rect 15561 7850 15627 7853
rect 19977 7850 20043 7853
rect 15561 7848 20043 7850
rect 15561 7792 15566 7848
rect 15622 7792 19982 7848
rect 20038 7792 20043 7848
rect 15561 7790 20043 7792
rect 15561 7787 15627 7790
rect 19977 7787 20043 7790
rect 20253 7850 20319 7853
rect 27061 7850 27127 7853
rect 20253 7848 27127 7850
rect 20253 7792 20258 7848
rect 20314 7792 27066 7848
rect 27122 7792 27127 7848
rect 20253 7790 27127 7792
rect 20253 7787 20319 7790
rect 27061 7787 27127 7790
rect 11838 7714 11898 7756
rect 11470 7654 11898 7714
rect 13629 7714 13695 7717
rect 20069 7714 20135 7717
rect 25129 7714 25195 7717
rect 13629 7712 18890 7714
rect 13629 7656 13634 7712
rect 13690 7656 18890 7712
rect 13629 7654 18890 7656
rect 6545 7651 6611 7654
rect 11329 7651 11395 7654
rect 13629 7651 13695 7654
rect 0 7578 800 7608
rect 3601 7578 3667 7581
rect 0 7576 3667 7578
rect 0 7520 3606 7576
rect 3662 7520 3667 7576
rect 0 7518 3667 7520
rect 0 7488 800 7518
rect 3601 7515 3667 7518
rect 3877 7578 3943 7581
rect 9489 7578 9555 7581
rect 14641 7578 14707 7581
rect 3877 7576 9555 7578
rect 3877 7520 3882 7576
rect 3938 7520 9494 7576
rect 9550 7520 9555 7576
rect 3877 7518 9555 7520
rect 3877 7515 3943 7518
rect 9489 7515 9555 7518
rect 9630 7576 14707 7578
rect 9630 7520 14646 7576
rect 14702 7520 14707 7576
rect 9630 7518 14707 7520
rect 2681 7442 2747 7445
rect 9489 7442 9555 7445
rect 2681 7440 9555 7442
rect 2681 7384 2686 7440
rect 2742 7384 9494 7440
rect 9550 7384 9555 7440
rect 2681 7382 9555 7384
rect 2681 7379 2747 7382
rect 9489 7379 9555 7382
rect 5073 7306 5139 7309
rect 6361 7306 6427 7309
rect 5073 7304 6427 7306
rect 5073 7248 5078 7304
rect 5134 7248 6366 7304
rect 6422 7248 6427 7304
rect 5073 7246 6427 7248
rect 5073 7243 5139 7246
rect 6361 7243 6427 7246
rect 0 7170 800 7200
rect 9630 7170 9690 7518
rect 14641 7515 14707 7518
rect 14825 7578 14891 7581
rect 18830 7578 18890 7654
rect 20069 7712 21650 7714
rect 20069 7656 20074 7712
rect 20130 7656 21650 7712
rect 20069 7654 21650 7656
rect 20069 7651 20135 7654
rect 21357 7578 21423 7581
rect 14825 7576 18706 7578
rect 14825 7520 14830 7576
rect 14886 7520 18706 7576
rect 14825 7518 18706 7520
rect 18830 7576 21423 7578
rect 18830 7520 21362 7576
rect 21418 7520 21423 7576
rect 18830 7518 21423 7520
rect 21590 7578 21650 7654
rect 22004 7712 25195 7714
rect 22004 7656 25134 7712
rect 25190 7656 25195 7712
rect 22004 7654 25195 7656
rect 22004 7578 22064 7654
rect 25129 7651 25195 7654
rect 21590 7518 22064 7578
rect 22645 7578 22711 7581
rect 26233 7578 26299 7581
rect 22645 7576 26299 7578
rect 22645 7520 22650 7576
rect 22706 7520 26238 7576
rect 26294 7520 26299 7576
rect 22645 7518 26299 7520
rect 14825 7515 14891 7518
rect 9857 7442 9923 7445
rect 18505 7442 18571 7445
rect 9857 7440 11898 7442
rect 9857 7384 9862 7440
rect 9918 7384 11898 7440
rect 9857 7382 11898 7384
rect 9857 7379 9923 7382
rect 11838 7340 11898 7382
rect 12022 7440 18571 7442
rect 12022 7384 18510 7440
rect 18566 7384 18571 7440
rect 12022 7382 18571 7384
rect 18646 7442 18706 7518
rect 21357 7515 21423 7518
rect 22645 7515 22711 7518
rect 26233 7515 26299 7518
rect 27613 7442 27679 7445
rect 18646 7440 27679 7442
rect 18646 7384 27618 7440
rect 27674 7384 27679 7440
rect 18646 7382 27679 7384
rect 12022 7340 12082 7382
rect 18505 7379 18571 7382
rect 27613 7379 27679 7382
rect 9765 7306 9831 7309
rect 9765 7304 11714 7306
rect 9765 7248 9770 7304
rect 9826 7248 11714 7304
rect 11838 7280 12082 7340
rect 12709 7306 12775 7309
rect 20805 7306 20871 7309
rect 23749 7306 23815 7309
rect 12709 7304 20871 7306
rect 9765 7246 11714 7248
rect 9765 7243 9831 7246
rect 0 7110 9690 7170
rect 9949 7170 10015 7173
rect 11654 7170 11714 7246
rect 12709 7248 12714 7304
rect 12770 7248 20810 7304
rect 20866 7248 20871 7304
rect 12709 7246 20871 7248
rect 12709 7243 12775 7246
rect 20805 7243 20871 7246
rect 21038 7304 23815 7306
rect 21038 7248 23754 7304
rect 23810 7248 23815 7304
rect 21038 7246 23815 7248
rect 12801 7170 12867 7173
rect 9949 7168 11530 7170
rect 9949 7112 9954 7168
rect 10010 7112 11530 7168
rect 9949 7110 11530 7112
rect 11654 7168 12867 7170
rect 11654 7112 12806 7168
rect 12862 7112 12867 7168
rect 11654 7110 12867 7112
rect 0 7080 800 7110
rect 9949 7107 10015 7110
rect 3969 7034 4035 7037
rect 11329 7034 11395 7037
rect 3969 7032 11395 7034
rect 3969 6976 3974 7032
rect 4030 6976 11334 7032
rect 11390 6976 11395 7032
rect 3969 6974 11395 6976
rect 3969 6971 4035 6974
rect 11329 6971 11395 6974
rect 3877 6898 3943 6901
rect 1948 6896 3943 6898
rect 1948 6840 3882 6896
rect 3938 6840 3943 6896
rect 1948 6838 3943 6840
rect 0 6762 800 6792
rect 1948 6762 2008 6838
rect 3877 6835 3943 6838
rect 4797 6898 4863 6901
rect 6085 6898 6151 6901
rect 4797 6896 6151 6898
rect 4797 6840 4802 6896
rect 4858 6840 6090 6896
rect 6146 6840 6151 6896
rect 4797 6838 6151 6840
rect 4797 6835 4863 6838
rect 6085 6835 6151 6838
rect 6269 6898 6335 6901
rect 9949 6898 10015 6901
rect 6269 6896 10015 6898
rect 6269 6840 6274 6896
rect 6330 6840 9954 6896
rect 10010 6840 10015 6896
rect 6269 6838 10015 6840
rect 6269 6835 6335 6838
rect 9949 6835 10015 6838
rect 10133 6898 10199 6901
rect 11329 6898 11395 6901
rect 10133 6896 11395 6898
rect 10133 6840 10138 6896
rect 10194 6840 11334 6896
rect 11390 6840 11395 6896
rect 10133 6838 11395 6840
rect 11470 6898 11530 7110
rect 12801 7107 12867 7110
rect 13169 7170 13235 7173
rect 18597 7170 18663 7173
rect 19241 7170 19307 7173
rect 13169 7168 19307 7170
rect 13169 7112 13174 7168
rect 13230 7112 18602 7168
rect 18658 7112 19246 7168
rect 19302 7112 19307 7168
rect 13169 7110 19307 7112
rect 13169 7107 13235 7110
rect 18597 7107 18663 7110
rect 19241 7107 19307 7110
rect 19425 7170 19491 7173
rect 21038 7170 21098 7246
rect 23749 7243 23815 7246
rect 19425 7168 21098 7170
rect 19425 7112 19430 7168
rect 19486 7112 21098 7168
rect 19425 7110 21098 7112
rect 21357 7170 21423 7173
rect 22369 7170 22435 7173
rect 21357 7168 22435 7170
rect 21357 7112 21362 7168
rect 21418 7112 22374 7168
rect 22430 7112 22435 7168
rect 21357 7110 22435 7112
rect 19425 7107 19491 7110
rect 21357 7107 21423 7110
rect 22369 7107 22435 7110
rect 12157 7034 12223 7037
rect 24761 7034 24827 7037
rect 12157 7032 24827 7034
rect 12157 6976 12162 7032
rect 12218 6976 24766 7032
rect 24822 6976 24827 7032
rect 12157 6974 24827 6976
rect 12157 6971 12223 6974
rect 24761 6971 24827 6974
rect 17217 6898 17283 6901
rect 11470 6896 17283 6898
rect 11470 6840 17222 6896
rect 17278 6840 17283 6896
rect 11470 6838 17283 6840
rect 10133 6835 10199 6838
rect 11329 6835 11395 6838
rect 17217 6835 17283 6838
rect 17401 6898 17467 6901
rect 20713 6898 20779 6901
rect 17401 6896 20779 6898
rect 17401 6840 17406 6896
rect 17462 6840 20718 6896
rect 20774 6840 20779 6896
rect 17401 6838 20779 6840
rect 17401 6835 17467 6838
rect 20713 6835 20779 6838
rect 21357 6898 21423 6901
rect 30649 6898 30715 6901
rect 21357 6896 30715 6898
rect 21357 6840 21362 6896
rect 21418 6840 30654 6896
rect 30710 6840 30715 6896
rect 21357 6838 30715 6840
rect 21357 6835 21423 6838
rect 30649 6835 30715 6838
rect 0 6702 2008 6762
rect 4429 6762 4495 6765
rect 8845 6762 8911 6765
rect 12525 6762 12591 6765
rect 29085 6762 29151 6765
rect 4429 6760 8911 6762
rect 4429 6704 4434 6760
rect 4490 6704 8850 6760
rect 8906 6704 8911 6760
rect 4429 6702 8911 6704
rect 0 6672 800 6702
rect 4429 6699 4495 6702
rect 8845 6699 8911 6702
rect 9446 6702 12450 6762
rect 4337 6626 4403 6629
rect 9446 6626 9506 6702
rect 4337 6624 9506 6626
rect 4337 6568 4342 6624
rect 4398 6568 9506 6624
rect 4337 6566 9506 6568
rect 9581 6626 9647 6629
rect 12249 6626 12315 6629
rect 9581 6624 12315 6626
rect 9581 6568 9586 6624
rect 9642 6568 12254 6624
rect 12310 6568 12315 6624
rect 9581 6566 12315 6568
rect 12390 6626 12450 6702
rect 12525 6760 29151 6762
rect 12525 6704 12530 6760
rect 12586 6704 29090 6760
rect 29146 6704 29151 6760
rect 12525 6702 29151 6704
rect 12525 6699 12591 6702
rect 29085 6699 29151 6702
rect 12709 6626 12775 6629
rect 12390 6624 12775 6626
rect 12390 6568 12714 6624
rect 12770 6568 12775 6624
rect 12390 6566 12775 6568
rect 4337 6563 4403 6566
rect 9581 6563 9647 6566
rect 12249 6563 12315 6566
rect 12709 6563 12775 6566
rect 13077 6626 13143 6629
rect 16573 6626 16639 6629
rect 13077 6624 16639 6626
rect 13077 6568 13082 6624
rect 13138 6568 16578 6624
rect 16634 6568 16639 6624
rect 13077 6566 16639 6568
rect 13077 6563 13143 6566
rect 16573 6563 16639 6566
rect 17033 6626 17099 6629
rect 17953 6626 18019 6629
rect 19241 6626 19307 6629
rect 17033 6624 19307 6626
rect 17033 6568 17038 6624
rect 17094 6568 17958 6624
rect 18014 6568 19246 6624
rect 19302 6568 19307 6624
rect 17033 6566 19307 6568
rect 17033 6563 17099 6566
rect 17953 6563 18019 6566
rect 19241 6563 19307 6566
rect 19425 6626 19491 6629
rect 21357 6626 21423 6629
rect 19425 6624 21423 6626
rect 19425 6568 19430 6624
rect 19486 6568 21362 6624
rect 21418 6568 21423 6624
rect 19425 6566 21423 6568
rect 19425 6563 19491 6566
rect 21357 6563 21423 6566
rect 22001 6626 22067 6629
rect 22829 6626 22895 6629
rect 22001 6624 22895 6626
rect 22001 6568 22006 6624
rect 22062 6568 22834 6624
rect 22890 6568 22895 6624
rect 22001 6566 22895 6568
rect 22001 6563 22067 6566
rect 22829 6563 22895 6566
rect 3877 6490 3943 6493
rect 6637 6490 6703 6493
rect 3877 6488 6703 6490
rect 3877 6432 3882 6488
rect 3938 6432 6642 6488
rect 6698 6432 6703 6488
rect 3877 6430 6703 6432
rect 3877 6427 3943 6430
rect 6637 6427 6703 6430
rect 6821 6490 6887 6493
rect 12249 6490 12315 6493
rect 6821 6488 12315 6490
rect 6821 6432 6826 6488
rect 6882 6432 12254 6488
rect 12310 6432 12315 6488
rect 6821 6430 12315 6432
rect 6821 6427 6887 6430
rect 12249 6427 12315 6430
rect 12893 6490 12959 6493
rect 17861 6490 17927 6493
rect 23289 6490 23355 6493
rect 12893 6488 17418 6490
rect 12893 6432 12898 6488
rect 12954 6432 17418 6488
rect 12893 6430 17418 6432
rect 12893 6427 12959 6430
rect 0 6354 800 6384
rect 0 6294 17234 6354
rect 0 6264 800 6294
rect 4245 6218 4311 6221
rect 12525 6218 12591 6221
rect 4245 6216 12591 6218
rect 4245 6160 4250 6216
rect 4306 6160 12530 6216
rect 12586 6160 12591 6216
rect 4245 6158 12591 6160
rect 4245 6155 4311 6158
rect 12525 6155 12591 6158
rect 12709 6218 12775 6221
rect 17033 6218 17099 6221
rect 12709 6216 17099 6218
rect 12709 6160 12714 6216
rect 12770 6160 17038 6216
rect 17094 6160 17099 6216
rect 12709 6158 17099 6160
rect 12709 6155 12775 6158
rect 17033 6155 17099 6158
rect 3417 6082 3483 6085
rect 7005 6082 7071 6085
rect 3417 6080 7071 6082
rect 3417 6024 3422 6080
rect 3478 6024 7010 6080
rect 7066 6024 7071 6080
rect 3417 6022 7071 6024
rect 3417 6019 3483 6022
rect 7005 6019 7071 6022
rect 7189 6082 7255 6085
rect 12525 6082 12591 6085
rect 15653 6082 15719 6085
rect 7189 6080 12450 6082
rect 7189 6024 7194 6080
rect 7250 6024 12450 6080
rect 7189 6022 12450 6024
rect 7189 6019 7255 6022
rect 0 5946 800 5976
rect 2957 5946 3023 5949
rect 0 5944 3023 5946
rect 0 5888 2962 5944
rect 3018 5888 3023 5944
rect 0 5886 3023 5888
rect 0 5856 800 5886
rect 2957 5883 3023 5886
rect 3601 5946 3667 5949
rect 12390 5946 12450 6022
rect 12525 6080 15719 6082
rect 12525 6024 12530 6080
rect 12586 6024 15658 6080
rect 15714 6024 15719 6080
rect 12525 6022 15719 6024
rect 17174 6082 17234 6294
rect 17358 6218 17418 6430
rect 17861 6488 23355 6490
rect 17861 6432 17866 6488
rect 17922 6432 23294 6488
rect 23350 6432 23355 6488
rect 17861 6430 23355 6432
rect 17861 6427 17927 6430
rect 23289 6427 23355 6430
rect 17861 6354 17927 6357
rect 20529 6354 20595 6357
rect 17861 6352 20595 6354
rect 17861 6296 17866 6352
rect 17922 6296 20534 6352
rect 20590 6296 20595 6352
rect 17861 6294 20595 6296
rect 17861 6291 17927 6294
rect 20529 6291 20595 6294
rect 20713 6354 20779 6357
rect 26877 6354 26943 6357
rect 20713 6352 26943 6354
rect 20713 6296 20718 6352
rect 20774 6296 26882 6352
rect 26938 6296 26943 6352
rect 20713 6294 26943 6296
rect 20713 6291 20779 6294
rect 26877 6291 26943 6294
rect 23197 6218 23263 6221
rect 17358 6216 23263 6218
rect 17358 6160 23202 6216
rect 23258 6160 23263 6216
rect 17358 6158 23263 6160
rect 23197 6155 23263 6158
rect 25865 6082 25931 6085
rect 17174 6080 25931 6082
rect 17174 6024 25870 6080
rect 25926 6024 25931 6080
rect 17174 6022 25931 6024
rect 12525 6019 12591 6022
rect 15653 6019 15719 6022
rect 25865 6019 25931 6022
rect 15285 5946 15351 5949
rect 3601 5944 12266 5946
rect 3601 5888 3606 5944
rect 3662 5888 12266 5944
rect 3601 5886 12266 5888
rect 12390 5944 15351 5946
rect 12390 5888 15290 5944
rect 15346 5888 15351 5944
rect 12390 5886 15351 5888
rect 3601 5883 3667 5886
rect 4797 5810 4863 5813
rect 6085 5810 6151 5813
rect 4797 5808 6151 5810
rect 4797 5752 4802 5808
rect 4858 5752 6090 5808
rect 6146 5752 6151 5808
rect 4797 5750 6151 5752
rect 4797 5747 4863 5750
rect 6085 5747 6151 5750
rect 7005 5810 7071 5813
rect 10225 5810 10291 5813
rect 7005 5808 10291 5810
rect 7005 5752 7010 5808
rect 7066 5752 10230 5808
rect 10286 5752 10291 5808
rect 7005 5750 10291 5752
rect 7005 5747 7071 5750
rect 10225 5747 10291 5750
rect 10501 5810 10567 5813
rect 12065 5810 12131 5813
rect 10501 5808 12131 5810
rect 10501 5752 10506 5808
rect 10562 5752 12070 5808
rect 12126 5752 12131 5808
rect 10501 5750 12131 5752
rect 12206 5810 12266 5886
rect 15285 5883 15351 5886
rect 17217 5946 17283 5949
rect 25221 5946 25287 5949
rect 17217 5944 25287 5946
rect 17217 5888 17222 5944
rect 17278 5888 25226 5944
rect 25282 5888 25287 5944
rect 17217 5886 25287 5888
rect 17217 5883 17283 5886
rect 25221 5883 25287 5886
rect 19609 5810 19675 5813
rect 12206 5808 19675 5810
rect 12206 5752 19614 5808
rect 19670 5752 19675 5808
rect 12206 5750 19675 5752
rect 10501 5747 10567 5750
rect 12065 5747 12131 5750
rect 19609 5747 19675 5750
rect 19885 5810 19951 5813
rect 22737 5810 22803 5813
rect 23197 5810 23263 5813
rect 19885 5808 23263 5810
rect 19885 5752 19890 5808
rect 19946 5752 22742 5808
rect 22798 5752 23202 5808
rect 23258 5752 23263 5808
rect 19885 5750 23263 5752
rect 19885 5747 19951 5750
rect 22737 5747 22803 5750
rect 23197 5747 23263 5750
rect 2405 5674 2471 5677
rect 5257 5674 5323 5677
rect 2405 5672 5323 5674
rect 2405 5616 2410 5672
rect 2466 5616 5262 5672
rect 5318 5616 5323 5672
rect 2405 5614 5323 5616
rect 2405 5611 2471 5614
rect 5257 5611 5323 5614
rect 5441 5674 5507 5677
rect 12985 5674 13051 5677
rect 18689 5674 18755 5677
rect 5441 5672 9874 5674
rect 5441 5616 5446 5672
rect 5502 5616 9874 5672
rect 5441 5614 9874 5616
rect 5441 5611 5507 5614
rect 0 5538 800 5568
rect 3141 5538 3207 5541
rect 0 5536 3207 5538
rect 0 5480 3146 5536
rect 3202 5480 3207 5536
rect 0 5478 3207 5480
rect 0 5448 800 5478
rect 3141 5475 3207 5478
rect 3325 5538 3391 5541
rect 9581 5538 9647 5541
rect 3325 5536 9647 5538
rect 3325 5480 3330 5536
rect 3386 5480 9586 5536
rect 9642 5480 9647 5536
rect 3325 5478 9647 5480
rect 9814 5538 9874 5614
rect 12985 5672 18755 5674
rect 12985 5616 12990 5672
rect 13046 5616 18694 5672
rect 18750 5616 18755 5672
rect 12985 5614 18755 5616
rect 12985 5611 13051 5614
rect 18689 5611 18755 5614
rect 19517 5674 19583 5677
rect 22001 5674 22067 5677
rect 19517 5672 22067 5674
rect 19517 5616 19522 5672
rect 19578 5616 22006 5672
rect 22062 5616 22067 5672
rect 19517 5614 22067 5616
rect 19517 5611 19583 5614
rect 22001 5611 22067 5614
rect 15193 5538 15259 5541
rect 9814 5536 15259 5538
rect 9814 5480 15198 5536
rect 15254 5480 15259 5536
rect 9814 5478 15259 5480
rect 3325 5475 3391 5478
rect 9581 5475 9647 5478
rect 15193 5475 15259 5478
rect 15377 5538 15443 5541
rect 20069 5538 20135 5541
rect 15377 5536 20135 5538
rect 15377 5480 15382 5536
rect 15438 5480 20074 5536
rect 20130 5480 20135 5536
rect 15377 5478 20135 5480
rect 15377 5475 15443 5478
rect 20069 5475 20135 5478
rect 20529 5538 20595 5541
rect 20805 5538 20871 5541
rect 27153 5538 27219 5541
rect 20529 5536 27219 5538
rect 20529 5480 20534 5536
rect 20590 5480 20810 5536
rect 20866 5480 27158 5536
rect 27214 5480 27219 5536
rect 20529 5478 27219 5480
rect 20529 5475 20595 5478
rect 20805 5475 20871 5478
rect 27153 5475 27219 5478
rect 1056 5352 33076 5364
rect 0 5130 800 5160
rect 0 5040 858 5130
rect 1056 5056 11616 5352
rect 11912 5056 21616 5352
rect 21912 5056 31616 5352
rect 31912 5056 33076 5352
rect 1056 5044 33076 5056
rect 798 4994 858 5040
rect 933 4994 999 4997
rect 798 4992 999 4994
rect 798 4936 938 4992
rect 994 4936 999 4992
rect 798 4934 999 4936
rect 933 4931 999 4934
rect 3785 4858 3851 4861
rect 798 4856 3851 4858
rect 798 4800 3790 4856
rect 3846 4800 3851 4856
rect 798 4798 3851 4800
rect 798 4752 858 4798
rect 3785 4795 3851 4798
rect 4521 4858 4587 4861
rect 7741 4858 7807 4861
rect 4521 4856 7807 4858
rect 4521 4800 4526 4856
rect 4582 4800 7746 4856
rect 7802 4800 7807 4856
rect 4521 4798 7807 4800
rect 4521 4795 4587 4798
rect 7741 4795 7807 4798
rect 7925 4858 7991 4861
rect 13813 4858 13879 4861
rect 7925 4856 13879 4858
rect 7925 4800 7930 4856
rect 7986 4800 13818 4856
rect 13874 4800 13879 4856
rect 7925 4798 13879 4800
rect 7925 4795 7991 4798
rect 13813 4795 13879 4798
rect 13997 4858 14063 4861
rect 15193 4858 15259 4861
rect 13997 4856 15259 4858
rect 13997 4800 14002 4856
rect 14058 4800 15198 4856
rect 15254 4800 15259 4856
rect 13997 4798 15259 4800
rect 13997 4795 14063 4798
rect 15193 4795 15259 4798
rect 18321 4858 18387 4861
rect 28441 4858 28507 4861
rect 18321 4856 28507 4858
rect 18321 4800 18326 4856
rect 18382 4800 28446 4856
rect 28502 4800 28507 4856
rect 18321 4798 28507 4800
rect 18321 4795 18387 4798
rect 28441 4795 28507 4798
rect 0 4662 858 4752
rect 1056 4692 33076 4704
rect 0 4632 800 4662
rect 1056 4396 10956 4692
rect 11252 4396 20956 4692
rect 21252 4396 30956 4692
rect 31252 4396 33076 4692
rect 1056 4384 33076 4396
rect 0 4314 800 4344
rect 5717 4314 5783 4317
rect 18137 4314 18203 4317
rect 0 4312 5783 4314
rect 0 4256 5722 4312
rect 5778 4256 5783 4312
rect 0 4254 5783 4256
rect 0 4224 800 4254
rect 5717 4251 5783 4254
rect 5950 4312 18203 4314
rect 5950 4256 18142 4312
rect 18198 4256 18203 4312
rect 5950 4254 18203 4256
rect 933 4178 999 4181
rect 3049 4178 3115 4181
rect 933 4176 3115 4178
rect 933 4120 938 4176
rect 994 4120 3054 4176
rect 3110 4120 3115 4176
rect 933 4118 3115 4120
rect 933 4115 999 4118
rect 3049 4115 3115 4118
rect 5533 4178 5599 4181
rect 5950 4178 6010 4254
rect 18137 4251 18203 4254
rect 20345 4314 20411 4317
rect 22093 4314 22159 4317
rect 20345 4312 22159 4314
rect 20345 4256 20350 4312
rect 20406 4256 22098 4312
rect 22154 4256 22159 4312
rect 20345 4254 22159 4256
rect 20345 4251 20411 4254
rect 22093 4251 22159 4254
rect 12065 4178 12131 4181
rect 5533 4176 6010 4178
rect 5533 4120 5538 4176
rect 5594 4120 6010 4176
rect 5533 4118 6010 4120
rect 6548 4176 12131 4178
rect 6548 4120 12070 4176
rect 12126 4120 12131 4176
rect 6548 4118 12131 4120
rect 5533 4115 5599 4118
rect 5625 4042 5691 4045
rect 6548 4042 6608 4118
rect 12065 4115 12131 4118
rect 12249 4178 12315 4181
rect 13629 4178 13695 4181
rect 12249 4176 13695 4178
rect 12249 4120 12254 4176
rect 12310 4120 13634 4176
rect 13690 4120 13695 4176
rect 12249 4118 13695 4120
rect 12249 4115 12315 4118
rect 13629 4115 13695 4118
rect 13813 4178 13879 4181
rect 16573 4178 16639 4181
rect 13813 4176 16639 4178
rect 13813 4120 13818 4176
rect 13874 4120 16578 4176
rect 16634 4120 16639 4176
rect 13813 4118 16639 4120
rect 13813 4115 13879 4118
rect 16573 4115 16639 4118
rect 17309 4178 17375 4181
rect 22185 4178 22251 4181
rect 17309 4176 22251 4178
rect 17309 4120 17314 4176
rect 17370 4120 22190 4176
rect 22246 4120 22251 4176
rect 17309 4118 22251 4120
rect 17309 4115 17375 4118
rect 22185 4115 22251 4118
rect 5625 4040 6608 4042
rect 5625 3984 5630 4040
rect 5686 3984 6608 4040
rect 5625 3982 6608 3984
rect 6913 4042 6979 4045
rect 18505 4042 18571 4045
rect 6913 4040 18571 4042
rect 6913 3984 6918 4040
rect 6974 3984 18510 4040
rect 18566 3984 18571 4040
rect 6913 3982 18571 3984
rect 5625 3979 5691 3982
rect 6913 3979 6979 3982
rect 18505 3979 18571 3982
rect 20621 4042 20687 4045
rect 26325 4042 26391 4045
rect 20621 4040 26391 4042
rect 20621 3984 20626 4040
rect 20682 3984 26330 4040
rect 26386 3984 26391 4040
rect 20621 3982 26391 3984
rect 20621 3979 20687 3982
rect 26325 3979 26391 3982
rect 0 3906 800 3936
rect 4981 3906 5047 3909
rect 12065 3906 12131 3909
rect 15377 3906 15443 3909
rect 0 3846 2790 3906
rect 0 3816 800 3846
rect 2730 3770 2790 3846
rect 4981 3904 12131 3906
rect 4981 3848 4986 3904
rect 5042 3848 12070 3904
rect 12126 3848 12131 3904
rect 4981 3846 12131 3848
rect 4981 3843 5047 3846
rect 12065 3843 12131 3846
rect 12252 3904 15443 3906
rect 12252 3848 15382 3904
rect 15438 3848 15443 3904
rect 12252 3846 15443 3848
rect 7557 3770 7623 3773
rect 2730 3768 7623 3770
rect 2730 3712 7562 3768
rect 7618 3712 7623 3768
rect 2730 3710 7623 3712
rect 7557 3707 7623 3710
rect 7741 3770 7807 3773
rect 12252 3770 12312 3846
rect 15377 3843 15443 3846
rect 7741 3768 12312 3770
rect 7741 3712 7746 3768
rect 7802 3712 12312 3768
rect 7741 3710 12312 3712
rect 14549 3770 14615 3773
rect 16205 3770 16271 3773
rect 14549 3768 16271 3770
rect 14549 3712 14554 3768
rect 14610 3712 16210 3768
rect 16266 3712 16271 3768
rect 14549 3710 16271 3712
rect 7741 3707 7807 3710
rect 14549 3707 14615 3710
rect 16205 3707 16271 3710
rect 16757 3770 16823 3773
rect 21357 3770 21423 3773
rect 22461 3770 22527 3773
rect 16757 3768 22527 3770
rect 16757 3712 16762 3768
rect 16818 3712 21362 3768
rect 21418 3712 22466 3768
rect 22522 3712 22527 3768
rect 16757 3710 22527 3712
rect 16757 3707 16823 3710
rect 21357 3707 21423 3710
rect 22461 3707 22527 3710
rect 4245 3634 4311 3637
rect 5441 3634 5507 3637
rect 4245 3632 5507 3634
rect 4245 3576 4250 3632
rect 4306 3576 5446 3632
rect 5502 3576 5507 3632
rect 4245 3574 5507 3576
rect 4245 3571 4311 3574
rect 5441 3571 5507 3574
rect 5809 3634 5875 3637
rect 13445 3634 13511 3637
rect 26877 3634 26943 3637
rect 5809 3632 12450 3634
rect 5809 3576 5814 3632
rect 5870 3576 12450 3632
rect 5809 3574 12450 3576
rect 5809 3571 5875 3574
rect 0 3498 800 3528
rect 4245 3498 4311 3501
rect 6085 3498 6151 3501
rect 0 3438 4170 3498
rect 0 3408 800 3438
rect 0 3090 800 3120
rect 3417 3090 3483 3093
rect 0 3088 3483 3090
rect 0 3032 3422 3088
rect 3478 3032 3483 3088
rect 0 3030 3483 3032
rect 4110 3090 4170 3438
rect 4245 3496 6151 3498
rect 4245 3440 4250 3496
rect 4306 3440 6090 3496
rect 6146 3440 6151 3496
rect 4245 3438 6151 3440
rect 4245 3435 4311 3438
rect 6085 3435 6151 3438
rect 7281 3498 7347 3501
rect 11973 3498 12039 3501
rect 7281 3496 12039 3498
rect 7281 3440 7286 3496
rect 7342 3440 11978 3496
rect 12034 3440 12039 3496
rect 7281 3438 12039 3440
rect 12390 3498 12450 3574
rect 13445 3632 26943 3634
rect 13445 3576 13450 3632
rect 13506 3576 26882 3632
rect 26938 3576 26943 3632
rect 13445 3574 26943 3576
rect 13445 3571 13511 3574
rect 26877 3571 26943 3574
rect 17953 3498 18019 3501
rect 12390 3496 18019 3498
rect 12390 3440 17958 3496
rect 18014 3440 18019 3496
rect 12390 3438 18019 3440
rect 7281 3435 7347 3438
rect 11973 3435 12039 3438
rect 17953 3435 18019 3438
rect 5441 3362 5507 3365
rect 8201 3362 8267 3365
rect 5441 3360 8267 3362
rect 5441 3304 5446 3360
rect 5502 3304 8206 3360
rect 8262 3304 8267 3360
rect 5441 3302 8267 3304
rect 5441 3299 5507 3302
rect 8201 3299 8267 3302
rect 8477 3362 8543 3365
rect 11329 3362 11395 3365
rect 14549 3362 14615 3365
rect 8477 3360 11395 3362
rect 8477 3304 8482 3360
rect 8538 3304 11334 3360
rect 11390 3304 11395 3360
rect 8477 3302 11395 3304
rect 8477 3299 8543 3302
rect 11329 3299 11395 3302
rect 12068 3360 14615 3362
rect 12068 3304 14554 3360
rect 14610 3304 14615 3360
rect 12068 3302 14615 3304
rect 4613 3226 4679 3229
rect 12068 3226 12128 3302
rect 14549 3299 14615 3302
rect 14917 3362 14983 3365
rect 27153 3362 27219 3365
rect 14917 3360 27219 3362
rect 14917 3304 14922 3360
rect 14978 3304 27158 3360
rect 27214 3304 27219 3360
rect 14917 3302 27219 3304
rect 14917 3299 14983 3302
rect 27153 3299 27219 3302
rect 4613 3224 12128 3226
rect 4613 3168 4618 3224
rect 4674 3168 12128 3224
rect 4613 3166 12128 3168
rect 12249 3226 12315 3229
rect 15929 3226 15995 3229
rect 12249 3224 15995 3226
rect 12249 3168 12254 3224
rect 12310 3168 15934 3224
rect 15990 3168 15995 3224
rect 12249 3166 15995 3168
rect 4613 3163 4679 3166
rect 12249 3163 12315 3166
rect 15929 3163 15995 3166
rect 17309 3226 17375 3229
rect 23933 3226 23999 3229
rect 17309 3224 23999 3226
rect 17309 3168 17314 3224
rect 17370 3168 23938 3224
rect 23994 3168 23999 3224
rect 17309 3166 23999 3168
rect 17309 3163 17375 3166
rect 23933 3163 23999 3166
rect 24577 3090 24643 3093
rect 4110 3088 24643 3090
rect 4110 3032 24582 3088
rect 24638 3032 24643 3088
rect 4110 3030 24643 3032
rect 0 3000 800 3030
rect 3417 3027 3483 3030
rect 24577 3027 24643 3030
rect 4429 2954 4495 2957
rect 7373 2954 7439 2957
rect 4429 2952 7439 2954
rect 4429 2896 4434 2952
rect 4490 2896 7378 2952
rect 7434 2896 7439 2952
rect 4429 2894 7439 2896
rect 4429 2891 4495 2894
rect 7373 2891 7439 2894
rect 7557 2954 7623 2957
rect 17309 2954 17375 2957
rect 7557 2952 17375 2954
rect 7557 2896 7562 2952
rect 7618 2896 17314 2952
rect 17370 2896 17375 2952
rect 7557 2894 17375 2896
rect 7557 2891 7623 2894
rect 17309 2891 17375 2894
rect 17769 2954 17835 2957
rect 20161 2954 20227 2957
rect 17769 2952 20227 2954
rect 17769 2896 17774 2952
rect 17830 2896 20166 2952
rect 20222 2896 20227 2952
rect 17769 2894 20227 2896
rect 17769 2891 17835 2894
rect 20161 2891 20227 2894
rect 20345 2954 20411 2957
rect 23289 2954 23355 2957
rect 20345 2952 23355 2954
rect 20345 2896 20350 2952
rect 20406 2896 23294 2952
rect 23350 2896 23355 2952
rect 20345 2894 23355 2896
rect 20345 2891 20411 2894
rect 23289 2891 23355 2894
rect 28993 2954 29059 2957
rect 33400 2954 34200 2984
rect 28993 2952 34200 2954
rect 28993 2896 28998 2952
rect 29054 2896 34200 2952
rect 28993 2894 34200 2896
rect 28993 2891 29059 2894
rect 33400 2864 34200 2894
rect 1669 2818 1735 2821
rect 27613 2818 27679 2821
rect 1669 2816 27679 2818
rect 1669 2760 1674 2816
rect 1730 2760 27618 2816
rect 27674 2760 27679 2816
rect 1669 2758 27679 2760
rect 1669 2755 1735 2758
rect 27613 2755 27679 2758
rect 0 2682 800 2712
rect 4061 2682 4127 2685
rect 9489 2682 9555 2685
rect 0 2680 4127 2682
rect 0 2624 4066 2680
rect 4122 2624 4127 2680
rect 0 2622 4127 2624
rect 0 2592 800 2622
rect 4061 2619 4127 2622
rect 4294 2680 9555 2682
rect 4294 2624 9494 2680
rect 9550 2624 9555 2680
rect 4294 2622 9555 2624
rect 4294 2546 4354 2622
rect 9489 2619 9555 2622
rect 9673 2682 9739 2685
rect 15009 2682 15075 2685
rect 9673 2680 15075 2682
rect 9673 2624 9678 2680
rect 9734 2624 15014 2680
rect 15070 2624 15075 2680
rect 9673 2622 15075 2624
rect 9673 2619 9739 2622
rect 15009 2619 15075 2622
rect 19241 2682 19307 2685
rect 20713 2682 20779 2685
rect 19241 2680 20779 2682
rect 19241 2624 19246 2680
rect 19302 2624 20718 2680
rect 20774 2624 20779 2680
rect 19241 2622 20779 2624
rect 19241 2619 19307 2622
rect 20713 2619 20779 2622
rect 2730 2486 4354 2546
rect 4797 2546 4863 2549
rect 6545 2546 6611 2549
rect 4797 2544 6611 2546
rect 4797 2488 4802 2544
rect 4858 2488 6550 2544
rect 6606 2488 6611 2544
rect 4797 2486 6611 2488
rect 0 2274 800 2304
rect 2730 2274 2790 2486
rect 4797 2483 4863 2486
rect 6545 2483 6611 2486
rect 6913 2546 6979 2549
rect 15653 2546 15719 2549
rect 6913 2544 15719 2546
rect 6913 2488 6918 2544
rect 6974 2488 15658 2544
rect 15714 2488 15719 2544
rect 6913 2486 15719 2488
rect 6913 2483 6979 2486
rect 15653 2483 15719 2486
rect 15837 2546 15903 2549
rect 20529 2546 20595 2549
rect 15837 2544 20595 2546
rect 15837 2488 15842 2544
rect 15898 2488 20534 2544
rect 20590 2488 20595 2544
rect 15837 2486 20595 2488
rect 15837 2483 15903 2486
rect 20529 2483 20595 2486
rect 3325 2410 3391 2413
rect 7005 2410 7071 2413
rect 3325 2408 7071 2410
rect 3325 2352 3330 2408
rect 3386 2352 7010 2408
rect 7066 2352 7071 2408
rect 3325 2350 7071 2352
rect 3325 2347 3391 2350
rect 7005 2347 7071 2350
rect 7373 2410 7439 2413
rect 12249 2410 12315 2413
rect 7373 2408 12315 2410
rect 7373 2352 7378 2408
rect 7434 2352 12254 2408
rect 12310 2352 12315 2408
rect 7373 2350 12315 2352
rect 7373 2347 7439 2350
rect 12249 2347 12315 2350
rect 12387 2410 12453 2413
rect 18597 2410 18663 2413
rect 20161 2410 20227 2413
rect 12387 2408 18522 2410
rect 12387 2352 12392 2408
rect 12448 2352 18522 2408
rect 12387 2350 18522 2352
rect 12387 2347 12453 2350
rect 0 2214 2790 2274
rect 5901 2274 5967 2277
rect 18462 2274 18522 2350
rect 18597 2408 20227 2410
rect 18597 2352 18602 2408
rect 18658 2352 20166 2408
rect 20222 2352 20227 2408
rect 18597 2350 20227 2352
rect 18597 2347 18663 2350
rect 20161 2347 20227 2350
rect 20529 2274 20595 2277
rect 5901 2272 18338 2274
rect 5901 2216 5906 2272
rect 5962 2216 18338 2272
rect 5901 2214 18338 2216
rect 18462 2272 20595 2274
rect 18462 2216 20534 2272
rect 20590 2216 20595 2272
rect 18462 2214 20595 2216
rect 0 2184 800 2214
rect 5901 2211 5967 2214
rect 4521 2138 4587 2141
rect 18045 2138 18111 2141
rect 4521 2136 18111 2138
rect 4521 2080 4526 2136
rect 4582 2080 18050 2136
rect 18106 2080 18111 2136
rect 4521 2078 18111 2080
rect 18278 2138 18338 2214
rect 20529 2211 20595 2214
rect 21357 2138 21423 2141
rect 18278 2136 21423 2138
rect 18278 2080 21362 2136
rect 21418 2080 21423 2136
rect 18278 2078 21423 2080
rect 4521 2075 4587 2078
rect 18045 2075 18111 2078
rect 21357 2075 21423 2078
rect 4705 2002 4771 2005
rect 22001 2002 22067 2005
rect 4705 2000 22067 2002
rect 4705 1944 4710 2000
rect 4766 1944 22006 2000
rect 22062 1944 22067 2000
rect 4705 1942 22067 1944
rect 4705 1939 4771 1942
rect 22001 1939 22067 1942
rect 0 1866 800 1896
rect 2773 1866 2839 1869
rect 0 1864 2839 1866
rect 0 1808 2778 1864
rect 2834 1808 2839 1864
rect 0 1806 2839 1808
rect 0 1776 800 1806
rect 2773 1803 2839 1806
rect 2957 1866 3023 1869
rect 12249 1866 12315 1869
rect 2957 1864 12315 1866
rect 2957 1808 2962 1864
rect 3018 1808 12254 1864
rect 12310 1808 12315 1864
rect 2957 1806 12315 1808
rect 2957 1803 3023 1806
rect 12249 1803 12315 1806
rect 13077 1866 13143 1869
rect 15837 1866 15903 1869
rect 13077 1864 15903 1866
rect 13077 1808 13082 1864
rect 13138 1808 15842 1864
rect 15898 1808 15903 1864
rect 13077 1806 15903 1808
rect 13077 1803 13143 1806
rect 15837 1803 15903 1806
rect 17861 1866 17927 1869
rect 19977 1866 20043 1869
rect 17861 1864 20043 1866
rect 17861 1808 17866 1864
rect 17922 1808 19982 1864
rect 20038 1808 20043 1864
rect 17861 1806 20043 1808
rect 17861 1803 17927 1806
rect 19977 1803 20043 1806
rect 4889 1730 4955 1733
rect 12157 1730 12223 1733
rect 4889 1728 12223 1730
rect 4889 1672 4894 1728
rect 4950 1672 12162 1728
rect 12218 1672 12223 1728
rect 4889 1670 12223 1672
rect 4889 1667 4955 1670
rect 12157 1667 12223 1670
rect 12985 1730 13051 1733
rect 16021 1730 16087 1733
rect 18413 1730 18479 1733
rect 12985 1728 18479 1730
rect 12985 1672 12990 1728
rect 13046 1672 16026 1728
rect 16082 1672 18418 1728
rect 18474 1672 18479 1728
rect 12985 1670 18479 1672
rect 12985 1667 13051 1670
rect 16021 1667 16087 1670
rect 18413 1667 18479 1670
rect 18597 1730 18663 1733
rect 22185 1730 22251 1733
rect 18597 1728 22251 1730
rect 18597 1672 18602 1728
rect 18658 1672 22190 1728
rect 22246 1672 22251 1728
rect 18597 1670 22251 1672
rect 18597 1667 18663 1670
rect 22185 1667 22251 1670
rect 20253 1594 20319 1597
rect 2730 1592 20319 1594
rect 2730 1536 20258 1592
rect 20314 1536 20319 1592
rect 2730 1534 20319 1536
rect 0 1458 800 1488
rect 2730 1458 2790 1534
rect 20253 1531 20319 1534
rect 0 1398 2790 1458
rect 10501 1458 10567 1461
rect 12341 1458 12407 1461
rect 10501 1456 12407 1458
rect 10501 1400 10506 1456
rect 10562 1400 12346 1456
rect 12402 1400 12407 1456
rect 10501 1398 12407 1400
rect 0 1368 800 1398
rect 10501 1395 10567 1398
rect 12341 1395 12407 1398
rect 15009 1458 15075 1461
rect 19793 1458 19859 1461
rect 15009 1456 19859 1458
rect 15009 1400 15014 1456
rect 15070 1400 19798 1456
rect 19854 1400 19859 1456
rect 15009 1398 19859 1400
rect 15009 1395 15075 1398
rect 19793 1395 19859 1398
rect 21357 1458 21423 1461
rect 24853 1458 24919 1461
rect 21357 1456 24919 1458
rect 21357 1400 21362 1456
rect 21418 1400 24858 1456
rect 24914 1400 24919 1456
rect 21357 1398 24919 1400
rect 21357 1395 21423 1398
rect 24853 1395 24919 1398
rect 3877 1322 3943 1325
rect 19885 1322 19951 1325
rect 3877 1320 19951 1322
rect 3877 1264 3882 1320
rect 3938 1264 19890 1320
rect 19946 1264 19951 1320
rect 3877 1262 19951 1264
rect 3877 1259 3943 1262
rect 19885 1259 19951 1262
rect 3969 1186 4035 1189
rect 15745 1186 15811 1189
rect 3969 1184 15811 1186
rect 3969 1128 3974 1184
rect 4030 1128 15750 1184
rect 15806 1128 15811 1184
rect 3969 1126 15811 1128
rect 3969 1123 4035 1126
rect 15745 1123 15811 1126
rect 20253 1186 20319 1189
rect 23473 1186 23539 1189
rect 20253 1184 23539 1186
rect 20253 1128 20258 1184
rect 20314 1128 23478 1184
rect 23534 1128 23539 1184
rect 20253 1126 23539 1128
rect 20253 1123 20319 1126
rect 23473 1123 23539 1126
rect 0 1050 800 1080
rect 22737 1050 22803 1053
rect 0 1048 22803 1050
rect 0 992 22742 1048
rect 22798 992 22803 1048
rect 0 990 22803 992
rect 0 960 800 990
rect 22737 987 22803 990
rect 4337 914 4403 917
rect 14917 914 14983 917
rect 24853 914 24919 917
rect 4337 912 24919 914
rect 4337 856 4342 912
rect 4398 856 14922 912
rect 14978 856 24858 912
rect 24914 856 24919 912
rect 4337 854 24919 856
rect 4337 851 4403 854
rect 14917 851 14983 854
rect 24853 851 24919 854
rect 3601 778 3667 781
rect 20345 778 20411 781
rect 3601 776 20411 778
rect 3601 720 3606 776
rect 3662 720 20350 776
rect 20406 720 20411 776
rect 3601 718 20411 720
rect 3601 715 3667 718
rect 20345 715 20411 718
rect 21357 778 21423 781
rect 24209 778 24275 781
rect 21357 776 24275 778
rect 21357 720 21362 776
rect 21418 720 24214 776
rect 24270 720 24275 776
rect 21357 718 24275 720
rect 21357 715 21423 718
rect 24209 715 24275 718
rect 0 642 800 672
rect 1393 642 1459 645
rect 0 640 1459 642
rect 0 584 1398 640
rect 1454 584 1459 640
rect 0 582 1459 584
rect 0 552 800 582
rect 1393 579 1459 582
rect 3049 642 3115 645
rect 20253 642 20319 645
rect 22093 642 22159 645
rect 3049 640 22159 642
rect 3049 584 3054 640
rect 3110 584 20258 640
rect 20314 584 22098 640
rect 22154 584 22159 640
rect 3049 582 22159 584
rect 3049 579 3115 582
rect 20253 579 20319 582
rect 22093 579 22159 582
rect 3417 506 3483 509
rect 23289 506 23355 509
rect 3417 504 23355 506
rect 3417 448 3422 504
rect 3478 448 23294 504
rect 23350 448 23355 504
rect 3417 446 23355 448
rect 3417 443 3483 446
rect 23289 443 23355 446
rect 3785 370 3851 373
rect 20713 370 20779 373
rect 3785 368 20779 370
rect 3785 312 3790 368
rect 3846 312 20718 368
rect 20774 312 20779 368
rect 3785 310 20779 312
rect 3785 307 3851 310
rect 20713 307 20779 310
rect 0 234 800 264
rect 1577 234 1643 237
rect 0 232 1643 234
rect 0 176 1582 232
rect 1638 176 1643 232
rect 0 174 1643 176
rect 0 144 800 174
rect 1577 171 1643 174
rect 9949 234 10015 237
rect 12065 234 12131 237
rect 15193 234 15259 237
rect 9949 232 12131 234
rect 9949 176 9954 232
rect 10010 176 12070 232
rect 12126 176 12131 232
rect 9949 174 12131 176
rect 9949 171 10015 174
rect 12065 171 12131 174
rect 12206 232 15259 234
rect 12206 176 15198 232
rect 15254 176 15259 232
rect 12206 174 15259 176
rect 9489 98 9555 101
rect 12206 98 12266 174
rect 15193 171 15259 174
rect 9489 96 12266 98
rect 9489 40 9494 96
rect 9550 40 12266 96
rect 9489 38 12266 40
rect 12341 98 12407 101
rect 17953 98 18019 101
rect 12341 96 18019 98
rect 12341 40 12346 96
rect 12402 40 17958 96
rect 18014 40 18019 96
rect 12341 38 18019 40
rect 9489 35 9555 38
rect 12341 35 12407 38
rect 17953 35 18019 38
use sky130_fd_sc_hd__diode_2  ANTENNA_clkgen.delay_155ns_1.enablebuffer_A
timestamp 1515178157
transform -1 0 24380 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkgen.delay_155ns_1.genblk1\[0\].control_invert_A
timestamp 1515178157
transform -1 0 24380 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkgen.delay_155ns_1.genblk1\[0\].dly_binary.and_bypass_switch_A_N
timestamp 1515178157
transform -1 0 27140 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkgen.delay_155ns_1.genblk1\[0\].dly_binary.out_mux_S
timestamp 1515178157
transform 1 0 25852 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkgen.delay_155ns_1.genblk1\[1\].control_invert_A
timestamp 1515178157
transform -1 0 25484 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkgen.delay_155ns_1.genblk1\[2\].control_invert_A
timestamp 1515178157
transform -1 0 26312 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkgen.delay_155ns_1.genblk1\[3\].control_invert_A
timestamp 1515178157
transform -1 0 24932 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkgen.delay_155ns_1.genblk1\[3\].dly_binary.and_bypass_switch_A_N
timestamp 1515178157
transform 1 0 23276 0 -1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkgen.delay_155ns_1.genblk1\[3\].dly_binary.out_mux_A0
timestamp 1515178157
transform -1 0 30820 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkgen.delay_155ns_1.genblk1\[3\].dly_binary.out_mux_S
timestamp 1515178157
transform -1 0 29992 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkgen.delay_155ns_1.genblk1\[4\].control_invert_A
timestamp 1515178157
transform -1 0 24932 0 -1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkgen.delay_155ns_1.genblk1\[4\].dly_binary.and_bypass_switch_B
timestamp 1515178157
transform 1 0 23828 0 1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkgen.delay_155ns_1.genblk1\[4\].dly_binary.out_mux_A1
timestamp 1515178157
transform -1 0 25484 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkgen.delay_155ns_2.enablebuffer_A
timestamp 1515178157
transform -1 0 23460 0 1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkgen.delay_155ns_2.genblk1\[0\].control_invert_A
timestamp 1515178157
transform -1 0 24380 0 -1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkgen.delay_155ns_2.genblk1\[0\].dly_binary.and_bypass_switch_B
timestamp 1515178157
transform 1 0 25024 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkgen.delay_155ns_2.genblk1\[0\].dly_binary.out_mux_A1
timestamp 1515178157
transform -1 0 22908 0 -1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkgen.delay_155ns_2.genblk1\[1\].control_invert_A
timestamp 1515178157
transform -1 0 23276 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkgen.delay_155ns_2.genblk1\[1\].dly_binary.and_bypass_switch_A_N
timestamp 1515178157
transform -1 0 22172 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkgen.delay_155ns_2.genblk1\[1\].dly_binary.and_bypass_switch_B
timestamp 1515178157
transform -1 0 22724 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkgen.delay_155ns_2.genblk1\[1\].dly_binary.out_mux_A1
timestamp 1515178157
transform -1 0 26588 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkgen.delay_155ns_2.genblk1\[1\].dly_binary.out_mux_S
timestamp 1515178157
transform -1 0 25668 0 1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkgen.delay_155ns_2.genblk1\[2\].control_invert_A
timestamp 1515178157
transform -1 0 25760 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkgen.delay_155ns_2.genblk1\[2\].dly_binary.and_bypass_switch_A_N
timestamp 1515178157
transform -1 0 22356 0 -1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkgen.delay_155ns_2.genblk1\[2\].dly_binary.out_mux_S
timestamp 1515178157
transform -1 0 27232 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkgen.delay_155ns_2.genblk1\[3\].control_invert_A
timestamp 1515178157
transform -1 0 24564 0 1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkgen.delay_155ns_2.genblk1\[3\].dly_binary.and_bypass_switch_A_N
timestamp 1515178157
transform -1 0 23736 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkgen.delay_155ns_2.genblk1\[3\].dly_binary.out_mux_S
timestamp 1515178157
transform -1 0 27784 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkgen.delay_155ns_2.genblk1\[4\].control_invert_A
timestamp 1515178157
transform -1 0 28704 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkgen.delay_155ns_2.genblk1\[4\].dly_binary.and_bypass_switch_A_N
timestamp 1515178157
transform 1 0 27048 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkgen.delay_155ns_2.genblk1\[4\].dly_binary.out_mux_A0
timestamp 1515178157
transform -1 0 29256 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkgen.delay_155ns_2.genblk1\[4\].dly_binary.out_mux_S
timestamp 1515178157
transform -1 0 28888 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkgen.delay_155ns_3.enablebuffer_A
timestamp 1515178157
transform 1 0 16836 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkgen.delay_155ns_3.genblk1\[0\].control_invert_A
timestamp 1515178157
transform -1 0 27784 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkgen.delay_155ns_3.genblk1\[1\].control_invert_A
timestamp 1515178157
transform -1 0 27048 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkgen.delay_155ns_3.genblk1\[2\].control_invert_A
timestamp 1515178157
transform -1 0 27232 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkgen.delay_155ns_3.genblk1\[3\].control_invert_A
timestamp 1515178157
transform -1 0 28152 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkgen.delay_155ns_3.genblk1\[4\].control_invert_A
timestamp 1515178157
transform -1 0 24932 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_delay_sample_n12_in
timestamp 1515178157
transform -1 0 27784 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_delay_sample_p11_in
timestamp 1515178157
transform -1 0 30912 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_edgedetect.dly_315ns_1.enablebuffer_A
timestamp 1515178157
transform 1 0 9292 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_edgedetect.dly_315ns_1.genblk1\[0\].control_invert_A
timestamp 1515178157
transform -1 0 28336 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_edgedetect.dly_315ns_1.genblk1\[0\].dly_binary.and_bypass_switch_A_N
timestamp 1515178157
transform 1 0 27416 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_edgedetect.dly_315ns_1.genblk1\[0\].dly_binary.and_bypass_switch_B
timestamp 1515178157
transform -1 0 12328 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_edgedetect.dly_315ns_1.genblk1\[0\].dly_binary.out_mux_A1
timestamp 1515178157
transform -1 0 29440 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_edgedetect.dly_315ns_1.genblk1\[0\].dly_binary.out_mux_S
timestamp 1515178157
transform -1 0 30084 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_edgedetect.dly_315ns_1.genblk1\[1\].control_invert_A
timestamp 1515178157
transform -1 0 29072 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_edgedetect.dly_315ns_1.genblk1\[1\].dly_binary.and_bypass_switch_B
timestamp 1515178157
transform -1 0 26496 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_edgedetect.dly_315ns_1.genblk1\[1\].dly_binary.out_mux_A1
timestamp 1515178157
transform -1 0 29256 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_edgedetect.dly_315ns_1.genblk1\[2\].control_invert_A
timestamp 1515178157
transform -1 0 28152 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_edgedetect.dly_315ns_1.genblk1\[3\].control_invert_A
timestamp 1515178157
transform -1 0 28520 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.genblk1\[0\].delay_unit_in
timestamp 1515178157
transform -1 0 30360 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_edgedetect.dly_315ns_1.genblk1\[4\].control_invert_A
timestamp 1515178157
transform -1 0 29072 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[0\].delay_unit_in
timestamp 1515178157
transform -1 0 30084 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_edgedetect.dly_315ns_1.genblk1\[5\].control_invert_A
timestamp 1515178157
transform -1 0 28704 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_edgedetect.nor1_B_N
timestamp 1515178157
transform -1 0 27600 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_edgedetect.or1_A
timestamp 1515178157
transform -1 0 30544 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_edgedetect.or1_B
timestamp 1515178157
transform -1 0 31096 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_inbuf_1_A
timestamp 1515178157
transform -1 0 25116 0 1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_inbuf_2_A
timestamp 1515178157
transform -1 0 27232 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_inbuf_3_A
timestamp 1515178157
transform -1 0 27232 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_outbuf_1_A
timestamp 1515178157
transform -1 0 26220 0 1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  clkgen.clkdig_inverter
timestamp 1515178157
transform 1 0 22816 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  clkgen.delay_155ns_1.enablebuffer
timestamp 1515178157
transform 1 0 21344 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  clkgen.delay_155ns_1.genblk1\[0\].bypass_enable
timestamp 1515178157
transform -1 0 18952 0 1 544
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  clkgen.delay_155ns_1.genblk1\[0\].control_invert
timestamp 1515178157
transform -1 0 21620 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  clkgen.delay_155ns_1.genblk1\[0\].dly_binary.and_bypass_switch
timestamp 1515178157
transform 1 0 1748 0 -1 3808
box -38 -48 590 592
use sky130_mm_sc_hd_dlyPoly5ns  clkgen.delay_155ns_1.genblk1\[0\].dly_binary.genblk1\[0\].delay_unit
timestamp 1515178157
transform 1 0 7268 0 1 2720
box -38 -48 2246 592
use sky130_fd_sc_hd__mux2_1  clkgen.delay_155ns_1.genblk1\[0\].dly_binary.out_mux
timestamp 1515178157
transform 1 0 7728 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  clkgen.delay_155ns_1.genblk1\[1\].bypass_enable
timestamp 1515178157
transform -1 0 22448 0 -1 2720
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  clkgen.delay_155ns_1.genblk1\[1\].control_invert
timestamp 1515178157
transform -1 0 23736 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  clkgen.delay_155ns_1.genblk1\[1\].dly_binary.and_bypass_switch
timestamp 1515178157
transform -1 0 18032 0 -1 3808
box -38 -48 590 592
use sky130_mm_sc_hd_dlyPoly5ns  clkgen.delay_155ns_1.genblk1\[1\].dly_binary.genblk1\[0\].delay_unit
timestamp 1515178157
transform -1 0 9476 0 1 1632
box -38 -48 2246 592
use sky130_mm_sc_hd_dlyPoly5ns  clkgen.delay_155ns_1.genblk1\[1\].dly_binary.genblk1\[1\].delay_unit
timestamp 1515178157
transform 1 0 9016 0 -1 3808
box -38 -48 2246 592
use sky130_fd_sc_hd__mux2_1  clkgen.delay_155ns_1.genblk1\[1\].dly_binary.out_mux
timestamp 1515178157
transform -1 0 6348 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  clkgen.delay_155ns_1.genblk1\[2\].bypass_enable
timestamp 1515178157
transform -1 0 22724 0 1 2720
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  clkgen.delay_155ns_1.genblk1\[2\].control_invert
timestamp 1515178157
transform -1 0 24656 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  clkgen.delay_155ns_1.genblk1\[2\].dly_binary.and_bypass_switch
timestamp 1515178157
transform -1 0 14536 0 1 544
box -38 -48 590 592
use sky130_mm_sc_hd_dlyPoly5ns  clkgen.delay_155ns_1.genblk1\[2\].dly_binary.genblk1\[0\].delay_unit
timestamp 1515178157
transform -1 0 6900 0 1 2720
box -38 -48 2246 592
use sky130_mm_sc_hd_dlyPoly5ns  clkgen.delay_155ns_1.genblk1\[2\].dly_binary.genblk1\[1\].delay_unit
timestamp 1515178157
transform 1 0 7544 0 -1 2720
box -38 -48 2246 592
use sky130_mm_sc_hd_dlyPoly5ns  clkgen.delay_155ns_1.genblk1\[2\].dly_binary.genblk1\[2\].delay_unit
timestamp 1515178157
transform 1 0 10120 0 -1 2720
box -38 -48 2246 592
use sky130_mm_sc_hd_dlyPoly5ns  clkgen.delay_155ns_1.genblk1\[2\].dly_binary.genblk1\[3\].delay_unit
timestamp 1515178157
transform -1 0 12604 0 1 2720
box -38 -48 2246 592
use sky130_fd_sc_hd__mux2_1  clkgen.delay_155ns_1.genblk1\[2\].dly_binary.out_mux
timestamp 1515178157
transform -1 0 9200 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  clkgen.delay_155ns_1.genblk1\[3\].bypass_enable
timestamp 1515178157
transform 1 0 19320 0 1 544
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  clkgen.delay_155ns_1.genblk1\[3\].control_invert
timestamp 1515178157
transform -1 0 24012 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  clkgen.delay_155ns_1.genblk1\[3\].dly_binary.and_bypass_switch
timestamp 1515178157
transform -1 0 16192 0 1 1632
box -38 -48 590 592
use sky130_mm_sc_hd_dlyPoly5ns  clkgen.delay_155ns_1.genblk1\[3\].dly_binary.genblk1\[0\].delay_unit
timestamp 1515178157
transform -1 0 6624 0 -1 2720
box -38 -48 2246 592
use sky130_mm_sc_hd_dlyPoly5ns  clkgen.delay_155ns_1.genblk1\[3\].dly_binary.genblk1\[1\].delay_unit
timestamp 1515178157
transform 1 0 7544 0 -1 1632
box -38 -48 2246 592
use sky130_mm_sc_hd_dlyPoly5ns  clkgen.delay_155ns_1.genblk1\[3\].dly_binary.genblk1\[2\].delay_unit
timestamp 1515178157
transform 1 0 10396 0 1 1632
box -38 -48 2246 592
use sky130_mm_sc_hd_dlyPoly5ns  clkgen.delay_155ns_1.genblk1\[3\].dly_binary.genblk1\[3\].delay_unit
timestamp 1515178157
transform 1 0 12788 0 -1 2720
box -38 -48 2246 592
use sky130_mm_sc_hd_dlyPoly5ns  clkgen.delay_155ns_1.genblk1\[3\].dly_binary.genblk1\[4\].delay_unit
timestamp 1515178157
transform 1 0 12972 0 1 2720
box -38 -48 2246 592
use sky130_mm_sc_hd_dlyPoly5ns  clkgen.delay_155ns_1.genblk1\[3\].dly_binary.genblk1\[5\].delay_unit
timestamp 1515178157
transform 1 0 15548 0 -1 2720
box -38 -48 2246 592
use sky130_mm_sc_hd_dlyPoly5ns  clkgen.delay_155ns_1.genblk1\[3\].dly_binary.genblk1\[6\].delay_unit
timestamp 1515178157
transform 1 0 18492 0 -1 3808
box -38 -48 2246 592
use sky130_mm_sc_hd_dlyPoly5ns  clkgen.delay_155ns_1.genblk1\[3\].dly_binary.genblk1\[7\].delay_unit
timestamp 1515178157
transform -1 0 20700 0 -1 2720
box -38 -48 2246 592
use sky130_fd_sc_hd__mux2_1  clkgen.delay_155ns_1.genblk1\[3\].dly_binary.out_mux
timestamp 1515178157
transform -1 0 2576 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  clkgen.delay_155ns_1.genblk1\[4\].bypass_enable
timestamp 1515178157
transform 1 0 20424 0 1 1632
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  clkgen.delay_155ns_1.genblk1\[4\].control_invert
timestamp 1515178157
transform -1 0 21804 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  clkgen.delay_155ns_1.genblk1\[4\].dly_binary.and_bypass_switch
timestamp 1515178157
transform -1 0 21620 0 -1 2720
box -38 -48 590 592
use sky130_mm_sc_hd_dlyPoly5ns  clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[0\].delay_unit
timestamp 1515178157
transform -1 0 3864 0 -1 2720
box -38 -48 2246 592
use sky130_mm_sc_hd_dlyPoly5ns  clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[1\].delay_unit
timestamp 1515178157
transform 1 0 1564 0 1 1632
box -38 -48 2246 592
use sky130_mm_sc_hd_dlyPoly5ns  clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[2\].delay_unit
timestamp 1515178157
transform -1 0 3772 0 1 544
box -38 -48 2246 592
use sky130_mm_sc_hd_dlyPoly5ns  clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[3\].delay_unit
timestamp 1515178157
transform 1 0 1840 0 -1 1632
box -38 -48 2246 592
use sky130_mm_sc_hd_dlyPoly5ns  clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[4\].delay_unit
timestamp 1515178157
transform 1 0 4416 0 1 544
box -38 -48 2246 592
use sky130_mm_sc_hd_dlyPoly5ns  clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[5\].delay_unit
timestamp 1515178157
transform -1 0 6900 0 1 1632
box -38 -48 2246 592
use sky130_mm_sc_hd_dlyPoly5ns  clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[6\].delay_unit
timestamp 1515178157
transform 1 0 4416 0 -1 1632
box -38 -48 2246 592
use sky130_mm_sc_hd_dlyPoly5ns  clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[7\].delay_unit
timestamp 1515178157
transform 1 0 7268 0 1 544
box -38 -48 2246 592
use sky130_mm_sc_hd_dlyPoly5ns  clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[8\].delay_unit
timestamp 1515178157
transform 1 0 10120 0 1 544
box -38 -48 2246 592
use sky130_mm_sc_hd_dlyPoly5ns  clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[9\].delay_unit
timestamp 1515178157
transform -1 0 12328 0 -1 1632
box -38 -48 2246 592
use sky130_mm_sc_hd_dlyPoly5ns  clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[10\].delay_unit
timestamp 1515178157
transform 1 0 12972 0 -1 1632
box -38 -48 2246 592
use sky130_mm_sc_hd_dlyPoly5ns  clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[11\].delay_unit
timestamp 1515178157
transform -1 0 15180 0 1 1632
box -38 -48 2246 592
use sky130_mm_sc_hd_dlyPoly5ns  clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[12\].delay_unit
timestamp 1515178157
transform 1 0 15640 0 1 544
box -38 -48 2246 592
use sky130_mm_sc_hd_dlyPoly5ns  clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[13\].delay_unit
timestamp 1515178157
transform 1 0 15824 0 -1 1632
box -38 -48 2246 592
use sky130_mm_sc_hd_dlyPoly5ns  clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[14\].delay_unit
timestamp 1515178157
transform 1 0 17848 0 1 1632
box -38 -48 2246 592
use sky130_mm_sc_hd_dlyPoly5ns  clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[15\].delay_unit
timestamp 1515178157
transform -1 0 21160 0 -1 1632
box -38 -48 2246 592
use sky130_fd_sc_hd__mux2_1  clkgen.delay_155ns_1.genblk1\[4\].dly_binary.out_mux
timestamp 1515178157
transform -1 0 13616 0 1 544
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  clkgen.delay_155ns_2.enablebuffer
timestamp 1515178157
transform -1 0 22540 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  clkgen.delay_155ns_2.genblk1\[0\].bypass_enable
timestamp 1515178157
transform -1 0 23184 0 -1 3808
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  clkgen.delay_155ns_2.genblk1\[0\].control_invert
timestamp 1515178157
transform 1 0 21988 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  clkgen.delay_155ns_2.genblk1\[0\].dly_binary.and_bypass_switch
timestamp 1515178157
transform -1 0 20516 0 1 2720
box -38 -48 590 592
use sky130_mm_sc_hd_dlyPoly5ns  clkgen.delay_155ns_2.genblk1\[0\].dly_binary.genblk1\[0\].delay_unit
timestamp 1515178157
transform -1 0 3772 0 1 3808
box -38 -48 2246 592
use sky130_fd_sc_hd__mux2_1  clkgen.delay_155ns_2.genblk1\[0\].dly_binary.out_mux
timestamp 1515178157
transform -1 0 16468 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  clkgen.delay_155ns_2.genblk1\[1\].bypass_enable
timestamp 1515178157
transform 1 0 23276 0 -1 4896
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  clkgen.delay_155ns_2.genblk1\[1\].control_invert
timestamp 1515178157
transform 1 0 20148 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  clkgen.delay_155ns_2.genblk1\[1\].dly_binary.and_bypass_switch
timestamp 1515178157
transform -1 0 17112 0 1 1632
box -38 -48 590 592
use sky130_mm_sc_hd_dlyPoly5ns  clkgen.delay_155ns_2.genblk1\[1\].dly_binary.genblk1\[0\].delay_unit
timestamp 1515178157
transform -1 0 4048 0 -1 4896
box -38 -48 2246 592
use sky130_mm_sc_hd_dlyPoly5ns  clkgen.delay_155ns_2.genblk1\[1\].dly_binary.genblk1\[1\].delay_unit
timestamp 1515178157
transform 1 0 4416 0 -1 4896
box -38 -48 2246 592
use sky130_fd_sc_hd__mux2_1  clkgen.delay_155ns_2.genblk1\[1\].dly_binary.out_mux
timestamp 1515178157
transform -1 0 2852 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  clkgen.delay_155ns_2.genblk1\[2\].bypass_enable
timestamp 1515178157
transform 1 0 21896 0 -1 3808
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  clkgen.delay_155ns_2.genblk1\[2\].control_invert
timestamp 1515178157
transform -1 0 23368 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  clkgen.delay_155ns_2.genblk1\[2\].dly_binary.and_bypass_switch
timestamp 1515178157
transform -1 0 19044 0 -1 4896
box -38 -48 590 592
use sky130_mm_sc_hd_dlyPoly5ns  clkgen.delay_155ns_2.genblk1\[2\].dly_binary.genblk1\[0\].delay_unit
timestamp 1515178157
transform -1 0 6624 0 -1 3808
box -38 -48 2246 592
use sky130_mm_sc_hd_dlyPoly5ns  clkgen.delay_155ns_2.genblk1\[2\].dly_binary.genblk1\[1\].delay_unit
timestamp 1515178157
transform 1 0 6716 0 1 3808
box -38 -48 2246 592
use sky130_mm_sc_hd_dlyPoly5ns  clkgen.delay_155ns_2.genblk1\[2\].dly_binary.genblk1\[2\].delay_unit
timestamp 1515178157
transform 1 0 7544 0 -1 4896
box -38 -48 2246 592
use sky130_mm_sc_hd_dlyPoly5ns  clkgen.delay_155ns_2.genblk1\[2\].dly_binary.genblk1\[3\].delay_unit
timestamp 1515178157
transform 1 0 9936 0 1 3808
box -38 -48 2246 592
use sky130_fd_sc_hd__mux2_1  clkgen.delay_155ns_2.genblk1\[2\].dly_binary.out_mux
timestamp 1515178157
transform -1 0 5060 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  clkgen.delay_155ns_2.genblk1\[3\].bypass_enable
timestamp 1515178157
transform -1 0 22908 0 -1 4896
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  clkgen.delay_155ns_2.genblk1\[3\].control_invert
timestamp 1515178157
transform 1 0 21344 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  clkgen.delay_155ns_2.genblk1\[3\].dly_binary.and_bypass_switch
timestamp 1515178157
transform -1 0 17388 0 1 4896
box -38 -48 590 592
use sky130_mm_sc_hd_dlyPoly5ns  clkgen.delay_155ns_2.genblk1\[3\].dly_binary.genblk1\[0\].delay_unit
timestamp 1515178157
transform -1 0 6624 0 -1 5984
box -38 -48 2246 592
use sky130_mm_sc_hd_dlyPoly5ns  clkgen.delay_155ns_2.genblk1\[3\].dly_binary.genblk1\[1\].delay_unit
timestamp 1515178157
transform 1 0 7268 0 -1 5984
box -38 -48 2246 592
use sky130_mm_sc_hd_dlyPoly5ns  clkgen.delay_155ns_2.genblk1\[3\].dly_binary.genblk1\[2\].delay_unit
timestamp 1515178157
transform 1 0 9936 0 1 4896
box -38 -48 2246 592
use sky130_mm_sc_hd_dlyPoly5ns  clkgen.delay_155ns_2.genblk1\[3\].dly_binary.genblk1\[3\].delay_unit
timestamp 1515178157
transform 1 0 10120 0 -1 5984
box -38 -48 2246 592
use sky130_mm_sc_hd_dlyPoly5ns  clkgen.delay_155ns_2.genblk1\[3\].dly_binary.genblk1\[4\].delay_unit
timestamp 1515178157
transform 1 0 12972 0 1 4896
box -38 -48 2246 592
use sky130_mm_sc_hd_dlyPoly5ns  clkgen.delay_155ns_2.genblk1\[3\].dly_binary.genblk1\[5\].delay_unit
timestamp 1515178157
transform 1 0 14904 0 -1 3808
box -38 -48 2246 592
use sky130_mm_sc_hd_dlyPoly5ns  clkgen.delay_155ns_2.genblk1\[3\].dly_binary.genblk1\[6\].delay_unit
timestamp 1515178157
transform 1 0 15824 0 -1 4896
box -38 -48 2246 592
use sky130_mm_sc_hd_dlyPoly5ns  clkgen.delay_155ns_2.genblk1\[3\].dly_binary.genblk1\[7\].delay_unit
timestamp 1515178157
transform 1 0 17848 0 1 4896
box -38 -48 2246 592
use sky130_fd_sc_hd__mux2_1  clkgen.delay_155ns_2.genblk1\[3\].dly_binary.out_mux
timestamp 1515178157
transform -1 0 4048 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  clkgen.delay_155ns_2.genblk1\[4\].bypass_enable
timestamp 1515178157
transform -1 0 21528 0 -1 3808
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  clkgen.delay_155ns_2.genblk1\[4\].control_invert
timestamp 1515178157
transform -1 0 25944 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  clkgen.delay_155ns_2.genblk1\[4\].dly_binary.and_bypass_switch
timestamp 1515178157
transform -1 0 17112 0 1 5984
box -38 -48 590 592
use sky130_mm_sc_hd_dlyPoly5ns  clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[0\].delay_unit
timestamp 1515178157
transform -1 0 8004 0 1 4896
box -38 -48 2246 592
use sky130_mm_sc_hd_dlyPoly5ns  clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[1\].delay_unit
timestamp 1515178157
transform 1 0 7268 0 1 5984
box -38 -48 2246 592
use sky130_mm_sc_hd_dlyPoly5ns  clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[2\].delay_unit
timestamp 1515178157
transform 1 0 10396 0 1 5984
box -38 -48 2246 592
use sky130_mm_sc_hd_dlyPoly5ns  clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[3\].delay_unit
timestamp 1515178157
transform 1 0 12788 0 -1 5984
box -38 -48 2246 592
use sky130_mm_sc_hd_dlyPoly5ns  clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[4\].delay_unit
timestamp 1515178157
transform 1 0 12972 0 1 5984
box -38 -48 2246 592
use sky130_mm_sc_hd_dlyPoly5ns  clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[5\].delay_unit
timestamp 1515178157
transform 1 0 15824 0 -1 5984
box -38 -48 2246 592
use sky130_mm_sc_hd_dlyPoly5ns  clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[6\].delay_unit
timestamp 1515178157
transform 1 0 17940 0 1 5984
box -38 -48 2246 592
use sky130_mm_sc_hd_dlyPoly5ns  clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[7\].delay_unit
timestamp 1515178157
transform 1 0 19412 0 -1 5984
box -38 -48 2246 592
use sky130_mm_sc_hd_dlyPoly5ns  clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[8\].delay_unit
timestamp 1515178157
transform 1 0 21344 0 1 4896
box -38 -48 2246 592
use sky130_mm_sc_hd_dlyPoly5ns  clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[9\].delay_unit
timestamp 1515178157
transform 1 0 24196 0 -1 5984
box -38 -48 2246 592
use sky130_mm_sc_hd_dlyPoly5ns  clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[10\].delay_unit
timestamp 1515178157
transform -1 0 26128 0 1 4896
box -38 -48 2246 592
use sky130_mm_sc_hd_dlyPoly5ns  clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[11\].delay_unit
timestamp 1515178157
transform 1 0 24380 0 1 5984
box -38 -48 2246 592
use sky130_mm_sc_hd_dlyPoly5ns  clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[12\].delay_unit
timestamp 1515178157
transform 1 0 26772 0 -1 5984
box -38 -48 2246 592
use sky130_mm_sc_hd_dlyPoly5ns  clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[13\].delay_unit
timestamp 1515178157
transform -1 0 29256 0 1 4896
box -38 -48 2246 592
use sky130_mm_sc_hd_dlyPoly5ns  clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[14\].delay_unit
timestamp 1515178157
transform 1 0 28060 0 1 5984
box -38 -48 2246 592
use sky130_mm_sc_hd_dlyPoly5ns  clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[15\].delay_unit
timestamp 1515178157
transform 1 0 29900 0 -1 5984
box -38 -48 2246 592
use sky130_fd_sc_hd__mux2_1  clkgen.delay_155ns_2.genblk1\[4\].dly_binary.out_mux
timestamp 1515178157
transform 1 0 2944 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  clkgen.delay_155ns_3.enablebuffer
timestamp 1515178157
transform 1 0 18492 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  clkgen.delay_155ns_3.genblk1\[0\].bypass_enable
timestamp 1515178157
transform -1 0 20884 0 1 4896
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  clkgen.delay_155ns_3.genblk1\[0\].control_invert
timestamp 1515178157
transform 1 0 14812 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  clkgen.delay_155ns_3.genblk1\[0\].dly_binary.and_bypass_switch
timestamp 1515178157
transform -1 0 16192 0 1 5984
box -38 -48 590 592
use sky130_mm_sc_hd_dlyPoly5ns  clkgen.delay_155ns_3.genblk1\[0\].dly_binary.genblk1\[0\].delay_unit
timestamp 1515178157
transform -1 0 6440 0 1 5984
box -38 -48 2246 592
use sky130_fd_sc_hd__mux2_1  clkgen.delay_155ns_3.genblk1\[0\].dly_binary.out_mux
timestamp 1515178157
transform -1 0 5152 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  clkgen.delay_155ns_3.genblk1\[1\].bypass_enable
timestamp 1515178157
transform -1 0 12328 0 -1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  clkgen.delay_155ns_3.genblk1\[1\].control_invert
timestamp 1515178157
transform -1 0 20792 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  clkgen.delay_155ns_3.genblk1\[1\].dly_binary.and_bypass_switch
timestamp 1515178157
transform -1 0 13340 0 -1 8160
box -38 -48 590 592
use sky130_mm_sc_hd_dlyPoly5ns  clkgen.delay_155ns_3.genblk1\[1\].dly_binary.genblk1\[0\].delay_unit
timestamp 1515178157
transform -1 0 6624 0 -1 7072
box -38 -48 2246 592
use sky130_mm_sc_hd_dlyPoly5ns  clkgen.delay_155ns_3.genblk1\[1\].dly_binary.genblk1\[1\].delay_unit
timestamp 1515178157
transform 1 0 7084 0 -1 7072
box -38 -48 2246 592
use sky130_fd_sc_hd__mux2_1  clkgen.delay_155ns_3.genblk1\[1\].dly_binary.out_mux
timestamp 1515178157
transform -1 0 4048 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  clkgen.delay_155ns_3.genblk1\[2\].bypass_enable
timestamp 1515178157
transform -1 0 23644 0 -1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  clkgen.delay_155ns_3.genblk1\[2\].control_invert
timestamp 1515178157
transform 1 0 20608 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  clkgen.delay_155ns_3.genblk1\[2\].dly_binary.and_bypass_switch
timestamp 1515178157
transform -1 0 8832 0 -1 8160
box -38 -48 590 592
use sky130_mm_sc_hd_dlyPoly5ns  clkgen.delay_155ns_3.genblk1\[2\].dly_binary.genblk1\[0\].delay_unit
timestamp 1515178157
transform -1 0 6900 0 1 7072
box -38 -48 2246 592
use sky130_mm_sc_hd_dlyPoly5ns  clkgen.delay_155ns_3.genblk1\[2\].dly_binary.genblk1\[1\].delay_unit
timestamp 1515178157
transform 1 0 7268 0 1 7072
box -38 -48 2246 592
use sky130_mm_sc_hd_dlyPoly5ns  clkgen.delay_155ns_3.genblk1\[2\].dly_binary.genblk1\[2\].delay_unit
timestamp 1515178157
transform 1 0 9292 0 -1 8160
box -38 -48 2246 592
use sky130_mm_sc_hd_dlyPoly5ns  clkgen.delay_155ns_3.genblk1\[2\].dly_binary.genblk1\[3\].delay_unit
timestamp 1515178157
transform -1 0 12328 0 -1 7072
box -38 -48 2246 592
use sky130_fd_sc_hd__mux2_1  clkgen.delay_155ns_3.genblk1\[2\].dly_binary.out_mux
timestamp 1515178157
transform -1 0 7912 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  clkgen.delay_155ns_3.genblk1\[3\].bypass_enable
timestamp 1515178157
transform -1 0 22816 0 -1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  clkgen.delay_155ns_3.genblk1\[3\].control_invert
timestamp 1515178157
transform -1 0 25300 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  clkgen.delay_155ns_3.genblk1\[3\].dly_binary.and_bypass_switch
timestamp 1515178157
transform 1 0 10120 0 1 7072
box -38 -48 590 592
use sky130_mm_sc_hd_dlyPoly5ns  clkgen.delay_155ns_3.genblk1\[3\].dly_binary.genblk1\[0\].delay_unit
timestamp 1515178157
transform 1 0 12788 0 -1 7072
box -38 -48 2246 592
use sky130_mm_sc_hd_dlyPoly5ns  clkgen.delay_155ns_3.genblk1\[3\].dly_binary.genblk1\[1\].delay_unit
timestamp 1515178157
transform 1 0 13708 0 -1 8160
box -38 -48 2246 592
use sky130_mm_sc_hd_dlyPoly5ns  clkgen.delay_155ns_3.genblk1\[3\].dly_binary.genblk1\[2\].delay_unit
timestamp 1515178157
transform 1 0 15364 0 -1 7072
box -38 -48 2246 592
use sky130_mm_sc_hd_dlyPoly5ns  clkgen.delay_155ns_3.genblk1\[3\].dly_binary.genblk1\[3\].delay_unit
timestamp 1515178157
transform 1 0 17020 0 1 7072
box -38 -48 2246 592
use sky130_mm_sc_hd_dlyPoly5ns  clkgen.delay_155ns_3.genblk1\[3\].dly_binary.genblk1\[4\].delay_unit
timestamp 1515178157
transform 1 0 18492 0 -1 7072
box -38 -48 2246 592
use sky130_mm_sc_hd_dlyPoly5ns  clkgen.delay_155ns_3.genblk1\[3\].dly_binary.genblk1\[5\].delay_unit
timestamp 1515178157
transform 1 0 21068 0 -1 7072
box -38 -48 2246 592
use sky130_mm_sc_hd_dlyPoly5ns  clkgen.delay_155ns_3.genblk1\[3\].dly_binary.genblk1\[6\].delay_unit
timestamp 1515178157
transform 1 0 21344 0 1 5984
box -38 -48 2246 592
use sky130_mm_sc_hd_dlyPoly5ns  clkgen.delay_155ns_3.genblk1\[3\].dly_binary.genblk1\[7\].delay_unit
timestamp 1515178157
transform -1 0 24748 0 1 7072
box -38 -48 2246 592
use sky130_fd_sc_hd__mux2_1  clkgen.delay_155ns_3.genblk1\[3\].dly_binary.out_mux
timestamp 1515178157
transform -1 0 11868 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  clkgen.delay_155ns_3.genblk1\[4\].bypass_enable
timestamp 1515178157
transform -1 0 23368 0 -1 5984
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  clkgen.delay_155ns_3.genblk1\[4\].control_invert
timestamp 1515178157
transform 1 0 14904 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  clkgen.delay_155ns_3.genblk1\[4\].dly_binary.and_bypass_switch
timestamp 1515178157
transform -1 0 12236 0 -1 3808
box -38 -48 590 592
use sky130_mm_sc_hd_dlyPoly5ns  clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[0\].delay_unit
timestamp 1515178157
transform 1 0 10120 0 -1 4896
box -38 -48 2246 592
use sky130_mm_sc_hd_dlyPoly5ns  clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[1\].delay_unit
timestamp 1515178157
transform 1 0 13248 0 -1 4896
box -38 -48 2246 592
use sky130_mm_sc_hd_dlyPoly5ns  clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[2\].delay_unit
timestamp 1515178157
transform -1 0 15180 0 1 3808
box -38 -48 2246 592
use sky130_mm_sc_hd_dlyPoly5ns  clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[3\].delay_unit
timestamp 1515178157
transform 1 0 16100 0 1 3808
box -38 -48 2246 592
use sky130_mm_sc_hd_dlyPoly5ns  clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[4\].delay_unit
timestamp 1515178157
transform 1 0 17388 0 1 2720
box -38 -48 2246 592
use sky130_mm_sc_hd_dlyPoly5ns  clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[5\].delay_unit
timestamp 1515178157
transform 1 0 18676 0 1 3808
box -38 -48 2246 592
use sky130_mm_sc_hd_dlyPoly5ns  clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[6\].delay_unit
timestamp 1515178157
transform 1 0 19872 0 -1 4896
box -38 -48 2246 592
use sky130_mm_sc_hd_dlyPoly5ns  clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[7\].delay_unit
timestamp 1515178157
transform 1 0 21344 0 1 3808
box -38 -48 2246 592
use sky130_mm_sc_hd_dlyPoly5ns  clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[8\].delay_unit
timestamp 1515178157
transform 1 0 24196 0 -1 4896
box -38 -48 2246 592
use sky130_mm_sc_hd_dlyPoly5ns  clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[9\].delay_unit
timestamp 1515178157
transform -1 0 26128 0 1 3808
box -38 -48 2246 592
use sky130_mm_sc_hd_dlyPoly5ns  clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[10\].delay_unit
timestamp 1515178157
transform 1 0 24472 0 -1 3808
box -38 -48 2246 592
use sky130_mm_sc_hd_dlyPoly5ns  clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[11\].delay_unit
timestamp 1515178157
transform 1 0 26772 0 -1 4896
box -38 -48 2246 592
use sky130_mm_sc_hd_dlyPoly5ns  clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[12\].delay_unit
timestamp 1515178157
transform 1 0 27048 0 1 3808
box -38 -48 2246 592
use sky130_mm_sc_hd_dlyPoly5ns  clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[13\].delay_unit
timestamp 1515178157
transform 1 0 29900 0 -1 4896
box -38 -48 2246 592
use sky130_mm_sc_hd_dlyPoly5ns  clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[14\].delay_unit
timestamp 1515178157
transform -1 0 31832 0 1 3808
box -38 -48 2246 592
use sky130_mm_sc_hd_dlyPoly5ns  clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[15\].delay_unit
timestamp 1515178157
transform -1 0 32292 0 1 4896
box -38 -48 2246 592
use sky130_fd_sc_hd__mux2_1  clkgen.delay_155ns_3.genblk1\[4\].dly_binary.out_mux
timestamp 1515178157
transform 1 0 15640 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__nor2b_1  clkgen.nor1
timestamp 1515178157
transform 1 0 1564 0 1 4896
box -38 -48 498 592
use sky130_mm_sc_hd_dlyPoly5ns  delay_sample_n12
timestamp 1515178157
transform 1 0 1564 0 1 2720
box -38 -48 2246 592
use sky130_mm_sc_hd_dlyPoly5ns  delay_sample_p11
timestamp 1515178157
transform -1 0 3772 0 -1 9248
box -38 -48 2246 592
use sky130_fd_sc_hd__buf_4  edgedetect.dly_315ns_1.enablebuffer
timestamp 1515178157
transform 1 0 15640 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  edgedetect.dly_315ns_1.genblk1\[0\].bypass_enable
timestamp 1515178157
transform 1 0 24196 0 -1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  edgedetect.dly_315ns_1.genblk1\[0\].control_invert
timestamp 1515178157
transform -1 0 26220 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  edgedetect.dly_315ns_1.genblk1\[0\].dly_binary.and_bypass_switch
timestamp 1515178157
transform -1 0 18032 0 -1 8160
box -38 -48 590 592
use sky130_mm_sc_hd_dlyPoly5ns  edgedetect.dly_315ns_1.genblk1\[0\].dly_binary.genblk1\[0\].delay_unit
timestamp 1515178157
transform -1 0 3956 0 -1 8160
box -38 -48 2246 592
use sky130_fd_sc_hd__mux2_1  edgedetect.dly_315ns_1.genblk1\[0\].dly_binary.out_mux
timestamp 1515178157
transform -1 0 2852 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  edgedetect.dly_315ns_1.genblk1\[1\].bypass_enable
timestamp 1515178157
transform -1 0 23736 0 -1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  edgedetect.dly_315ns_1.genblk1\[1\].control_invert
timestamp 1515178157
transform -1 0 27876 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  edgedetect.dly_315ns_1.genblk1\[1\].dly_binary.and_bypass_switch
timestamp 1515178157
transform -1 0 19044 0 -1 8160
box -38 -48 590 592
use sky130_mm_sc_hd_dlyPoly5ns  edgedetect.dly_315ns_1.genblk1\[1\].dly_binary.genblk1\[0\].delay_unit
timestamp 1515178157
transform -1 0 3772 0 1 8160
box -38 -48 2246 592
use sky130_mm_sc_hd_dlyPoly5ns  edgedetect.dly_315ns_1.genblk1\[1\].dly_binary.genblk1\[1\].delay_unit
timestamp 1515178157
transform 1 0 4324 0 -1 8160
box -38 -48 2246 592
use sky130_fd_sc_hd__mux2_1  edgedetect.dly_315ns_1.genblk1\[1\].dly_binary.out_mux
timestamp 1515178157
transform -1 0 7912 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  edgedetect.dly_315ns_1.genblk1\[2\].bypass_enable
timestamp 1515178157
transform -1 0 24656 0 -1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  edgedetect.dly_315ns_1.genblk1\[2\].control_invert
timestamp 1515178157
transform -1 0 27048 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.and_bypass_switch
timestamp 1515178157
transform -1 0 20240 0 1 9248
box -38 -48 590 592
use sky130_mm_sc_hd_dlyPoly5ns  edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.genblk1\[0\].delay_unit
timestamp 1515178157
transform -1 0 3772 0 1 9248
box -38 -48 2246 592
use sky130_mm_sc_hd_dlyPoly5ns  edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.genblk1\[1\].delay_unit
timestamp 1515178157
transform 1 0 4692 0 1 9248
box -38 -48 2246 592
use sky130_mm_sc_hd_dlyPoly5ns  edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.genblk1\[2\].delay_unit
timestamp 1515178157
transform 1 0 7544 0 -1 10336
box -38 -48 2246 592
use sky130_mm_sc_hd_dlyPoly5ns  edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.genblk1\[3\].delay_unit
timestamp 1515178157
transform 1 0 9936 0 -1 11424
box -38 -48 2246 592
use sky130_fd_sc_hd__mux2_1  edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.out_mux
timestamp 1515178157
transform -1 0 9108 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  edgedetect.dly_315ns_1.genblk1\[3\].bypass_enable
timestamp 1515178157
transform -1 0 25484 0 -1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  edgedetect.dly_315ns_1.genblk1\[3\].control_invert
timestamp 1515178157
transform -1 0 27324 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.and_bypass_switch
timestamp 1515178157
transform -1 0 22908 0 -1 10336
box -38 -48 590 592
use sky130_mm_sc_hd_dlyPoly5ns  edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.genblk1\[0\].delay_unit
timestamp 1515178157
transform -1 0 4048 0 -1 10336
box -38 -48 2246 592
use sky130_mm_sc_hd_dlyPoly5ns  edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.genblk1\[1\].delay_unit
timestamp 1515178157
transform 1 0 4416 0 -1 10336
box -38 -48 2246 592
use sky130_mm_sc_hd_dlyPoly5ns  edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.genblk1\[2\].delay_unit
timestamp 1515178157
transform 1 0 7268 0 1 9248
box -38 -48 2246 592
use sky130_mm_sc_hd_dlyPoly5ns  edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.genblk1\[3\].delay_unit
timestamp 1515178157
transform 1 0 10396 0 1 9248
box -38 -48 2246 592
use sky130_mm_sc_hd_dlyPoly5ns  edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.genblk1\[4\].delay_unit
timestamp 1515178157
transform 1 0 12788 0 -1 11424
box -38 -48 2246 592
use sky130_mm_sc_hd_dlyPoly5ns  edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.genblk1\[5\].delay_unit
timestamp 1515178157
transform 1 0 12972 0 1 9248
box -38 -48 2246 592
use sky130_mm_sc_hd_dlyPoly5ns  edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.genblk1\[6\].delay_unit
timestamp 1515178157
transform 1 0 15640 0 -1 11424
box -38 -48 2246 592
use sky130_mm_sc_hd_dlyPoly5ns  edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.genblk1\[7\].delay_unit
timestamp 1515178157
transform 1 0 15824 0 -1 10336
box -38 -48 2246 592
use sky130_fd_sc_hd__mux2_1  edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.out_mux
timestamp 1515178157
transform -1 0 19320 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  edgedetect.dly_315ns_1.genblk1\[4\].bypass_enable
timestamp 1515178157
transform -1 0 26312 0 -1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  edgedetect.dly_315ns_1.genblk1\[4\].control_invert
timestamp 1515178157
transform -1 0 27968 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.and_bypass_switch
timestamp 1515178157
transform -1 0 21896 0 1 7072
box -38 -48 590 592
use sky130_mm_sc_hd_dlyPoly5ns  edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[0\].delay_unit
timestamp 1515178157
transform -1 0 3772 0 -1 11424
box -38 -48 2246 592
use sky130_mm_sc_hd_dlyPoly5ns  edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[1\].delay_unit
timestamp 1515178157
transform 1 0 1564 0 1 10336
box -38 -48 2246 592
use sky130_mm_sc_hd_dlyPoly5ns  edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[2\].delay_unit
timestamp 1515178157
transform 1 0 4692 0 1 10336
box -38 -48 2246 592
use sky130_mm_sc_hd_dlyPoly5ns  edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[3\].delay_unit
timestamp 1515178157
transform -1 0 6624 0 -1 11424
box -38 -48 2246 592
use sky130_mm_sc_hd_dlyPoly5ns  edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[4\].delay_unit
timestamp 1515178157
transform 1 0 7268 0 -1 11424
box -38 -48 2246 592
use sky130_mm_sc_hd_dlyPoly5ns  edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[5\].delay_unit
timestamp 1515178157
transform -1 0 9476 0 1 10336
box -38 -48 2246 592
use sky130_mm_sc_hd_dlyPoly5ns  edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[6\].delay_unit
timestamp 1515178157
transform 1 0 10120 0 -1 10336
box -38 -48 2246 592
use sky130_mm_sc_hd_dlyPoly5ns  edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[7\].delay_unit
timestamp 1515178157
transform 1 0 10396 0 1 10336
box -38 -48 2246 592
use sky130_mm_sc_hd_dlyPoly5ns  edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[8\].delay_unit
timestamp 1515178157
transform 1 0 13248 0 -1 10336
box -38 -48 2246 592
use sky130_mm_sc_hd_dlyPoly5ns  edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[9\].delay_unit
timestamp 1515178157
transform -1 0 15180 0 1 10336
box -38 -48 2246 592
use sky130_mm_sc_hd_dlyPoly5ns  edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[10\].delay_unit
timestamp 1515178157
transform 1 0 18492 0 -1 11424
box -38 -48 2246 592
use sky130_mm_sc_hd_dlyPoly5ns  edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[11\].delay_unit
timestamp 1515178157
transform -1 0 18124 0 1 10336
box -38 -48 2246 592
use sky130_mm_sc_hd_dlyPoly5ns  edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[12\].delay_unit
timestamp 1515178157
transform 1 0 18492 0 1 10336
box -38 -48 2246 592
use sky130_mm_sc_hd_dlyPoly5ns  edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[13\].delay_unit
timestamp 1515178157
transform 1 0 21344 0 1 10336
box -38 -48 2246 592
use sky130_mm_sc_hd_dlyPoly5ns  edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[14\].delay_unit
timestamp 1515178157
transform -1 0 23552 0 -1 11424
box -38 -48 2246 592
use sky130_mm_sc_hd_dlyPoly5ns  edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[15\].delay_unit
timestamp 1515178157
transform 1 0 23920 0 1 10336
box -38 -48 2246 592
use sky130_fd_sc_hd__mux2_1  edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.out_mux
timestamp 1515178157
transform 1 0 16284 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  edgedetect.dly_315ns_1.genblk1\[5\].bypass_enable
timestamp 1515178157
transform -1 0 25576 0 1 7072
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  edgedetect.dly_315ns_1.genblk1\[5\].control_invert
timestamp 1515178157
transform -1 0 28520 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.and_bypass_switch
timestamp 1515178157
transform -1 0 20148 0 1 7072
box -38 -48 590 592
use sky130_mm_sc_hd_dlyPoly5ns  edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[0\].delay_unit
timestamp 1515178157
transform -1 0 6532 0 -1 9248
box -38 -48 2246 592
use sky130_mm_sc_hd_dlyPoly5ns  edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[1\].delay_unit
timestamp 1515178157
transform 1 0 4692 0 1 8160
box -38 -48 2246 592
use sky130_mm_sc_hd_dlyPoly5ns  edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[2\].delay_unit
timestamp 1515178157
transform 1 0 7268 0 1 8160
box -38 -48 2246 592
use sky130_mm_sc_hd_dlyPoly5ns  edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[3\].delay_unit
timestamp 1515178157
transform 1 0 9568 0 -1 9248
box -38 -48 2246 592
use sky130_mm_sc_hd_dlyPoly5ns  edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[4\].delay_unit
timestamp 1515178157
transform 1 0 10396 0 1 8160
box -38 -48 2246 592
use sky130_mm_sc_hd_dlyPoly5ns  edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[5\].delay_unit
timestamp 1515178157
transform 1 0 12236 0 1 7072
box -38 -48 2246 592
use sky130_mm_sc_hd_dlyPoly5ns  edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[6\].delay_unit
timestamp 1515178157
transform 1 0 13248 0 -1 9248
box -38 -48 2246 592
use sky130_mm_sc_hd_dlyPoly5ns  edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[7\].delay_unit
timestamp 1515178157
transform -1 0 15180 0 1 8160
box -38 -48 2246 592
use sky130_mm_sc_hd_dlyPoly5ns  edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[8\].delay_unit
timestamp 1515178157
transform 1 0 15916 0 1 8160
box -38 -48 2246 592
use sky130_mm_sc_hd_dlyPoly5ns  edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[9\].delay_unit
timestamp 1515178157
transform 1 0 17112 0 1 9248
box -38 -48 2246 592
use sky130_mm_sc_hd_dlyPoly5ns  edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[10\].delay_unit
timestamp 1515178157
transform 1 0 18492 0 1 8160
box -38 -48 2246 592
use sky130_mm_sc_hd_dlyPoly5ns  edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[11\].delay_unit
timestamp 1515178157
transform 1 0 19780 0 -1 8160
box -38 -48 2246 592
use sky130_mm_sc_hd_dlyPoly5ns  edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[12\].delay_unit
timestamp 1515178157
transform 1 0 21344 0 1 8160
box -38 -48 2246 592
use sky130_mm_sc_hd_dlyPoly5ns  edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[13\].delay_unit
timestamp 1515178157
transform 1 0 23920 0 1 8160
box -38 -48 2246 592
use sky130_mm_sc_hd_dlyPoly5ns  edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[14\].delay_unit
timestamp 1515178157
transform -1 0 26404 0 -1 8160
box -38 -48 2246 592
use sky130_mm_sc_hd_dlyPoly5ns  edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[15\].delay_unit
timestamp 1515178157
transform 1 0 25024 0 -1 9248
box -38 -48 2246 592
use sky130_mm_sc_hd_dlyPoly5ns  edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[16\].delay_unit
timestamp 1515178157
transform 1 0 27048 0 1 8160
box -38 -48 2246 592
use sky130_mm_sc_hd_dlyPoly5ns  edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[17\].delay_unit
timestamp 1515178157
transform -1 0 18032 0 -1 9248
box -38 -48 2246 592
use sky130_mm_sc_hd_dlyPoly5ns  edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[18\].delay_unit
timestamp 1515178157
transform 1 0 18768 0 -1 9248
box -38 -48 2246 592
use sky130_mm_sc_hd_dlyPoly5ns  edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[19\].delay_unit
timestamp 1515178157
transform 1 0 19780 0 -1 10336
box -38 -48 2246 592
use sky130_mm_sc_hd_dlyPoly5ns  edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[20\].delay_unit
timestamp 1515178157
transform 1 0 21344 0 1 9248
box -38 -48 2246 592
use sky130_mm_sc_hd_dlyPoly5ns  edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[21\].delay_unit
timestamp 1515178157
transform 1 0 21528 0 -1 9248
box -38 -48 2246 592
use sky130_mm_sc_hd_dlyPoly5ns  edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[22\].delay_unit
timestamp 1515178157
transform 1 0 24196 0 -1 10336
box -38 -48 2246 592
use sky130_mm_sc_hd_dlyPoly5ns  edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[23\].delay_unit
timestamp 1515178157
transform 1 0 24380 0 1 9248
box -38 -48 2246 592
use sky130_mm_sc_hd_dlyPoly5ns  edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[24\].delay_unit
timestamp 1515178157
transform 1 0 26772 0 -1 10336
box -38 -48 2246 592
use sky130_mm_sc_hd_dlyPoly5ns  edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[25\].delay_unit
timestamp 1515178157
transform 1 0 27600 0 1 10336
box -38 -48 2246 592
use sky130_mm_sc_hd_dlyPoly5ns  edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[26\].delay_unit
timestamp 1515178157
transform 1 0 29900 0 -1 10336
box -38 -48 2246 592
use sky130_mm_sc_hd_dlyPoly5ns  edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[27\].delay_unit
timestamp 1515178157
transform -1 0 32568 0 -1 8160
box -38 -48 2246 592
use sky130_mm_sc_hd_dlyPoly5ns  edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[28\].delay_unit
timestamp 1515178157
transform -1 0 29256 0 1 9248
box -38 -48 2246 592
use sky130_mm_sc_hd_dlyPoly5ns  edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[29\].delay_unit
timestamp 1515178157
transform 1 0 29624 0 1 9248
box -38 -48 2246 592
use sky130_mm_sc_hd_dlyPoly5ns  edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[30\].delay_unit
timestamp 1515178157
transform 1 0 29900 0 -1 9248
box -38 -48 2246 592
use sky130_mm_sc_hd_dlyPoly5ns  edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[31\].delay_unit
timestamp 1515178157
transform -1 0 32292 0 1 8160
box -38 -48 2246 592
use sky130_fd_sc_hd__mux2_1  edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.out_mux
timestamp 1515178157
transform -1 0 16468 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__nor2b_1  edgedetect.nor1
timestamp 1515178157
transform 1 0 24196 0 -1 7072
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  edgedetect.or1
timestamp 1515178157
transform -1 0 2024 0 1 7072
box -38 -48 498 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3
timestamp 1515178157
transform 1 0 1380 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29
timestamp 1515178157
transform 1 0 3772 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32
timestamp 1515178157
transform 1 0 4048 0 1 544
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_60
timestamp 1515178157
transform 1 0 6624 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_63
timestamp 1515178157
transform 1 0 6900 0 1 544
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_91
timestamp 1515178157
transform 1 0 9476 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_94
timestamp 1515178157
transform 1 0 9752 0 1 544
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_122
timestamp 1515178157
transform 1 0 12328 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_125
timestamp 1515178157
transform 1 0 12604 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_136
timestamp 1515178157
transform 1 0 13616 0 1 544
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_146
timestamp 1515178157
transform 1 0 14536 0 1 544
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_153
timestamp 1515178157
transform 1 0 15180 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_156
timestamp 1515178157
transform 1 0 15456 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_182
timestamp 1515178157
transform 1 0 17848 0 1 544
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_187
timestamp 1515178157
transform 1 0 18308 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_194
timestamp 1515178157
transform 1 0 18952 0 1 544
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_203
timestamp 1515178157
transform 1 0 19780 0 1 544
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_210
timestamp 1515178157
transform 1 0 20424 0 1 544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_216
timestamp 1515178157
transform 1 0 20976 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_218
timestamp 1515178157
transform 1 0 21160 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_223
timestamp 1515178157
transform 1 0 21620 0 1 544
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_229
timestamp 1515178157
transform 1 0 22172 0 1 544
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_235
timestamp 1515178157
transform 1 0 22724 0 1 544
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_241
timestamp 1515178157
transform 1 0 23276 0 1 544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_247
timestamp 1515178157
transform 1 0 23828 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_249
timestamp 1515178157
transform 1 0 24012 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_253
timestamp 1515178157
transform 1 0 24380 0 1 544
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_259
timestamp 1515178157
transform 1 0 24932 0 1 544
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_265
timestamp 1515178157
transform 1 0 25484 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_277
timestamp 1515178157
transform 1 0 26588 0 1 544
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_280
timestamp 1515178157
transform 1 0 26864 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_292
timestamp 1515178157
transform 1 0 27968 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_304
timestamp 1515178157
transform 1 0 29072 0 1 544
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_311
timestamp 1515178157
transform 1 0 29716 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_323
timestamp 1515178157
transform 1 0 30820 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_335
timestamp 1515178157
transform 1 0 31924 0 1 544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_342
timestamp 1515178157
transform 1 0 32568 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_3
timestamp 1515178157
transform 1 0 1380 0 -1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_7
timestamp 1515178157
transform 1 0 1748 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_32
timestamp 1515178157
transform 1 0 4048 0 -1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_60
timestamp 1515178157
transform 1 0 6624 0 -1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_1_63
timestamp 1515178157
transform 1 0 6900 0 -1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_69
timestamp 1515178157
transform 1 0 7452 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_94
timestamp 1515178157
transform 1 0 9752 0 -1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_122
timestamp 1515178157
transform 1 0 12328 0 -1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_125
timestamp 1515178157
transform 1 0 12604 0 -1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_153
timestamp 1515178157
transform 1 0 15180 0 -1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_159
timestamp 1515178157
transform 1 0 15732 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_184
timestamp 1515178157
transform 1 0 18032 0 -1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_1_187
timestamp 1515178157
transform 1 0 18308 0 -1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_193
timestamp 1515178157
transform 1 0 18860 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_218
timestamp 1515178157
transform 1 0 21160 0 -1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_225
timestamp 1515178157
transform 1 0 21804 0 -1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_231
timestamp 1515178157
transform 1 0 22356 0 -1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_237
timestamp 1515178157
transform 1 0 22908 0 -1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_243
timestamp 1515178157
transform 1 0 23460 0 -1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_247
timestamp 1515178157
transform 1 0 23828 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_249
timestamp 1515178157
transform 1 0 24012 0 -1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_253
timestamp 1515178157
transform 1 0 24380 0 -1 1632
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_259
timestamp 1515178157
transform 1 0 24932 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_271
timestamp 1515178157
transform 1 0 26036 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_283
timestamp 1515178157
transform 1 0 27140 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_295
timestamp 1515178157
transform 1 0 28244 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_1_307
timestamp 1515178157
transform 1 0 29348 0 -1 1632
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_1_311
timestamp 1515178157
transform 1 0 29716 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_323
timestamp 1515178157
transform 1 0 30820 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_335
timestamp 1515178157
transform 1 0 31924 0 -1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_343
timestamp 1515178157
transform 1 0 32660 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_3
timestamp 1515178157
transform 1 0 1380 0 1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_29
timestamp 1515178157
transform 1 0 3772 0 1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_2_32
timestamp 1515178157
transform 1 0 4048 0 1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_38
timestamp 1515178157
transform 1 0 4600 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_63
timestamp 1515178157
transform 1 0 6900 0 1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_91
timestamp 1515178157
transform 1 0 9476 0 1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_2_94
timestamp 1515178157
transform 1 0 9752 0 1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_100
timestamp 1515178157
transform 1 0 10304 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_125
timestamp 1515178157
transform 1 0 12604 0 1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_153
timestamp 1515178157
transform 1 0 15180 0 1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_156
timestamp 1515178157
transform 1 0 15456 0 1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_164
timestamp 1515178157
transform 1 0 16192 0 1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_174
timestamp 1515178157
transform 1 0 17112 0 1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_2_206
timestamp 1515178157
transform 1 0 20056 0 1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_215
timestamp 1515178157
transform 1 0 20884 0 1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_218
timestamp 1515178157
transform 1 0 21160 0 1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_223
timestamp 1515178157
transform 1 0 21620 0 1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_230
timestamp 1515178157
transform 1 0 22264 0 1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_237
timestamp 1515178157
transform 1 0 22908 0 1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_243
timestamp 1515178157
transform 1 0 23460 0 1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_249
timestamp 1515178157
transform 1 0 24012 0 1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_255
timestamp 1515178157
transform 1 0 24564 0 1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_261
timestamp 1515178157
transform 1 0 25116 0 1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_267
timestamp 1515178157
transform 1 0 25668 0 1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_273
timestamp 1515178157
transform 1 0 26220 0 1 1632
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_2_280
timestamp 1515178157
transform 1 0 26864 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_292
timestamp 1515178157
transform 1 0 27968 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_304
timestamp 1515178157
transform 1 0 29072 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_316
timestamp 1515178157
transform 1 0 30176 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_328
timestamp 1515178157
transform 1 0 31280 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_340
timestamp 1515178157
transform 1 0 32384 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_342
timestamp 1515178157
transform 1 0 32568 0 1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_3
timestamp 1515178157
transform 1 0 1380 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_3_30
timestamp 1515178157
transform 1 0 3864 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_3_60
timestamp 1515178157
transform 1 0 6624 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_3_63
timestamp 1515178157
transform 1 0 6900 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_69
timestamp 1515178157
transform 1 0 7452 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_94
timestamp 1515178157
transform 1 0 9752 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_122
timestamp 1515178157
transform 1 0 12328 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_125
timestamp 1515178157
transform 1 0 12604 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_3_151
timestamp 1515178157
transform 1 0 14996 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_3_181
timestamp 1515178157
transform 1 0 17756 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_185
timestamp 1515178157
transform 1 0 18124 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_187
timestamp 1515178157
transform 1 0 18308 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_213
timestamp 1515178157
transform 1 0 20700 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_223
timestamp 1515178157
transform 1 0 21620 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_232
timestamp 1515178157
transform 1 0 22448 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_239
timestamp 1515178157
transform 1 0 23092 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_246
timestamp 1515178157
transform 1 0 23736 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_249
timestamp 1515178157
transform 1 0 24012 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_253
timestamp 1515178157
transform 1 0 24380 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_259
timestamp 1515178157
transform 1 0 24932 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_265
timestamp 1515178157
transform 1 0 25484 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_271
timestamp 1515178157
transform 1 0 26036 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_277
timestamp 1515178157
transform 1 0 26588 0 -1 2720
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_3_283
timestamp 1515178157
transform 1 0 27140 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_295
timestamp 1515178157
transform 1 0 28244 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_3_307
timestamp 1515178157
transform 1 0 29348 0 -1 2720
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_3_311
timestamp 1515178157
transform 1 0 29716 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_323
timestamp 1515178157
transform 1 0 30820 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_335
timestamp 1515178157
transform 1 0 31924 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_343
timestamp 1515178157
transform 1 0 32660 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_3
timestamp 1515178157
transform 1 0 1380 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_29
timestamp 1515178157
transform 1 0 3772 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_4_32
timestamp 1515178157
transform 1 0 4048 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_38
timestamp 1515178157
transform 1 0 4600 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_63
timestamp 1515178157
transform 1 0 6900 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_91
timestamp 1515178157
transform 1 0 9476 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_4_94
timestamp 1515178157
transform 1 0 9752 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_100
timestamp 1515178157
transform 1 0 10304 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_125
timestamp 1515178157
transform 1 0 12604 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_153
timestamp 1515178157
transform 1 0 15180 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_156
timestamp 1515178157
transform 1 0 15456 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_167
timestamp 1515178157
transform 1 0 16468 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_173
timestamp 1515178157
transform 1 0 17020 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_201
timestamp 1515178157
transform 1 0 19596 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_4_211
timestamp 1515178157
transform 1 0 20516 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_4_218
timestamp 1515178157
transform 1 0 21160 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_226
timestamp 1515178157
transform 1 0 21896 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_235
timestamp 1515178157
transform 1 0 22724 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_242
timestamp 1515178157
transform 1 0 23368 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_249
timestamp 1515178157
transform 1 0 24012 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_256
timestamp 1515178157
transform 1 0 24656 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_262
timestamp 1515178157
transform 1 0 25208 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_268
timestamp 1515178157
transform 1 0 25760 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_274
timestamp 1515178157
transform 1 0 26312 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_278
timestamp 1515178157
transform 1 0 26680 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_280
timestamp 1515178157
transform 1 0 26864 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_284
timestamp 1515178157
transform 1 0 27232 0 1 2720
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_4_290
timestamp 1515178157
transform 1 0 27784 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_302
timestamp 1515178157
transform 1 0 28888 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_314
timestamp 1515178157
transform 1 0 29992 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_326
timestamp 1515178157
transform 1 0 31096 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_338
timestamp 1515178157
transform 1 0 32200 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_342
timestamp 1515178157
transform 1 0 32568 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_3
timestamp 1515178157
transform 1 0 1380 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_13
timestamp 1515178157
transform 1 0 2300 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_32
timestamp 1515178157
transform 1 0 4048 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_60
timestamp 1515178157
transform 1 0 6624 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_63
timestamp 1515178157
transform 1 0 6900 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_68
timestamp 1515178157
transform 1 0 7360 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_81
timestamp 1515178157
transform 1 0 8556 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_85
timestamp 1515178157
transform 1 0 8924 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_110
timestamp 1515178157
transform 1 0 11224 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_114
timestamp 1515178157
transform 1 0 11592 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_5_121
timestamp 1515178157
transform 1 0 12236 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_125
timestamp 1515178157
transform 1 0 12604 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_5_142
timestamp 1515178157
transform 1 0 14168 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_5_174
timestamp 1515178157
transform 1 0 17112 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_184
timestamp 1515178157
transform 1 0 18032 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_187
timestamp 1515178157
transform 1 0 18308 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_213
timestamp 1515178157
transform 1 0 20700 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_222
timestamp 1515178157
transform 1 0 21528 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_231
timestamp 1515178157
transform 1 0 22356 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_240
timestamp 1515178157
transform 1 0 23184 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_246
timestamp 1515178157
transform 1 0 23736 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_249
timestamp 1515178157
transform 1 0 24012 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_253
timestamp 1515178157
transform 1 0 24380 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_278
timestamp 1515178157
transform 1 0 26680 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_284
timestamp 1515178157
transform 1 0 27232 0 -1 3808
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_5_290
timestamp 1515178157
transform 1 0 27784 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_302
timestamp 1515178157
transform 1 0 28888 0 -1 3808
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_5_311
timestamp 1515178157
transform 1 0 29716 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_323
timestamp 1515178157
transform 1 0 30820 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_335
timestamp 1515178157
transform 1 0 31924 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_343
timestamp 1515178157
transform 1 0 32660 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_3
timestamp 1515178157
transform 1 0 1380 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_29
timestamp 1515178157
transform 1 0 3772 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_32
timestamp 1515178157
transform 1 0 4048 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_43
timestamp 1515178157
transform 1 0 5060 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_47
timestamp 1515178157
transform 1 0 5428 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_57
timestamp 1515178157
transform 1 0 6348 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_85
timestamp 1515178157
transform 1 0 8924 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_91
timestamp 1515178157
transform 1 0 9476 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_94
timestamp 1515178157
transform 1 0 9752 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_6_120
timestamp 1515178157
transform 1 0 12144 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_128
timestamp 1515178157
transform 1 0 12880 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_153
timestamp 1515178157
transform 1 0 15180 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_6_156
timestamp 1515178157
transform 1 0 15456 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_162
timestamp 1515178157
transform 1 0 16008 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_187
timestamp 1515178157
transform 1 0 18308 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_215
timestamp 1515178157
transform 1 0 20884 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_218
timestamp 1515178157
transform 1 0 21160 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_244
timestamp 1515178157
transform 1 0 23552 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_6_272
timestamp 1515178157
transform 1 0 26128 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_278
timestamp 1515178157
transform 1 0 26680 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_280
timestamp 1515178157
transform 1 0 26864 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_306
timestamp 1515178157
transform 1 0 29256 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_6_334
timestamp 1515178157
transform 1 0 31832 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_340
timestamp 1515178157
transform 1 0 32384 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_342
timestamp 1515178157
transform 1 0 32568 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_3
timestamp 1515178157
transform 1 0 1380 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_7
timestamp 1515178157
transform 1 0 1748 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_32
timestamp 1515178157
transform 1 0 4048 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_60
timestamp 1515178157
transform 1 0 6624 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_7_63
timestamp 1515178157
transform 1 0 6900 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_69
timestamp 1515178157
transform 1 0 7452 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_94
timestamp 1515178157
transform 1 0 9752 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_122
timestamp 1515178157
transform 1 0 12328 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_7_125
timestamp 1515178157
transform 1 0 12604 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_131
timestamp 1515178157
transform 1 0 13156 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_156
timestamp 1515178157
transform 1 0 15456 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_184
timestamp 1515178157
transform 1 0 18032 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_187
timestamp 1515178157
transform 1 0 18308 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_7_195
timestamp 1515178157
transform 1 0 19044 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_203
timestamp 1515178157
transform 1 0 19780 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_228
timestamp 1515178157
transform 1 0 22080 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_237
timestamp 1515178157
transform 1 0 22908 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_246
timestamp 1515178157
transform 1 0 23736 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_249
timestamp 1515178157
transform 1 0 24012 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_275
timestamp 1515178157
transform 1 0 26404 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_7_303
timestamp 1515178157
transform 1 0 28980 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_309
timestamp 1515178157
transform 1 0 29532 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_311
timestamp 1515178157
transform 1 0 29716 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_7_337
timestamp 1515178157
transform 1 0 32108 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_343
timestamp 1515178157
transform 1 0 32660 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_3
timestamp 1515178157
transform 1 0 1380 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_10
timestamp 1515178157
transform 1 0 2024 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_29
timestamp 1515178157
transform 1 0 3772 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_8_32
timestamp 1515178157
transform 1 0 4048 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_8_44
timestamp 1515178157
transform 1 0 5152 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_50
timestamp 1515178157
transform 1 0 5704 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_75
timestamp 1515178157
transform 1 0 8004 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_88
timestamp 1515178157
transform 1 0 9200 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_92
timestamp 1515178157
transform 1 0 9568 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_94
timestamp 1515178157
transform 1 0 9752 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_8_120
timestamp 1515178157
transform 1 0 12144 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_128
timestamp 1515178157
transform 1 0 12880 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_153
timestamp 1515178157
transform 1 0 15180 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_156
timestamp 1515178157
transform 1 0 15456 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_167
timestamp 1515178157
transform 1 0 16468 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_177
timestamp 1515178157
transform 1 0 17388 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_181
timestamp 1515178157
transform 1 0 17756 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_206
timestamp 1515178157
transform 1 0 20056 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_215
timestamp 1515178157
transform 1 0 20884 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_218
timestamp 1515178157
transform 1 0 21160 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_244
timestamp 1515178157
transform 1 0 23552 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_8_272
timestamp 1515178157
transform 1 0 26128 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_278
timestamp 1515178157
transform 1 0 26680 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_280
timestamp 1515178157
transform 1 0 26864 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_8_306
timestamp 1515178157
transform 1 0 29256 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_314
timestamp 1515178157
transform 1 0 29992 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_339
timestamp 1515178157
transform 1 0 32292 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_342
timestamp 1515178157
transform 1 0 32568 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_9_3
timestamp 1515178157
transform 1 0 1380 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_9
timestamp 1515178157
transform 1 0 1932 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_19
timestamp 1515178157
transform 1 0 2852 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_32
timestamp 1515178157
transform 1 0 4048 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_60
timestamp 1515178157
transform 1 0 6624 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_63
timestamp 1515178157
transform 1 0 6900 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_9_91
timestamp 1515178157
transform 1 0 9476 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_97
timestamp 1515178157
transform 1 0 10028 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_122
timestamp 1515178157
transform 1 0 12328 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_125
timestamp 1515178157
transform 1 0 12604 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_9_151
timestamp 1515178157
transform 1 0 14996 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_159
timestamp 1515178157
transform 1 0 15732 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_184
timestamp 1515178157
transform 1 0 18032 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_187
timestamp 1515178157
transform 1 0 18308 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_195
timestamp 1515178157
transform 1 0 19044 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_223
timestamp 1515178157
transform 1 0 21620 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_233
timestamp 1515178157
transform 1 0 22540 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_9_242
timestamp 1515178157
transform 1 0 23368 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_9_249
timestamp 1515178157
transform 1 0 24012 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_275
timestamp 1515178157
transform 1 0 26404 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_9_303
timestamp 1515178157
transform 1 0 28980 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_309
timestamp 1515178157
transform 1 0 29532 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_311
timestamp 1515178157
transform 1 0 29716 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_9_337
timestamp 1515178157
transform 1 0 32108 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_343
timestamp 1515178157
transform 1 0 32660 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_3
timestamp 1515178157
transform 1 0 1380 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_16
timestamp 1515178157
transform 1 0 2576 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_29
timestamp 1515178157
transform 1 0 3772 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_32
timestamp 1515178157
transform 1 0 4048 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_10_58
timestamp 1515178157
transform 1 0 6440 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_66
timestamp 1515178157
transform 1 0 7176 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_91
timestamp 1515178157
transform 1 0 9476 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_10_94
timestamp 1515178157
transform 1 0 9752 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_100
timestamp 1515178157
transform 1 0 10304 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_125
timestamp 1515178157
transform 1 0 12604 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_153
timestamp 1515178157
transform 1 0 15180 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_156
timestamp 1515178157
transform 1 0 15456 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_164
timestamp 1515178157
transform 1 0 16192 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_10_174
timestamp 1515178157
transform 1 0 17112 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_182
timestamp 1515178157
transform 1 0 17848 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_207
timestamp 1515178157
transform 1 0 20148 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_10_214
timestamp 1515178157
transform 1 0 20792 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_218
timestamp 1515178157
transform 1 0 21160 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_10_244
timestamp 1515178157
transform 1 0 23552 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_252
timestamp 1515178157
transform 1 0 24288 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_277
timestamp 1515178157
transform 1 0 26588 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_280
timestamp 1515178157
transform 1 0 26864 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_10_284
timestamp 1515178157
transform 1 0 27232 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_292
timestamp 1515178157
transform 1 0 27968 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_317
timestamp 1515178157
transform 1 0 30268 0 1 5984
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_10_323
timestamp 1515178157
transform 1 0 30820 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_335
timestamp 1515178157
transform 1 0 31924 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_10_342
timestamp 1515178157
transform 1 0 32568 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_11_3
timestamp 1515178157
transform 1 0 1380 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_9
timestamp 1515178157
transform 1 0 1932 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_19
timestamp 1515178157
transform 1 0 2852 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_32
timestamp 1515178157
transform 1 0 4048 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_60
timestamp 1515178157
transform 1 0 6624 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_63
timestamp 1515178157
transform 1 0 6900 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_11_89
timestamp 1515178157
transform 1 0 9292 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_97
timestamp 1515178157
transform 1 0 10028 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_122
timestamp 1515178157
transform 1 0 12328 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_125
timestamp 1515178157
transform 1 0 12604 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_151
timestamp 1515178157
transform 1 0 14996 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_11_179
timestamp 1515178157
transform 1 0 17572 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_185
timestamp 1515178157
transform 1 0 18124 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_187
timestamp 1515178157
transform 1 0 18308 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_213
timestamp 1515178157
transform 1 0 20700 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_11_241
timestamp 1515178157
transform 1 0 23276 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_247
timestamp 1515178157
transform 1 0 23828 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_249
timestamp 1515178157
transform 1 0 24012 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_256
timestamp 1515178157
transform 1 0 24656 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_263
timestamp 1515178157
transform 1 0 25300 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_270
timestamp 1515178157
transform 1 0 25944 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_276
timestamp 1515178157
transform 1 0 26496 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_282
timestamp 1515178157
transform 1 0 27048 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_288
timestamp 1515178157
transform 1 0 27600 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_294
timestamp 1515178157
transform 1 0 28152 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_300
timestamp 1515178157
transform 1 0 28704 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_306
timestamp 1515178157
transform 1 0 29256 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_311
timestamp 1515178157
transform 1 0 29716 0 -1 7072
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_11_315
timestamp 1515178157
transform 1 0 30084 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_327
timestamp 1515178157
transform 1 0 31188 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_339
timestamp 1515178157
transform 1 0 32292 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_343
timestamp 1515178157
transform 1 0 32660 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_3
timestamp 1515178157
transform 1 0 1380 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_10
timestamp 1515178157
transform 1 0 2024 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_29
timestamp 1515178157
transform 1 0 3772 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_12_32
timestamp 1515178157
transform 1 0 4048 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_38
timestamp 1515178157
transform 1 0 4600 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_63
timestamp 1515178157
transform 1 0 6900 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_91
timestamp 1515178157
transform 1 0 9476 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_94
timestamp 1515178157
transform 1 0 9752 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_104
timestamp 1515178157
transform 1 0 10672 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_117
timestamp 1515178157
transform 1 0 11868 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_145
timestamp 1515178157
transform 1 0 14444 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_12_152
timestamp 1515178157
transform 1 0 15088 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_156
timestamp 1515178157
transform 1 0 15456 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_12_164
timestamp 1515178157
transform 1 0 16192 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_172
timestamp 1515178157
transform 1 0 16928 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_197
timestamp 1515178157
transform 1 0 19228 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_207
timestamp 1515178157
transform 1 0 20148 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_12_214
timestamp 1515178157
transform 1 0 20792 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_218
timestamp 1515178157
transform 1 0 21160 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_12_226
timestamp 1515178157
transform 1 0 21896 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_232
timestamp 1515178157
transform 1 0 22448 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_257
timestamp 1515178157
transform 1 0 24748 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_266
timestamp 1515178157
transform 1 0 25576 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_12_273
timestamp 1515178157
transform 1 0 26220 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_12_280
timestamp 1515178157
transform 1 0 26864 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_284
timestamp 1515178157
transform 1 0 27232 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_290
timestamp 1515178157
transform 1 0 27784 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_296
timestamp 1515178157
transform 1 0 28336 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_302
timestamp 1515178157
transform 1 0 28888 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_308
timestamp 1515178157
transform 1 0 29440 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_314
timestamp 1515178157
transform 1 0 29992 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_320
timestamp 1515178157
transform 1 0 30544 0 1 7072
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_12_326
timestamp 1515178157
transform 1 0 31096 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_12_338
timestamp 1515178157
transform 1 0 32200 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_342
timestamp 1515178157
transform 1 0 32568 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_3
timestamp 1515178157
transform 1 0 1380 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_31
timestamp 1515178157
transform 1 0 3956 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_13_59
timestamp 1515178157
transform 1 0 6532 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_63
timestamp 1515178157
transform 1 0 6900 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_74
timestamp 1515178157
transform 1 0 7912 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_84
timestamp 1515178157
transform 1 0 8832 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_88
timestamp 1515178157
transform 1 0 9200 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_113
timestamp 1515178157
transform 1 0 11500 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_122
timestamp 1515178157
transform 1 0 12328 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_125
timestamp 1515178157
transform 1 0 12604 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_133
timestamp 1515178157
transform 1 0 13340 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_161
timestamp 1515178157
transform 1 0 15916 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_174
timestamp 1515178157
transform 1 0 17112 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_184
timestamp 1515178157
transform 1 0 18032 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_187
timestamp 1515178157
transform 1 0 18308 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_13_195
timestamp 1515178157
transform 1 0 19044 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_13_227
timestamp 1515178157
transform 1 0 21988 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_236
timestamp 1515178157
transform 1 0 22816 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_13_245
timestamp 1515178157
transform 1 0 23644 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_249
timestamp 1515178157
transform 1 0 24012 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_275
timestamp 1515178157
transform 1 0 26404 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_282
timestamp 1515178157
transform 1 0 27048 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_288
timestamp 1515178157
transform 1 0 27600 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_294
timestamp 1515178157
transform 1 0 28152 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_300
timestamp 1515178157
transform 1 0 28704 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_306
timestamp 1515178157
transform 1 0 29256 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_13_311
timestamp 1515178157
transform 1 0 29716 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_317
timestamp 1515178157
transform 1 0 30268 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_342
timestamp 1515178157
transform 1 0 32568 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_3
timestamp 1515178157
transform 1 0 1380 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_29
timestamp 1515178157
transform 1 0 3772 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_14_32
timestamp 1515178157
transform 1 0 4048 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_38
timestamp 1515178157
transform 1 0 4600 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_63
timestamp 1515178157
transform 1 0 6900 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_91
timestamp 1515178157
transform 1 0 9476 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_14_94
timestamp 1515178157
transform 1 0 9752 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_100
timestamp 1515178157
transform 1 0 10304 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_125
timestamp 1515178157
transform 1 0 12604 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_153
timestamp 1515178157
transform 1 0 15180 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_156
timestamp 1515178157
transform 1 0 15456 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_160
timestamp 1515178157
transform 1 0 15824 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_185
timestamp 1515178157
transform 1 0 18124 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_213
timestamp 1515178157
transform 1 0 20700 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_218
timestamp 1515178157
transform 1 0 21160 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_244
timestamp 1515178157
transform 1 0 23552 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_14_272
timestamp 1515178157
transform 1 0 26128 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_278
timestamp 1515178157
transform 1 0 26680 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_280
timestamp 1515178157
transform 1 0 26864 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_14_306
timestamp 1515178157
transform 1 0 29256 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_314
timestamp 1515178157
transform 1 0 29992 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_339
timestamp 1515178157
transform 1 0 32292 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_342
timestamp 1515178157
transform 1 0 32568 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_3
timestamp 1515178157
transform 1 0 1380 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_15_29
timestamp 1515178157
transform 1 0 3772 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_15_59
timestamp 1515178157
transform 1 0 6532 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_63
timestamp 1515178157
transform 1 0 6900 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_74
timestamp 1515178157
transform 1 0 7912 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_87
timestamp 1515178157
transform 1 0 9108 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_91
timestamp 1515178157
transform 1 0 9476 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_116
timestamp 1515178157
transform 1 0 11776 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_122
timestamp 1515178157
transform 1 0 12328 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_15_125
timestamp 1515178157
transform 1 0 12604 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_131
timestamp 1515178157
transform 1 0 13156 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_156
timestamp 1515178157
transform 1 0 15456 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_184
timestamp 1515178157
transform 1 0 18032 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_187
timestamp 1515178157
transform 1 0 18308 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_191
timestamp 1515178157
transform 1 0 18676 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_15_216
timestamp 1515178157
transform 1 0 20976 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_15_246
timestamp 1515178157
transform 1 0 23736 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_249
timestamp 1515178157
transform 1 0 24012 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_256
timestamp 1515178157
transform 1 0 24656 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_284
timestamp 1515178157
transform 1 0 27232 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_291
timestamp 1515178157
transform 1 0 27876 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_298
timestamp 1515178157
transform 1 0 28520 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_15_304
timestamp 1515178157
transform 1 0 29072 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_15_311
timestamp 1515178157
transform 1 0 29716 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_15_337
timestamp 1515178157
transform 1 0 32108 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_343
timestamp 1515178157
transform 1 0 32660 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_3
timestamp 1515178157
transform 1 0 1380 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_29
timestamp 1515178157
transform 1 0 3772 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_16_32
timestamp 1515178157
transform 1 0 4048 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_38
timestamp 1515178157
transform 1 0 4600 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_63
timestamp 1515178157
transform 1 0 6900 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_91
timestamp 1515178157
transform 1 0 9476 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_16_94
timestamp 1515178157
transform 1 0 9752 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_100
timestamp 1515178157
transform 1 0 10304 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_125
timestamp 1515178157
transform 1 0 12604 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_153
timestamp 1515178157
transform 1 0 15180 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_156
timestamp 1515178157
transform 1 0 15456 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_16_167
timestamp 1515178157
transform 1 0 16468 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_173
timestamp 1515178157
transform 1 0 17020 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_198
timestamp 1515178157
transform 1 0 19320 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_208
timestamp 1515178157
transform 1 0 20240 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_215
timestamp 1515178157
transform 1 0 20884 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_218
timestamp 1515178157
transform 1 0 21160 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_16_244
timestamp 1515178157
transform 1 0 23552 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_252
timestamp 1515178157
transform 1 0 24288 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_277
timestamp 1515178157
transform 1 0 26588 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_280
timestamp 1515178157
transform 1 0 26864 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_306
timestamp 1515178157
transform 1 0 29256 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_16_334
timestamp 1515178157
transform 1 0 31832 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_340
timestamp 1515178157
transform 1 0 32384 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_342
timestamp 1515178157
transform 1 0 32568 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_3
timestamp 1515178157
transform 1 0 1380 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_7
timestamp 1515178157
transform 1 0 1748 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_32
timestamp 1515178157
transform 1 0 4048 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_60
timestamp 1515178157
transform 1 0 6624 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_17_63
timestamp 1515178157
transform 1 0 6900 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_69
timestamp 1515178157
transform 1 0 7452 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_94
timestamp 1515178157
transform 1 0 9752 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_122
timestamp 1515178157
transform 1 0 12328 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_17_125
timestamp 1515178157
transform 1 0 12604 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_131
timestamp 1515178157
transform 1 0 13156 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_156
timestamp 1515178157
transform 1 0 15456 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_184
timestamp 1515178157
transform 1 0 18032 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_187
timestamp 1515178157
transform 1 0 18308 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_198
timestamp 1515178157
transform 1 0 19320 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_202
timestamp 1515178157
transform 1 0 19688 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_227
timestamp 1515178157
transform 1 0 21988 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_237
timestamp 1515178157
transform 1 0 22908 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_246
timestamp 1515178157
transform 1 0 23736 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_249
timestamp 1515178157
transform 1 0 24012 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_275
timestamp 1515178157
transform 1 0 26404 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_17_303
timestamp 1515178157
transform 1 0 28980 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_309
timestamp 1515178157
transform 1 0 29532 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_311
timestamp 1515178157
transform 1 0 29716 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_17_337
timestamp 1515178157
transform 1 0 32108 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_343
timestamp 1515178157
transform 1 0 32660 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_3
timestamp 1515178157
transform 1 0 1380 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_29
timestamp 1515178157
transform 1 0 3772 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_18_32
timestamp 1515178157
transform 1 0 4048 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_38
timestamp 1515178157
transform 1 0 4600 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_63
timestamp 1515178157
transform 1 0 6900 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_91
timestamp 1515178157
transform 1 0 9476 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_18_94
timestamp 1515178157
transform 1 0 9752 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_100
timestamp 1515178157
transform 1 0 10304 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_125
timestamp 1515178157
transform 1 0 12604 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_153
timestamp 1515178157
transform 1 0 15180 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_156
timestamp 1515178157
transform 1 0 15456 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_160
timestamp 1515178157
transform 1 0 15824 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_185
timestamp 1515178157
transform 1 0 18124 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_213
timestamp 1515178157
transform 1 0 20700 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_218
timestamp 1515178157
transform 1 0 21160 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_244
timestamp 1515178157
transform 1 0 23552 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_18_272
timestamp 1515178157
transform 1 0 26128 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_278
timestamp 1515178157
transform 1 0 26680 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_280
timestamp 1515178157
transform 1 0 26864 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_284
timestamp 1515178157
transform 1 0 27232 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_312
timestamp 1515178157
transform 1 0 29808 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_318
timestamp 1515178157
transform 1 0 30360 0 1 10336
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_18_324
timestamp 1515178157
transform 1 0 30912 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_336
timestamp 1515178157
transform 1 0 32016 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_340
timestamp 1515178157
transform 1 0 32384 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_342
timestamp 1515178157
transform 1 0 32568 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_3
timestamp 1515178157
transform 1 0 1380 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_29
timestamp 1515178157
transform 1 0 3772 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_32
timestamp 1515178157
transform 1 0 4048 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_60
timestamp 1515178157
transform 1 0 6624 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_63
timestamp 1515178157
transform 1 0 6900 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_91
timestamp 1515178157
transform 1 0 9476 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_94
timestamp 1515178157
transform 1 0 9752 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_120
timestamp 1515178157
transform 1 0 12144 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_125
timestamp 1515178157
transform 1 0 12604 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_151
timestamp 1515178157
transform 1 0 14996 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_156
timestamp 1515178157
transform 1 0 15456 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_182
timestamp 1515178157
transform 1 0 17848 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_187
timestamp 1515178157
transform 1 0 18308 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_213
timestamp 1515178157
transform 1 0 20700 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_218
timestamp 1515178157
transform 1 0 21160 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_244
timestamp 1515178157
transform 1 0 23552 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_249
timestamp 1515178157
transform 1 0 24012 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_256
timestamp 1515178157
transform 1 0 24656 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_265
timestamp 1515178157
transform 1 0 25484 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_274
timestamp 1515178157
transform 1 0 26312 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_278
timestamp 1515178157
transform 1 0 26680 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_280
timestamp 1515178157
transform 1 0 26864 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_285
timestamp 1515178157
transform 1 0 27324 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_292
timestamp 1515178157
transform 1 0 27968 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_298
timestamp 1515178157
transform 1 0 28520 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_19_304
timestamp 1515178157
transform 1 0 29072 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_19_311
timestamp 1515178157
transform 1 0 29716 0 -1 11424
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_19_315
timestamp 1515178157
transform 1 0 30084 0 -1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_327
timestamp 1515178157
transform 1 0 31188 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_19_339
timestamp 1515178157
transform 1 0 32292 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_342
timestamp 1515178157
transform 1 0 32568 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  inbuf_1
timestamp 1515178157
transform -1 0 22908 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  inbuf_2
timestamp 1515178157
transform 1 0 20516 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  inbuf_3
timestamp 1515178157
transform -1 0 7360 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__bufbuf_8  outbuf_1
timestamp 1515178157
transform -1 0 4048 0 -1 3808
box -38 -48 1418 592
use sky130_fd_sc_hd__bufbuf_8  outbuf_2
timestamp 1515178157
transform -1 0 14168 0 -1 3808
box -38 -48 1418 592
use sky130_fd_sc_hd__bufbuf_8  outbuf_3
timestamp 1515178157
transform 1 0 2392 0 1 7072
box -38 -48 1418 592
use sky130_fd_sc_hd__bufbuf_8  outbuf_4
timestamp 1515178157
transform -1 0 3772 0 1 4896
box -38 -48 1418 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1515178157
transform 1 0 1104 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1515178157
transform -1 0 33028 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1515178157
transform 1 0 1104 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1515178157
transform -1 0 33028 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1515178157
transform 1 0 1104 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1515178157
transform -1 0 33028 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1515178157
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1515178157
transform -1 0 33028 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1515178157
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1515178157
transform -1 0 33028 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1515178157
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1515178157
transform -1 0 33028 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1515178157
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1515178157
transform -1 0 33028 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1515178157
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1515178157
transform -1 0 33028 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1515178157
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1515178157
transform -1 0 33028 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1515178157
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1515178157
transform -1 0 33028 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1515178157
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1515178157
transform -1 0 33028 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1515178157
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1515178157
transform -1 0 33028 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1515178157
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1515178157
transform -1 0 33028 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1515178157
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1515178157
transform -1 0 33028 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1515178157
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1515178157
transform -1 0 33028 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1515178157
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1515178157
transform -1 0 33028 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1515178157
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1515178157
transform -1 0 33028 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1515178157
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1515178157
transform -1 0 33028 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1515178157
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1515178157
transform -1 0 33028 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1515178157
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1515178157
transform -1 0 33028 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_40
timestamp 1515178157
transform 1 0 3956 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_41
timestamp 1515178157
transform 1 0 6808 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_42
timestamp 1515178157
transform 1 0 9660 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_43
timestamp 1515178157
transform 1 0 12512 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_44
timestamp 1515178157
transform 1 0 15364 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_45
timestamp 1515178157
transform 1 0 18216 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_46
timestamp 1515178157
transform 1 0 21068 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_47
timestamp 1515178157
transform 1 0 23920 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_48
timestamp 1515178157
transform 1 0 26772 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_49
timestamp 1515178157
transform 1 0 29624 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_50
timestamp 1515178157
transform 1 0 32476 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_51
timestamp 1515178157
transform 1 0 6808 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_52
timestamp 1515178157
transform 1 0 12512 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_53
timestamp 1515178157
transform 1 0 18216 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_54
timestamp 1515178157
transform 1 0 23920 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_55
timestamp 1515178157
transform 1 0 29624 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_56
timestamp 1515178157
transform 1 0 3956 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_57
timestamp 1515178157
transform 1 0 9660 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_58
timestamp 1515178157
transform 1 0 15364 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_59
timestamp 1515178157
transform 1 0 21068 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_60
timestamp 1515178157
transform 1 0 26772 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_61
timestamp 1515178157
transform 1 0 32476 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_62
timestamp 1515178157
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_63
timestamp 1515178157
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_64
timestamp 1515178157
transform 1 0 18216 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_65
timestamp 1515178157
transform 1 0 23920 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_66
timestamp 1515178157
transform 1 0 29624 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_67
timestamp 1515178157
transform 1 0 3956 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_68
timestamp 1515178157
transform 1 0 9660 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_69
timestamp 1515178157
transform 1 0 15364 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_70
timestamp 1515178157
transform 1 0 21068 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_71
timestamp 1515178157
transform 1 0 26772 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_72
timestamp 1515178157
transform 1 0 32476 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_73
timestamp 1515178157
transform 1 0 6808 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_74
timestamp 1515178157
transform 1 0 12512 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_75
timestamp 1515178157
transform 1 0 18216 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_76
timestamp 1515178157
transform 1 0 23920 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_77
timestamp 1515178157
transform 1 0 29624 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_78
timestamp 1515178157
transform 1 0 3956 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_79
timestamp 1515178157
transform 1 0 9660 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_80
timestamp 1515178157
transform 1 0 15364 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_81
timestamp 1515178157
transform 1 0 21068 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_82
timestamp 1515178157
transform 1 0 26772 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_83
timestamp 1515178157
transform 1 0 32476 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_84
timestamp 1515178157
transform 1 0 6808 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_85
timestamp 1515178157
transform 1 0 12512 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_86
timestamp 1515178157
transform 1 0 18216 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_87
timestamp 1515178157
transform 1 0 23920 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_88
timestamp 1515178157
transform 1 0 29624 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_89
timestamp 1515178157
transform 1 0 3956 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_90
timestamp 1515178157
transform 1 0 9660 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_91
timestamp 1515178157
transform 1 0 15364 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_92
timestamp 1515178157
transform 1 0 21068 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_93
timestamp 1515178157
transform 1 0 26772 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_94
timestamp 1515178157
transform 1 0 32476 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_95
timestamp 1515178157
transform 1 0 6808 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_96
timestamp 1515178157
transform 1 0 12512 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_97
timestamp 1515178157
transform 1 0 18216 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_98
timestamp 1515178157
transform 1 0 23920 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_99
timestamp 1515178157
transform 1 0 29624 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_100
timestamp 1515178157
transform 1 0 3956 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_101
timestamp 1515178157
transform 1 0 9660 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_102
timestamp 1515178157
transform 1 0 15364 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_103
timestamp 1515178157
transform 1 0 21068 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_104
timestamp 1515178157
transform 1 0 26772 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_105
timestamp 1515178157
transform 1 0 32476 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_106
timestamp 1515178157
transform 1 0 6808 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_107
timestamp 1515178157
transform 1 0 12512 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_108
timestamp 1515178157
transform 1 0 18216 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_109
timestamp 1515178157
transform 1 0 23920 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_110
timestamp 1515178157
transform 1 0 29624 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_111
timestamp 1515178157
transform 1 0 3956 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_112
timestamp 1515178157
transform 1 0 9660 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_113
timestamp 1515178157
transform 1 0 15364 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_114
timestamp 1515178157
transform 1 0 21068 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_115
timestamp 1515178157
transform 1 0 26772 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_116
timestamp 1515178157
transform 1 0 32476 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_117
timestamp 1515178157
transform 1 0 6808 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_118
timestamp 1515178157
transform 1 0 12512 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_119
timestamp 1515178157
transform 1 0 18216 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_120
timestamp 1515178157
transform 1 0 23920 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_121
timestamp 1515178157
transform 1 0 29624 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_122
timestamp 1515178157
transform 1 0 3956 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_123
timestamp 1515178157
transform 1 0 9660 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_124
timestamp 1515178157
transform 1 0 15364 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_125
timestamp 1515178157
transform 1 0 21068 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_126
timestamp 1515178157
transform 1 0 26772 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_127
timestamp 1515178157
transform 1 0 32476 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_128
timestamp 1515178157
transform 1 0 6808 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_129
timestamp 1515178157
transform 1 0 12512 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130
timestamp 1515178157
transform 1 0 18216 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 1515178157
transform 1 0 23920 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 1515178157
transform 1 0 29624 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 1515178157
transform 1 0 3956 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 1515178157
transform 1 0 9660 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 1515178157
transform 1 0 15364 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 1515178157
transform 1 0 21068 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1515178157
transform 1 0 26772 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1515178157
transform 1 0 32476 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1515178157
transform 1 0 6808 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1515178157
transform 1 0 12512 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1515178157
transform 1 0 18216 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1515178157
transform 1 0 23920 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1515178157
transform 1 0 29624 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1515178157
transform 1 0 3956 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1515178157
transform 1 0 9660 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1515178157
transform 1 0 15364 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1515178157
transform 1 0 21068 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1515178157
transform 1 0 26772 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1515178157
transform 1 0 32476 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1515178157
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1515178157
transform 1 0 6808 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1515178157
transform 1 0 9660 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1515178157
transform 1 0 12512 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1515178157
transform 1 0 15364 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1515178157
transform 1 0 18216 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1515178157
transform 1 0 21068 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1515178157
transform 1 0 23920 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1515178157
transform 1 0 26772 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1515178157
transform 1 0 29624 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1515178157
transform 1 0 32476 0 -1 11424
box -38 -48 130 592
<< labels >>
rlabel metal1 s 17066 10880 17066 10880 4 VDD
rlabel metal1 s 17066 11424 17066 11424 4 VSS
rlabel metal1 s 24380 6222 24380 6222 4 clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[11\]
rlabel metal1 s 26381 6188 26381 6188 4 clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[12\]
rlabel metal1 s 27876 6222 27876 6222 4 clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[14\]
rlabel metal1 s 24242 6970 24242 6970 4 clkgen.delay_155ns_3.bypass_enable_w\[3\]
rlabel metal1 s 20884 6834 20884 6834 4 clkgen.delay_155ns_3.genblk1\[3\].dly_binary.signal_w\[5\]
rlabel metal1 s 21666 6222 21666 6222 4 clkgen.delay_155ns_3.genblk1\[3\].dly_binary.signal_w\[6\]
rlabel metal1 s 24426 7310 24426 7310 4 clkgen.delay_155ns_3.genblk1\[3\].dly_binary.signal_w\[7\]
rlabel metal1 s 25254 7378 25254 7378 4 edgedetect.dly_315ns_1.bypass_enable_w\[0\]
rlabel metal1 s 25254 11152 25254 11152 4 edgedetect.dly_315ns_1.bypass_enable_w\[3\]
rlabel metal1 s 26082 11220 26082 11220 4 edgedetect.dly_315ns_1.bypass_enable_w\[4\]
rlabel metal1 s 25346 7276 25346 7276 4 edgedetect.dly_315ns_1.bypass_enable_w\[5\]
rlabel metal1 s 19734 9418 19734 9418 4 edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.bypass_in
rlabel metal1 s 18446 10166 18446 10166 4 edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.out
rlabel metal1 s 18722 9996 18722 9996 4 edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.bypass_in
rlabel metal1 s 19228 9894 19228 9894 4 edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.out
rlabel metal1 s 17825 10132 17825 10132 4 edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.signal_w\[8\]
rlabel metal1 s 17434 7854 17434 7854 4 edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.bypass_in
rlabel metal1 s 18032 7718 18032 7718 4 edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.out
rlabel metal1 s 18170 11186 18170 11186 4 edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[10\]
rlabel metal1 s 20493 10540 20493 10540 4 edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[13\]
rlabel metal1 s 23276 11186 23276 11186 4 edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[14\]
rlabel metal1 s 21551 11220 21551 11220 4 edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[15\]
rlabel metal1 s 18768 8398 18768 8398 4 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[10\]
rlabel metal1 s 21781 7956 21781 7956 4 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[12\]
rlabel metal1 s 23345 8364 23345 8364 4 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[13\]
rlabel metal1 s 25921 8364 25921 8364 4 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[14\]
rlabel metal1 s 18308 9010 18308 9010 4 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[17\]
rlabel metal1 s 18814 8976 18814 8976 4 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[18\]
rlabel metal1 s 21528 9486 21528 9486 4 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[20\]
rlabel metal1 s 21850 9078 21850 9078 4 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[21\]
rlabel metal1 s 23529 9044 23529 9044 4 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[22\]
rlabel metal1 s 24702 9486 24702 9486 4 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[23\]
rlabel metal1 s 29601 10540 29601 10540 4 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[26\]
rlabel metal1 s 32246 7922 32246 7922 4 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[27\]
rlabel metal1 s 30567 7956 30567 7956 4 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[28\]
rlabel metal1 s 17342 9486 17342 9486 4 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[9\]
rlabel metal1 s 4094 10098 4094 10098 4 edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.signal_w\[0\]
rlabel metal1 s 4462 10064 4462 10064 4 edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.signal_w\[1\]
rlabel metal1 s 7314 9520 7314 9520 4 edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.signal_w\[2\]
rlabel metal1 s 9246 9452 9246 9452 4 edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.signal_w\[3\]
rlabel metal1 s 12972 6834 12972 6834 4 clkgen.delay_155ns_3.genblk1\[3\].dly_binary.signal_w\[0\]
rlabel metal1 s 7130 6222 7130 6222 4 clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[1\]
rlabel metal1 s 9246 6188 9246 6188 4 clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[2\]
rlabel metal1 s 14973 6188 14973 6188 4 clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[5\]
rlabel metal1 s 15134 11696 15134 11696 4 dlycontrol4_in[3]
rlabel metal1 s 16928 6222 16928 6222 4 clkgen.delay_155ns_2.genblk1\[4\].dly_binary.bypass_in
rlabel metal1 s 15778 6222 15778 6222 4 clkgen.delay_155ns_3.genblk1\[0\].dly_binary.bypass_in
rlabel metal1 s 16790 7922 16790 7922 4 edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[16\]
rlabel metal1 s 3565 10540 3565 10540 4 edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[2\]
rlabel metal1 s 11960 10132 11960 10132 4 edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[7\]
rlabel metal1 s 12926 10098 12926 10098 4 edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[8\]
rlabel metal1 s 6624 6222 6624 6222 4 clkgen.delay_155ns_3.genblk1\[0\].dly_binary.signal_w\[0\]
rlabel metal1 s 6992 7922 6992 7922 4 clkgen.delay_155ns_3.genblk1\[1\].dly_binary.out
rlabel metal1 s 16284 7310 16284 7310 4 edgedetect.dly_315ns_1.enable_dlycontrol_w
rlabel metal1 s 2254 6732 2254 6732 4 edgedetect.dly_315ns_1.genblk1\[0\].dly_binary.bypass_in
rlabel metal1 s 2254 6970 2254 6970 4 edgedetect.dly_315ns_1.genblk1\[0\].dly_binary.signal_w\[1\]
rlabel metal1 s 1863 8364 1863 8364 4 edgedetect.dly_315ns_1.genblk1\[1\].dly_binary.signal_w\[1\]
rlabel metal1 s 6325 7956 6325 7956 4 edgedetect.dly_315ns_1.genblk1\[1\].dly_binary.signal_w\[2\]
rlabel metal1 s 7130 6800 7130 6800 4 clkgen.delay_155ns_3.genblk1\[1\].dly_binary.signal_w\[1\]
rlabel metal1 s 10120 7446 10120 7446 4 clkgen.delay_155ns_3.genblk1\[2\].dly_binary.out
rlabel metal1 s 7406 10098 7406 10098 4 edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.signal_w\[2\]
rlabel metal1 s 9545 10132 9545 10132 4 edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.signal_w\[3\]
rlabel metal1 s 9108 9146 9108 9146 4 edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.signal_w\[4\]
rlabel metal1 s 12328 6834 12328 6834 4 clkgen.delay_155ns_3.genblk1\[2\].dly_binary.signal_w\[3\]
rlabel metal1 s 6693 8364 6693 8364 4 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[2\]
rlabel metal1 s 10810 8280 10810 8280 4 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[4\]
rlabel metal1 s 12236 8364 12236 8364 4 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[5\]
rlabel metal1 s 10327 6868 10327 6868 4 clkgen.delay_155ns_3.genblk1\[2\].dly_binary.signal_w\[4\]
rlabel metal1 s 2162 7310 2162 7310 4 sample_p_1
rlabel metal1 s 9936 2482 9936 2482 4 clkgen.delay_155ns_1.genblk1\[2\].dly_binary.signal_w\[2\]
rlabel metal1 s 9108 5066 9108 5066 4 clkgen.delay_155ns_1.genblk1\[2\].dly_binary.signal_w\[4\]
rlabel metal1 s 16100 1802 16100 1802 4 clkgen.delay_155ns_1.genblk1\[3\].dly_binary.bypass_in
rlabel metal1 s 7268 1394 7268 1394 4 clkgen.delay_155ns_1.genblk1\[3\].dly_binary.signal_w\[1\]
rlabel metal1 s 9545 1428 9545 1428 4 clkgen.delay_155ns_1.genblk1\[3\].dly_binary.signal_w\[2\]
rlabel metal1 s 15364 2482 15364 2482 4 clkgen.delay_155ns_1.genblk1\[3\].dly_binary.signal_w\[5\]
rlabel metal1 s 13754 4692 13754 4692 4 clkgen.delay_155ns_3.genblk1\[3\].dly_binary.out
rlabel metal1 s 14973 1428 14973 1428 4 clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[11\]
rlabel metal1 s 16146 1394 16146 1394 4 clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[13\]
rlabel metal1 s 4899 1836 4899 1836 4 clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[6\]
rlabel metal1 s 7084 782 7084 782 4 clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[7\]
rlabel metal1 s 11454 3502 11454 3502 4 clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[0\]
rlabel metal1 s 12282 4675 12282 4675 4 clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[1\]
rlabel metal1 s 13110 306 13110 306 4 dlycontrol1_in[0]
rlabel metal1 s 9269 748 9269 748 4 clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[8\]
rlabel metal1 s 2346 5644 2346 5644 4 clkgen.delay_155ns_2.genblk1\[0\].dly_binary.out
rlabel metal1 s 7866 4658 7866 4658 4 clkgen.delay_155ns_2.genblk1\[2\].dly_binary.signal_w\[2\]
rlabel metal1 s 9660 4046 9660 4046 4 clkgen.delay_155ns_2.genblk1\[2\].dly_binary.signal_w\[3\]
rlabel metal1 s 11937 4012 11937 4012 4 clkgen.delay_155ns_2.genblk1\[2\].dly_binary.signal_w\[4\]
rlabel metal1 s 7314 5712 7314 5712 4 clkgen.delay_155ns_2.genblk1\[3\].dly_binary.signal_w\[1\]
rlabel metal1 s 9752 5134 9752 5134 4 clkgen.delay_155ns_2.genblk1\[3\].dly_binary.signal_w\[2\]
rlabel metal1 s 10396 5746 10396 5746 4 clkgen.delay_155ns_2.genblk1\[3\].dly_binary.signal_w\[3\]
rlabel metal1 s 14122 3536 14122 3536 4 clkgen.clk_comp_out
rlabel metal1 s 2254 5134 2254 5134 4 clkgen.clk_dig_delayed_w
rlabel metal1 s 7130 3468 7130 3468 4 clkgen.delay_155ns_1.genblk1\[0\].dly_binary.in
rlabel metal1 s 7176 2958 7176 2958 4 clkgen.delay_155ns_1.genblk1\[0\].dly_binary.signal_w\[0\]
rlabel metal1 s 8602 3570 8602 3570 4 clkgen.delay_155ns_1.genblk1\[0\].dly_binary.signal_w\[1\]
rlabel metal1 s 8188 2618 8188 2618 4 clkgen.delay_155ns_1.genblk1\[1\].dly_binary.signal_w\[1\]
rlabel metal1 s 5980 3978 5980 3978 4 clkgen.delay_155ns_1.genblk1\[1\].dly_binary.signal_w\[2\]
rlabel metal1 s 14766 714 14766 714 4 clkgen.delay_155ns_1.genblk1\[2\].dly_binary.bypass_in
rlabel metal1 s 7590 2448 7590 2448 4 clkgen.delay_155ns_1.genblk1\[2\].dly_binary.signal_w\[1\]
rlabel metal1 s 5428 4998 5428 4998 4 clkgen.delay_155ns_3.genblk1\[0\].dly_binary.out
rlabel metal1 s 18722 748 18722 748 4 clkgen.delay_155ns_1.bypass_enable_w\[0\]
rlabel metal1 s 18354 4522 18354 4522 4 clkgen.delay_155ns_2.genblk1\[1\].dly_binary.out
rlabel metal1 s 18584 4590 18584 4590 4 clkgen.delay_155ns_2.genblk1\[2\].dly_binary.bypass_in
rlabel metal1 s 21298 2312 21298 2312 4 clkgen.delay_155ns_1.genblk1\[3\].dly_binary.out
rlabel metal1 s 22218 2516 22218 2516 4 clkgen.delay_155ns_1.bypass_enable_w\[1\]
rlabel metal1 s 21390 2550 21390 2550 4 clkgen.delay_155ns_1.genblk1\[1\].dly_binary.bypass_in
rlabel metal1 s 22494 2992 22494 2992 4 clkgen.delay_155ns_1.bypass_enable_w\[2\]
rlabel metal1 s 17549 2516 17549 2516 4 clkgen.delay_155ns_1.genblk1\[3\].dly_binary.signal_w\[6\]
rlabel metal1 s 21574 952 21574 952 4 clkgen.delay_155ns_1.bypass_enable_w\[3\]
rlabel metal1 s 17986 5135 17986 5135 4 clkgen.delay_155ns_2.genblk1\[3\].dly_binary.signal_w\[7\]
rlabel metal1 s 17066 5270 17066 5270 4 clkgen.delay_155ns_3.genblk1\[4\].dly_binary.bypass_in
rlabel metal1 s 21574 1530 21574 1530 4 clkgen.delay_155ns_1.bypass_enable_w\[4\]
rlabel metal1 s 24426 3570 24426 3570 4 clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[10\]
rlabel metal1 s 26473 3604 26473 3604 4 clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[11\]
rlabel metal1 s 27370 4046 27370 4046 4 clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[12\]
rlabel metal1 s 29578 4658 29578 4658 4 clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[13\]
rlabel metal1 s 31970 5134 31970 5134 4 clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[15\]
rlabel metal1 s 17894 5168 17894 5168 4 clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[16\]
rlabel metal1 s 17825 1428 17825 1428 4 clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[14\]
rlabel metal1 s 18998 4046 18998 4046 4 clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[5\]
rlabel metal1 s 20194 4658 20194 4658 4 clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[6\]
rlabel metal1 s 21528 4046 21528 4046 4 clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[7\]
rlabel metal1 s 24104 4658 24104 4658 4 clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[8\]
rlabel metal1 s 19849 1836 19849 1836 4 clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[15\]
rlabel metal1 s 23506 2482 23506 2482 4 dlycontrol1_in[1]
rlabel metal1 s 21390 1904 21390 1904 4 dlycontrol2_in[3]
rlabel metal1 s 29026 5134 29026 5134 4 clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[13\]
rlabel metal1 s 20332 1870 20332 1870 4 clkgen.delay_155ns_1.enable_dlycontrol_w
rlabel metal1 s 18262 646 18262 646 4 clkgen.delay_155ns_1.genblk1\[0\].dly_binary.bypass_in
rlabel metal1 s 19872 3094 19872 3094 4 clkgen.clk_dig_out
rlabel metal1 s 22172 2074 22172 2074 4 clkgen.delay_155ns_2.bypass_enable_w\[0\]
rlabel metal1 s 17825 5780 17825 5780 4 clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[6\]
rlabel metal1 s 23874 5746 23874 5746 4 clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[9\]
rlabel metal1 s 20332 5134 20332 5134 4 clkgen.delay_155ns_3.bypass_enable_w\[0\]
rlabel metal1 s 22678 3162 22678 3162 4 clkgen.delay_155ns_2.bypass_enable_w\[2\]
rlabel metal1 s 21896 2006 21896 2006 4 clkgen.delay_155ns_2.bypass_enable_w\[3\]
rlabel metal1 s 21298 3502 21298 3502 4 clkgen.delay_155ns_2.bypass_enable_w\[4\]
rlabel metal1 s 23920 1870 23920 1870 4 ena_in
rlabel metal1 s 21712 3502 21712 3502 4 clkgen.delay_155ns_2.enable_dlycontrol_w
rlabel metal3 s 1740 1836 1740 1836 4 clk_dig_out
rlabel metal3 s 12374 1411 12374 1411 4 clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[10\]
rlabel metal3 s 18722 5661 18722 5661 4 clkgen.delay_155ns_3.enable_dlycontrol_w
rlabel metal3 s 17388 6324 17388 6324 4 clkgen.delay_155ns_3.genblk1\[2\].dly_binary.bypass_in
rlabel metal3 s 5750 7276 5750 7276 4 clkgen.delay_155ns_3.genblk1\[2\].dly_binary.signal_w\[1\]
rlabel metal3 s 4140 3264 4140 3264 4 dlycontrol1_in[2]
rlabel metal3 s 0 4632 800 4752 4 dlycontrol2_in[0]
port 10 nsew
rlabel metal3 s 0 5040 800 5160 4 dlycontrol2_in[1]
port 11 nsew
rlabel metal3 s 17204 6188 17204 6188 4 dlycontrol2_in[4]
rlabel metal3 s 1326 6732 1326 6732 4 dlycontrol3_in[0]
rlabel metal3 s 22034 10421 22034 10421 4 dlycontrol3_in[2]
rlabel metal3 s 0 8304 800 8424 4 dlycontrol3_in[4]
port 19 nsew
rlabel metal3 s 820 8772 820 8772 4 dlycontrol4_in[0]
rlabel metal3 s 0 9120 800 9240 4 dlycontrol4_in[1]
port 21 nsew
rlabel metal3 s 11040 8228 11040 8228 4 edgedetect.dly_315ns_1.genblk1\[1\].dly_binary.out
rlabel metal3 s 12466 11883 12466 11883 4 edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[0\]
rlabel metal3 s 16974 10540 16974 10540 4 edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[12\]
rlabel metal3 s 8740 10540 8740 10540 4 edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[6\]
rlabel metal3 s 17894 6443 17894 6443 4 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.out
rlabel metal3 s 2714 7395 2714 7395 4 edgedetect.start_conv_edge_w
rlabel metal3 s 1717 2244 1717 2244 4 enable_dlycontrol_in
rlabel metal3 s 1050 612 1050 612 4 sample_n_out
rlabel metal3 s 866 11220 866 11220 4 sample_p_in
rlabel metal3 s 820 11628 820 11628 4 sample_p_out
rlabel metal3 s 1717 1428 1717 1428 4 start_conv_in
flabel metal3 s 1056 4384 33076 4704 0 FreeSans 2400 0 0 0 VDD
port 1 nsew
flabel metal3 s 1056 8384 33076 8704 0 FreeSans 2400 0 0 0 VDD
port 1 nsew
flabel metal3 s 1056 5044 33076 5364 0 FreeSans 2400 0 0 0 VSS
port 2 nsew
flabel metal3 s 1056 9044 33076 9364 0 FreeSans 2400 0 0 0 VSS
port 2 nsew
flabel metal3 s 33400 2864 34200 2984 0 FreeSans 600 0 0 0 clk_comp_out
port 3 nsew
flabel metal3 s 0 1776 800 1896 0 FreeSans 600 0 0 0 clk_dig_out
port 4 nsew
flabel metal3 s 0 2592 800 2712 0 FreeSans 600 0 0 0 dlycontrol1_in[0]
port 5 nsew
flabel metal3 s 0 3000 800 3120 0 FreeSans 600 0 0 0 dlycontrol1_in[1]
port 6 nsew
flabel metal3 s 0 3408 800 3528 0 FreeSans 600 0 0 0 dlycontrol1_in[2]
port 7 nsew
flabel metal3 s 0 3816 800 3936 0 FreeSans 600 0 0 0 dlycontrol1_in[3]
port 8 nsew
flabel metal3 s 0 4224 800 4344 0 FreeSans 600 0 0 0 dlycontrol1_in[4]
port 9 nsew
flabel metal3 s 400 4692 400 4692 0 FreeSans 600 0 0 0 dlycontrol2_in[0]
flabel metal3 s 400 5100 400 5100 0 FreeSans 600 0 0 0 dlycontrol2_in[1]
flabel metal3 s 0 5448 800 5568 0 FreeSans 600 0 0 0 dlycontrol2_in[2]
port 12 nsew
flabel metal3 s 0 5856 800 5976 0 FreeSans 600 0 0 0 dlycontrol2_in[3]
port 13 nsew
flabel metal3 s 0 6264 800 6384 0 FreeSans 600 0 0 0 dlycontrol2_in[4]
port 14 nsew
flabel metal3 s 0 6672 800 6792 0 FreeSans 600 0 0 0 dlycontrol3_in[0]
port 15 nsew
flabel metal3 s 0 7080 800 7200 0 FreeSans 600 0 0 0 dlycontrol3_in[1]
port 16 nsew
flabel metal3 s 0 7488 800 7608 0 FreeSans 600 0 0 0 dlycontrol3_in[2]
port 17 nsew
flabel metal3 s 0 7896 800 8016 0 FreeSans 600 0 0 0 dlycontrol3_in[3]
port 18 nsew
flabel metal3 s 400 8364 400 8364 0 FreeSans 600 0 0 0 dlycontrol3_in[4]
flabel metal3 s 0 8712 800 8832 0 FreeSans 600 0 0 0 dlycontrol4_in[0]
port 20 nsew
flabel metal3 s 400 9180 400 9180 0 FreeSans 600 0 0 0 dlycontrol4_in[1]
flabel metal3 s 0 9528 800 9648 0 FreeSans 600 0 0 0 dlycontrol4_in[2]
port 22 nsew
flabel metal3 s 0 9936 800 10056 0 FreeSans 600 0 0 0 dlycontrol4_in[3]
port 23 nsew
flabel metal3 s 0 10344 800 10464 0 FreeSans 600 0 0 0 dlycontrol4_in[4]
port 24 nsew
flabel metal3 s 0 10752 800 10872 0 FreeSans 600 0 0 0 dlycontrol4_in[5]
port 25 nsew
flabel metal3 s 0 960 800 1080 0 FreeSans 600 0 0 0 ena_in
port 26 nsew
flabel metal3 s 0 2184 800 2304 0 FreeSans 600 0 0 0 enable_dlycontrol_in
port 27 nsew
flabel metal3 s 33400 8848 34200 8968 0 FreeSans 600 0 0 0 ndecision_finish_in
port 28 nsew
flabel metal3 s 0 144 800 264 0 FreeSans 600 0 0 0 sample_n_in
port 29 nsew
flabel metal3 s 0 552 800 672 0 FreeSans 600 0 0 0 sample_n_out
port 30 nsew
flabel metal3 s 0 11160 800 11280 0 FreeSans 600 0 0 0 sample_p_in
port 31 nsew
flabel metal3 s 0 11568 800 11688 0 FreeSans 600 0 0 0 sample_p_out
port 32 nsew
flabel metal3 s 0 1368 800 1488 0 FreeSans 600 0 0 0 start_conv_in
port 33 nsew
rlabel metal2 s 29854 5967 29854 5967 4 clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[15\]
rlabel metal2 s 19734 5967 19734 5967 4 clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[7\]
rlabel metal2 s 22034 8653 22034 8653 4 clkgen.delay_155ns_3.bypass_enable_w\[2\]
rlabel metal2 s 17158 7718 17158 7718 4 clkgen.delay_155ns_3.genblk1\[3\].dly_binary.bypass_in
rlabel metal2 s 17158 7089 17158 7089 4 clkgen.delay_155ns_3.genblk1\[3\].dly_binary.signal_w\[3\]
rlabel metal2 s 18814 7055 18814 7055 4 clkgen.delay_155ns_3.genblk1\[3\].dly_binary.signal_w\[4\]
rlabel metal2 s 20838 7225 20838 7225 4 clkgen.delay_155ns_3.genblk1\[3\].dly_binary.signal_w\[8\]
rlabel metal2 s 20746 6545 20746 6545 4 dlycontrol3_in[1]
rlabel metal2 s 17250 6392 17250 6392 4 dlycontrol3_in[3]
rlabel metal2 s 27002 8755 27002 8755 4 dlycontrol4_in[2]
rlabel metal2 s 27738 10200 27738 10200 4 edgedetect.dly_315ns_1.bypass_enable_w\[1\]
rlabel metal2 s 26910 9622 26910 9622 4 edgedetect.dly_315ns_1.bypass_enable_w\[2\]
rlabel metal2 s 17618 7735 17618 7735 4 edgedetect.dly_315ns_1.genblk1\[0\].dly_binary.in
rlabel metal2 s 18630 7463 18630 7463 4 edgedetect.dly_315ns_1.genblk1\[0\].dly_binary.out
rlabel metal2 s 18998 8874 18998 8874 4 edgedetect.dly_315ns_1.genblk1\[1\].dly_binary.bypass_in
rlabel metal2 s 18538 7599 18538 7599 4 edgedetect.dly_315ns_1.genblk1\[1\].dly_binary.signal_w\[0\]
rlabel metal2 s 18078 11050 18078 11050 4 edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[11\]
rlabel metal2 s 17986 8891 17986 8891 4 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.bypass_in
rlabel metal2 s 19642 7769 19642 7769 4 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[0\]
rlabel metal2 s 20286 8143 20286 8143 4 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[11\]
rlabel metal2 s 24610 8483 24610 8483 4 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[15\]
rlabel metal2 s 27186 8704 27186 8704 4 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[16\]
rlabel metal2 s 20562 9639 20562 9639 4 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[19\]
rlabel metal2 s 26818 9792 26818 9792 4 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[24\]
rlabel metal2 s 28566 10285 28566 10285 4 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[25\]
rlabel metal2 s 27462 9299 27462 9299 4 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[29\]
rlabel metal2 s 31418 9520 31418 9520 4 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[30\]
rlabel metal2 s 32154 8704 32154 8704 4 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[31\]
rlabel metal2 s 17066 9163 17066 9163 4 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[32\]
flabel metal2 s 20944 496 21264 11472 0 FreeSans 2240 90 0 0 VDD
port 1 nsew
flabel metal2 s 30944 496 31264 11472 0 FreeSans 2240 90 0 0 VDD
port 1 nsew
flabel metal2 s 21604 496 21924 11472 0 FreeSans 2240 90 0 0 VSS
port 2 nsew
flabel metal2 s 31604 496 31924 11472 0 FreeSans 2240 90 0 0 VSS
port 2 nsew
rlabel metal2 s 6854 7548 6854 7548 4 clkgen.delay_155ns_3.genblk1\[2\].dly_binary.signal_w\[0\]
rlabel metal2 s 9430 7616 9430 7616 4 clkgen.delay_155ns_3.genblk1\[2\].dly_binary.signal_w\[2\]
rlabel metal2 s 16882 9316 16882 9316 4 edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.signal_w\[0\]
rlabel metal2 s 1978 8483 1978 8483 4 edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.signal_w\[1\]
rlabel metal2 s 12190 10319 12190 10319 4 edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.signal_w\[4\]
rlabel metal2 s 13110 10506 13110 10506 4 edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.signal_w\[5\]
rlabel metal2 s 15686 10336 15686 10336 4 edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.signal_w\[6\]
rlabel metal2 s 15962 10812 15962 10812 4 edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.signal_w\[7\]
rlabel metal2 s 16606 6477 16606 6477 4 clkgen.delay_155ns_2.genblk1\[3\].dly_binary.out
rlabel metal2 s 1610 10880 1610 10880 4 edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[1\]
rlabel metal2 s 6486 10863 6486 10863 4 edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[3\]
rlabel metal2 s 7314 11356 7314 11356 4 edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[4\]
rlabel metal2 s 9430 10880 9430 10880 4 edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[5\]
rlabel metal2 s 15042 10353 15042 10353 4 edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[9\]
rlabel metal2 s 14582 7463 14582 7463 4 clkgen.delay_155ns_3.genblk1\[3\].dly_binary.signal_w\[1\]
rlabel metal2 s 15502 7395 15502 7395 4 clkgen.delay_155ns_3.genblk1\[3\].dly_binary.signal_w\[2\]
rlabel metal2 s 7222 5899 7222 5899 4 clkgen.delay_155ns_2.genblk1\[3\].dly_binary.signal_w\[0\]
rlabel metal2 s 2162 8942 2162 8942 4 clkgen.delay_155ns_1.genblk1\[3\].dly_binary.signal_w\[8\]
rlabel metal2 s 12834 5950 12834 5950 4 clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[3\]
rlabel metal2 s 1610 6154 1610 6154 4 clkgen.enable_loop_in
rlabel metal2 s 4738 8721 4738 8721 4 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[1\]
rlabel metal2 s 14582 5916 14582 5916 4 clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[4\]
rlabel metal2 s 2254 7769 2254 7769 4 clkgen.delay_155ns_2.genblk1\[1\].dly_binary.bypass_in
rlabel metal2 s 14398 7344 14398 7344 4 clkgen.delay_155ns_3.bypass_enable_w\[1\]
rlabel metal2 s 4002 11101 4002 11101 4 dlycontrol4_in[4]
rlabel metal2 s 4094 11203 4094 11203 4 dlycontrol4_in[5]
rlabel metal2 s 16514 7871 16514 7871 4 clkgen.delay_155ns_2.genblk1\[3\].dly_binary.bypass_in
rlabel metal2 s 9614 8704 9614 8704 4 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[3\]
rlabel metal2 s 13294 8364 13294 8364 4 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[6\]
rlabel metal2 s 15042 8721 15042 8721 4 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[7\]
rlabel metal2 s 14030 8364 14030 8364 4 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[8\]
rlabel metal2 s 2622 7667 2622 7667 4 edgedetect.ena_in
flabel metal2 s 10944 496 11264 11472 0 FreeSans 2240 90 0 0 VDD
port 1 nsew
rlabel metal2 s 3450 6409 3450 6409 4 clkgen.delay_155ns_3.genblk1\[1\].dly_binary.bypass_in
rlabel metal2 s 6578 7259 6578 7259 4 clkgen.delay_155ns_3.genblk1\[1\].dly_binary.signal_w\[0\]
flabel metal2 s 11604 496 11924 11472 0 FreeSans 2240 90 0 0 VSS
port 2 nsew
rlabel metal2 s 8878 6800 8878 6800 4 clkgen.delay_155ns_3.genblk1\[1\].dly_binary.signal_w\[2\]
rlabel metal2 s 15870 8007 15870 8007 4 edgedetect.dly_315ns_1.genblk1\[0\].dly_binary.signal_w\[0\]
rlabel metal2 s 15042 544 15042 544 4 clkgen.delay_155ns_3.bypass_enable_w\[4\]
rlabel metal2 s 13662 4080 13662 4080 4 clkgen.delay_155ns_3.genblk1\[0\].dly_binary.in
rlabel metal2 s 4646 5695 4646 5695 4 clkgen.delay_155ns_3.genblk1\[0\].dly_binary.signal_w\[1\]
rlabel metal2 s 13202 510 13202 510 4 clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[16\]
rlabel metal2 s 1702 2176 1702 2176 4 clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[1\]
rlabel metal2 s 3358 1309 3358 1309 4 clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[2\]
rlabel metal2 s 1978 1071 1978 1071 4 clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[3\]
rlabel metal2 s 4462 1088 4462 1088 4 clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[4\]
rlabel metal2 s 6762 1326 6762 1326 4 clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[5\]
rlabel metal2 s 12282 1088 12282 1088 4 clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[9\]
rlabel metal2 s 1978 3859 1978 3859 4 clkgen.delay_155ns_2.genblk1\[0\].dly_binary.signal_w\[1\]
rlabel metal2 s 14122 510 14122 510 4 clkgen.delay_155ns_1.genblk1\[1\].dly_binary.out
rlabel metal2 s 15778 1445 15778 1445 4 clkgen.delay_155ns_2.genblk1\[1\].dly_binary.signal_w\[0\]
rlabel metal2 s 2254 4845 2254 4845 4 clkgen.delay_155ns_2.genblk1\[1\].dly_binary.signal_w\[1\]
rlabel metal2 s 15042 4369 15042 4369 4 clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[2\]
rlabel metal2 s 13386 3859 13386 3859 4 clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[3\]
rlabel metal2 s 6210 4845 6210 4845 4 clkgen.delay_155ns_2.genblk1\[1\].dly_binary.signal_w\[2\]
rlabel metal2 s 3634 1754 3634 1754 4 dlycontrol2_in[2]
rlabel metal2 s 15226 5389 15226 5389 4 clkgen.delay_155ns_2.genblk1\[2\].dly_binary.out
rlabel metal2 s 4830 3859 4830 3859 4 clkgen.delay_155ns_2.genblk1\[2\].dly_binary.signal_w\[1\]
rlabel metal2 s 15042 2329 15042 2329 4 clkgen.delay_155ns_1.genblk1\[2\].dly_binary.out
rlabel metal2 s 14030 408 14030 408 4 clkgen.delay_155ns_1.genblk1\[2\].dly_binary.signal_w\[0\]
rlabel metal2 s 12466 2754 12466 2754 4 clkgen.delay_155ns_1.genblk1\[2\].dly_binary.signal_w\[3\]
rlabel metal2 s 12282 5440 12282 5440 4 clkgen.delay_155ns_2.genblk1\[3\].dly_binary.signal_w\[4\]
rlabel metal2 s 14766 4335 14766 4335 4 clkgen.delay_155ns_2.genblk1\[3\].dly_binary.signal_w\[5\]
rlabel metal2 s 16606 3604 16606 3604 4 clkgen.delay_155ns_2.genblk1\[3\].dly_binary.signal_w\[6\]
rlabel metal2 s 13846 4488 13846 4488 4 clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[0\]
rlabel metal2 s 14950 3383 14950 3383 4 ndecision_finish_in
rlabel metal2 s 3726 4046 3726 4046 4 sample_n_1
rlabel metal2 s 1702 2873 1702 2873 4 sample_n_in
rlabel metal2 s 15686 2295 15686 2295 4 clkgen.delay_155ns_1.genblk1\[3\].dly_binary.signal_w\[0\]
rlabel metal2 s 12834 2176 12834 2176 4 clkgen.delay_155ns_1.genblk1\[3\].dly_binary.signal_w\[3\]
rlabel metal2 s 14168 2516 14168 2516 4 clkgen.delay_155ns_1.genblk1\[3\].dly_binary.signal_w\[4\]
rlabel metal2 s 13478 3553 13478 3553 4 clk_comp_out
rlabel metal2 s 13570 476 13570 476 4 clkgen.delay_155ns_1.genblk1\[4\].dly_binary.out
rlabel metal2 s 13386 1343 13386 1343 4 clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[12\]
rlabel metal2 s 17342 3060 17342 3060 4 dlycontrol1_in[3]
rlabel metal2 s 21390 1768 21390 1768 4 dlycontrol1_in[4]
rlabel metal2 s 25990 5457 25990 5457 4 clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[10\]
rlabel metal2 s 18538 4233 18538 4233 4 clkgen.delay_155ns_2.genblk1\[2\].dly_binary.signal_w\[0\]
rlabel metal2 s 32062 5797 32062 5797 4 clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[16\]
rlabel metal2 s 17802 2975 17802 2975 4 clkgen.delay_155ns_2.genblk1\[0\].dly_binary.bypass_in
rlabel metal2 s 19918 1632 19918 1632 4 clkgen.delay_155ns_2.genblk1\[0\].dly_binary.signal_w\[0\]
rlabel metal2 s 17250 3162 17250 3162 4 clkgen.delay_155ns_1.genblk1\[1\].dly_binary.signal_w\[0\]
rlabel metal2 s 21482 5457 21482 5457 4 clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[8\]
rlabel metal2 s 20746 816 20746 816 4 clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[0\]
rlabel metal2 s 20654 3587 20654 3587 4 clkgen.delay_155ns_1.genblk1\[3\].dly_binary.signal_w\[7\]
rlabel metal2 s 17158 3298 17158 3298 4 clkgen.delay_155ns_1.genblk1\[0\].dly_binary.out
rlabel metal2 s 32062 4352 32062 4352 4 clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[14\]
rlabel metal2 s 20838 1088 20838 1088 4 clkgen.delay_155ns_1.genblk1\[4\].dly_binary.bypass_in
rlabel metal2 s 19642 5440 19642 5440 4 clkgen.delay_155ns_2.genblk1\[3\].dly_binary.signal_w\[8\]
rlabel metal2 s 17894 3485 17894 3485 4 clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[4\]
rlabel metal2 s 25990 4369 25990 4369 4 clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[9\]
rlabel metal2 s 20286 1071 20286 1071 4 clkgen.delay_155ns_2.bypass_enable_w\[1\]
<< properties >>
string FIXED_BBOX 0 0 34200 12000
string GDS_END 1667446
string GDS_FILE adc_top.gds.gz
string GDS_START 927278
<< end >>
