magic
tech sky130A
magscale 1 2
timestamp 1695640753
<< metal3 >>
rect -7128 5932 -5556 5960
rect -7128 4708 -5640 5932
rect -5576 4708 -5556 5932
rect -7128 4680 -5556 4708
rect -5316 5932 -3744 5960
rect -5316 4708 -3828 5932
rect -3764 4708 -3744 5932
rect -5316 4680 -3744 4708
rect -3504 5932 -1932 5960
rect -3504 4708 -2016 5932
rect -1952 4708 -1932 5932
rect -3504 4680 -1932 4708
rect -1692 5932 -120 5960
rect -1692 4708 -204 5932
rect -140 4708 -120 5932
rect -1692 4680 -120 4708
rect 120 5932 1692 5960
rect 120 4708 1608 5932
rect 1672 4708 1692 5932
rect 120 4680 1692 4708
rect 1932 5932 3504 5960
rect 1932 4708 3420 5932
rect 3484 4708 3504 5932
rect 1932 4680 3504 4708
rect 3744 5932 5316 5960
rect 3744 4708 5232 5932
rect 5296 4708 5316 5932
rect 3744 4680 5316 4708
rect 5556 5932 7128 5960
rect 5556 4708 7044 5932
rect 7108 4708 7128 5932
rect 5556 4680 7128 4708
rect -7128 4412 -5556 4440
rect -7128 3188 -5640 4412
rect -5576 3188 -5556 4412
rect -7128 3160 -5556 3188
rect -5316 4412 -3744 4440
rect -5316 3188 -3828 4412
rect -3764 3188 -3744 4412
rect -5316 3160 -3744 3188
rect -3504 4412 -1932 4440
rect -3504 3188 -2016 4412
rect -1952 3188 -1932 4412
rect -3504 3160 -1932 3188
rect -1692 4412 -120 4440
rect -1692 3188 -204 4412
rect -140 3188 -120 4412
rect -1692 3160 -120 3188
rect 120 4412 1692 4440
rect 120 3188 1608 4412
rect 1672 3188 1692 4412
rect 120 3160 1692 3188
rect 1932 4412 3504 4440
rect 1932 3188 3420 4412
rect 3484 3188 3504 4412
rect 1932 3160 3504 3188
rect 3744 4412 5316 4440
rect 3744 3188 5232 4412
rect 5296 3188 5316 4412
rect 3744 3160 5316 3188
rect 5556 4412 7128 4440
rect 5556 3188 7044 4412
rect 7108 3188 7128 4412
rect 5556 3160 7128 3188
rect -7128 2892 -5556 2920
rect -7128 1668 -5640 2892
rect -5576 1668 -5556 2892
rect -7128 1640 -5556 1668
rect -5316 2892 -3744 2920
rect -5316 1668 -3828 2892
rect -3764 1668 -3744 2892
rect -5316 1640 -3744 1668
rect -3504 2892 -1932 2920
rect -3504 1668 -2016 2892
rect -1952 1668 -1932 2892
rect -3504 1640 -1932 1668
rect -1692 2892 -120 2920
rect -1692 1668 -204 2892
rect -140 1668 -120 2892
rect -1692 1640 -120 1668
rect 120 2892 1692 2920
rect 120 1668 1608 2892
rect 1672 1668 1692 2892
rect 120 1640 1692 1668
rect 1932 2892 3504 2920
rect 1932 1668 3420 2892
rect 3484 1668 3504 2892
rect 1932 1640 3504 1668
rect 3744 2892 5316 2920
rect 3744 1668 5232 2892
rect 5296 1668 5316 2892
rect 3744 1640 5316 1668
rect 5556 2892 7128 2920
rect 5556 1668 7044 2892
rect 7108 1668 7128 2892
rect 5556 1640 7128 1668
rect -7128 1372 -5556 1400
rect -7128 148 -5640 1372
rect -5576 148 -5556 1372
rect -7128 120 -5556 148
rect -5316 1372 -3744 1400
rect -5316 148 -3828 1372
rect -3764 148 -3744 1372
rect -5316 120 -3744 148
rect -3504 1372 -1932 1400
rect -3504 148 -2016 1372
rect -1952 148 -1932 1372
rect -3504 120 -1932 148
rect -1692 1372 -120 1400
rect -1692 148 -204 1372
rect -140 148 -120 1372
rect -1692 120 -120 148
rect 120 1372 1692 1400
rect 120 148 1608 1372
rect 1672 148 1692 1372
rect 120 120 1692 148
rect 1932 1372 3504 1400
rect 1932 148 3420 1372
rect 3484 148 3504 1372
rect 1932 120 3504 148
rect 3744 1372 5316 1400
rect 3744 148 5232 1372
rect 5296 148 5316 1372
rect 3744 120 5316 148
rect 5556 1372 7128 1400
rect 5556 148 7044 1372
rect 7108 148 7128 1372
rect 5556 120 7128 148
rect -7128 -148 -5556 -120
rect -7128 -1372 -5640 -148
rect -5576 -1372 -5556 -148
rect -7128 -1400 -5556 -1372
rect -5316 -148 -3744 -120
rect -5316 -1372 -3828 -148
rect -3764 -1372 -3744 -148
rect -5316 -1400 -3744 -1372
rect -3504 -148 -1932 -120
rect -3504 -1372 -2016 -148
rect -1952 -1372 -1932 -148
rect -3504 -1400 -1932 -1372
rect -1692 -148 -120 -120
rect -1692 -1372 -204 -148
rect -140 -1372 -120 -148
rect -1692 -1400 -120 -1372
rect 120 -148 1692 -120
rect 120 -1372 1608 -148
rect 1672 -1372 1692 -148
rect 120 -1400 1692 -1372
rect 1932 -148 3504 -120
rect 1932 -1372 3420 -148
rect 3484 -1372 3504 -148
rect 1932 -1400 3504 -1372
rect 3744 -148 5316 -120
rect 3744 -1372 5232 -148
rect 5296 -1372 5316 -148
rect 3744 -1400 5316 -1372
rect 5556 -148 7128 -120
rect 5556 -1372 7044 -148
rect 7108 -1372 7128 -148
rect 5556 -1400 7128 -1372
rect -7128 -1668 -5556 -1640
rect -7128 -2892 -5640 -1668
rect -5576 -2892 -5556 -1668
rect -7128 -2920 -5556 -2892
rect -5316 -1668 -3744 -1640
rect -5316 -2892 -3828 -1668
rect -3764 -2892 -3744 -1668
rect -5316 -2920 -3744 -2892
rect -3504 -1668 -1932 -1640
rect -3504 -2892 -2016 -1668
rect -1952 -2892 -1932 -1668
rect -3504 -2920 -1932 -2892
rect -1692 -1668 -120 -1640
rect -1692 -2892 -204 -1668
rect -140 -2892 -120 -1668
rect -1692 -2920 -120 -2892
rect 120 -1668 1692 -1640
rect 120 -2892 1608 -1668
rect 1672 -2892 1692 -1668
rect 120 -2920 1692 -2892
rect 1932 -1668 3504 -1640
rect 1932 -2892 3420 -1668
rect 3484 -2892 3504 -1668
rect 1932 -2920 3504 -2892
rect 3744 -1668 5316 -1640
rect 3744 -2892 5232 -1668
rect 5296 -2892 5316 -1668
rect 3744 -2920 5316 -2892
rect 5556 -1668 7128 -1640
rect 5556 -2892 7044 -1668
rect 7108 -2892 7128 -1668
rect 5556 -2920 7128 -2892
rect -7128 -3188 -5556 -3160
rect -7128 -4412 -5640 -3188
rect -5576 -4412 -5556 -3188
rect -7128 -4440 -5556 -4412
rect -5316 -3188 -3744 -3160
rect -5316 -4412 -3828 -3188
rect -3764 -4412 -3744 -3188
rect -5316 -4440 -3744 -4412
rect -3504 -3188 -1932 -3160
rect -3504 -4412 -2016 -3188
rect -1952 -4412 -1932 -3188
rect -3504 -4440 -1932 -4412
rect -1692 -3188 -120 -3160
rect -1692 -4412 -204 -3188
rect -140 -4412 -120 -3188
rect -1692 -4440 -120 -4412
rect 120 -3188 1692 -3160
rect 120 -4412 1608 -3188
rect 1672 -4412 1692 -3188
rect 120 -4440 1692 -4412
rect 1932 -3188 3504 -3160
rect 1932 -4412 3420 -3188
rect 3484 -4412 3504 -3188
rect 1932 -4440 3504 -4412
rect 3744 -3188 5316 -3160
rect 3744 -4412 5232 -3188
rect 5296 -4412 5316 -3188
rect 3744 -4440 5316 -4412
rect 5556 -3188 7128 -3160
rect 5556 -4412 7044 -3188
rect 7108 -4412 7128 -3188
rect 5556 -4440 7128 -4412
rect -7128 -4708 -5556 -4680
rect -7128 -5932 -5640 -4708
rect -5576 -5932 -5556 -4708
rect -7128 -5960 -5556 -5932
rect -5316 -4708 -3744 -4680
rect -5316 -5932 -3828 -4708
rect -3764 -5932 -3744 -4708
rect -5316 -5960 -3744 -5932
rect -3504 -4708 -1932 -4680
rect -3504 -5932 -2016 -4708
rect -1952 -5932 -1932 -4708
rect -3504 -5960 -1932 -5932
rect -1692 -4708 -120 -4680
rect -1692 -5932 -204 -4708
rect -140 -5932 -120 -4708
rect -1692 -5960 -120 -5932
rect 120 -4708 1692 -4680
rect 120 -5932 1608 -4708
rect 1672 -5932 1692 -4708
rect 120 -5960 1692 -5932
rect 1932 -4708 3504 -4680
rect 1932 -5932 3420 -4708
rect 3484 -5932 3504 -4708
rect 1932 -5960 3504 -5932
rect 3744 -4708 5316 -4680
rect 3744 -5932 5232 -4708
rect 5296 -5932 5316 -4708
rect 3744 -5960 5316 -5932
rect 5556 -4708 7128 -4680
rect 5556 -5932 7044 -4708
rect 7108 -5932 7128 -4708
rect 5556 -5960 7128 -5932
<< via3 >>
rect -5640 4708 -5576 5932
rect -3828 4708 -3764 5932
rect -2016 4708 -1952 5932
rect -204 4708 -140 5932
rect 1608 4708 1672 5932
rect 3420 4708 3484 5932
rect 5232 4708 5296 5932
rect 7044 4708 7108 5932
rect -5640 3188 -5576 4412
rect -3828 3188 -3764 4412
rect -2016 3188 -1952 4412
rect -204 3188 -140 4412
rect 1608 3188 1672 4412
rect 3420 3188 3484 4412
rect 5232 3188 5296 4412
rect 7044 3188 7108 4412
rect -5640 1668 -5576 2892
rect -3828 1668 -3764 2892
rect -2016 1668 -1952 2892
rect -204 1668 -140 2892
rect 1608 1668 1672 2892
rect 3420 1668 3484 2892
rect 5232 1668 5296 2892
rect 7044 1668 7108 2892
rect -5640 148 -5576 1372
rect -3828 148 -3764 1372
rect -2016 148 -1952 1372
rect -204 148 -140 1372
rect 1608 148 1672 1372
rect 3420 148 3484 1372
rect 5232 148 5296 1372
rect 7044 148 7108 1372
rect -5640 -1372 -5576 -148
rect -3828 -1372 -3764 -148
rect -2016 -1372 -1952 -148
rect -204 -1372 -140 -148
rect 1608 -1372 1672 -148
rect 3420 -1372 3484 -148
rect 5232 -1372 5296 -148
rect 7044 -1372 7108 -148
rect -5640 -2892 -5576 -1668
rect -3828 -2892 -3764 -1668
rect -2016 -2892 -1952 -1668
rect -204 -2892 -140 -1668
rect 1608 -2892 1672 -1668
rect 3420 -2892 3484 -1668
rect 5232 -2892 5296 -1668
rect 7044 -2892 7108 -1668
rect -5640 -4412 -5576 -3188
rect -3828 -4412 -3764 -3188
rect -2016 -4412 -1952 -3188
rect -204 -4412 -140 -3188
rect 1608 -4412 1672 -3188
rect 3420 -4412 3484 -3188
rect 5232 -4412 5296 -3188
rect 7044 -4412 7108 -3188
rect -5640 -5932 -5576 -4708
rect -3828 -5932 -3764 -4708
rect -2016 -5932 -1952 -4708
rect -204 -5932 -140 -4708
rect 1608 -5932 1672 -4708
rect 3420 -5932 3484 -4708
rect 5232 -5932 5296 -4708
rect 7044 -5932 7108 -4708
<< mimcap >>
rect -7088 5880 -5888 5920
rect -7088 4760 -7048 5880
rect -5928 4760 -5888 5880
rect -7088 4720 -5888 4760
rect -5276 5880 -4076 5920
rect -5276 4760 -5236 5880
rect -4116 4760 -4076 5880
rect -5276 4720 -4076 4760
rect -3464 5880 -2264 5920
rect -3464 4760 -3424 5880
rect -2304 4760 -2264 5880
rect -3464 4720 -2264 4760
rect -1652 5880 -452 5920
rect -1652 4760 -1612 5880
rect -492 4760 -452 5880
rect -1652 4720 -452 4760
rect 160 5880 1360 5920
rect 160 4760 200 5880
rect 1320 4760 1360 5880
rect 160 4720 1360 4760
rect 1972 5880 3172 5920
rect 1972 4760 2012 5880
rect 3132 4760 3172 5880
rect 1972 4720 3172 4760
rect 3784 5880 4984 5920
rect 3784 4760 3824 5880
rect 4944 4760 4984 5880
rect 3784 4720 4984 4760
rect 5596 5880 6796 5920
rect 5596 4760 5636 5880
rect 6756 4760 6796 5880
rect 5596 4720 6796 4760
rect -7088 4360 -5888 4400
rect -7088 3240 -7048 4360
rect -5928 3240 -5888 4360
rect -7088 3200 -5888 3240
rect -5276 4360 -4076 4400
rect -5276 3240 -5236 4360
rect -4116 3240 -4076 4360
rect -5276 3200 -4076 3240
rect -3464 4360 -2264 4400
rect -3464 3240 -3424 4360
rect -2304 3240 -2264 4360
rect -3464 3200 -2264 3240
rect -1652 4360 -452 4400
rect -1652 3240 -1612 4360
rect -492 3240 -452 4360
rect -1652 3200 -452 3240
rect 160 4360 1360 4400
rect 160 3240 200 4360
rect 1320 3240 1360 4360
rect 160 3200 1360 3240
rect 1972 4360 3172 4400
rect 1972 3240 2012 4360
rect 3132 3240 3172 4360
rect 1972 3200 3172 3240
rect 3784 4360 4984 4400
rect 3784 3240 3824 4360
rect 4944 3240 4984 4360
rect 3784 3200 4984 3240
rect 5596 4360 6796 4400
rect 5596 3240 5636 4360
rect 6756 3240 6796 4360
rect 5596 3200 6796 3240
rect -7088 2840 -5888 2880
rect -7088 1720 -7048 2840
rect -5928 1720 -5888 2840
rect -7088 1680 -5888 1720
rect -5276 2840 -4076 2880
rect -5276 1720 -5236 2840
rect -4116 1720 -4076 2840
rect -5276 1680 -4076 1720
rect -3464 2840 -2264 2880
rect -3464 1720 -3424 2840
rect -2304 1720 -2264 2840
rect -3464 1680 -2264 1720
rect -1652 2840 -452 2880
rect -1652 1720 -1612 2840
rect -492 1720 -452 2840
rect -1652 1680 -452 1720
rect 160 2840 1360 2880
rect 160 1720 200 2840
rect 1320 1720 1360 2840
rect 160 1680 1360 1720
rect 1972 2840 3172 2880
rect 1972 1720 2012 2840
rect 3132 1720 3172 2840
rect 1972 1680 3172 1720
rect 3784 2840 4984 2880
rect 3784 1720 3824 2840
rect 4944 1720 4984 2840
rect 3784 1680 4984 1720
rect 5596 2840 6796 2880
rect 5596 1720 5636 2840
rect 6756 1720 6796 2840
rect 5596 1680 6796 1720
rect -7088 1320 -5888 1360
rect -7088 200 -7048 1320
rect -5928 200 -5888 1320
rect -7088 160 -5888 200
rect -5276 1320 -4076 1360
rect -5276 200 -5236 1320
rect -4116 200 -4076 1320
rect -5276 160 -4076 200
rect -3464 1320 -2264 1360
rect -3464 200 -3424 1320
rect -2304 200 -2264 1320
rect -3464 160 -2264 200
rect -1652 1320 -452 1360
rect -1652 200 -1612 1320
rect -492 200 -452 1320
rect -1652 160 -452 200
rect 160 1320 1360 1360
rect 160 200 200 1320
rect 1320 200 1360 1320
rect 160 160 1360 200
rect 1972 1320 3172 1360
rect 1972 200 2012 1320
rect 3132 200 3172 1320
rect 1972 160 3172 200
rect 3784 1320 4984 1360
rect 3784 200 3824 1320
rect 4944 200 4984 1320
rect 3784 160 4984 200
rect 5596 1320 6796 1360
rect 5596 200 5636 1320
rect 6756 200 6796 1320
rect 5596 160 6796 200
rect -7088 -200 -5888 -160
rect -7088 -1320 -7048 -200
rect -5928 -1320 -5888 -200
rect -7088 -1360 -5888 -1320
rect -5276 -200 -4076 -160
rect -5276 -1320 -5236 -200
rect -4116 -1320 -4076 -200
rect -5276 -1360 -4076 -1320
rect -3464 -200 -2264 -160
rect -3464 -1320 -3424 -200
rect -2304 -1320 -2264 -200
rect -3464 -1360 -2264 -1320
rect -1652 -200 -452 -160
rect -1652 -1320 -1612 -200
rect -492 -1320 -452 -200
rect -1652 -1360 -452 -1320
rect 160 -200 1360 -160
rect 160 -1320 200 -200
rect 1320 -1320 1360 -200
rect 160 -1360 1360 -1320
rect 1972 -200 3172 -160
rect 1972 -1320 2012 -200
rect 3132 -1320 3172 -200
rect 1972 -1360 3172 -1320
rect 3784 -200 4984 -160
rect 3784 -1320 3824 -200
rect 4944 -1320 4984 -200
rect 3784 -1360 4984 -1320
rect 5596 -200 6796 -160
rect 5596 -1320 5636 -200
rect 6756 -1320 6796 -200
rect 5596 -1360 6796 -1320
rect -7088 -1720 -5888 -1680
rect -7088 -2840 -7048 -1720
rect -5928 -2840 -5888 -1720
rect -7088 -2880 -5888 -2840
rect -5276 -1720 -4076 -1680
rect -5276 -2840 -5236 -1720
rect -4116 -2840 -4076 -1720
rect -5276 -2880 -4076 -2840
rect -3464 -1720 -2264 -1680
rect -3464 -2840 -3424 -1720
rect -2304 -2840 -2264 -1720
rect -3464 -2880 -2264 -2840
rect -1652 -1720 -452 -1680
rect -1652 -2840 -1612 -1720
rect -492 -2840 -452 -1720
rect -1652 -2880 -452 -2840
rect 160 -1720 1360 -1680
rect 160 -2840 200 -1720
rect 1320 -2840 1360 -1720
rect 160 -2880 1360 -2840
rect 1972 -1720 3172 -1680
rect 1972 -2840 2012 -1720
rect 3132 -2840 3172 -1720
rect 1972 -2880 3172 -2840
rect 3784 -1720 4984 -1680
rect 3784 -2840 3824 -1720
rect 4944 -2840 4984 -1720
rect 3784 -2880 4984 -2840
rect 5596 -1720 6796 -1680
rect 5596 -2840 5636 -1720
rect 6756 -2840 6796 -1720
rect 5596 -2880 6796 -2840
rect -7088 -3240 -5888 -3200
rect -7088 -4360 -7048 -3240
rect -5928 -4360 -5888 -3240
rect -7088 -4400 -5888 -4360
rect -5276 -3240 -4076 -3200
rect -5276 -4360 -5236 -3240
rect -4116 -4360 -4076 -3240
rect -5276 -4400 -4076 -4360
rect -3464 -3240 -2264 -3200
rect -3464 -4360 -3424 -3240
rect -2304 -4360 -2264 -3240
rect -3464 -4400 -2264 -4360
rect -1652 -3240 -452 -3200
rect -1652 -4360 -1612 -3240
rect -492 -4360 -452 -3240
rect -1652 -4400 -452 -4360
rect 160 -3240 1360 -3200
rect 160 -4360 200 -3240
rect 1320 -4360 1360 -3240
rect 160 -4400 1360 -4360
rect 1972 -3240 3172 -3200
rect 1972 -4360 2012 -3240
rect 3132 -4360 3172 -3240
rect 1972 -4400 3172 -4360
rect 3784 -3240 4984 -3200
rect 3784 -4360 3824 -3240
rect 4944 -4360 4984 -3240
rect 3784 -4400 4984 -4360
rect 5596 -3240 6796 -3200
rect 5596 -4360 5636 -3240
rect 6756 -4360 6796 -3240
rect 5596 -4400 6796 -4360
rect -7088 -4760 -5888 -4720
rect -7088 -5880 -7048 -4760
rect -5928 -5880 -5888 -4760
rect -7088 -5920 -5888 -5880
rect -5276 -4760 -4076 -4720
rect -5276 -5880 -5236 -4760
rect -4116 -5880 -4076 -4760
rect -5276 -5920 -4076 -5880
rect -3464 -4760 -2264 -4720
rect -3464 -5880 -3424 -4760
rect -2304 -5880 -2264 -4760
rect -3464 -5920 -2264 -5880
rect -1652 -4760 -452 -4720
rect -1652 -5880 -1612 -4760
rect -492 -5880 -452 -4760
rect -1652 -5920 -452 -5880
rect 160 -4760 1360 -4720
rect 160 -5880 200 -4760
rect 1320 -5880 1360 -4760
rect 160 -5920 1360 -5880
rect 1972 -4760 3172 -4720
rect 1972 -5880 2012 -4760
rect 3132 -5880 3172 -4760
rect 1972 -5920 3172 -5880
rect 3784 -4760 4984 -4720
rect 3784 -5880 3824 -4760
rect 4944 -5880 4984 -4760
rect 3784 -5920 4984 -5880
rect 5596 -4760 6796 -4720
rect 5596 -5880 5636 -4760
rect 6756 -5880 6796 -4760
rect 5596 -5920 6796 -5880
<< mimcapcontact >>
rect -7048 4760 -5928 5880
rect -5236 4760 -4116 5880
rect -3424 4760 -2304 5880
rect -1612 4760 -492 5880
rect 200 4760 1320 5880
rect 2012 4760 3132 5880
rect 3824 4760 4944 5880
rect 5636 4760 6756 5880
rect -7048 3240 -5928 4360
rect -5236 3240 -4116 4360
rect -3424 3240 -2304 4360
rect -1612 3240 -492 4360
rect 200 3240 1320 4360
rect 2012 3240 3132 4360
rect 3824 3240 4944 4360
rect 5636 3240 6756 4360
rect -7048 1720 -5928 2840
rect -5236 1720 -4116 2840
rect -3424 1720 -2304 2840
rect -1612 1720 -492 2840
rect 200 1720 1320 2840
rect 2012 1720 3132 2840
rect 3824 1720 4944 2840
rect 5636 1720 6756 2840
rect -7048 200 -5928 1320
rect -5236 200 -4116 1320
rect -3424 200 -2304 1320
rect -1612 200 -492 1320
rect 200 200 1320 1320
rect 2012 200 3132 1320
rect 3824 200 4944 1320
rect 5636 200 6756 1320
rect -7048 -1320 -5928 -200
rect -5236 -1320 -4116 -200
rect -3424 -1320 -2304 -200
rect -1612 -1320 -492 -200
rect 200 -1320 1320 -200
rect 2012 -1320 3132 -200
rect 3824 -1320 4944 -200
rect 5636 -1320 6756 -200
rect -7048 -2840 -5928 -1720
rect -5236 -2840 -4116 -1720
rect -3424 -2840 -2304 -1720
rect -1612 -2840 -492 -1720
rect 200 -2840 1320 -1720
rect 2012 -2840 3132 -1720
rect 3824 -2840 4944 -1720
rect 5636 -2840 6756 -1720
rect -7048 -4360 -5928 -3240
rect -5236 -4360 -4116 -3240
rect -3424 -4360 -2304 -3240
rect -1612 -4360 -492 -3240
rect 200 -4360 1320 -3240
rect 2012 -4360 3132 -3240
rect 3824 -4360 4944 -3240
rect 5636 -4360 6756 -3240
rect -7048 -5880 -5928 -4760
rect -5236 -5880 -4116 -4760
rect -3424 -5880 -2304 -4760
rect -1612 -5880 -492 -4760
rect 200 -5880 1320 -4760
rect 2012 -5880 3132 -4760
rect 3824 -5880 4944 -4760
rect 5636 -5880 6756 -4760
<< metal4 >>
rect -6540 5881 -6436 6080
rect -5660 5932 -5556 6080
rect -7049 5880 -5927 5881
rect -7049 4760 -7048 5880
rect -5928 4760 -5927 5880
rect -7049 4759 -5927 4760
rect -6540 4361 -6436 4759
rect -5660 4708 -5640 5932
rect -5576 4708 -5556 5932
rect -4728 5881 -4624 6080
rect -3848 5932 -3744 6080
rect -5237 5880 -4115 5881
rect -5237 4760 -5236 5880
rect -4116 4760 -4115 5880
rect -5237 4759 -4115 4760
rect -5660 4412 -5556 4708
rect -7049 4360 -5927 4361
rect -7049 3240 -7048 4360
rect -5928 3240 -5927 4360
rect -7049 3239 -5927 3240
rect -6540 2841 -6436 3239
rect -5660 3188 -5640 4412
rect -5576 3188 -5556 4412
rect -4728 4361 -4624 4759
rect -3848 4708 -3828 5932
rect -3764 4708 -3744 5932
rect -2916 5881 -2812 6080
rect -2036 5932 -1932 6080
rect -3425 5880 -2303 5881
rect -3425 4760 -3424 5880
rect -2304 4760 -2303 5880
rect -3425 4759 -2303 4760
rect -3848 4412 -3744 4708
rect -5237 4360 -4115 4361
rect -5237 3240 -5236 4360
rect -4116 3240 -4115 4360
rect -5237 3239 -4115 3240
rect -5660 2892 -5556 3188
rect -7049 2840 -5927 2841
rect -7049 1720 -7048 2840
rect -5928 1720 -5927 2840
rect -7049 1719 -5927 1720
rect -6540 1321 -6436 1719
rect -5660 1668 -5640 2892
rect -5576 1668 -5556 2892
rect -4728 2841 -4624 3239
rect -3848 3188 -3828 4412
rect -3764 3188 -3744 4412
rect -2916 4361 -2812 4759
rect -2036 4708 -2016 5932
rect -1952 4708 -1932 5932
rect -1104 5881 -1000 6080
rect -224 5932 -120 6080
rect -1613 5880 -491 5881
rect -1613 4760 -1612 5880
rect -492 4760 -491 5880
rect -1613 4759 -491 4760
rect -2036 4412 -1932 4708
rect -3425 4360 -2303 4361
rect -3425 3240 -3424 4360
rect -2304 3240 -2303 4360
rect -3425 3239 -2303 3240
rect -3848 2892 -3744 3188
rect -5237 2840 -4115 2841
rect -5237 1720 -5236 2840
rect -4116 1720 -4115 2840
rect -5237 1719 -4115 1720
rect -5660 1372 -5556 1668
rect -7049 1320 -5927 1321
rect -7049 200 -7048 1320
rect -5928 200 -5927 1320
rect -7049 199 -5927 200
rect -6540 -199 -6436 199
rect -5660 148 -5640 1372
rect -5576 148 -5556 1372
rect -4728 1321 -4624 1719
rect -3848 1668 -3828 2892
rect -3764 1668 -3744 2892
rect -2916 2841 -2812 3239
rect -2036 3188 -2016 4412
rect -1952 3188 -1932 4412
rect -1104 4361 -1000 4759
rect -224 4708 -204 5932
rect -140 4708 -120 5932
rect 708 5881 812 6080
rect 1588 5932 1692 6080
rect 199 5880 1321 5881
rect 199 4760 200 5880
rect 1320 4760 1321 5880
rect 199 4759 1321 4760
rect -224 4412 -120 4708
rect -1613 4360 -491 4361
rect -1613 3240 -1612 4360
rect -492 3240 -491 4360
rect -1613 3239 -491 3240
rect -2036 2892 -1932 3188
rect -3425 2840 -2303 2841
rect -3425 1720 -3424 2840
rect -2304 1720 -2303 2840
rect -3425 1719 -2303 1720
rect -3848 1372 -3744 1668
rect -5237 1320 -4115 1321
rect -5237 200 -5236 1320
rect -4116 200 -4115 1320
rect -5237 199 -4115 200
rect -5660 -148 -5556 148
rect -7049 -200 -5927 -199
rect -7049 -1320 -7048 -200
rect -5928 -1320 -5927 -200
rect -7049 -1321 -5927 -1320
rect -6540 -1719 -6436 -1321
rect -5660 -1372 -5640 -148
rect -5576 -1372 -5556 -148
rect -4728 -199 -4624 199
rect -3848 148 -3828 1372
rect -3764 148 -3744 1372
rect -2916 1321 -2812 1719
rect -2036 1668 -2016 2892
rect -1952 1668 -1932 2892
rect -1104 2841 -1000 3239
rect -224 3188 -204 4412
rect -140 3188 -120 4412
rect 708 4361 812 4759
rect 1588 4708 1608 5932
rect 1672 4708 1692 5932
rect 2520 5881 2624 6080
rect 3400 5932 3504 6080
rect 2011 5880 3133 5881
rect 2011 4760 2012 5880
rect 3132 4760 3133 5880
rect 2011 4759 3133 4760
rect 1588 4412 1692 4708
rect 199 4360 1321 4361
rect 199 3240 200 4360
rect 1320 3240 1321 4360
rect 199 3239 1321 3240
rect -224 2892 -120 3188
rect -1613 2840 -491 2841
rect -1613 1720 -1612 2840
rect -492 1720 -491 2840
rect -1613 1719 -491 1720
rect -2036 1372 -1932 1668
rect -3425 1320 -2303 1321
rect -3425 200 -3424 1320
rect -2304 200 -2303 1320
rect -3425 199 -2303 200
rect -3848 -148 -3744 148
rect -5237 -200 -4115 -199
rect -5237 -1320 -5236 -200
rect -4116 -1320 -4115 -200
rect -5237 -1321 -4115 -1320
rect -5660 -1668 -5556 -1372
rect -7049 -1720 -5927 -1719
rect -7049 -2840 -7048 -1720
rect -5928 -2840 -5927 -1720
rect -7049 -2841 -5927 -2840
rect -6540 -3239 -6436 -2841
rect -5660 -2892 -5640 -1668
rect -5576 -2892 -5556 -1668
rect -4728 -1719 -4624 -1321
rect -3848 -1372 -3828 -148
rect -3764 -1372 -3744 -148
rect -2916 -199 -2812 199
rect -2036 148 -2016 1372
rect -1952 148 -1932 1372
rect -1104 1321 -1000 1719
rect -224 1668 -204 2892
rect -140 1668 -120 2892
rect 708 2841 812 3239
rect 1588 3188 1608 4412
rect 1672 3188 1692 4412
rect 2520 4361 2624 4759
rect 3400 4708 3420 5932
rect 3484 4708 3504 5932
rect 4332 5881 4436 6080
rect 5212 5932 5316 6080
rect 3823 5880 4945 5881
rect 3823 4760 3824 5880
rect 4944 4760 4945 5880
rect 3823 4759 4945 4760
rect 3400 4412 3504 4708
rect 2011 4360 3133 4361
rect 2011 3240 2012 4360
rect 3132 3240 3133 4360
rect 2011 3239 3133 3240
rect 1588 2892 1692 3188
rect 199 2840 1321 2841
rect 199 1720 200 2840
rect 1320 1720 1321 2840
rect 199 1719 1321 1720
rect -224 1372 -120 1668
rect -1613 1320 -491 1321
rect -1613 200 -1612 1320
rect -492 200 -491 1320
rect -1613 199 -491 200
rect -2036 -148 -1932 148
rect -3425 -200 -2303 -199
rect -3425 -1320 -3424 -200
rect -2304 -1320 -2303 -200
rect -3425 -1321 -2303 -1320
rect -3848 -1668 -3744 -1372
rect -5237 -1720 -4115 -1719
rect -5237 -2840 -5236 -1720
rect -4116 -2840 -4115 -1720
rect -5237 -2841 -4115 -2840
rect -5660 -3188 -5556 -2892
rect -7049 -3240 -5927 -3239
rect -7049 -4360 -7048 -3240
rect -5928 -4360 -5927 -3240
rect -7049 -4361 -5927 -4360
rect -6540 -4759 -6436 -4361
rect -5660 -4412 -5640 -3188
rect -5576 -4412 -5556 -3188
rect -4728 -3239 -4624 -2841
rect -3848 -2892 -3828 -1668
rect -3764 -2892 -3744 -1668
rect -2916 -1719 -2812 -1321
rect -2036 -1372 -2016 -148
rect -1952 -1372 -1932 -148
rect -1104 -199 -1000 199
rect -224 148 -204 1372
rect -140 148 -120 1372
rect 708 1321 812 1719
rect 1588 1668 1608 2892
rect 1672 1668 1692 2892
rect 2520 2841 2624 3239
rect 3400 3188 3420 4412
rect 3484 3188 3504 4412
rect 4332 4361 4436 4759
rect 5212 4708 5232 5932
rect 5296 4708 5316 5932
rect 6144 5881 6248 6080
rect 7024 5932 7128 6080
rect 5635 5880 6757 5881
rect 5635 4760 5636 5880
rect 6756 4760 6757 5880
rect 5635 4759 6757 4760
rect 5212 4412 5316 4708
rect 3823 4360 4945 4361
rect 3823 3240 3824 4360
rect 4944 3240 4945 4360
rect 3823 3239 4945 3240
rect 3400 2892 3504 3188
rect 2011 2840 3133 2841
rect 2011 1720 2012 2840
rect 3132 1720 3133 2840
rect 2011 1719 3133 1720
rect 1588 1372 1692 1668
rect 199 1320 1321 1321
rect 199 200 200 1320
rect 1320 200 1321 1320
rect 199 199 1321 200
rect -224 -148 -120 148
rect -1613 -200 -491 -199
rect -1613 -1320 -1612 -200
rect -492 -1320 -491 -200
rect -1613 -1321 -491 -1320
rect -2036 -1668 -1932 -1372
rect -3425 -1720 -2303 -1719
rect -3425 -2840 -3424 -1720
rect -2304 -2840 -2303 -1720
rect -3425 -2841 -2303 -2840
rect -3848 -3188 -3744 -2892
rect -5237 -3240 -4115 -3239
rect -5237 -4360 -5236 -3240
rect -4116 -4360 -4115 -3240
rect -5237 -4361 -4115 -4360
rect -5660 -4708 -5556 -4412
rect -7049 -4760 -5927 -4759
rect -7049 -5880 -7048 -4760
rect -5928 -5880 -5927 -4760
rect -7049 -5881 -5927 -5880
rect -6540 -6080 -6436 -5881
rect -5660 -5932 -5640 -4708
rect -5576 -5932 -5556 -4708
rect -4728 -4759 -4624 -4361
rect -3848 -4412 -3828 -3188
rect -3764 -4412 -3744 -3188
rect -2916 -3239 -2812 -2841
rect -2036 -2892 -2016 -1668
rect -1952 -2892 -1932 -1668
rect -1104 -1719 -1000 -1321
rect -224 -1372 -204 -148
rect -140 -1372 -120 -148
rect 708 -199 812 199
rect 1588 148 1608 1372
rect 1672 148 1692 1372
rect 2520 1321 2624 1719
rect 3400 1668 3420 2892
rect 3484 1668 3504 2892
rect 4332 2841 4436 3239
rect 5212 3188 5232 4412
rect 5296 3188 5316 4412
rect 6144 4361 6248 4759
rect 7024 4708 7044 5932
rect 7108 4708 7128 5932
rect 7024 4412 7128 4708
rect 5635 4360 6757 4361
rect 5635 3240 5636 4360
rect 6756 3240 6757 4360
rect 5635 3239 6757 3240
rect 5212 2892 5316 3188
rect 3823 2840 4945 2841
rect 3823 1720 3824 2840
rect 4944 1720 4945 2840
rect 3823 1719 4945 1720
rect 3400 1372 3504 1668
rect 2011 1320 3133 1321
rect 2011 200 2012 1320
rect 3132 200 3133 1320
rect 2011 199 3133 200
rect 1588 -148 1692 148
rect 199 -200 1321 -199
rect 199 -1320 200 -200
rect 1320 -1320 1321 -200
rect 199 -1321 1321 -1320
rect -224 -1668 -120 -1372
rect -1613 -1720 -491 -1719
rect -1613 -2840 -1612 -1720
rect -492 -2840 -491 -1720
rect -1613 -2841 -491 -2840
rect -2036 -3188 -1932 -2892
rect -3425 -3240 -2303 -3239
rect -3425 -4360 -3424 -3240
rect -2304 -4360 -2303 -3240
rect -3425 -4361 -2303 -4360
rect -3848 -4708 -3744 -4412
rect -5237 -4760 -4115 -4759
rect -5237 -5880 -5236 -4760
rect -4116 -5880 -4115 -4760
rect -5237 -5881 -4115 -5880
rect -5660 -6080 -5556 -5932
rect -4728 -6080 -4624 -5881
rect -3848 -5932 -3828 -4708
rect -3764 -5932 -3744 -4708
rect -2916 -4759 -2812 -4361
rect -2036 -4412 -2016 -3188
rect -1952 -4412 -1932 -3188
rect -1104 -3239 -1000 -2841
rect -224 -2892 -204 -1668
rect -140 -2892 -120 -1668
rect 708 -1719 812 -1321
rect 1588 -1372 1608 -148
rect 1672 -1372 1692 -148
rect 2520 -199 2624 199
rect 3400 148 3420 1372
rect 3484 148 3504 1372
rect 4332 1321 4436 1719
rect 5212 1668 5232 2892
rect 5296 1668 5316 2892
rect 6144 2841 6248 3239
rect 7024 3188 7044 4412
rect 7108 3188 7128 4412
rect 7024 2892 7128 3188
rect 5635 2840 6757 2841
rect 5635 1720 5636 2840
rect 6756 1720 6757 2840
rect 5635 1719 6757 1720
rect 5212 1372 5316 1668
rect 3823 1320 4945 1321
rect 3823 200 3824 1320
rect 4944 200 4945 1320
rect 3823 199 4945 200
rect 3400 -148 3504 148
rect 2011 -200 3133 -199
rect 2011 -1320 2012 -200
rect 3132 -1320 3133 -200
rect 2011 -1321 3133 -1320
rect 1588 -1668 1692 -1372
rect 199 -1720 1321 -1719
rect 199 -2840 200 -1720
rect 1320 -2840 1321 -1720
rect 199 -2841 1321 -2840
rect -224 -3188 -120 -2892
rect -1613 -3240 -491 -3239
rect -1613 -4360 -1612 -3240
rect -492 -4360 -491 -3240
rect -1613 -4361 -491 -4360
rect -2036 -4708 -1932 -4412
rect -3425 -4760 -2303 -4759
rect -3425 -5880 -3424 -4760
rect -2304 -5880 -2303 -4760
rect -3425 -5881 -2303 -5880
rect -3848 -6080 -3744 -5932
rect -2916 -6080 -2812 -5881
rect -2036 -5932 -2016 -4708
rect -1952 -5932 -1932 -4708
rect -1104 -4759 -1000 -4361
rect -224 -4412 -204 -3188
rect -140 -4412 -120 -3188
rect 708 -3239 812 -2841
rect 1588 -2892 1608 -1668
rect 1672 -2892 1692 -1668
rect 2520 -1719 2624 -1321
rect 3400 -1372 3420 -148
rect 3484 -1372 3504 -148
rect 4332 -199 4436 199
rect 5212 148 5232 1372
rect 5296 148 5316 1372
rect 6144 1321 6248 1719
rect 7024 1668 7044 2892
rect 7108 1668 7128 2892
rect 7024 1372 7128 1668
rect 5635 1320 6757 1321
rect 5635 200 5636 1320
rect 6756 200 6757 1320
rect 5635 199 6757 200
rect 5212 -148 5316 148
rect 3823 -200 4945 -199
rect 3823 -1320 3824 -200
rect 4944 -1320 4945 -200
rect 3823 -1321 4945 -1320
rect 3400 -1668 3504 -1372
rect 2011 -1720 3133 -1719
rect 2011 -2840 2012 -1720
rect 3132 -2840 3133 -1720
rect 2011 -2841 3133 -2840
rect 1588 -3188 1692 -2892
rect 199 -3240 1321 -3239
rect 199 -4360 200 -3240
rect 1320 -4360 1321 -3240
rect 199 -4361 1321 -4360
rect -224 -4708 -120 -4412
rect -1613 -4760 -491 -4759
rect -1613 -5880 -1612 -4760
rect -492 -5880 -491 -4760
rect -1613 -5881 -491 -5880
rect -2036 -6080 -1932 -5932
rect -1104 -6080 -1000 -5881
rect -224 -5932 -204 -4708
rect -140 -5932 -120 -4708
rect 708 -4759 812 -4361
rect 1588 -4412 1608 -3188
rect 1672 -4412 1692 -3188
rect 2520 -3239 2624 -2841
rect 3400 -2892 3420 -1668
rect 3484 -2892 3504 -1668
rect 4332 -1719 4436 -1321
rect 5212 -1372 5232 -148
rect 5296 -1372 5316 -148
rect 6144 -199 6248 199
rect 7024 148 7044 1372
rect 7108 148 7128 1372
rect 7024 -148 7128 148
rect 5635 -200 6757 -199
rect 5635 -1320 5636 -200
rect 6756 -1320 6757 -200
rect 5635 -1321 6757 -1320
rect 5212 -1668 5316 -1372
rect 3823 -1720 4945 -1719
rect 3823 -2840 3824 -1720
rect 4944 -2840 4945 -1720
rect 3823 -2841 4945 -2840
rect 3400 -3188 3504 -2892
rect 2011 -3240 3133 -3239
rect 2011 -4360 2012 -3240
rect 3132 -4360 3133 -3240
rect 2011 -4361 3133 -4360
rect 1588 -4708 1692 -4412
rect 199 -4760 1321 -4759
rect 199 -5880 200 -4760
rect 1320 -5880 1321 -4760
rect 199 -5881 1321 -5880
rect -224 -6080 -120 -5932
rect 708 -6080 812 -5881
rect 1588 -5932 1608 -4708
rect 1672 -5932 1692 -4708
rect 2520 -4759 2624 -4361
rect 3400 -4412 3420 -3188
rect 3484 -4412 3504 -3188
rect 4332 -3239 4436 -2841
rect 5212 -2892 5232 -1668
rect 5296 -2892 5316 -1668
rect 6144 -1719 6248 -1321
rect 7024 -1372 7044 -148
rect 7108 -1372 7128 -148
rect 7024 -1668 7128 -1372
rect 5635 -1720 6757 -1719
rect 5635 -2840 5636 -1720
rect 6756 -2840 6757 -1720
rect 5635 -2841 6757 -2840
rect 5212 -3188 5316 -2892
rect 3823 -3240 4945 -3239
rect 3823 -4360 3824 -3240
rect 4944 -4360 4945 -3240
rect 3823 -4361 4945 -4360
rect 3400 -4708 3504 -4412
rect 2011 -4760 3133 -4759
rect 2011 -5880 2012 -4760
rect 3132 -5880 3133 -4760
rect 2011 -5881 3133 -5880
rect 1588 -6080 1692 -5932
rect 2520 -6080 2624 -5881
rect 3400 -5932 3420 -4708
rect 3484 -5932 3504 -4708
rect 4332 -4759 4436 -4361
rect 5212 -4412 5232 -3188
rect 5296 -4412 5316 -3188
rect 6144 -3239 6248 -2841
rect 7024 -2892 7044 -1668
rect 7108 -2892 7128 -1668
rect 7024 -3188 7128 -2892
rect 5635 -3240 6757 -3239
rect 5635 -4360 5636 -3240
rect 6756 -4360 6757 -3240
rect 5635 -4361 6757 -4360
rect 5212 -4708 5316 -4412
rect 3823 -4760 4945 -4759
rect 3823 -5880 3824 -4760
rect 4944 -5880 4945 -4760
rect 3823 -5881 4945 -5880
rect 3400 -6080 3504 -5932
rect 4332 -6080 4436 -5881
rect 5212 -5932 5232 -4708
rect 5296 -5932 5316 -4708
rect 6144 -4759 6248 -4361
rect 7024 -4412 7044 -3188
rect 7108 -4412 7128 -3188
rect 7024 -4708 7128 -4412
rect 5635 -4760 6757 -4759
rect 5635 -5880 5636 -4760
rect 6756 -5880 6757 -4760
rect 5635 -5881 6757 -5880
rect 5212 -6080 5316 -5932
rect 6144 -6080 6248 -5881
rect 7024 -5932 7044 -4708
rect 7108 -5932 7128 -4708
rect 7024 -6080 7128 -5932
<< properties >>
string FIXED_BBOX 5556 4680 6836 5960
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 6 l 6 val 76.56 carea 2.00 cperi 0.19 nx 8 ny 8 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
