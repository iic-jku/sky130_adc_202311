magic
tech sky130A
magscale 1 2
timestamp 1699972208
<< nwell >>
rect -42 962 872 1260
rect 876 964 992 1036
rect 1726 964 1842 1036
rect -42 943 686 962
rect 102 857 686 943
rect 102 842 722 857
rect 836 842 872 962
rect 102 622 872 842
rect 1846 962 2760 1260
rect 1846 842 1882 962
rect 2032 943 2760 962
rect 2032 857 2616 943
rect 1996 842 2616 857
rect 1846 622 2616 842
rect 102 -381 2760 -334
rect 102 -431 2616 -381
rect 102 -666 2452 -431
<< pwell >>
rect -42 286 690 622
rect 2028 286 2760 622
rect -42 176 2760 286
rect -42 156 1576 176
rect -42 90 1642 156
rect -42 58 1576 90
rect -42 -14 1642 58
rect 1654 -14 2760 176
rect -42 -334 2760 -14
<< pdiff >>
rect 924 970 976 1030
rect 1742 970 1794 1030
<< nsubdiff >>
rect 839 -398 961 -373
rect 839 -619 961 -592
rect 1755 -398 1877 -373
rect 1755 -619 1877 -592
<< nsubdiffcont >>
rect 839 -592 961 -398
rect 1755 -592 1877 -398
<< locali >>
rect 686 953 836 1040
rect 526 857 836 953
rect 1882 953 2032 1040
rect 722 842 836 857
rect 1226 840 1492 922
rect 1882 908 2192 953
rect 1882 866 1944 908
rect 2012 866 2192 908
rect 1882 857 2192 866
rect 1882 842 1996 857
rect 722 756 930 798
rect 1788 756 1996 798
rect 60 378 206 576
rect 722 450 922 492
rect 1796 450 1996 492
rect 526 312 836 412
rect 722 212 836 312
rect 1164 212 1554 412
rect 1882 312 2192 412
rect 2512 378 2658 576
rect 1882 212 1996 312
rect 1128 -57 1559 38
rect 60 -289 206 -91
rect 2512 -289 2658 -91
rect 839 -398 961 -364
rect 1755 -398 1877 -364
rect 839 -601 961 -592
rect 1755 -601 1877 -592
rect 528 -635 2219 -601
<< viali >>
rect 1944 866 2012 908
rect 414 740 488 778
rect 2230 740 2304 778
rect 330 578 364 612
rect 2356 576 2390 610
rect 978 120 1012 154
rect 1086 120 1120 154
rect 1598 120 1632 154
rect 1706 120 1740 154
rect 332 -324 366 -290
rect 1202 -324 1236 -290
rect 1342 -328 1378 -292
rect 2352 -324 2386 -290
rect 412 -424 446 -388
rect 1494 -492 1530 -456
rect 2272 -424 2306 -388
<< metal1 >>
rect 310 1590 382 1744
rect 310 1506 316 1590
rect 376 1506 382 1590
rect 310 1077 382 1506
rect 686 1734 758 1744
rect 686 1650 692 1734
rect 752 1650 758 1734
rect 310 1025 319 1077
rect 371 1025 382 1077
rect 564 1134 638 1140
rect 564 1078 570 1134
rect 632 1078 638 1134
rect 564 1072 638 1078
rect 310 1019 382 1025
rect 570 784 638 1072
rect 686 1026 758 1650
rect 1014 1134 1082 1140
rect 1014 1078 1020 1134
rect 1076 1078 1082 1134
rect 1014 1072 1082 1078
rect 686 974 696 1026
rect 748 974 758 1026
rect 686 964 758 974
rect 918 1030 982 1036
rect 918 970 924 1030
rect 976 970 982 1030
rect 918 964 982 970
rect 1114 1030 1178 1036
rect 1114 970 1120 1030
rect 1172 970 1178 1030
rect 1114 964 1178 970
rect 1026 912 1090 918
rect 1026 852 1032 912
rect 1084 852 1090 912
rect 1026 846 1090 852
rect 1323 908 1395 1668
rect 1960 1302 2032 1744
rect 1960 1218 1966 1302
rect 2026 1218 2032 1302
rect 1636 1134 1704 1140
rect 1636 1078 1642 1134
rect 1698 1078 1704 1134
rect 1636 1072 1704 1078
rect 1540 1030 1604 1036
rect 1540 970 1546 1030
rect 1598 970 1604 1030
rect 1540 964 1604 970
rect 1736 1030 1800 1036
rect 1736 970 1742 1030
rect 1794 970 1800 1030
rect 1736 964 1800 970
rect 1960 1026 2032 1218
rect 2340 1446 2412 1744
rect 2340 1362 2346 1446
rect 2406 1362 2412 1446
rect 1960 974 1970 1026
rect 2022 974 2032 1026
rect 1960 964 2032 974
rect 2080 1134 2154 1140
rect 2080 1078 2086 1134
rect 2148 1078 2154 1134
rect 2080 1072 2154 1078
rect 2340 1073 2412 1362
rect 1323 856 1333 908
rect 1385 856 1395 908
rect 1323 846 1395 856
rect 1628 912 1692 918
rect 1628 852 1634 912
rect 1686 852 1692 912
rect 1930 914 2026 922
rect 1930 860 1938 914
rect 2018 860 2026 914
rect 1930 854 2026 860
rect 1628 846 1692 852
rect 1026 842 1072 846
rect 402 778 638 784
rect 402 740 414 778
rect 488 740 638 778
rect 402 734 638 740
rect 310 621 382 627
rect 310 569 321 621
rect 373 569 382 621
rect 310 560 382 569
rect 928 412 976 842
rect 1024 410 1072 842
rect 1646 842 1692 846
rect 1646 410 1694 842
rect 1742 412 1790 842
rect 2080 784 2148 1072
rect 2340 1021 2349 1073
rect 2401 1021 2412 1073
rect 2340 1015 2412 1021
rect 2722 857 2760 953
rect 2080 778 2316 784
rect 2080 740 2230 778
rect 2304 740 2316 778
rect 2080 734 2316 740
rect 2340 617 2411 623
rect 2340 565 2351 617
rect 2403 565 2411 617
rect 2340 559 2411 565
rect 2722 313 2760 409
rect 310 181 382 187
rect 310 97 316 181
rect 376 166 382 181
rect 2340 177 2412 183
rect 2340 166 2346 177
rect 376 154 1026 166
rect 376 120 978 154
rect 1012 120 1026 154
rect 376 108 1026 120
rect 1076 160 1642 166
rect 1076 154 1578 160
rect 1076 120 1086 154
rect 1120 120 1578 154
rect 1076 108 1578 120
rect 376 97 382 108
rect 310 91 382 97
rect 1572 96 1578 108
rect 1636 96 1642 160
rect 1692 154 2346 166
rect 1692 120 1706 154
rect 1740 120 2346 154
rect 1692 108 2346 120
rect 1572 90 1642 96
rect 2340 93 2346 108
rect 2406 93 2412 177
rect 2340 87 2412 93
rect 514 -122 1254 -26
rect 1559 -122 2304 -26
rect 1930 -210 2026 -204
rect 310 -280 382 -273
rect 310 -334 316 -280
rect 376 -334 382 -280
rect 310 -339 382 -334
rect 1184 -280 1248 -274
rect 1930 -276 1936 -210
rect 2020 -276 2026 -210
rect 1184 -336 1190 -280
rect 1242 -336 1248 -280
rect 1184 -342 1248 -336
rect 1328 -282 1394 -276
rect 1328 -342 1334 -282
rect 1388 -342 1394 -282
rect 1328 -348 1394 -342
rect 406 -380 482 -374
rect 406 -434 412 -380
rect 476 -434 482 -380
rect 406 -440 482 -434
rect 1482 -450 1556 -442
rect 1482 -502 1492 -450
rect 1550 -502 1556 -450
rect 1482 -508 1556 -502
rect 1930 -570 2026 -276
rect 2340 -284 2412 -278
rect 2340 -338 2346 -284
rect 2406 -338 2412 -284
rect 2340 -344 2412 -338
rect 2244 -382 2314 -376
rect 2244 -434 2250 -382
rect 2308 -434 2314 -382
rect 2244 -440 2314 -434
rect 102 -666 2452 -570
<< via1 >>
rect 316 1506 376 1590
rect 692 1650 752 1734
rect 319 1025 371 1077
rect 570 1078 632 1134
rect 1020 1078 1076 1134
rect 696 974 748 1026
rect 924 970 976 1030
rect 1120 970 1172 1030
rect 1032 852 1084 912
rect 1966 1218 2026 1302
rect 1642 1078 1698 1134
rect 1546 970 1598 1030
rect 1742 970 1794 1030
rect 2346 1362 2406 1446
rect 1970 974 2022 1026
rect 2086 1078 2148 1134
rect 1333 856 1385 908
rect 1634 852 1686 912
rect 1938 908 2018 914
rect 1938 866 1944 908
rect 1944 866 2012 908
rect 2012 866 2018 908
rect 1938 860 2018 866
rect 321 612 373 621
rect 321 578 330 612
rect 330 578 364 612
rect 364 578 373 612
rect 321 569 373 578
rect 2349 1021 2401 1073
rect 2351 610 2403 617
rect 2351 576 2356 610
rect 2356 576 2390 610
rect 2390 576 2403 610
rect 2351 565 2403 576
rect 316 97 376 181
rect 1578 154 1636 160
rect 1578 120 1598 154
rect 1598 120 1632 154
rect 1632 120 1636 154
rect 1578 96 1636 120
rect 2346 93 2406 177
rect 316 -290 376 -280
rect 316 -324 332 -290
rect 332 -324 366 -290
rect 366 -324 376 -290
rect 316 -334 376 -324
rect 1936 -276 2020 -210
rect 1190 -290 1242 -280
rect 1190 -324 1202 -290
rect 1202 -324 1236 -290
rect 1236 -324 1242 -290
rect 1190 -336 1242 -324
rect 1334 -292 1388 -282
rect 1334 -328 1342 -292
rect 1342 -328 1378 -292
rect 1378 -328 1388 -292
rect 1334 -342 1388 -328
rect 412 -388 476 -380
rect 412 -424 446 -388
rect 446 -424 476 -388
rect 412 -434 476 -424
rect 1492 -456 1550 -450
rect 1492 -492 1494 -456
rect 1494 -492 1530 -456
rect 1530 -492 1550 -456
rect 1492 -502 1550 -492
rect 2346 -290 2406 -284
rect 2346 -324 2352 -290
rect 2352 -324 2386 -290
rect 2386 -324 2406 -290
rect 2346 -338 2406 -324
rect 2250 -388 2308 -382
rect 2250 -424 2272 -388
rect 2272 -424 2306 -388
rect 2306 -424 2308 -388
rect 2250 -434 2308 -424
<< metal2 >>
rect -42 1734 2760 1740
rect -42 1650 692 1734
rect 752 1650 2760 1734
rect -42 1644 2760 1650
rect -42 1590 2760 1596
rect -42 1506 316 1590
rect 376 1506 2760 1590
rect -42 1500 2760 1506
rect -42 1446 2760 1452
rect -42 1362 2346 1446
rect 2406 1362 2760 1446
rect -42 1356 2760 1362
rect -42 1302 2760 1308
rect -42 1218 1966 1302
rect 2026 1218 2760 1302
rect -42 1212 2760 1218
rect 562 1134 1082 1140
rect 310 1077 382 1083
rect 310 1025 319 1077
rect 371 1025 382 1077
rect 562 1078 570 1134
rect 632 1078 1020 1134
rect 1076 1078 1082 1134
rect 562 1072 1082 1078
rect 1636 1134 2156 1140
rect 1636 1078 1642 1134
rect 1698 1078 2086 1134
rect 2148 1078 2156 1134
rect 1636 1072 2156 1078
rect 2340 1073 2412 1079
rect 310 621 382 1025
rect 686 1030 1178 1036
rect 686 1026 924 1030
rect 686 974 696 1026
rect 748 974 924 1026
rect 686 970 924 974
rect 976 970 1120 1030
rect 1172 970 1178 1030
rect 686 964 1178 970
rect 1540 1030 2032 1036
rect 1540 970 1546 1030
rect 1598 970 1742 1030
rect 1794 1026 2032 1030
rect 1794 974 1970 1026
rect 2022 974 2032 1026
rect 1794 970 2032 974
rect 1540 964 2032 970
rect 2340 1021 2349 1073
rect 2401 1021 2412 1073
rect 1026 912 1692 918
rect 1026 852 1032 912
rect 1084 908 1634 912
rect 1084 856 1333 908
rect 1385 856 1634 908
rect 1084 852 1634 856
rect 1686 852 1692 912
rect 1026 846 1692 852
rect 1930 914 2026 922
rect 1930 860 1938 914
rect 2018 860 2026 914
rect 310 569 321 621
rect 373 569 382 621
rect 310 181 382 569
rect 310 97 316 181
rect 376 97 382 181
rect 310 -280 382 97
rect 1572 160 1642 166
rect 1572 96 1578 160
rect 1636 96 1642 160
rect 310 -334 316 -280
rect 376 -334 382 -280
rect 310 -339 382 -334
rect 1184 -280 1248 -274
rect 1184 -336 1190 -280
rect 1242 -336 1248 -280
rect 1184 -374 1248 -336
rect 406 -380 1248 -374
rect 406 -434 412 -380
rect 476 -434 1248 -380
rect 406 -440 1248 -434
rect 1328 -282 1394 -276
rect 1328 -342 1334 -282
rect 1388 -342 1394 -282
rect 1328 -574 1394 -342
rect 1572 -442 1642 96
rect 1930 -210 2026 860
rect 1930 -276 1936 -210
rect 2020 -276 2026 -210
rect 1930 -282 2026 -276
rect 2340 617 2412 1021
rect 2340 565 2351 617
rect 2403 565 2412 617
rect 2340 177 2412 565
rect 2340 93 2346 177
rect 2406 93 2412 177
rect 2340 -284 2412 93
rect 2340 -338 2346 -284
rect 2406 -338 2412 -284
rect 2340 -344 2412 -338
rect 1482 -450 1642 -442
rect 1482 -502 1492 -450
rect 1550 -502 1642 -450
rect 1482 -508 1642 -502
rect 2244 -382 2314 -376
rect 2244 -434 2250 -382
rect 2308 -434 2314 -382
rect 2244 -574 2314 -434
rect 1328 -644 2314 -574
use sky130_fd_pr__nfet_01v8_ZRZL87  sky130_fd_pr__nfet_01v8_ZRZL87_0
timestamp 1695375165
transform -1 0 1669 0 -1 312
box -363 -310 363 310
use sky130_fd_pr__nfet_01v8_ZRZL87  sky130_fd_pr__nfet_01v8_ZRZL87_1
timestamp 1695375165
transform 1 0 1049 0 -1 312
box -363 -310 363 310
use sky130_fd_pr__pfet_01v8_3HMKL2  sky130_fd_pr__pfet_01v8_3HMKL2_0
timestamp 1695375165
transform -1 0 1669 0 1 941
box -363 -319 363 319
use sky130_fd_pr__pfet_01v8_3HMKL2  sky130_fd_pr__pfet_01v8_3HMKL2_1
timestamp 1695375165
transform 1 0 1049 0 1 941
box -363 -319 363 319
use sky130_fd_sc_hd__and2_1  sky130_fd_sc_hd__and2_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 1128 0 -1 -74
box -38 -48 498 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 -4 0 1 361
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_1
timestamp 1694700623
transform 1 0 252 0 1 361
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_2
timestamp 1694700623
transform -1 0 2722 0 -1 -74
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_3
timestamp 1694700623
transform -1 0 2466 0 -1 -74
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_4
timestamp 1694700623
transform 1 0 252 0 -1 -74
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_5
timestamp 1694700623
transform 1 0 -4 0 -1 -74
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_6
timestamp 1694700623
transform -1 0 2722 0 1 361
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_7
timestamp 1694700623
transform -1 0 2466 0 1 361
box -38 -48 314 592
<< labels >>
flabel metal1 2722 857 2760 953 0 FreeSans 160 0 0 0 vdd_mux21
port 11 nsew
flabel metal1 2722 313 2760 409 0 FreeSans 160 0 0 0 vss_mux21
port 0 nsew
flabel metal1 686 1026 758 1668 0 FreeSans 320 90 0 0 in1_mux21
port 8 nsew
flabel metal1 1323 908 1395 1668 0 FreeSans 320 90 0 0 out_mux21
port 7 nsew
flabel metal1 2340 1073 2412 1668 0 FreeSans 320 90 0 0 s0_mux21
port 10 nsew
flabel metal1 1960 1026 2032 1668 0 FreeSans 320 90 0 0 in0_mux21
port 9 nsew
flabel metal1 310 1077 382 1661 0 FreeSans 320 90 0 0 s1_mux21
port 2 nsew
<< end >>
