magic
tech sky130A
magscale 1 2
timestamp 1698999411
<< pwell >>
rect -213 -76 213 76
<< nmos >>
rect -129 -50 -29 50
rect 29 -50 129 50
<< ndiff >>
rect -187 17 -129 50
rect -187 -17 -175 17
rect -141 -17 -129 17
rect -187 -50 -129 -17
rect -29 17 29 50
rect -29 -17 -17 17
rect 17 -17 29 17
rect -29 -50 29 -17
rect 129 17 187 50
rect 129 -17 141 17
rect 175 -17 187 17
rect 129 -50 187 -17
<< ndiffc >>
rect -175 -17 -141 17
rect -17 -17 17 17
rect 141 -17 175 17
<< poly >>
rect -129 50 -29 76
rect 29 50 129 76
rect -129 -76 -29 -50
rect 29 -76 129 -50
<< locali >>
rect -175 17 -141 54
rect -175 -54 -141 -17
rect -17 17 17 54
rect -17 -54 17 -17
rect 141 17 175 54
rect 141 -54 175 -17
<< end >>
