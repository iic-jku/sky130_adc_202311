magic
tech sky130A
magscale 1 2
timestamp 1699000694
<< metal3 >>
rect 93510 59508 99838 59620
rect 93510 44417 93622 59508
rect 84476 44297 93622 44417
rect 93510 44296 93622 44297
rect 93512 43296 93624 43298
rect 84414 43176 93624 43296
rect 93512 13198 93624 43176
rect 93512 13086 100078 13198
use adc_top  adc_top_0
timestamp 1698999411
transform 1 0 0 0 1 0
box -1076 -4 85624 80516
<< end >>
