magic
tech sky130A
magscale 1 2
timestamp 1697443107
<< locali >>
rect -3890 1913 -3644 2113
rect -3130 1913 -2980 2113
rect -3717 1764 -3669 1866
rect -3201 1764 -3153 1866
rect -3890 504 -3644 604
rect -3130 590 -2980 604
rect -3130 514 -3055 590
rect -2995 514 -2980 590
rect -3130 504 -2980 514
rect -3717 364 -3669 466
rect -3201 364 -3153 466
<< viali >>
rect -3055 514 -2995 590
<< metal1 >>
rect -3843 2113 -3795 2770
rect -3747 2113 -3699 2770
rect -3890 2104 -3699 2113
rect -3651 2104 -3603 2770
rect -3557 2764 -3505 2770
rect -3557 2662 -3505 2668
rect -3555 2104 -3507 2662
rect -3459 2482 -3411 2770
rect -3365 2764 -3313 2770
rect -3365 2662 -3313 2668
rect -3461 2476 -3409 2482
rect -3461 2374 -3409 2380
rect -3459 2104 -3411 2374
rect -3363 2104 -3315 2662
rect -3267 2626 -3219 2770
rect -3269 2620 -3217 2626
rect -3269 2518 -3217 2524
rect -3267 2104 -3219 2518
rect -3171 2104 -3123 2770
rect -3075 2626 -3027 2770
rect -3077 2620 -3025 2626
rect -3077 2518 -3025 2524
rect -3890 2060 -3714 2104
rect -3891 2051 -3714 2060
rect -3891 1975 -3881 2051
rect -3757 1975 -3714 2051
rect -3891 1966 -3714 1975
rect -3890 1913 -3714 1966
rect -3843 1400 -3795 1913
rect -3651 1652 -3603 1872
rect -3653 1646 -3601 1652
rect -3653 1544 -3601 1550
rect -3651 1400 -3603 1544
rect -3459 1508 -3411 1872
rect -3267 1652 -3219 1872
rect -3269 1646 -3217 1652
rect -3269 1544 -3217 1550
rect -3461 1502 -3409 1508
rect -3461 1400 -3409 1406
rect -3267 1400 -3219 1544
rect -3075 1508 -3027 2518
rect -3077 1502 -3025 1508
rect -3077 1400 -3025 1406
rect -3843 1108 -3795 1252
rect -3845 1102 -3793 1108
rect -3845 1000 -3793 1006
rect -3843 108 -3795 1000
rect -3747 604 -3699 1252
rect -3651 604 -3603 1252
rect -3557 1246 -3505 1252
rect -3557 1144 -3505 1150
rect -3555 604 -3507 1144
rect -3459 964 -3411 1252
rect -3365 1246 -3313 1252
rect -3365 1144 -3313 1150
rect -3461 958 -3409 964
rect -3461 856 -3409 862
rect -3459 604 -3411 856
rect -3363 604 -3315 1144
rect -3267 1108 -3219 1252
rect -3269 1102 -3217 1108
rect -3269 1000 -3217 1006
rect -3267 604 -3219 1000
rect -3171 604 -3123 1252
rect -3075 604 -3027 1252
rect -3125 590 -2980 604
rect -3125 514 -3113 590
rect -2990 514 -2980 590
rect -3125 504 -2980 514
rect -3651 252 -3603 472
rect -3653 246 -3601 252
rect -3653 144 -3601 150
rect -3845 102 -3793 108
rect -3845 0 -3793 6
rect -3651 0 -3603 144
rect -3459 108 -3411 472
rect -3267 252 -3219 472
rect -3269 246 -3217 252
rect -3269 144 -3217 150
rect -3461 102 -3409 108
rect -3461 0 -3409 6
rect -3267 0 -3219 144
rect -3075 0 -3027 504
<< via1 >>
rect -3557 2668 -3505 2764
rect -3365 2668 -3313 2764
rect -3461 2380 -3409 2476
rect -3269 2524 -3217 2620
rect -3077 2524 -3025 2620
rect -3881 1975 -3757 2051
rect -3653 1550 -3601 1646
rect -3269 1550 -3217 1646
rect -3461 1406 -3409 1502
rect -3077 1406 -3025 1502
rect -3845 1006 -3793 1102
rect -3557 1150 -3505 1246
rect -3365 1150 -3313 1246
rect -3461 862 -3409 958
rect -3269 1006 -3217 1102
rect -3113 514 -3055 590
rect -3055 514 -2995 590
rect -2995 514 -2990 590
rect -3653 150 -3601 246
rect -3845 6 -3793 102
rect -3269 150 -3217 246
rect -3461 6 -3409 102
<< metal2 >>
rect -3557 2764 -3505 2770
rect -3365 2764 -3313 2770
rect -3890 2668 -3557 2764
rect -3505 2668 -3365 2764
rect -3313 2668 -2980 2764
rect -3557 2662 -3505 2668
rect -3365 2662 -3313 2668
rect -3269 2620 -3217 2626
rect -3077 2620 -3025 2626
rect -3890 2524 -3269 2620
rect -3217 2524 -3077 2620
rect -3025 2524 -2980 2620
rect -3269 2518 -3217 2524
rect -3461 2476 -3409 2482
rect -3890 2380 -3461 2476
rect -3409 2466 -2981 2476
rect -3409 2390 -3113 2466
rect -2989 2452 -2981 2466
rect -2989 2390 -2980 2452
rect -3409 2380 -2980 2390
rect -3461 2374 -3409 2380
rect -3891 2051 -3747 2060
rect -3891 1975 -3881 2051
rect -3757 1975 -3747 2051
rect -3891 1966 -3747 1975
rect -3653 1646 -3601 1652
rect -3269 1646 -3217 1652
rect -3890 1550 -3653 1646
rect -3601 1636 -3269 1646
rect -3601 1560 -3369 1636
rect -3601 1550 -3269 1560
rect -3217 1550 -2980 1646
rect -3653 1544 -3601 1550
rect -3269 1544 -3217 1550
rect -3461 1502 -3409 1508
rect -3077 1502 -3025 1508
rect -3890 1492 -3461 1502
rect -3890 1416 -3625 1492
rect -3501 1416 -3461 1492
rect -3890 1406 -3461 1416
rect -3409 1406 -3077 1502
rect -3025 1406 -2980 1502
rect -3461 1400 -3409 1406
rect -3077 1400 -3025 1406
rect -3557 1246 -3505 1252
rect -3365 1246 -3313 1252
rect -3890 1150 -3557 1246
rect -3505 1150 -3365 1246
rect -3313 1150 -2980 1246
rect -3557 1144 -3505 1150
rect -3365 1144 -3313 1150
rect -3845 1102 -3793 1108
rect -3269 1102 -3217 1108
rect -3890 1006 -3845 1102
rect -3793 1006 -3269 1102
rect -3217 1006 -2980 1102
rect -3845 1000 -3793 1006
rect -3269 1000 -3217 1006
rect -3461 958 -3409 964
rect -3890 948 -3461 958
rect -3890 872 -3881 948
rect -3757 872 -3461 948
rect -3890 862 -3461 872
rect -3409 862 -2980 958
rect -3461 856 -3409 862
rect -3123 590 -2980 604
rect -3123 514 -3113 590
rect -2989 514 -2980 590
rect -3123 504 -2980 514
rect -3653 246 -3601 252
rect -3269 246 -3217 252
rect -3890 150 -3653 246
rect -3601 236 -3269 246
rect -3601 160 -3369 236
rect -3601 150 -3269 160
rect -3217 150 -2980 246
rect -3653 144 -3601 150
rect -3269 144 -3217 150
rect -3845 102 -3793 108
rect -3461 102 -3409 108
rect -3890 6 -3845 102
rect -3793 92 -3461 102
rect -3793 16 -3625 92
rect -3501 16 -3461 92
rect -3793 6 -3461 16
rect -3409 6 -2980 102
rect -3845 0 -3793 6
rect -3461 0 -3409 6
<< via2 >>
rect -3113 2390 -2989 2466
rect -3881 1975 -3757 2051
rect -3369 1560 -3269 1636
rect -3269 1560 -3245 1636
rect -3625 1416 -3501 1492
rect -3881 872 -3757 948
rect -3113 514 -2990 590
rect -2990 514 -2989 590
rect -3369 160 -3269 236
rect -3269 160 -3245 236
rect -3625 16 -3501 92
<< metal3 >>
rect -3891 2051 -3747 2764
rect -3891 1975 -3881 2051
rect -3757 1975 -3747 2051
rect -3891 948 -3747 1975
rect -3891 872 -3881 948
rect -3757 872 -3747 948
rect -3891 6 -3747 872
rect -3635 1492 -3491 2764
rect -3635 1416 -3625 1492
rect -3501 1416 -3491 1492
rect -3635 92 -3491 1416
rect -3635 16 -3625 92
rect -3501 16 -3491 92
rect -3635 6 -3491 16
rect -3379 1636 -3235 2764
rect -3379 1560 -3369 1636
rect -3245 1560 -3235 1636
rect -3379 236 -3235 1560
rect -3379 160 -3369 236
rect -3245 160 -3235 236
rect -3379 6 -3235 160
rect -3123 2466 -2979 2764
rect -3123 2390 -3113 2466
rect -2989 2390 -2979 2466
rect -3123 590 -2979 2390
rect -3123 514 -3113 590
rect -2989 514 -2979 590
rect -3123 6 -2979 514
use sky130_fd_pr__nfet_01v8_QWA63T  sky130_fd_pr__nfet_01v8_QWA63T_1
timestamp 1696930192
transform 1 0 -3435 0 1 554
box -455 -260 455 260
use sky130_fd_pr__pfet_01v8_UAU7GH  sky130_fd_pr__pfet_01v8_UAU7GH_1
timestamp 1696931086
transform 1 0 -3435 0 1 2013
box -455 -319 455 319
<< end >>
