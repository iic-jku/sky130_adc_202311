magic
tech sky130A
magscale 1 2
timestamp 1699263546
<< locali >>
rect -293 6162 -2 6394
rect -293 5822 -272 6162
rect -32 5822 -2 6162
rect -293 5644 -2 5822
rect 89 5644 98 6394
rect 20702 6162 21002 6394
rect 20702 5822 20732 6162
rect 20972 5822 21002 6162
rect 7462 -1126 7762 -894
rect 7462 -1466 7492 -1126
rect 7732 -1466 7762 -1126
rect 7462 -1644 7762 -1466
rect 8021 -4558 9206 -4538
rect 8021 -5268 8041 -4558
rect 8529 -4770 9206 -4558
rect 8529 -5110 8786 -4770
rect 9026 -5110 9206 -4770
rect 8529 -5268 9206 -5110
rect 8021 -5288 9206 -5268
rect 10280 -6994 10420 5654
rect 20702 5644 21002 5822
rect 12938 -1126 13238 -894
rect 12938 -1466 12968 -1126
rect 13208 -1466 13238 -1126
rect 12938 -1644 13238 -1466
rect 11644 -4770 11944 -4538
rect 11644 -5110 11674 -4770
rect 11914 -5110 11944 -4770
rect 11644 -5288 11944 -5110
<< viali >>
rect -272 5822 -32 6162
rect 20732 5822 20972 6162
rect 7492 -1466 7732 -1126
rect 8041 -5268 8529 -4558
rect 8786 -5110 9026 -4770
rect 12968 -1466 13208 -1126
rect 11674 -5110 11914 -4770
<< metal1 >>
rect 10100 39020 10600 39050
rect 10100 38780 10130 39020
rect 10570 38780 10600 39020
rect 10100 38750 10600 38780
rect -293 6162 -2 6192
rect -293 5822 -272 6162
rect -32 5822 -2 6162
rect -293 5792 -2 5822
rect 89 5792 98 6192
rect 20702 6162 21002 6192
rect 20702 5822 20732 6162
rect 20972 5822 21002 6162
rect 20702 5792 21002 5822
rect 7462 -1126 7762 -1096
rect 7462 -1466 7492 -1126
rect 7732 -1466 7762 -1126
rect 7462 -1496 7762 -1466
rect 12938 -1126 13238 -1096
rect 12938 -1466 12968 -1126
rect 13208 -1466 13238 -1126
rect 12938 -1496 13238 -1466
rect 8021 -4558 8549 -4538
rect 8021 -5268 8041 -4558
rect 8529 -5268 8549 -4558
rect 8756 -4770 9056 -4740
rect 8756 -5110 8786 -4770
rect 9026 -5110 9056 -4770
rect 8756 -5140 9056 -5110
rect 11644 -4770 11944 -4740
rect 11644 -5110 11674 -4770
rect 11914 -5110 11944 -4770
rect 11644 -5140 11944 -5110
rect 8021 -5288 8549 -5268
<< via1 >>
rect 10130 38780 10570 39020
rect -272 5822 -32 6162
rect 20732 5822 20972 6162
rect 7492 -1466 7732 -1126
rect 12968 -1466 13208 -1126
rect 8786 -5110 9026 -4770
rect 11674 -5110 11914 -4770
<< metal2 >>
rect 8021 37768 8549 39050
rect 10100 39020 10600 39050
rect 10100 38780 10130 39020
rect 10570 38780 10600 39020
rect 10100 38750 10600 38780
rect 8021 37428 8051 37768
rect 8519 37428 8549 37768
rect 8021 37310 8549 37428
rect 6624 7858 7058 7878
rect 6624 7698 6644 7858
rect 7038 7698 7058 7858
rect 6624 7180 7058 7698
rect 13080 7858 13514 7878
rect 13080 7698 13100 7858
rect 13494 7698 13514 7858
rect 13080 7180 13514 7698
rect 140 7016 574 7036
rect 140 6816 160 7016
rect 554 6816 574 7016
rect 140 6796 574 6816
rect 1434 7016 1868 7036
rect 1434 6816 1454 7016
rect 1848 6816 1868 7016
rect 1434 6796 1868 6816
rect 2728 7016 3162 7036
rect 2728 6816 2748 7016
rect 3142 6816 3162 7016
rect 2728 6796 3162 6816
rect 4022 7016 4456 7036
rect 4022 6816 4042 7016
rect 4436 6816 4456 7016
rect 4022 6796 4456 6816
rect 5316 7016 5750 7036
rect 5316 6816 5336 7016
rect 5730 6816 5750 7016
rect 5316 6796 5750 6816
rect 6610 7016 7044 7036
rect 6610 6816 6630 7016
rect 7024 6816 7044 7016
rect 6610 6796 7044 6816
rect 7904 7016 8338 7036
rect 7904 6816 7924 7016
rect 8318 6816 8338 7016
rect 7904 6796 8338 6816
rect 9198 7016 9632 7036
rect 9198 6816 9218 7016
rect 9612 6816 9632 7016
rect 9198 6796 9632 6816
rect 10492 7016 10926 7036
rect 10492 6816 10512 7016
rect 10906 6816 10926 7016
rect 10492 6796 10926 6816
rect 11786 7016 12220 7036
rect 11786 6816 11806 7016
rect 12200 6816 12220 7016
rect 11786 6796 12220 6816
rect 13080 7016 13514 7036
rect 13080 6816 13100 7016
rect 13494 6816 13514 7016
rect 13080 6796 13514 6816
rect 14374 7016 14808 7036
rect 14374 6816 14394 7016
rect 14788 6816 14808 7016
rect 14374 6796 14808 6816
rect 15668 7016 16102 7036
rect 15668 6816 15688 7016
rect 16082 6816 16102 7016
rect 15668 6796 16102 6816
rect 16962 7016 17396 7036
rect 16962 6816 16982 7016
rect 17376 6816 17396 7016
rect 16962 6796 17396 6816
rect 18256 7016 18690 7036
rect 18256 6816 18276 7016
rect 18670 6816 18690 7016
rect 18256 6796 18690 6816
rect 19550 7016 19984 7036
rect 19550 6816 19570 7016
rect 19964 6816 19984 7016
rect 19550 6796 19984 6816
rect -293 6162 21002 6192
rect -293 5822 -272 6162
rect -32 5822 8051 6162
rect 8519 5822 20732 6162
rect 20972 5822 21002 6162
rect -293 5792 21002 5822
rect 20655 5146 20702 5242
rect 20655 5002 20702 5098
rect 6624 4214 7058 4234
rect 6624 4054 6644 4214
rect 7038 4054 7058 4214
rect 6624 3486 7058 4054
rect 13080 4214 13514 4234
rect 13080 4054 13100 4214
rect 13494 4054 13514 4214
rect 13080 3486 13514 4054
rect 5316 3372 5750 3392
rect 5316 3172 5336 3372
rect 5730 3172 5750 3372
rect 5316 3152 5750 3172
rect 6610 3372 7044 3392
rect 6610 3172 6630 3372
rect 7024 3172 7044 3372
rect 6610 3152 7044 3172
rect 7904 3372 8338 3392
rect 7904 3172 7924 3372
rect 8318 3172 8338 3372
rect 7904 3152 8338 3172
rect 9198 3372 9632 3392
rect 9198 3172 9218 3372
rect 9612 3172 9632 3372
rect 9198 3152 9632 3172
rect 10492 3372 10926 3392
rect 10492 3172 10512 3372
rect 10906 3172 10926 3372
rect 10492 3152 10926 3172
rect 11786 3372 12220 3392
rect 11786 3172 11806 3372
rect 12200 3172 12220 3372
rect 11786 3152 12220 3172
rect 13080 3372 13514 3392
rect 13080 3172 13100 3372
rect 13494 3172 13514 3372
rect 13080 3152 13514 3172
rect 14374 3372 14808 3392
rect 14374 3172 14394 3372
rect 14788 3172 14808 3372
rect 14374 3152 14808 3172
rect 8021 2518 8549 2548
rect 8021 2178 8051 2518
rect 8519 2178 8549 2518
rect 8021 2148 8549 2178
rect 15481 1502 15528 1598
rect 15481 1358 15528 1454
rect 6624 570 7058 590
rect 6624 410 6644 570
rect 7038 410 7058 570
rect 6624 -252 7058 410
rect 13080 570 13514 590
rect 13080 410 13100 570
rect 13494 410 13514 570
rect 13080 -108 13514 410
rect 12937 -204 13514 -108
rect 6624 -348 7762 -252
rect 7904 -272 8338 -252
rect 7904 -472 7924 -272
rect 8318 -472 8338 -272
rect 7904 -492 8338 -472
rect 9198 -272 9632 -252
rect 9198 -472 9218 -272
rect 9612 -472 9632 -272
rect 9198 -492 9632 -472
rect 10492 -272 10926 -252
rect 10492 -472 10512 -272
rect 10906 -472 10926 -272
rect 10492 -492 10926 -472
rect 11786 -272 12220 -252
rect 11786 -472 11806 -272
rect 12200 -472 12220 -272
rect 11786 -492 12220 -472
rect 7462 -1126 13238 -1096
rect 7462 -1466 7492 -1126
rect 7732 -1466 8051 -1126
rect 8519 -1466 12968 -1126
rect 13208 -1466 13238 -1126
rect 7462 -1496 13238 -1466
rect 12891 -2142 12938 -2046
rect 12891 -2286 12938 -2190
rect 6624 -3074 7058 -3054
rect 6624 -3234 6644 -3074
rect 7038 -3234 7058 -3074
rect 6624 -3896 7058 -3234
rect 13080 -3074 13514 -3054
rect 13080 -3234 13100 -3074
rect 13494 -3234 13514 -3074
rect 13080 -3348 13514 -3234
rect 13078 -3752 13514 -3348
rect 11621 -3848 13514 -3752
rect 13078 -3896 13514 -3848
rect 6622 -3992 9065 -3896
rect 9197 -3916 9631 -3896
rect 9197 -4116 9217 -3916
rect 9611 -4116 9631 -3916
rect 9197 -4136 9631 -4116
rect 10492 -3916 10926 -3896
rect 10492 -4116 10512 -3916
rect 10906 -4116 10926 -3916
rect 10492 -4136 10926 -4116
rect 8021 -4770 11944 -4740
rect 8021 -5110 8051 -4770
rect 8519 -5110 8786 -4770
rect 9026 -5110 11674 -4770
rect 11914 -5110 11944 -4770
rect 8021 -5140 11944 -5110
rect 11597 -5786 11644 -5690
rect 11597 -5930 11644 -5834
<< via2 >>
rect 10130 38780 10570 39020
rect 8051 37428 8519 37768
rect 6644 7698 7038 7858
rect 13100 7698 13494 7858
rect 160 6816 554 7016
rect 1454 6816 1848 7016
rect 2748 6816 3142 7016
rect 4042 6816 4436 7016
rect 5336 6816 5730 7016
rect 6630 6816 7024 7016
rect 7924 6816 8318 7016
rect 9218 6816 9612 7016
rect 10512 6816 10906 7016
rect 11806 6816 12200 7016
rect 13100 6816 13494 7016
rect 14394 6816 14788 7016
rect 15688 6816 16082 7016
rect 16982 6816 17376 7016
rect 18276 6816 18670 7016
rect 19570 6816 19964 7016
rect 8051 5822 8519 6162
rect 6644 4054 7038 4214
rect 13100 4054 13494 4214
rect 5336 3172 5730 3372
rect 6630 3172 7024 3372
rect 7924 3172 8318 3372
rect 9218 3172 9612 3372
rect 10512 3172 10906 3372
rect 11806 3172 12200 3372
rect 13100 3172 13494 3372
rect 14394 3172 14788 3372
rect 8051 2178 8519 2518
rect 6644 410 7038 570
rect 13100 410 13494 570
rect 7924 -472 8318 -272
rect 9218 -472 9612 -272
rect 10512 -472 10906 -272
rect 11806 -472 12200 -272
rect 8051 -1466 8519 -1126
rect 6644 -3234 7038 -3074
rect 13100 -3234 13494 -3074
rect 9217 -4116 9611 -3916
rect 10512 -4116 10906 -3916
rect 8051 -5110 8519 -4770
<< metal3 >>
rect 10100 39020 10600 39050
rect 10100 38780 10130 39020
rect 10570 38780 10600 39020
rect 10100 38750 10600 38780
rect 8021 37768 8549 37798
rect 8021 37428 8051 37768
rect 8519 37428 8549 37768
rect 8021 37398 8549 37428
rect 6624 8228 7058 8248
rect 6624 7698 6644 8228
rect 7038 7698 7058 8228
rect 6624 7678 7058 7698
rect 13080 8228 13514 8248
rect 13080 7698 13100 8228
rect 13494 7698 13514 8228
rect 13080 7678 13514 7698
rect 140 7160 574 7180
rect 140 6816 160 7160
rect 554 6816 574 7160
rect 140 6652 574 6816
rect 1434 7016 1868 7180
rect 1434 6672 1454 7016
rect 1848 6672 1868 7016
rect 1434 6652 1868 6672
rect 2728 7160 3162 7180
rect 2728 6816 2748 7160
rect 3142 6816 3162 7160
rect 2728 6652 3162 6816
rect 4022 7016 4456 7180
rect 4022 6672 4042 7016
rect 4436 6672 4456 7016
rect 4022 6652 4456 6672
rect 5316 7160 5750 7180
rect 5316 6816 5336 7160
rect 5730 6816 5750 7160
rect 5316 6652 5750 6816
rect 6610 7016 7044 7180
rect 6610 6672 6630 7016
rect 7024 6672 7044 7016
rect 6610 6652 7044 6672
rect 7904 7160 8338 7180
rect 7904 6816 7924 7160
rect 8318 6816 8338 7160
rect 7904 6652 8338 6816
rect 9198 7016 9632 7180
rect 9198 6672 9218 7016
rect 9612 6672 9632 7016
rect 9198 6652 9632 6672
rect 10492 7160 10926 7180
rect 10492 6816 10512 7160
rect 10906 6816 10926 7160
rect 10492 6652 10926 6816
rect 11786 7016 12220 7180
rect 11786 6672 11806 7016
rect 12200 6672 12220 7016
rect 11786 6652 12220 6672
rect 13080 7160 13514 7180
rect 13080 6816 13100 7160
rect 13494 6816 13514 7160
rect 13080 6652 13514 6816
rect 14374 7016 14808 7180
rect 14374 6672 14394 7016
rect 14788 6672 14808 7016
rect 14374 6652 14808 6672
rect 15668 7160 16102 7180
rect 15668 6816 15688 7160
rect 16082 6816 16102 7160
rect 15668 6652 16102 6816
rect 16962 7016 17396 7180
rect 16962 6672 16982 7016
rect 17376 6672 17396 7016
rect 16962 6652 17396 6672
rect 18256 7160 18690 7180
rect 18256 6816 18276 7160
rect 18670 6816 18690 7160
rect 18256 6652 18690 6816
rect 19550 7016 19984 7180
rect 19550 6672 19570 7016
rect 19964 6672 19984 7016
rect 19550 6652 19984 6672
rect 8021 6162 8549 6192
rect 8021 5822 8051 6162
rect 8519 5822 8549 6162
rect 8021 5792 8549 5822
rect 6624 4584 7058 4604
rect 6624 4054 6644 4584
rect 7038 4054 7058 4584
rect 6624 4034 7058 4054
rect 13080 4584 13514 4604
rect 13080 4054 13100 4584
rect 13494 4054 13514 4584
rect 13080 4034 13514 4054
rect 5316 3516 5750 3536
rect 5316 3172 5336 3516
rect 5730 3172 5750 3516
rect 5316 3008 5750 3172
rect 6610 3372 7044 3536
rect 6610 3028 6630 3372
rect 7024 3028 7044 3372
rect 6610 3008 7044 3028
rect 7904 3516 8338 3536
rect 7904 3172 7924 3516
rect 8318 3172 8338 3516
rect 7904 3008 8338 3172
rect 9198 3372 9632 3536
rect 9198 3028 9218 3372
rect 9612 3028 9632 3372
rect 9198 3008 9632 3028
rect 10492 3516 10926 3536
rect 10492 3172 10512 3516
rect 10906 3172 10926 3516
rect 10492 3008 10926 3172
rect 11786 3372 12220 3536
rect 11786 3028 11806 3372
rect 12200 3028 12220 3372
rect 11786 3008 12220 3028
rect 13080 3516 13514 3536
rect 13080 3172 13100 3516
rect 13494 3172 13514 3516
rect 13080 3008 13514 3172
rect 14374 3372 14808 3536
rect 14374 3028 14394 3372
rect 14788 3028 14808 3372
rect 14374 3008 14808 3028
rect 8021 2518 8549 2548
rect 8021 2178 8051 2518
rect 8519 2178 8549 2518
rect 8021 2148 8549 2178
rect 6624 940 7058 960
rect 6624 410 6644 940
rect 7038 410 7058 940
rect 6624 390 7058 410
rect 13080 940 13514 960
rect 13080 410 13100 940
rect 13494 410 13514 940
rect 13080 390 13514 410
rect 7904 -128 8338 -108
rect 7904 -472 7924 -128
rect 8318 -472 8338 -128
rect 7904 -636 8338 -472
rect 9198 -272 9632 -108
rect 9198 -616 9218 -272
rect 9612 -616 9632 -272
rect 9198 -636 9632 -616
rect 10492 -128 10926 -108
rect 10492 -472 10512 -128
rect 10906 -472 10926 -128
rect 10492 -636 10926 -472
rect 11786 -272 12220 -108
rect 11786 -616 11806 -272
rect 12200 -616 12220 -272
rect 11786 -636 12220 -616
rect 8021 -1126 8549 -1096
rect 8021 -1466 8051 -1126
rect 8519 -1466 8549 -1126
rect 8021 -1496 8549 -1466
rect 6624 -2704 7058 -2684
rect 6624 -3234 6644 -2704
rect 7038 -3234 7058 -2704
rect 6624 -3254 7058 -3234
rect 13080 -2704 13514 -2684
rect 13080 -3234 13100 -2704
rect 13494 -3234 13514 -2704
rect 13080 -3254 13514 -3234
rect 9197 -3772 9631 -3752
rect 9197 -4116 9217 -3772
rect 9611 -4116 9631 -3772
rect 9197 -4280 9631 -4116
rect 10492 -3916 10926 -3752
rect 10492 -4260 10512 -3916
rect 10906 -4260 10926 -3916
rect 10492 -4280 10926 -4260
rect 8021 -4770 8549 -4740
rect 8021 -5110 8051 -4770
rect 8519 -5110 8549 -4770
rect 8021 -5140 8549 -5110
<< via3 >>
rect 10130 38780 10570 39020
rect 8051 37428 8519 37768
rect 6644 7858 7038 8228
rect 6644 7698 7038 7858
rect 13100 7858 13494 8228
rect 13100 7698 13494 7858
rect 160 7016 554 7160
rect 160 7000 554 7016
rect 1454 6816 1848 6832
rect 1454 6672 1848 6816
rect 2748 7016 3142 7160
rect 2748 7000 3142 7016
rect 4042 6816 4436 6832
rect 4042 6672 4436 6816
rect 5336 7016 5730 7160
rect 5336 7000 5730 7016
rect 6630 6816 7024 6832
rect 6630 6672 7024 6816
rect 7924 7016 8318 7160
rect 7924 7000 8318 7016
rect 9218 6816 9612 6832
rect 9218 6672 9612 6816
rect 10512 7016 10906 7160
rect 10512 7000 10906 7016
rect 11806 6816 12200 6832
rect 11806 6672 12200 6816
rect 13100 7016 13494 7160
rect 13100 7000 13494 7016
rect 14394 6816 14788 6832
rect 14394 6672 14788 6816
rect 15688 7016 16082 7160
rect 15688 7000 16082 7016
rect 16982 6816 17376 6832
rect 16982 6672 17376 6816
rect 18276 7016 18670 7160
rect 18276 7000 18670 7016
rect 19570 6816 19964 6832
rect 19570 6672 19964 6816
rect 8051 5822 8519 6162
rect 6644 4214 7038 4584
rect 6644 4054 7038 4214
rect 13100 4214 13494 4584
rect 13100 4054 13494 4214
rect 5336 3372 5730 3516
rect 5336 3356 5730 3372
rect 6630 3172 7024 3188
rect 6630 3028 7024 3172
rect 7924 3372 8318 3516
rect 7924 3356 8318 3372
rect 9218 3172 9612 3188
rect 9218 3028 9612 3172
rect 10512 3372 10906 3516
rect 10512 3356 10906 3372
rect 11806 3172 12200 3188
rect 11806 3028 12200 3172
rect 13100 3372 13494 3516
rect 13100 3356 13494 3372
rect 14394 3172 14788 3188
rect 14394 3028 14788 3172
rect 8051 2178 8519 2518
rect 6644 570 7038 940
rect 6644 410 7038 570
rect 13100 570 13494 940
rect 13100 410 13494 570
rect 7924 -272 8318 -128
rect 7924 -288 8318 -272
rect 9218 -472 9612 -456
rect 9218 -616 9612 -472
rect 10512 -272 10906 -128
rect 10512 -288 10906 -272
rect 11806 -472 12200 -456
rect 11806 -616 12200 -472
rect 8051 -1466 8519 -1126
rect 6644 -3074 7038 -2704
rect 6644 -3234 7038 -3074
rect 13100 -3074 13494 -2704
rect 13100 -3234 13494 -3074
rect 9217 -3916 9611 -3772
rect 9217 -3932 9611 -3916
rect 10512 -4116 10906 -4100
rect 10512 -4260 10906 -4116
rect 8051 -5110 8519 -4770
<< metal4 >>
rect 8021 39020 12606 39050
rect 8021 38780 8051 39020
rect 8519 38780 10130 39020
rect 10570 38780 12606 39020
rect 8021 38750 12606 38780
rect 8021 38520 12606 38550
rect 8021 38280 9880 38520
rect 10820 38280 12108 38520
rect 12576 38280 12606 38520
rect 8021 38250 12606 38280
rect 8021 37768 8549 37798
rect 8021 37428 8051 37768
rect 8519 37428 8549 37768
rect 8021 37398 8549 37428
rect -2821 22066 -9 22126
rect -2821 21616 -950 22066
rect -69 21616 -9 22066
rect -2821 21556 -9 21616
rect 20113 22066 22925 22126
rect 20113 21616 20173 22066
rect 21054 21616 22925 22066
rect 20113 21556 22925 21616
rect -2821 20244 -9 20304
rect -2821 19794 -2762 20244
rect -1881 19794 -9 20244
rect -2821 19734 -9 19794
rect 20113 20244 22925 20304
rect 20113 19794 21985 20244
rect 22866 19794 22925 20244
rect 20113 19734 22925 19794
rect -2821 18422 -9 18482
rect -2821 17972 -950 18422
rect -69 17972 -9 18422
rect -2821 17912 -9 17972
rect 20113 18422 22925 18482
rect 20113 17972 20173 18422
rect 21054 17972 22925 18422
rect 20113 17912 22925 17972
rect -2821 16600 -9 16660
rect -2821 16150 -2762 16600
rect -1881 16150 -9 16600
rect -2821 16090 -9 16150
rect 20113 16600 22925 16660
rect 20113 16150 21985 16600
rect 22866 16150 22925 16600
rect 20113 16090 22925 16150
rect -2821 14778 -9 14838
rect -2821 14328 -950 14778
rect -69 14328 -9 14778
rect -2821 14268 -9 14328
rect 20113 14778 22925 14838
rect 20113 14328 20173 14778
rect 21054 14328 22925 14778
rect 20113 14268 22925 14328
rect -2821 12956 -9 13016
rect -2821 12506 -2762 12956
rect -1881 12506 -9 12956
rect -2821 12446 -9 12506
rect 20113 12956 22925 13016
rect 20113 12506 21985 12956
rect 22866 12506 22925 12956
rect 20113 12446 22925 12506
rect -2821 11134 -9 11194
rect -2821 10684 -950 11134
rect -69 10684 -9 11134
rect -2821 10624 -9 10684
rect 20113 11134 22925 11194
rect 20113 10684 20173 11134
rect 21054 10684 22925 11134
rect 20113 10624 22925 10684
rect -2821 9312 -9 9372
rect -2821 8862 -2762 9312
rect -1881 8862 -9 9312
rect -2821 8802 -9 8862
rect 20113 9312 22925 9372
rect 20113 8862 21985 9312
rect 22866 8862 22925 9312
rect 20113 8802 22925 8862
rect 6622 8228 7622 8248
rect 6622 7698 6644 8228
rect 7038 8188 7622 8228
rect 7563 7738 7622 8188
rect 7038 7698 7622 7738
rect 6622 7678 7622 7698
rect 13078 8228 14078 8248
rect 13078 7698 13100 8228
rect 13494 8188 14078 8228
rect 14019 7738 14078 8188
rect 13494 7698 14078 7738
rect 13078 7678 14078 7698
rect -2821 7490 22925 7550
rect -2821 7040 -950 7490
rect -69 7160 20173 7490
rect -69 7040 160 7160
rect -2821 7000 160 7040
rect 554 7000 2748 7160
rect 3142 7000 5336 7160
rect 5730 7000 7924 7160
rect 8318 7000 10512 7160
rect 10906 7000 13100 7160
rect 13494 7000 15688 7160
rect 16082 7000 18276 7160
rect 18670 7040 20173 7160
rect 21054 7040 22925 7490
rect 18670 7000 22925 7040
rect -2821 6980 22925 7000
rect -1291 6832 21393 6852
rect -1291 6672 1454 6832
rect 1848 6672 4042 6832
rect 4436 6672 6630 6832
rect 7024 6672 9218 6832
rect 9612 6672 11806 6832
rect 12200 6672 14394 6832
rect 14788 6672 16982 6832
rect 17376 6672 19570 6832
rect 19964 6672 21393 6832
rect -1291 6282 21393 6672
rect 8021 6162 8549 6192
rect 8021 5822 8051 6162
rect 8519 5822 8549 6162
rect 8021 5792 8549 5822
rect -2821 5668 -9 5728
rect -2821 5218 -2762 5668
rect -1881 5218 -9 5668
rect -2821 5158 -9 5218
rect 20113 5668 22925 5728
rect 20113 5218 21985 5668
rect 22866 5218 22925 5668
rect 20113 5158 22925 5218
rect 6622 4584 7622 4604
rect 6622 4054 6644 4584
rect 7038 4544 7622 4584
rect 7563 4094 7622 4544
rect 7038 4054 7622 4094
rect 6622 4034 7622 4054
rect 13078 4584 14078 4604
rect 13078 4054 13100 4584
rect 13494 4544 14078 4584
rect 14019 4094 14078 4544
rect 13494 4054 14078 4094
rect 13078 4034 14078 4054
rect -2821 3846 22925 3906
rect -2821 3396 -950 3846
rect -69 3516 20173 3846
rect -69 3396 5336 3516
rect -2821 3356 5336 3396
rect 5730 3356 7924 3516
rect 8318 3356 10512 3516
rect 10906 3356 13100 3516
rect 13494 3396 20173 3516
rect 21054 3396 22925 3846
rect 13494 3356 22925 3396
rect -2821 3336 22925 3356
rect -1291 3188 21393 3208
rect -1291 3028 6630 3188
rect 7024 3028 9218 3188
rect 9612 3028 11806 3188
rect 12200 3028 14394 3188
rect 14788 3028 21393 3188
rect -1291 2638 21393 3028
rect 8021 2518 8549 2548
rect 8021 2178 8051 2518
rect 8519 2178 8549 2518
rect 8021 2148 8549 2178
rect -2821 2024 -9 2084
rect -2821 1574 -2762 2024
rect -1881 1574 -9 2024
rect -2821 1514 -9 1574
rect 20113 2024 22925 2084
rect 20113 1574 21985 2024
rect 22866 1574 22925 2024
rect 20113 1514 22925 1574
rect 6622 940 7622 960
rect 6622 410 6644 940
rect 7038 900 7622 940
rect 7563 450 7622 900
rect 7038 410 7622 450
rect 6622 390 7622 410
rect 13078 940 14078 960
rect 13078 410 13100 940
rect 13494 900 14078 940
rect 14019 450 14078 900
rect 13494 410 14078 450
rect 13078 390 14078 410
rect -2821 202 22925 262
rect -2821 -248 -950 202
rect -69 -128 20173 202
rect -69 -248 7924 -128
rect -2821 -288 7924 -248
rect 8318 -288 10512 -128
rect 10906 -248 20173 -128
rect 21054 -248 22925 202
rect 10906 -288 22925 -248
rect -2821 -308 22925 -288
rect -1291 -456 21393 -436
rect -1291 -616 9218 -456
rect 9612 -616 11806 -456
rect 12200 -616 21393 -456
rect -1291 -1006 21393 -616
rect 8021 -1126 8549 -1096
rect 8021 -1466 8051 -1126
rect 8519 -1466 8549 -1126
rect 8021 -1496 8549 -1466
rect -2821 -1620 -9 -1560
rect -2821 -2070 -2762 -1620
rect -1881 -2070 -9 -1620
rect -2821 -2130 -9 -2070
rect 20113 -1620 22925 -1560
rect 20113 -2070 21985 -1620
rect 22866 -2070 22925 -1620
rect 20113 -2130 22925 -2070
rect 6622 -2704 7622 -2684
rect 6622 -3234 6644 -2704
rect 7038 -2744 7622 -2704
rect 7563 -3194 7622 -2744
rect 7038 -3234 7622 -3194
rect 6622 -3254 7622 -3234
rect 13078 -2704 14078 -2684
rect 13078 -3234 13100 -2704
rect 13494 -2744 14078 -2704
rect 14019 -3194 14078 -2744
rect 13494 -3234 14078 -3194
rect 13078 -3254 14078 -3234
rect -2821 -3442 22925 -3382
rect -2821 -3892 -950 -3442
rect -69 -3772 20173 -3442
rect -69 -3892 9217 -3772
rect -2821 -3932 9217 -3892
rect 9611 -3892 20173 -3772
rect 21054 -3892 22925 -3442
rect 9611 -3932 22925 -3892
rect -2821 -3952 22925 -3932
rect -1291 -4100 21393 -4080
rect -1291 -4260 10512 -4100
rect 10906 -4260 21393 -4100
rect -1291 -4650 21393 -4260
rect 8021 -4770 8549 -4740
rect 8021 -5110 8051 -4770
rect 8519 -5110 8549 -4770
rect 8021 -5140 8549 -5110
rect -2821 -5264 -9 -5204
rect -2821 -5714 -2762 -5264
rect -1881 -5714 -9 -5264
rect -2821 -5774 -9 -5714
rect 20113 -5264 22925 -5204
rect 20113 -5714 21985 -5264
rect 22866 -5714 22925 -5264
rect 20113 -5774 22925 -5714
rect -2821 -7086 -9 -7026
rect -2821 -7536 -950 -7086
rect -69 -7536 -9 -7086
rect -2821 -7596 -9 -7536
rect 20113 -7086 22925 -7026
rect 20113 -7536 20173 -7086
rect 21054 -7536 22925 -7086
rect 20113 -7596 22925 -7536
<< via4 >>
rect 8051 38780 8519 39020
rect 9880 38280 10820 38520
rect 12108 38280 12576 38520
rect 8051 37428 8519 37768
rect -950 21616 -69 22066
rect 20173 21616 21054 22066
rect -2762 19794 -1881 20244
rect 21985 19794 22866 20244
rect -950 17972 -69 18422
rect 20173 17972 21054 18422
rect -2762 16150 -1881 16600
rect 21985 16150 22866 16600
rect -950 14328 -69 14778
rect 20173 14328 21054 14778
rect -2762 12506 -1881 12956
rect 21985 12506 22866 12956
rect -950 10684 -69 11134
rect 20173 10684 21054 11134
rect -2762 8862 -1881 9312
rect 21985 8862 22866 9312
rect 6682 7738 7038 8188
rect 7038 7738 7563 8188
rect 13138 7738 13494 8188
rect 13494 7738 14019 8188
rect -950 7040 -69 7490
rect 20173 7040 21054 7490
rect 8051 5822 8519 6162
rect -2762 5218 -1881 5668
rect 21985 5218 22866 5668
rect 6682 4094 7038 4544
rect 7038 4094 7563 4544
rect 13138 4094 13494 4544
rect 13494 4094 14019 4544
rect -950 3396 -69 3846
rect 20173 3396 21054 3846
rect 8051 2178 8519 2518
rect -2762 1574 -1881 2024
rect 21985 1574 22866 2024
rect 6682 450 7038 900
rect 7038 450 7563 900
rect 13138 450 13494 900
rect 13494 450 14019 900
rect -950 -248 -69 202
rect 20173 -248 21054 202
rect 8051 -1466 8519 -1126
rect -2762 -2070 -1881 -1620
rect 21985 -2070 22866 -1620
rect 6682 -3194 7038 -2744
rect 7038 -3194 7563 -2744
rect 13138 -3194 13494 -2744
rect 13494 -3194 14019 -2744
rect -950 -3892 -69 -3442
rect 20173 -3892 21054 -3442
rect 8051 -5110 8519 -4770
rect -2762 -5714 -1881 -5264
rect 21985 -5714 22866 -5264
rect -950 -7536 -69 -7086
rect 20173 -7536 21054 -7086
<< metal5 >>
rect 8021 39020 8549 39050
rect 8021 38780 8051 39020
rect 8519 38780 8549 39020
rect -2821 20244 -1821 22126
rect -2821 19794 -2762 20244
rect -1881 19794 -1821 20244
rect -2821 16600 -1821 19794
rect -2821 16150 -2762 16600
rect -1881 16150 -1821 16600
rect -2821 12956 -1821 16150
rect -2821 12506 -2762 12956
rect -1881 12506 -1821 12956
rect -2821 9312 -1821 12506
rect -2821 8862 -2762 9312
rect -1881 8862 -1821 9312
rect -2821 5668 -1821 8862
rect -2821 5218 -2762 5668
rect -1881 5218 -1821 5668
rect -2821 2024 -1821 5218
rect -2821 1574 -2762 2024
rect -1881 1574 -1821 2024
rect -2821 -1620 -1821 1574
rect -2821 -2070 -2762 -1620
rect -1881 -2070 -1821 -1620
rect -2821 -5264 -1821 -2070
rect -2821 -5714 -2762 -5264
rect -1881 -5714 -1821 -5264
rect -2821 -7596 -1821 -5714
rect -1009 22066 -9 22126
rect -1009 21616 -950 22066
rect -69 21616 -9 22066
rect -1009 18422 -9 21616
rect -1009 17972 -950 18422
rect -69 17972 -9 18422
rect -1009 14778 -9 17972
rect -1009 14328 -950 14778
rect -69 14328 -9 14778
rect -1009 11134 -9 14328
rect -1009 10684 -950 11134
rect -69 10684 -9 11134
rect -1009 7490 -9 10684
rect -1009 7040 -950 7490
rect -69 7040 -9 7490
rect -1009 3846 -9 7040
rect -1009 3396 -950 3846
rect -69 3396 -9 3846
rect -1009 202 -9 3396
rect -1009 -248 -950 202
rect -69 -248 -9 202
rect -1009 -3442 -9 -248
rect -1009 -3892 -950 -3442
rect -69 -3892 -9 -3442
rect -1009 -7086 -9 -3892
rect -1009 -7536 -950 -7086
rect -69 -7536 -9 -7086
rect 6622 8188 7622 38136
rect 6622 7738 6682 8188
rect 7563 7738 7622 8188
rect 6622 4544 7622 7738
rect 6622 4094 6682 4544
rect 7563 4094 7622 4544
rect 6622 900 7622 4094
rect 6622 450 6682 900
rect 7563 450 7622 900
rect 6622 -2744 7622 450
rect 6622 -3194 6682 -2744
rect 7563 -3194 7622 -2744
rect 6622 -7264 7622 -3194
rect 8021 37768 8549 38780
rect 9850 38520 10850 38750
rect 9850 38280 9880 38520
rect 10820 38280 10850 38520
rect 9850 38250 10850 38280
rect 12078 38520 12606 39050
rect 12078 38280 12108 38520
rect 12576 38280 12606 38520
rect 8021 37428 8051 37768
rect 8519 37428 8549 37768
rect 8021 6162 8549 37428
rect 12078 37310 12606 38280
rect 8021 5822 8051 6162
rect 8519 5822 8549 6162
rect 8021 2518 8549 5822
rect 8021 2178 8051 2518
rect 8519 2178 8549 2518
rect 8021 -1126 8549 2178
rect 8021 -1466 8051 -1126
rect 8519 -1466 8549 -1126
rect 8021 -4770 8549 -1466
rect 8021 -5110 8051 -4770
rect 8519 -5110 8549 -4770
rect 8021 -5418 8549 -5110
rect 13078 8188 14078 38136
rect 13078 7738 13138 8188
rect 14019 7738 14078 8188
rect 13078 4544 14078 7738
rect 13078 4094 13138 4544
rect 14019 4094 14078 4544
rect 13078 900 14078 4094
rect 13078 450 13138 900
rect 14019 450 14078 900
rect 13078 -2744 14078 450
rect 13078 -3194 13138 -2744
rect 14019 -3194 14078 -2744
rect 13078 -7264 14078 -3194
rect 20113 22066 21113 22126
rect 20113 21616 20173 22066
rect 21054 21616 21113 22066
rect 20113 18422 21113 21616
rect 20113 17972 20173 18422
rect 21054 17972 21113 18422
rect 20113 14778 21113 17972
rect 20113 14328 20173 14778
rect 21054 14328 21113 14778
rect 20113 11134 21113 14328
rect 20113 10684 20173 11134
rect 21054 10684 21113 11134
rect 20113 7490 21113 10684
rect 20113 7040 20173 7490
rect 21054 7040 21113 7490
rect 20113 3846 21113 7040
rect 20113 3396 20173 3846
rect 21054 3396 21113 3846
rect 20113 202 21113 3396
rect 20113 -248 20173 202
rect 21054 -248 21113 202
rect 20113 -3442 21113 -248
rect 20113 -3892 20173 -3442
rect 21054 -3892 21113 -3442
rect 20113 -7086 21113 -3892
rect -1009 -7596 -9 -7536
rect 20113 -7536 20173 -7086
rect 21054 -7536 21113 -7086
rect 20113 -7596 21113 -7536
rect 21925 20244 22925 22126
rect 21925 19794 21985 20244
rect 22866 19794 22925 20244
rect 21925 16600 22925 19794
rect 21925 16150 21985 16600
rect 22866 16150 22925 16600
rect 21925 12956 22925 16150
rect 21925 12506 21985 12956
rect 22866 12506 22925 12956
rect 21925 9312 22925 12506
rect 21925 8862 21985 9312
rect 22866 8862 22925 9312
rect 21925 5668 22925 8862
rect 21925 5218 21985 5668
rect 22866 5218 22925 5668
rect 21925 2024 22925 5218
rect 21925 1574 21985 2024
rect 22866 1574 22925 2024
rect 21925 -1620 22925 1574
rect 21925 -2070 21985 -1620
rect 22866 -2070 22925 -1620
rect 21925 -5264 22925 -2070
rect 21925 -5714 21985 -5264
rect 22866 -5714 22925 -5264
rect 21925 -7596 22925 -5714
use osc_nfet_w15_nf4_cc  osc_nfet_w15_nf4_cc_0
timestamp 1697705955
transform 1 0 9060 0 1 -5703
box -4 -238 2584 1959
use osc_nfet_w30_nf4_cc  osc_nfet_w30_nf4_cc_0
timestamp 1698146509
transform 1 0 7762 0 1 -2057
box 0 -240 5176 1957
use osc_nfet_w60_nf4_cc  osc_nfet_w60_nf4_cc_0
timestamp 1698146509
transform 1 0 4 0 1 1587
box 5172 -240 15524 1957
use osc_nfet_w120_nf4_cc  osc_nfet_w120_nf4_cc_0
timestamp 1698146509
transform 1 0 2 0 1 5229
box -4 -238 20700 1959
use sky130_fd_pr__cap_mim_m3_1_RX9LCP  sky130_fd_pr__cap_mim_m3_1_RX9LCP_0
timestamp 1696346236
transform 0 -1 20753 -1 0 -6400
box -786 -640 786 640
use sky130_fd_pr__cap_mim_m3_1_RX9LCP  sky130_fd_pr__cap_mim_m3_1_RX9LCP_1
timestamp 1696346236
transform 0 -1 22285 1 0 -6398
box -786 -640 786 640
use sky130_fd_pr__cap_mim_m3_1_RX9LCP  sky130_fd_pr__cap_mim_m3_1_RX9LCP_2
timestamp 1696346236
transform 0 -1 22285 -1 0 -4576
box -786 -640 786 640
use sky130_fd_pr__cap_mim_m3_1_RX9LCP  sky130_fd_pr__cap_mim_m3_1_RX9LCP_3
timestamp 1696346236
transform 0 -1 20753 1 0 -4578
box -786 -640 786 640
use sky130_fd_pr__cap_mim_m3_1_RX9LCP  sky130_fd_pr__cap_mim_m3_1_RX9LCP_4
timestamp 1696346236
transform 0 -1 20753 -1 0 -2756
box -786 -640 786 640
use sky130_fd_pr__cap_mim_m3_1_RX9LCP  sky130_fd_pr__cap_mim_m3_1_RX9LCP_5
timestamp 1696346236
transform 0 -1 22285 1 0 -2754
box -786 -640 786 640
use sky130_fd_pr__cap_mim_m3_1_RX9LCP  sky130_fd_pr__cap_mim_m3_1_RX9LCP_6
timestamp 1696346236
transform 0 -1 20753 1 0 -934
box -786 -640 786 640
use sky130_fd_pr__cap_mim_m3_1_RX9LCP  sky130_fd_pr__cap_mim_m3_1_RX9LCP_7
timestamp 1696346236
transform 0 -1 22285 -1 0 -932
box -786 -640 786 640
use sky130_fd_pr__cap_mim_m3_1_RX9LCP  sky130_fd_pr__cap_mim_m3_1_RX9LCP_8
timestamp 1696346236
transform 0 -1 20753 -1 0 888
box -786 -640 786 640
use sky130_fd_pr__cap_mim_m3_1_RX9LCP  sky130_fd_pr__cap_mim_m3_1_RX9LCP_9
timestamp 1696346236
transform 0 -1 22283 1 0 888
box -786 -640 786 640
use sky130_fd_pr__cap_mim_m3_1_RX9LCP  sky130_fd_pr__cap_mim_m3_1_RX9LCP_10
timestamp 1696346236
transform 0 -1 22283 -1 0 2710
box -786 -640 786 640
use sky130_fd_pr__cap_mim_m3_1_RX9LCP  sky130_fd_pr__cap_mim_m3_1_RX9LCP_11
timestamp 1696346236
transform 0 -1 20753 1 0 2710
box -786 -640 786 640
use sky130_fd_pr__cap_mim_m3_1_RX9LCP  sky130_fd_pr__cap_mim_m3_1_RX9LCP_12
timestamp 1696346236
transform 0 -1 20753 -1 0 4532
box -786 -640 786 640
use sky130_fd_pr__cap_mim_m3_1_RX9LCP  sky130_fd_pr__cap_mim_m3_1_RX9LCP_13
timestamp 1696346236
transform 0 -1 22283 1 0 4532
box -786 -640 786 640
use sky130_fd_pr__cap_mim_m3_1_RX9LCP  sky130_fd_pr__cap_mim_m3_1_RX9LCP_14
timestamp 1696346236
transform 0 -1 22283 -1 0 6354
box -786 -640 786 640
use sky130_fd_pr__cap_mim_m3_1_RX9LCP  sky130_fd_pr__cap_mim_m3_1_RX9LCP_15
timestamp 1696346236
transform 0 -1 20753 1 0 6354
box -786 -640 786 640
use sky130_fd_pr__cap_mim_m3_1_RX9LCP  sky130_fd_pr__cap_mim_m3_1_RX9LCP_16
timestamp 1696346236
transform 0 -1 20753 -1 0 8176
box -786 -640 786 640
use sky130_fd_pr__cap_mim_m3_1_RX9LCP  sky130_fd_pr__cap_mim_m3_1_RX9LCP_17
timestamp 1696346236
transform 0 -1 22283 1 0 8176
box -786 -640 786 640
use sky130_fd_pr__cap_mim_m3_1_RX9LCP  sky130_fd_pr__cap_mim_m3_1_RX9LCP_18
timestamp 1696346236
transform 0 -1 22283 -1 0 9998
box -786 -640 786 640
use sky130_fd_pr__cap_mim_m3_1_RX9LCP  sky130_fd_pr__cap_mim_m3_1_RX9LCP_19
timestamp 1696346236
transform 0 -1 20753 1 0 9998
box -786 -640 786 640
use sky130_fd_pr__cap_mim_m3_1_RX9LCP  sky130_fd_pr__cap_mim_m3_1_RX9LCP_20
timestamp 1696346236
transform 0 -1 20753 1 0 13642
box -786 -640 786 640
use sky130_fd_pr__cap_mim_m3_1_RX9LCP  sky130_fd_pr__cap_mim_m3_1_RX9LCP_21
timestamp 1696346236
transform 0 -1 20753 -1 0 11820
box -786 -640 786 640
use sky130_fd_pr__cap_mim_m3_1_RX9LCP  sky130_fd_pr__cap_mim_m3_1_RX9LCP_22
timestamp 1696346236
transform 0 -1 20753 -1 0 15464
box -786 -640 786 640
use sky130_fd_pr__cap_mim_m3_1_RX9LCP  sky130_fd_pr__cap_mim_m3_1_RX9LCP_23
timestamp 1696346236
transform 0 -1 22283 -1 0 13642
box -786 -640 786 640
use sky130_fd_pr__cap_mim_m3_1_RX9LCP  sky130_fd_pr__cap_mim_m3_1_RX9LCP_24
timestamp 1696346236
transform 0 -1 22283 1 0 11820
box -786 -640 786 640
use sky130_fd_pr__cap_mim_m3_1_RX9LCP  sky130_fd_pr__cap_mim_m3_1_RX9LCP_25
timestamp 1696346236
transform 0 -1 22283 1 0 15464
box -786 -640 786 640
use sky130_fd_pr__cap_mim_m3_1_RX9LCP  sky130_fd_pr__cap_mim_m3_1_RX9LCP_26
timestamp 1696346236
transform 0 -1 20753 1 0 20930
box -786 -640 786 640
use sky130_fd_pr__cap_mim_m3_1_RX9LCP  sky130_fd_pr__cap_mim_m3_1_RX9LCP_27
timestamp 1696346236
transform 0 -1 20753 1 0 17286
box -786 -640 786 640
use sky130_fd_pr__cap_mim_m3_1_RX9LCP  sky130_fd_pr__cap_mim_m3_1_RX9LCP_28
timestamp 1696346236
transform 0 -1 20753 -1 0 19108
box -786 -640 786 640
use sky130_fd_pr__cap_mim_m3_1_RX9LCP  sky130_fd_pr__cap_mim_m3_1_RX9LCP_29
timestamp 1696346236
transform 0 -1 22283 -1 0 20930
box -786 -640 786 640
use sky130_fd_pr__cap_mim_m3_1_RX9LCP  sky130_fd_pr__cap_mim_m3_1_RX9LCP_30
timestamp 1696346236
transform 0 -1 22283 -1 0 17286
box -786 -640 786 640
use sky130_fd_pr__cap_mim_m3_1_RX9LCP  sky130_fd_pr__cap_mim_m3_1_RX9LCP_31
timestamp 1696346236
transform 0 -1 22283 1 0 19108
box -786 -640 786 640
use sky130_fd_pr__cap_mim_m3_1_RX9LCP  sky130_fd_pr__cap_mim_m3_1_RX9LCP_32
timestamp 1696346236
transform 0 1 -649 1 0 20930
box -786 -640 786 640
use sky130_fd_pr__cap_mim_m3_1_RX9LCP  sky130_fd_pr__cap_mim_m3_1_RX9LCP_33
timestamp 1696346236
transform 0 1 -2181 -1 0 20928
box -786 -640 786 640
use sky130_fd_pr__cap_mim_m3_1_RX9LCP  sky130_fd_pr__cap_mim_m3_1_RX9LCP_34
timestamp 1696346236
transform 0 1 -2181 1 0 19106
box -786 -640 786 640
use sky130_fd_pr__cap_mim_m3_1_RX9LCP  sky130_fd_pr__cap_mim_m3_1_RX9LCP_35
timestamp 1696346236
transform 0 1 -649 -1 0 19108
box -786 -640 786 640
use sky130_fd_pr__cap_mim_m3_1_RX9LCP  sky130_fd_pr__cap_mim_m3_1_RX9LCP_36
timestamp 1696346236
transform 0 1 -649 1 0 17286
box -786 -640 786 640
use sky130_fd_pr__cap_mim_m3_1_RX9LCP  sky130_fd_pr__cap_mim_m3_1_RX9LCP_37
timestamp 1696346236
transform 0 1 -2181 -1 0 17284
box -786 -640 786 640
use sky130_fd_pr__cap_mim_m3_1_RX9LCP  sky130_fd_pr__cap_mim_m3_1_RX9LCP_38
timestamp 1696346236
transform 0 1 -649 -1 0 15464
box -786 -640 786 640
use sky130_fd_pr__cap_mim_m3_1_RX9LCP  sky130_fd_pr__cap_mim_m3_1_RX9LCP_39
timestamp 1696346236
transform 0 1 -2181 1 0 15462
box -786 -640 786 640
use sky130_fd_pr__cap_mim_m3_1_RX9LCP  sky130_fd_pr__cap_mim_m3_1_RX9LCP_40
timestamp 1696346236
transform 0 1 -649 1 0 13642
box -786 -640 786 640
use sky130_fd_pr__cap_mim_m3_1_RX9LCP  sky130_fd_pr__cap_mim_m3_1_RX9LCP_41
timestamp 1696346236
transform 0 1 -2179 -1 0 13642
box -786 -640 786 640
use sky130_fd_pr__cap_mim_m3_1_RX9LCP  sky130_fd_pr__cap_mim_m3_1_RX9LCP_42
timestamp 1696346236
transform 0 1 -2179 1 0 11820
box -786 -640 786 640
use sky130_fd_pr__cap_mim_m3_1_RX9LCP  sky130_fd_pr__cap_mim_m3_1_RX9LCP_43
timestamp 1696346236
transform 0 1 -649 -1 0 11820
box -786 -640 786 640
use sky130_fd_pr__cap_mim_m3_1_RX9LCP  sky130_fd_pr__cap_mim_m3_1_RX9LCP_44
timestamp 1696346236
transform 0 1 -649 1 0 9998
box -786 -640 786 640
use sky130_fd_pr__cap_mim_m3_1_RX9LCP  sky130_fd_pr__cap_mim_m3_1_RX9LCP_45
timestamp 1696346236
transform 0 1 -2179 -1 0 9998
box -786 -640 786 640
use sky130_fd_pr__cap_mim_m3_1_RX9LCP  sky130_fd_pr__cap_mim_m3_1_RX9LCP_46
timestamp 1696346236
transform 0 1 -2179 1 0 8176
box -786 -640 786 640
use sky130_fd_pr__cap_mim_m3_1_RX9LCP  sky130_fd_pr__cap_mim_m3_1_RX9LCP_47
timestamp 1696346236
transform 0 1 -649 -1 0 8176
box -786 -640 786 640
use sky130_fd_pr__cap_mim_m3_1_RX9LCP  sky130_fd_pr__cap_mim_m3_1_RX9LCP_48
timestamp 1696346236
transform 0 1 -649 1 0 6354
box -786 -640 786 640
use sky130_fd_pr__cap_mim_m3_1_RX9LCP  sky130_fd_pr__cap_mim_m3_1_RX9LCP_49
timestamp 1696346236
transform 0 1 -2179 -1 0 6354
box -786 -640 786 640
use sky130_fd_pr__cap_mim_m3_1_RX9LCP  sky130_fd_pr__cap_mim_m3_1_RX9LCP_50
timestamp 1696346236
transform 0 1 -2179 1 0 4532
box -786 -640 786 640
use sky130_fd_pr__cap_mim_m3_1_RX9LCP  sky130_fd_pr__cap_mim_m3_1_RX9LCP_51
timestamp 1696346236
transform 0 1 -649 -1 0 4532
box -786 -640 786 640
use sky130_fd_pr__cap_mim_m3_1_RX9LCP  sky130_fd_pr__cap_mim_m3_1_RX9LCP_52
timestamp 1696346236
transform 0 1 -649 -1 0 888
box -786 -640 786 640
use sky130_fd_pr__cap_mim_m3_1_RX9LCP  sky130_fd_pr__cap_mim_m3_1_RX9LCP_53
timestamp 1696346236
transform 0 1 -649 1 0 2710
box -786 -640 786 640
use sky130_fd_pr__cap_mim_m3_1_RX9LCP  sky130_fd_pr__cap_mim_m3_1_RX9LCP_54
timestamp 1696346236
transform 0 1 -649 1 0 -934
box -786 -640 786 640
use sky130_fd_pr__cap_mim_m3_1_RX9LCP  sky130_fd_pr__cap_mim_m3_1_RX9LCP_55
timestamp 1696346236
transform 0 1 -2179 1 0 888
box -786 -640 786 640
use sky130_fd_pr__cap_mim_m3_1_RX9LCP  sky130_fd_pr__cap_mim_m3_1_RX9LCP_56
timestamp 1696346236
transform 0 1 -2179 -1 0 2710
box -786 -640 786 640
use sky130_fd_pr__cap_mim_m3_1_RX9LCP  sky130_fd_pr__cap_mim_m3_1_RX9LCP_57
timestamp 1696346236
transform 0 1 -2179 -1 0 -934
box -786 -640 786 640
use sky130_fd_pr__cap_mim_m3_1_RX9LCP  sky130_fd_pr__cap_mim_m3_1_RX9LCP_58
timestamp 1696346236
transform 0 1 -649 -1 0 -6400
box -786 -640 786 640
use sky130_fd_pr__cap_mim_m3_1_RX9LCP  sky130_fd_pr__cap_mim_m3_1_RX9LCP_59
timestamp 1696346236
transform 0 1 -649 -1 0 -2756
box -786 -640 786 640
use sky130_fd_pr__cap_mim_m3_1_RX9LCP  sky130_fd_pr__cap_mim_m3_1_RX9LCP_60
timestamp 1696346236
transform 0 1 -649 1 0 -4578
box -786 -640 786 640
use sky130_fd_pr__cap_mim_m3_1_RX9LCP  sky130_fd_pr__cap_mim_m3_1_RX9LCP_61
timestamp 1696346236
transform 0 1 -2179 1 0 -6400
box -786 -640 786 640
use sky130_fd_pr__cap_mim_m3_1_RX9LCP  sky130_fd_pr__cap_mim_m3_1_RX9LCP_62
timestamp 1696346236
transform 0 1 -2179 1 0 -2756
box -786 -640 786 640
use sky130_fd_pr__cap_mim_m3_1_RX9LCP  sky130_fd_pr__cap_mim_m3_1_RX9LCP_63
timestamp 1696346236
transform 0 1 -2179 -1 0 -4578
box -786 -640 786 640
use uwb_inductor  uwb_inductor_0
timestamp 1698153454
transform 1 0 10350 0 1 40250
box -9750 -2114 9700 18700
<< labels >>
flabel locali 10280 -6994 10420 -6948 0 FreeSans 240 0 0 0 vss_osc
port 0 nsew
flabel metal2 20655 5146 20702 5242 0 FreeSans 240 0 0 0 en1_osc[3]
port 3 nsew
flabel metal2 15481 1502 15528 1598 0 FreeSans 240 0 0 0 en1_osc[2]
port 4 nsew
flabel metal2 12891 -2142 12938 -2046 0 FreeSans 240 0 0 0 en1_osc[1]
port 5 nsew
flabel metal2 11597 -5786 11644 -5690 0 FreeSans 240 0 0 0 en1_osc[0]
port 6 nsew
flabel metal2 20655 5002 20702 5098 0 FreeSans 240 0 0 0 en2_osc[3]
port 7 nsew
flabel metal2 15481 1358 15528 1454 0 FreeSans 240 0 0 0 en2_osc[2]
port 8 nsew
flabel metal2 12891 -2286 12938 -2190 0 FreeSans 240 0 0 0 en2_osc[1]
port 9 nsew
flabel metal2 11597 -5930 11644 -5834 0 FreeSans 240 0 0 0 en2_osc[0]
port 10 nsew
flabel metal5 6622 8248 7622 8736 0 FreeSans 800 0 0 0 outp_osc
port 2 nsew
flabel metal5 13078 8248 14078 8736 0 FreeSans 800 0 0 0 outn_osc
port 1 nsew
flabel metal5 9850 38550 10850 38650 0 FreeSans 1600 0 0 0 vdd_osc
port 11 nsew
<< end >>
