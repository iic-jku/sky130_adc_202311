magic
tech sky130A
magscale 1 2
timestamp 1696337182
<< metal3 >>
rect -1692 12012 -120 12040
rect -1692 10788 -204 12012
rect -140 10788 -120 12012
rect -1692 10760 -120 10788
rect 120 12012 1692 12040
rect 120 10788 1608 12012
rect 1672 10788 1692 12012
rect 120 10760 1692 10788
rect -1692 10492 -120 10520
rect -1692 9268 -204 10492
rect -140 9268 -120 10492
rect -1692 9240 -120 9268
rect 120 10492 1692 10520
rect 120 9268 1608 10492
rect 1672 9268 1692 10492
rect 120 9240 1692 9268
rect -1692 8972 -120 9000
rect -1692 7748 -204 8972
rect -140 7748 -120 8972
rect -1692 7720 -120 7748
rect 120 8972 1692 9000
rect 120 7748 1608 8972
rect 1672 7748 1692 8972
rect 120 7720 1692 7748
rect -1692 7452 -120 7480
rect -1692 6228 -204 7452
rect -140 6228 -120 7452
rect -1692 6200 -120 6228
rect 120 7452 1692 7480
rect 120 6228 1608 7452
rect 1672 6228 1692 7452
rect 120 6200 1692 6228
rect -1692 5932 -120 5960
rect -1692 4708 -204 5932
rect -140 4708 -120 5932
rect -1692 4680 -120 4708
rect 120 5932 1692 5960
rect 120 4708 1608 5932
rect 1672 4708 1692 5932
rect 120 4680 1692 4708
rect -1692 4412 -120 4440
rect -1692 3188 -204 4412
rect -140 3188 -120 4412
rect -1692 3160 -120 3188
rect 120 4412 1692 4440
rect 120 3188 1608 4412
rect 1672 3188 1692 4412
rect 120 3160 1692 3188
rect -1692 2892 -120 2920
rect -1692 1668 -204 2892
rect -140 1668 -120 2892
rect -1692 1640 -120 1668
rect 120 2892 1692 2920
rect 120 1668 1608 2892
rect 1672 1668 1692 2892
rect 120 1640 1692 1668
rect -1692 1372 -120 1400
rect -1692 148 -204 1372
rect -140 148 -120 1372
rect -1692 120 -120 148
rect 120 1372 1692 1400
rect 120 148 1608 1372
rect 1672 148 1692 1372
rect 120 120 1692 148
rect -1692 -148 -120 -120
rect -1692 -1372 -204 -148
rect -140 -1372 -120 -148
rect -1692 -1400 -120 -1372
rect 120 -148 1692 -120
rect 120 -1372 1608 -148
rect 1672 -1372 1692 -148
rect 120 -1400 1692 -1372
rect -1692 -1668 -120 -1640
rect -1692 -2892 -204 -1668
rect -140 -2892 -120 -1668
rect -1692 -2920 -120 -2892
rect 120 -1668 1692 -1640
rect 120 -2892 1608 -1668
rect 1672 -2892 1692 -1668
rect 120 -2920 1692 -2892
rect -1692 -3188 -120 -3160
rect -1692 -4412 -204 -3188
rect -140 -4412 -120 -3188
rect -1692 -4440 -120 -4412
rect 120 -3188 1692 -3160
rect 120 -4412 1608 -3188
rect 1672 -4412 1692 -3188
rect 120 -4440 1692 -4412
rect -1692 -4708 -120 -4680
rect -1692 -5932 -204 -4708
rect -140 -5932 -120 -4708
rect -1692 -5960 -120 -5932
rect 120 -4708 1692 -4680
rect 120 -5932 1608 -4708
rect 1672 -5932 1692 -4708
rect 120 -5960 1692 -5932
rect -1692 -6228 -120 -6200
rect -1692 -7452 -204 -6228
rect -140 -7452 -120 -6228
rect -1692 -7480 -120 -7452
rect 120 -6228 1692 -6200
rect 120 -7452 1608 -6228
rect 1672 -7452 1692 -6228
rect 120 -7480 1692 -7452
rect -1692 -7748 -120 -7720
rect -1692 -8972 -204 -7748
rect -140 -8972 -120 -7748
rect -1692 -9000 -120 -8972
rect 120 -7748 1692 -7720
rect 120 -8972 1608 -7748
rect 1672 -8972 1692 -7748
rect 120 -9000 1692 -8972
rect -1692 -9268 -120 -9240
rect -1692 -10492 -204 -9268
rect -140 -10492 -120 -9268
rect -1692 -10520 -120 -10492
rect 120 -9268 1692 -9240
rect 120 -10492 1608 -9268
rect 1672 -10492 1692 -9268
rect 120 -10520 1692 -10492
rect -1692 -10788 -120 -10760
rect -1692 -12012 -204 -10788
rect -140 -12012 -120 -10788
rect -1692 -12040 -120 -12012
rect 120 -10788 1692 -10760
rect 120 -12012 1608 -10788
rect 1672 -12012 1692 -10788
rect 120 -12040 1692 -12012
<< via3 >>
rect -204 10788 -140 12012
rect 1608 10788 1672 12012
rect -204 9268 -140 10492
rect 1608 9268 1672 10492
rect -204 7748 -140 8972
rect 1608 7748 1672 8972
rect -204 6228 -140 7452
rect 1608 6228 1672 7452
rect -204 4708 -140 5932
rect 1608 4708 1672 5932
rect -204 3188 -140 4412
rect 1608 3188 1672 4412
rect -204 1668 -140 2892
rect 1608 1668 1672 2892
rect -204 148 -140 1372
rect 1608 148 1672 1372
rect -204 -1372 -140 -148
rect 1608 -1372 1672 -148
rect -204 -2892 -140 -1668
rect 1608 -2892 1672 -1668
rect -204 -4412 -140 -3188
rect 1608 -4412 1672 -3188
rect -204 -5932 -140 -4708
rect 1608 -5932 1672 -4708
rect -204 -7452 -140 -6228
rect 1608 -7452 1672 -6228
rect -204 -8972 -140 -7748
rect 1608 -8972 1672 -7748
rect -204 -10492 -140 -9268
rect 1608 -10492 1672 -9268
rect -204 -12012 -140 -10788
rect 1608 -12012 1672 -10788
<< mimcap >>
rect -1652 11960 -452 12000
rect -1652 10840 -1612 11960
rect -492 10840 -452 11960
rect -1652 10800 -452 10840
rect 160 11960 1360 12000
rect 160 10840 200 11960
rect 1320 10840 1360 11960
rect 160 10800 1360 10840
rect -1652 10440 -452 10480
rect -1652 9320 -1612 10440
rect -492 9320 -452 10440
rect -1652 9280 -452 9320
rect 160 10440 1360 10480
rect 160 9320 200 10440
rect 1320 9320 1360 10440
rect 160 9280 1360 9320
rect -1652 8920 -452 8960
rect -1652 7800 -1612 8920
rect -492 7800 -452 8920
rect -1652 7760 -452 7800
rect 160 8920 1360 8960
rect 160 7800 200 8920
rect 1320 7800 1360 8920
rect 160 7760 1360 7800
rect -1652 7400 -452 7440
rect -1652 6280 -1612 7400
rect -492 6280 -452 7400
rect -1652 6240 -452 6280
rect 160 7400 1360 7440
rect 160 6280 200 7400
rect 1320 6280 1360 7400
rect 160 6240 1360 6280
rect -1652 5880 -452 5920
rect -1652 4760 -1612 5880
rect -492 4760 -452 5880
rect -1652 4720 -452 4760
rect 160 5880 1360 5920
rect 160 4760 200 5880
rect 1320 4760 1360 5880
rect 160 4720 1360 4760
rect -1652 4360 -452 4400
rect -1652 3240 -1612 4360
rect -492 3240 -452 4360
rect -1652 3200 -452 3240
rect 160 4360 1360 4400
rect 160 3240 200 4360
rect 1320 3240 1360 4360
rect 160 3200 1360 3240
rect -1652 2840 -452 2880
rect -1652 1720 -1612 2840
rect -492 1720 -452 2840
rect -1652 1680 -452 1720
rect 160 2840 1360 2880
rect 160 1720 200 2840
rect 1320 1720 1360 2840
rect 160 1680 1360 1720
rect -1652 1320 -452 1360
rect -1652 200 -1612 1320
rect -492 200 -452 1320
rect -1652 160 -452 200
rect 160 1320 1360 1360
rect 160 200 200 1320
rect 1320 200 1360 1320
rect 160 160 1360 200
rect -1652 -200 -452 -160
rect -1652 -1320 -1612 -200
rect -492 -1320 -452 -200
rect -1652 -1360 -452 -1320
rect 160 -200 1360 -160
rect 160 -1320 200 -200
rect 1320 -1320 1360 -200
rect 160 -1360 1360 -1320
rect -1652 -1720 -452 -1680
rect -1652 -2840 -1612 -1720
rect -492 -2840 -452 -1720
rect -1652 -2880 -452 -2840
rect 160 -1720 1360 -1680
rect 160 -2840 200 -1720
rect 1320 -2840 1360 -1720
rect 160 -2880 1360 -2840
rect -1652 -3240 -452 -3200
rect -1652 -4360 -1612 -3240
rect -492 -4360 -452 -3240
rect -1652 -4400 -452 -4360
rect 160 -3240 1360 -3200
rect 160 -4360 200 -3240
rect 1320 -4360 1360 -3240
rect 160 -4400 1360 -4360
rect -1652 -4760 -452 -4720
rect -1652 -5880 -1612 -4760
rect -492 -5880 -452 -4760
rect -1652 -5920 -452 -5880
rect 160 -4760 1360 -4720
rect 160 -5880 200 -4760
rect 1320 -5880 1360 -4760
rect 160 -5920 1360 -5880
rect -1652 -6280 -452 -6240
rect -1652 -7400 -1612 -6280
rect -492 -7400 -452 -6280
rect -1652 -7440 -452 -7400
rect 160 -6280 1360 -6240
rect 160 -7400 200 -6280
rect 1320 -7400 1360 -6280
rect 160 -7440 1360 -7400
rect -1652 -7800 -452 -7760
rect -1652 -8920 -1612 -7800
rect -492 -8920 -452 -7800
rect -1652 -8960 -452 -8920
rect 160 -7800 1360 -7760
rect 160 -8920 200 -7800
rect 1320 -8920 1360 -7800
rect 160 -8960 1360 -8920
rect -1652 -9320 -452 -9280
rect -1652 -10440 -1612 -9320
rect -492 -10440 -452 -9320
rect -1652 -10480 -452 -10440
rect 160 -9320 1360 -9280
rect 160 -10440 200 -9320
rect 1320 -10440 1360 -9320
rect 160 -10480 1360 -10440
rect -1652 -10840 -452 -10800
rect -1652 -11960 -1612 -10840
rect -492 -11960 -452 -10840
rect -1652 -12000 -452 -11960
rect 160 -10840 1360 -10800
rect 160 -11960 200 -10840
rect 1320 -11960 1360 -10840
rect 160 -12000 1360 -11960
<< mimcapcontact >>
rect -1612 10840 -492 11960
rect 200 10840 1320 11960
rect -1612 9320 -492 10440
rect 200 9320 1320 10440
rect -1612 7800 -492 8920
rect 200 7800 1320 8920
rect -1612 6280 -492 7400
rect 200 6280 1320 7400
rect -1612 4760 -492 5880
rect 200 4760 1320 5880
rect -1612 3240 -492 4360
rect 200 3240 1320 4360
rect -1612 1720 -492 2840
rect 200 1720 1320 2840
rect -1612 200 -492 1320
rect 200 200 1320 1320
rect -1612 -1320 -492 -200
rect 200 -1320 1320 -200
rect -1612 -2840 -492 -1720
rect 200 -2840 1320 -1720
rect -1612 -4360 -492 -3240
rect 200 -4360 1320 -3240
rect -1612 -5880 -492 -4760
rect 200 -5880 1320 -4760
rect -1612 -7400 -492 -6280
rect 200 -7400 1320 -6280
rect -1612 -8920 -492 -7800
rect 200 -8920 1320 -7800
rect -1612 -10440 -492 -9320
rect 200 -10440 1320 -9320
rect -1612 -11960 -492 -10840
rect 200 -11960 1320 -10840
<< metal4 >>
rect -1104 11961 -1000 12160
rect -224 12012 -120 12160
rect -1613 11960 -491 11961
rect -1613 10840 -1612 11960
rect -492 10840 -491 11960
rect -1613 10839 -491 10840
rect -1104 10441 -1000 10839
rect -224 10788 -204 12012
rect -140 10788 -120 12012
rect 708 11961 812 12160
rect 1588 12012 1692 12160
rect 199 11960 1321 11961
rect 199 10840 200 11960
rect 1320 10840 1321 11960
rect 199 10839 1321 10840
rect -224 10492 -120 10788
rect -1613 10440 -491 10441
rect -1613 9320 -1612 10440
rect -492 9320 -491 10440
rect -1613 9319 -491 9320
rect -1104 8921 -1000 9319
rect -224 9268 -204 10492
rect -140 9268 -120 10492
rect 708 10441 812 10839
rect 1588 10788 1608 12012
rect 1672 10788 1692 12012
rect 1588 10492 1692 10788
rect 199 10440 1321 10441
rect 199 9320 200 10440
rect 1320 9320 1321 10440
rect 199 9319 1321 9320
rect -224 8972 -120 9268
rect -1613 8920 -491 8921
rect -1613 7800 -1612 8920
rect -492 7800 -491 8920
rect -1613 7799 -491 7800
rect -1104 7401 -1000 7799
rect -224 7748 -204 8972
rect -140 7748 -120 8972
rect 708 8921 812 9319
rect 1588 9268 1608 10492
rect 1672 9268 1692 10492
rect 1588 8972 1692 9268
rect 199 8920 1321 8921
rect 199 7800 200 8920
rect 1320 7800 1321 8920
rect 199 7799 1321 7800
rect -224 7452 -120 7748
rect -1613 7400 -491 7401
rect -1613 6280 -1612 7400
rect -492 6280 -491 7400
rect -1613 6279 -491 6280
rect -1104 5881 -1000 6279
rect -224 6228 -204 7452
rect -140 6228 -120 7452
rect 708 7401 812 7799
rect 1588 7748 1608 8972
rect 1672 7748 1692 8972
rect 1588 7452 1692 7748
rect 199 7400 1321 7401
rect 199 6280 200 7400
rect 1320 6280 1321 7400
rect 199 6279 1321 6280
rect -224 5932 -120 6228
rect -1613 5880 -491 5881
rect -1613 4760 -1612 5880
rect -492 4760 -491 5880
rect -1613 4759 -491 4760
rect -1104 4361 -1000 4759
rect -224 4708 -204 5932
rect -140 4708 -120 5932
rect 708 5881 812 6279
rect 1588 6228 1608 7452
rect 1672 6228 1692 7452
rect 1588 5932 1692 6228
rect 199 5880 1321 5881
rect 199 4760 200 5880
rect 1320 4760 1321 5880
rect 199 4759 1321 4760
rect -224 4412 -120 4708
rect -1613 4360 -491 4361
rect -1613 3240 -1612 4360
rect -492 3240 -491 4360
rect -1613 3239 -491 3240
rect -1104 2841 -1000 3239
rect -224 3188 -204 4412
rect -140 3188 -120 4412
rect 708 4361 812 4759
rect 1588 4708 1608 5932
rect 1672 4708 1692 5932
rect 1588 4412 1692 4708
rect 199 4360 1321 4361
rect 199 3240 200 4360
rect 1320 3240 1321 4360
rect 199 3239 1321 3240
rect -224 2892 -120 3188
rect -1613 2840 -491 2841
rect -1613 1720 -1612 2840
rect -492 1720 -491 2840
rect -1613 1719 -491 1720
rect -1104 1321 -1000 1719
rect -224 1668 -204 2892
rect -140 1668 -120 2892
rect 708 2841 812 3239
rect 1588 3188 1608 4412
rect 1672 3188 1692 4412
rect 1588 2892 1692 3188
rect 199 2840 1321 2841
rect 199 1720 200 2840
rect 1320 1720 1321 2840
rect 199 1719 1321 1720
rect -224 1372 -120 1668
rect -1613 1320 -491 1321
rect -1613 200 -1612 1320
rect -492 200 -491 1320
rect -1613 199 -491 200
rect -1104 -199 -1000 199
rect -224 148 -204 1372
rect -140 148 -120 1372
rect 708 1321 812 1719
rect 1588 1668 1608 2892
rect 1672 1668 1692 2892
rect 1588 1372 1692 1668
rect 199 1320 1321 1321
rect 199 200 200 1320
rect 1320 200 1321 1320
rect 199 199 1321 200
rect -224 -148 -120 148
rect -1613 -200 -491 -199
rect -1613 -1320 -1612 -200
rect -492 -1320 -491 -200
rect -1613 -1321 -491 -1320
rect -1104 -1719 -1000 -1321
rect -224 -1372 -204 -148
rect -140 -1372 -120 -148
rect 708 -199 812 199
rect 1588 148 1608 1372
rect 1672 148 1692 1372
rect 1588 -148 1692 148
rect 199 -200 1321 -199
rect 199 -1320 200 -200
rect 1320 -1320 1321 -200
rect 199 -1321 1321 -1320
rect -224 -1668 -120 -1372
rect -1613 -1720 -491 -1719
rect -1613 -2840 -1612 -1720
rect -492 -2840 -491 -1720
rect -1613 -2841 -491 -2840
rect -1104 -3239 -1000 -2841
rect -224 -2892 -204 -1668
rect -140 -2892 -120 -1668
rect 708 -1719 812 -1321
rect 1588 -1372 1608 -148
rect 1672 -1372 1692 -148
rect 1588 -1668 1692 -1372
rect 199 -1720 1321 -1719
rect 199 -2840 200 -1720
rect 1320 -2840 1321 -1720
rect 199 -2841 1321 -2840
rect -224 -3188 -120 -2892
rect -1613 -3240 -491 -3239
rect -1613 -4360 -1612 -3240
rect -492 -4360 -491 -3240
rect -1613 -4361 -491 -4360
rect -1104 -4759 -1000 -4361
rect -224 -4412 -204 -3188
rect -140 -4412 -120 -3188
rect 708 -3239 812 -2841
rect 1588 -2892 1608 -1668
rect 1672 -2892 1692 -1668
rect 1588 -3188 1692 -2892
rect 199 -3240 1321 -3239
rect 199 -4360 200 -3240
rect 1320 -4360 1321 -3240
rect 199 -4361 1321 -4360
rect -224 -4708 -120 -4412
rect -1613 -4760 -491 -4759
rect -1613 -5880 -1612 -4760
rect -492 -5880 -491 -4760
rect -1613 -5881 -491 -5880
rect -1104 -6279 -1000 -5881
rect -224 -5932 -204 -4708
rect -140 -5932 -120 -4708
rect 708 -4759 812 -4361
rect 1588 -4412 1608 -3188
rect 1672 -4412 1692 -3188
rect 1588 -4708 1692 -4412
rect 199 -4760 1321 -4759
rect 199 -5880 200 -4760
rect 1320 -5880 1321 -4760
rect 199 -5881 1321 -5880
rect -224 -6228 -120 -5932
rect -1613 -6280 -491 -6279
rect -1613 -7400 -1612 -6280
rect -492 -7400 -491 -6280
rect -1613 -7401 -491 -7400
rect -1104 -7799 -1000 -7401
rect -224 -7452 -204 -6228
rect -140 -7452 -120 -6228
rect 708 -6279 812 -5881
rect 1588 -5932 1608 -4708
rect 1672 -5932 1692 -4708
rect 1588 -6228 1692 -5932
rect 199 -6280 1321 -6279
rect 199 -7400 200 -6280
rect 1320 -7400 1321 -6280
rect 199 -7401 1321 -7400
rect -224 -7748 -120 -7452
rect -1613 -7800 -491 -7799
rect -1613 -8920 -1612 -7800
rect -492 -8920 -491 -7800
rect -1613 -8921 -491 -8920
rect -1104 -9319 -1000 -8921
rect -224 -8972 -204 -7748
rect -140 -8972 -120 -7748
rect 708 -7799 812 -7401
rect 1588 -7452 1608 -6228
rect 1672 -7452 1692 -6228
rect 1588 -7748 1692 -7452
rect 199 -7800 1321 -7799
rect 199 -8920 200 -7800
rect 1320 -8920 1321 -7800
rect 199 -8921 1321 -8920
rect -224 -9268 -120 -8972
rect -1613 -9320 -491 -9319
rect -1613 -10440 -1612 -9320
rect -492 -10440 -491 -9320
rect -1613 -10441 -491 -10440
rect -1104 -10839 -1000 -10441
rect -224 -10492 -204 -9268
rect -140 -10492 -120 -9268
rect 708 -9319 812 -8921
rect 1588 -8972 1608 -7748
rect 1672 -8972 1692 -7748
rect 1588 -9268 1692 -8972
rect 199 -9320 1321 -9319
rect 199 -10440 200 -9320
rect 1320 -10440 1321 -9320
rect 199 -10441 1321 -10440
rect -224 -10788 -120 -10492
rect -1613 -10840 -491 -10839
rect -1613 -11960 -1612 -10840
rect -492 -11960 -491 -10840
rect -1613 -11961 -491 -11960
rect -1104 -12160 -1000 -11961
rect -224 -12012 -204 -10788
rect -140 -12012 -120 -10788
rect 708 -10839 812 -10441
rect 1588 -10492 1608 -9268
rect 1672 -10492 1692 -9268
rect 1588 -10788 1692 -10492
rect 199 -10840 1321 -10839
rect 199 -11960 200 -10840
rect 1320 -11960 1321 -10840
rect 199 -11961 1321 -11960
rect -224 -12160 -120 -12012
rect 708 -12160 812 -11961
rect 1588 -12012 1608 -10788
rect 1672 -12012 1692 -10788
rect 1588 -12160 1692 -12012
<< properties >>
string FIXED_BBOX 120 10760 1400 12040
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 6 l 6 val 76.56 carea 2.00 cperi 0.19 nx 2 ny 16 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
