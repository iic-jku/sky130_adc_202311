magic
tech sky130A
magscale 1 2
timestamp 1696930192
<< error_p >>
rect -365 -88 -307 -82
rect -173 -88 -115 -82
rect 211 -88 269 -82
rect -365 -122 -353 -88
rect -173 -122 -161 -88
rect 211 -122 223 -88
rect -365 -128 -307 -122
rect -173 -128 -115 -122
rect 211 -128 269 -122
<< pwell >>
rect -551 -260 551 260
<< nmos >>
rect -351 -50 -321 50
rect -255 -50 -225 50
rect -159 -50 -129 50
rect -63 -50 -33 50
rect 33 -50 63 50
rect 129 -50 159 50
rect 225 -50 255 50
rect 321 -50 351 50
<< ndiff >>
rect -413 38 -351 50
rect -413 -38 -401 38
rect -367 -38 -351 38
rect -413 -50 -351 -38
rect -321 38 -255 50
rect -321 -38 -305 38
rect -271 -38 -255 38
rect -321 -50 -255 -38
rect -225 38 -159 50
rect -225 -38 -209 38
rect -175 -38 -159 38
rect -225 -50 -159 -38
rect -129 38 -63 50
rect -129 -38 -113 38
rect -79 -38 -63 38
rect -129 -50 -63 -38
rect -33 38 33 50
rect -33 -38 -17 38
rect 17 -38 33 38
rect -33 -50 33 -38
rect 63 38 129 50
rect 63 -38 79 38
rect 113 -38 129 38
rect 63 -50 129 -38
rect 159 38 225 50
rect 159 -38 175 38
rect 209 -38 225 38
rect 159 -50 225 -38
rect 255 38 321 50
rect 255 -38 271 38
rect 305 -38 321 38
rect 255 -50 321 -38
rect 351 38 413 50
rect 351 -38 367 38
rect 401 -38 413 38
rect 351 -50 413 -38
<< ndiffc >>
rect -401 -38 -367 38
rect -305 -38 -271 38
rect -209 -38 -175 38
rect -113 -38 -79 38
rect -17 -38 17 38
rect 79 -38 113 38
rect 175 -38 209 38
rect 271 -38 305 38
rect 367 -38 401 38
<< psubdiff >>
rect -515 190 -419 224
rect 419 190 515 224
rect -515 128 -481 190
rect 481 128 515 190
rect -515 -190 -481 -128
rect 481 -190 515 -128
rect -515 -224 -419 -190
rect 419 -224 515 -190
<< psubdiffcont >>
rect -419 190 419 224
rect -515 -128 -481 128
rect 481 -128 515 128
rect -419 -224 419 -190
<< poly >>
rect -351 50 -321 76
rect -255 50 -225 76
rect -159 50 -129 76
rect -63 50 -33 76
rect 33 50 63 76
rect 129 50 159 76
rect 225 50 255 76
rect 321 50 351 76
rect -351 -72 -321 -50
rect -369 -88 -303 -72
rect -255 -76 -225 -50
rect -159 -72 -129 -50
rect -63 -72 -33 -50
rect 33 -72 63 -50
rect -369 -122 -353 -88
rect -319 -122 -303 -88
rect -369 -138 -303 -122
rect -177 -88 -111 -72
rect -177 -122 -161 -88
rect -127 -122 -111 -88
rect -177 -138 -111 -122
rect -63 -88 63 -72
rect 129 -76 159 -50
rect 225 -72 255 -50
rect -63 -122 -47 -88
rect 47 -122 63 -88
rect -63 -138 63 -122
rect 207 -88 273 -72
rect 321 -76 351 -50
rect 207 -122 223 -88
rect 257 -122 273 -88
rect 207 -138 273 -122
<< polycont >>
rect -353 -122 -319 -88
rect -161 -122 -127 -88
rect -47 -122 47 -88
rect 223 -122 257 -88
<< locali >>
rect -515 190 -419 224
rect 419 190 515 224
rect -515 128 -481 190
rect 481 128 515 190
rect -401 38 -367 54
rect -401 -54 -367 -38
rect -305 38 -271 54
rect -305 -54 -271 -38
rect -209 38 -175 54
rect -209 -54 -175 -38
rect -113 38 -79 54
rect -113 -54 -79 -38
rect -17 38 17 54
rect -17 -54 17 -38
rect 79 38 113 54
rect 79 -54 113 -38
rect 175 38 209 54
rect 175 -54 209 -38
rect 271 38 305 54
rect 271 -54 305 -38
rect 367 38 401 54
rect 367 -54 401 -38
rect -369 -122 -353 -88
rect -319 -122 -303 -88
rect -177 -122 -161 -88
rect -127 -122 -111 -88
rect -63 -122 -47 -88
rect 47 -122 63 -88
rect 207 -122 223 -88
rect 257 -122 273 -88
rect -515 -190 -481 -128
rect 481 -190 515 -128
rect -515 -224 -419 -190
rect 419 -224 515 -190
<< viali >>
rect -401 -38 -367 38
rect -305 -38 -271 38
rect -209 -38 -175 38
rect -113 -38 -79 38
rect -17 -38 17 38
rect 79 -38 113 38
rect 175 -38 209 38
rect 271 -38 305 38
rect 367 -38 401 38
rect -353 -122 -319 -88
rect -161 -122 -127 -88
rect -47 -122 47 -88
rect 223 -122 257 -88
<< metal1 >>
rect -407 38 -361 50
rect -407 -38 -401 38
rect -367 -38 -361 38
rect -407 -50 -361 -38
rect -311 38 -265 50
rect -311 -38 -305 38
rect -271 -38 -265 38
rect -311 -50 -265 -38
rect -215 38 -169 50
rect -215 -38 -209 38
rect -175 -38 -169 38
rect -215 -50 -169 -38
rect -119 38 -73 50
rect -119 -38 -113 38
rect -79 -38 -73 38
rect -119 -50 -73 -38
rect -23 38 23 50
rect -23 -38 -17 38
rect 17 -38 23 38
rect -23 -50 23 -38
rect 73 38 119 50
rect 73 -38 79 38
rect 113 -38 119 38
rect 73 -50 119 -38
rect 169 38 215 50
rect 169 -38 175 38
rect 209 -38 215 38
rect 169 -50 215 -38
rect 265 38 311 50
rect 265 -38 271 38
rect 305 -38 311 38
rect 265 -50 311 -38
rect 361 38 407 50
rect 361 -38 367 38
rect 401 -38 407 38
rect 361 -50 407 -38
rect -365 -88 -307 -82
rect -365 -122 -353 -88
rect -319 -122 -307 -88
rect -365 -128 -307 -122
rect -173 -88 -115 -82
rect -173 -122 -161 -88
rect -127 -122 -115 -88
rect -173 -128 -115 -122
rect -59 -88 59 -82
rect -59 -122 -47 -88
rect 47 -122 59 -88
rect -59 -128 59 -122
rect 211 -88 269 -82
rect 211 -122 223 -88
rect 257 -122 269 -88
rect 211 -128 269 -122
<< properties >>
string FIXED_BBOX -498 -207 498 207
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 0.5 l 0.150 m 1 nf 8 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
