magic
tech sky130A
magscale 1 2
timestamp 1699972208
<< nwell >>
rect 2877 38830 2941 38831
rect 1279 38265 3154 38830
rect 1279 38264 1569 38265
rect 1629 37421 3020 37437
rect 1463 37186 3020 37421
rect 1463 37177 2960 37186
rect 1463 37176 1925 37177
<< pwell >>
rect 898 39450 5230 39753
rect 898 36676 1213 39450
rect 4889 36758 5229 39450
rect 4889 36676 5230 36758
rect 898 36423 5230 36676
rect 898 36385 5229 36423
<< psubdiff >>
rect 924 39650 5204 39727
rect 924 39548 1335 39650
rect 1437 39548 1735 39650
rect 1837 39548 2135 39650
rect 2237 39548 2535 39650
rect 2637 39548 2935 39650
rect 3037 39548 3335 39650
rect 3437 39548 3735 39650
rect 3837 39548 4135 39650
rect 4237 39548 4535 39650
rect 4637 39548 5204 39650
rect 924 39476 5204 39548
rect 924 39467 1187 39476
rect 924 39365 1009 39467
rect 1111 39365 1187 39467
rect 924 39067 1187 39365
rect 924 38965 1009 39067
rect 1111 38965 1187 39067
rect 4915 39467 5203 39476
rect 4915 39365 5012 39467
rect 5114 39365 5203 39467
rect 4915 39067 5203 39365
rect 924 38667 1187 38965
rect 4915 38965 5012 39067
rect 5114 38965 5203 39067
rect 924 38565 1009 38667
rect 1111 38565 1187 38667
rect 924 38267 1187 38565
rect 924 38165 1009 38267
rect 1111 38165 1187 38267
rect 924 37867 1187 38165
rect 924 37765 1009 37867
rect 1111 37765 1187 37867
rect 924 37467 1187 37765
rect 924 37365 1009 37467
rect 1111 37365 1187 37467
rect 924 37067 1187 37365
rect 4915 38667 5203 38965
rect 4915 38565 5012 38667
rect 5114 38565 5203 38667
rect 4915 38267 5203 38565
rect 4915 38165 5012 38267
rect 5114 38165 5203 38267
rect 4915 37867 5203 38165
rect 4915 37765 5012 37867
rect 5114 37765 5203 37867
rect 4915 37467 5203 37765
rect 4915 37365 5012 37467
rect 5114 37365 5203 37467
rect 924 36965 1009 37067
rect 1111 36965 1187 37067
rect 4915 37067 5203 37365
rect 924 36650 1187 36965
rect 4915 36965 5012 37067
rect 5114 36965 5203 37067
rect 4915 36732 5203 36965
rect 4915 36650 5204 36732
rect 924 36649 2538 36650
rect 2685 36649 5204 36650
rect 924 36585 5204 36649
rect 924 36483 1009 36585
rect 1111 36483 1437 36585
rect 1539 36483 1837 36585
rect 1939 36483 2237 36585
rect 2339 36580 3437 36585
rect 2339 36483 2771 36580
rect 924 36478 2771 36483
rect 2873 36478 3098 36580
rect 3200 36483 3437 36580
rect 3539 36483 3837 36585
rect 3939 36483 4237 36585
rect 4339 36483 4637 36585
rect 4739 36483 5012 36585
rect 5114 36483 5204 36585
rect 3200 36478 5204 36483
rect 924 36449 5204 36478
rect 924 36411 5203 36449
<< psubdiffcont >>
rect 1335 39548 1437 39650
rect 1735 39548 1837 39650
rect 2135 39548 2237 39650
rect 2535 39548 2637 39650
rect 2935 39548 3037 39650
rect 3335 39548 3437 39650
rect 3735 39548 3837 39650
rect 4135 39548 4237 39650
rect 4535 39548 4637 39650
rect 1009 39365 1111 39467
rect 1009 38965 1111 39067
rect 5012 39365 5114 39467
rect 5012 38965 5114 39067
rect 1009 38565 1111 38667
rect 1009 38165 1111 38267
rect 1009 37765 1111 37867
rect 1009 37365 1111 37467
rect 5012 38565 5114 38667
rect 5012 38165 5114 38267
rect 5012 37765 5114 37867
rect 5012 37365 5114 37467
rect 1009 36965 1111 37067
rect 5012 36965 5114 37067
rect 1009 36483 1111 36585
rect 1437 36483 1539 36585
rect 1837 36483 1939 36585
rect 2237 36483 2339 36585
rect 2771 36478 2873 36580
rect 3098 36478 3200 36580
rect 3437 36483 3539 36585
rect 3837 36483 3939 36585
rect 4237 36483 4339 36585
rect 4637 36483 4739 36585
rect 5012 36483 5114 36585
<< poly >>
rect 2885 38981 2951 38994
rect 2885 38966 2901 38981
rect 2039 38964 2901 38966
rect 1650 38947 2901 38964
rect 2935 38947 2951 38981
rect 1650 38934 2951 38947
rect 1650 38870 2965 38892
rect 1650 38862 2921 38870
rect 1650 38819 1750 38862
rect 1808 38819 1908 38862
rect 2081 38816 2181 38862
rect 2239 38817 2339 38862
rect 2526 38817 2626 38862
rect 2684 38817 2784 38862
rect 2911 38836 2921 38862
rect 2955 38836 2965 38870
rect 2911 38820 2965 38836
rect 2526 38816 2538 38817
rect 2003 37144 2103 37197
rect 2161 37144 2261 37198
rect 2483 37144 2583 37198
rect 2641 37144 2741 37197
rect 2884 37172 2952 37182
rect 2884 37144 2902 37172
rect 2003 37138 2902 37144
rect 2936 37138 2952 37172
rect 2003 37114 2952 37138
rect 2003 37040 2969 37070
rect 2900 37037 2969 37040
rect 2900 37003 2917 37037
rect 2951 37003 2969 37037
rect 2900 36992 2969 37003
<< polycont >>
rect 2901 38947 2935 38981
rect 2921 38836 2955 38870
rect 2902 37138 2936 37172
rect 2917 37003 2951 37037
<< locali >>
rect 21068 75471 21140 75492
rect 503 75431 575 75452
rect 503 75397 522 75431
rect 556 75397 575 75431
rect 503 75376 575 75397
rect 629 75431 701 75452
rect 629 75397 648 75431
rect 682 75397 701 75431
rect 629 75376 701 75397
rect 749 75431 821 75452
rect 749 75397 768 75431
rect 802 75397 821 75431
rect 21068 75437 21087 75471
rect 21121 75437 21140 75471
rect 21068 75416 21140 75437
rect 21194 75471 21266 75492
rect 21194 75437 21213 75471
rect 21247 75437 21266 75471
rect 21194 75416 21266 75437
rect 21314 75471 21386 75492
rect 21314 75437 21333 75471
rect 21367 75437 21386 75471
rect 21314 75416 21386 75437
rect 749 75376 821 75397
rect 21068 75353 21140 75374
rect 503 75313 575 75334
rect 503 75279 522 75313
rect 556 75279 575 75313
rect 503 75258 575 75279
rect 629 75313 701 75334
rect 629 75279 648 75313
rect 682 75279 701 75313
rect 629 75258 701 75279
rect 749 75313 821 75334
rect 749 75279 768 75313
rect 802 75279 821 75313
rect 21068 75319 21087 75353
rect 21121 75319 21140 75353
rect 21068 75298 21140 75319
rect 21194 75353 21266 75374
rect 21194 75319 21213 75353
rect 21247 75319 21266 75353
rect 21194 75298 21266 75319
rect 21314 75353 21386 75374
rect 21314 75319 21333 75353
rect 21367 75319 21386 75353
rect 21314 75298 21386 75319
rect 749 75258 821 75279
rect 463 75039 946 75109
rect 463 75005 523 75039
rect 557 75005 645 75039
rect 679 75005 771 75039
rect 805 75005 946 75039
rect 463 74892 946 75005
rect 463 74858 523 74892
rect 557 74858 645 74892
rect 679 74858 771 74892
rect 805 74858 946 74892
rect 463 74755 946 74858
rect 463 74721 523 74755
rect 557 74721 645 74755
rect 679 74721 771 74755
rect 805 74721 946 74755
rect 463 74650 946 74721
rect 22010 74050 22082 74071
rect 22010 74016 22029 74050
rect 22063 74016 22082 74050
rect 22010 73995 22082 74016
rect 22136 74050 22208 74071
rect 22136 74016 22155 74050
rect 22189 74016 22208 74050
rect 22136 73995 22208 74016
rect 22256 74050 22328 74071
rect 22256 74016 22275 74050
rect 22309 74016 22328 74050
rect 22256 73995 22328 74016
rect 22010 73932 22082 73953
rect 22010 73898 22029 73932
rect 22063 73898 22082 73932
rect 22010 73877 22082 73898
rect 22136 73932 22208 73953
rect 22136 73898 22155 73932
rect 22189 73898 22208 73932
rect 22136 73877 22208 73898
rect 22256 73932 22328 73953
rect 22256 73898 22275 73932
rect 22309 73898 22328 73932
rect 22256 73877 22328 73898
rect 463 73279 946 73349
rect 463 73245 523 73279
rect 557 73245 645 73279
rect 679 73245 771 73279
rect 805 73245 946 73279
rect 463 73132 946 73245
rect 463 73098 523 73132
rect 557 73098 645 73132
rect 679 73098 771 73132
rect 805 73098 946 73132
rect 463 72995 946 73098
rect 463 72961 523 72995
rect 557 72961 645 72995
rect 679 72961 771 72995
rect 805 72961 946 72995
rect 463 72890 946 72961
rect 503 72758 575 72779
rect 503 72724 522 72758
rect 556 72724 575 72758
rect 503 72703 575 72724
rect 629 72758 701 72779
rect 629 72724 648 72758
rect 682 72724 701 72758
rect 629 72703 701 72724
rect 749 72758 821 72779
rect 749 72724 768 72758
rect 802 72724 821 72758
rect 749 72703 821 72724
rect 21068 72674 21140 72695
rect 503 72640 575 72661
rect 503 72606 522 72640
rect 556 72606 575 72640
rect 503 72585 575 72606
rect 629 72640 701 72661
rect 629 72606 648 72640
rect 682 72606 701 72640
rect 629 72585 701 72606
rect 749 72640 821 72661
rect 749 72606 768 72640
rect 802 72606 821 72640
rect 21068 72640 21087 72674
rect 21121 72640 21140 72674
rect 21068 72619 21140 72640
rect 21194 72674 21266 72695
rect 21194 72640 21213 72674
rect 21247 72640 21266 72674
rect 21194 72619 21266 72640
rect 21314 72674 21386 72695
rect 21314 72640 21333 72674
rect 21367 72640 21386 72674
rect 21314 72619 21386 72640
rect 749 72585 821 72606
rect 21068 72556 21140 72577
rect 21068 72522 21087 72556
rect 21121 72522 21140 72556
rect 21068 72501 21140 72522
rect 21194 72556 21266 72577
rect 21194 72522 21213 72556
rect 21247 72522 21266 72556
rect 21194 72501 21266 72522
rect 21314 72556 21386 72577
rect 21314 72522 21333 72556
rect 21367 72522 21386 72556
rect 21314 72501 21386 72522
rect 21068 71471 21140 71492
rect 503 71431 575 71452
rect 503 71397 522 71431
rect 556 71397 575 71431
rect 503 71376 575 71397
rect 629 71431 701 71452
rect 629 71397 648 71431
rect 682 71397 701 71431
rect 629 71376 701 71397
rect 749 71431 821 71452
rect 749 71397 768 71431
rect 802 71397 821 71431
rect 21068 71437 21087 71471
rect 21121 71437 21140 71471
rect 21068 71416 21140 71437
rect 21194 71471 21266 71492
rect 21194 71437 21213 71471
rect 21247 71437 21266 71471
rect 21194 71416 21266 71437
rect 21314 71471 21386 71492
rect 21314 71437 21333 71471
rect 21367 71437 21386 71471
rect 21314 71416 21386 71437
rect 749 71376 821 71397
rect 21068 71353 21140 71374
rect 503 71313 575 71334
rect 503 71279 522 71313
rect 556 71279 575 71313
rect 503 71258 575 71279
rect 629 71313 701 71334
rect 629 71279 648 71313
rect 682 71279 701 71313
rect 629 71258 701 71279
rect 749 71313 821 71334
rect 749 71279 768 71313
rect 802 71279 821 71313
rect 21068 71319 21087 71353
rect 21121 71319 21140 71353
rect 21068 71298 21140 71319
rect 21194 71353 21266 71374
rect 21194 71319 21213 71353
rect 21247 71319 21266 71353
rect 21194 71298 21266 71319
rect 21314 71353 21386 71374
rect 21314 71319 21333 71353
rect 21367 71319 21386 71353
rect 21314 71298 21386 71319
rect 749 71258 821 71279
rect 463 71039 946 71109
rect 463 71005 523 71039
rect 557 71005 645 71039
rect 679 71005 771 71039
rect 805 71005 946 71039
rect 463 70892 946 71005
rect 463 70858 523 70892
rect 557 70858 645 70892
rect 679 70858 771 70892
rect 805 70858 946 70892
rect 463 70755 946 70858
rect 463 70721 523 70755
rect 557 70721 645 70755
rect 679 70721 771 70755
rect 805 70721 946 70755
rect 463 70650 946 70721
rect 22010 70050 22082 70071
rect 22010 70016 22029 70050
rect 22063 70016 22082 70050
rect 22010 69995 22082 70016
rect 22136 70050 22208 70071
rect 22136 70016 22155 70050
rect 22189 70016 22208 70050
rect 22136 69995 22208 70016
rect 22256 70050 22328 70071
rect 22256 70016 22275 70050
rect 22309 70016 22328 70050
rect 22256 69995 22328 70016
rect 22010 69932 22082 69953
rect 22010 69898 22029 69932
rect 22063 69898 22082 69932
rect 22010 69877 22082 69898
rect 22136 69932 22208 69953
rect 22136 69898 22155 69932
rect 22189 69898 22208 69932
rect 22136 69877 22208 69898
rect 22256 69932 22328 69953
rect 22256 69898 22275 69932
rect 22309 69898 22328 69932
rect 22256 69877 22328 69898
rect 463 69279 946 69349
rect 463 69245 523 69279
rect 557 69245 645 69279
rect 679 69245 771 69279
rect 805 69245 946 69279
rect 463 69132 946 69245
rect 463 69098 523 69132
rect 557 69098 645 69132
rect 679 69098 771 69132
rect 805 69098 946 69132
rect 463 68995 946 69098
rect 463 68961 523 68995
rect 557 68961 645 68995
rect 679 68961 771 68995
rect 805 68961 946 68995
rect 463 68890 946 68961
rect 503 68758 575 68779
rect 503 68724 522 68758
rect 556 68724 575 68758
rect 503 68703 575 68724
rect 629 68758 701 68779
rect 629 68724 648 68758
rect 682 68724 701 68758
rect 629 68703 701 68724
rect 749 68758 821 68779
rect 749 68724 768 68758
rect 802 68724 821 68758
rect 749 68703 821 68724
rect 21068 68674 21140 68695
rect 503 68640 575 68661
rect 503 68606 522 68640
rect 556 68606 575 68640
rect 503 68585 575 68606
rect 629 68640 701 68661
rect 629 68606 648 68640
rect 682 68606 701 68640
rect 629 68585 701 68606
rect 749 68640 821 68661
rect 749 68606 768 68640
rect 802 68606 821 68640
rect 21068 68640 21087 68674
rect 21121 68640 21140 68674
rect 21068 68619 21140 68640
rect 21194 68674 21266 68695
rect 21194 68640 21213 68674
rect 21247 68640 21266 68674
rect 21194 68619 21266 68640
rect 21314 68674 21386 68695
rect 21314 68640 21333 68674
rect 21367 68640 21386 68674
rect 21314 68619 21386 68640
rect 749 68585 821 68606
rect 21068 68556 21140 68577
rect 21068 68522 21087 68556
rect 21121 68522 21140 68556
rect 21068 68501 21140 68522
rect 21194 68556 21266 68577
rect 21194 68522 21213 68556
rect 21247 68522 21266 68556
rect 21194 68501 21266 68522
rect 21314 68556 21386 68577
rect 21314 68522 21333 68556
rect 21367 68522 21386 68556
rect 21314 68501 21386 68522
rect 21068 67471 21140 67492
rect 503 67429 575 67450
rect 503 67395 522 67429
rect 556 67395 575 67429
rect 503 67374 575 67395
rect 629 67429 701 67450
rect 629 67395 648 67429
rect 682 67395 701 67429
rect 629 67374 701 67395
rect 749 67429 821 67450
rect 749 67395 768 67429
rect 802 67395 821 67429
rect 21068 67437 21087 67471
rect 21121 67437 21140 67471
rect 21068 67416 21140 67437
rect 21194 67471 21266 67492
rect 21194 67437 21213 67471
rect 21247 67437 21266 67471
rect 21194 67416 21266 67437
rect 21314 67471 21386 67492
rect 21314 67437 21333 67471
rect 21367 67437 21386 67471
rect 21314 67416 21386 67437
rect 749 67374 821 67395
rect 21068 67353 21140 67374
rect 503 67311 575 67332
rect 503 67277 522 67311
rect 556 67277 575 67311
rect 503 67256 575 67277
rect 629 67311 701 67332
rect 629 67277 648 67311
rect 682 67277 701 67311
rect 629 67256 701 67277
rect 749 67311 821 67332
rect 749 67277 768 67311
rect 802 67277 821 67311
rect 21068 67319 21087 67353
rect 21121 67319 21140 67353
rect 21068 67298 21140 67319
rect 21194 67353 21266 67374
rect 21194 67319 21213 67353
rect 21247 67319 21266 67353
rect 21194 67298 21266 67319
rect 21314 67353 21386 67374
rect 21314 67319 21333 67353
rect 21367 67319 21386 67353
rect 21314 67298 21386 67319
rect 749 67256 821 67277
rect 463 67039 946 67109
rect 463 67005 523 67039
rect 557 67005 645 67039
rect 679 67005 771 67039
rect 805 67005 946 67039
rect 463 66892 946 67005
rect 463 66858 523 66892
rect 557 66858 645 66892
rect 679 66858 771 66892
rect 805 66858 946 66892
rect 463 66755 946 66858
rect 463 66721 523 66755
rect 557 66721 645 66755
rect 679 66721 771 66755
rect 805 66721 946 66755
rect 463 66650 946 66721
rect 22010 66037 22082 66058
rect 22010 66003 22029 66037
rect 22063 66003 22082 66037
rect 22010 65982 22082 66003
rect 22136 66037 22208 66058
rect 22136 66003 22155 66037
rect 22189 66003 22208 66037
rect 22136 65982 22208 66003
rect 22256 66037 22328 66058
rect 22256 66003 22275 66037
rect 22309 66003 22328 66037
rect 22256 65982 22328 66003
rect 22010 65919 22082 65940
rect 22010 65885 22029 65919
rect 22063 65885 22082 65919
rect 22010 65864 22082 65885
rect 22136 65919 22208 65940
rect 22136 65885 22155 65919
rect 22189 65885 22208 65919
rect 22136 65864 22208 65885
rect 22256 65919 22328 65940
rect 22256 65885 22275 65919
rect 22309 65885 22328 65919
rect 22256 65864 22328 65885
rect 463 65280 946 65350
rect 463 65246 523 65280
rect 557 65246 645 65280
rect 679 65246 771 65280
rect 805 65246 946 65280
rect 463 65133 946 65246
rect 463 65099 523 65133
rect 557 65099 645 65133
rect 679 65099 771 65133
rect 805 65099 946 65133
rect 463 64996 946 65099
rect 463 64962 523 64996
rect 557 64962 645 64996
rect 679 64962 771 64996
rect 805 64962 946 64996
rect 463 64891 946 64962
rect 503 64689 575 64710
rect 503 64655 522 64689
rect 556 64655 575 64689
rect 503 64634 575 64655
rect 629 64689 701 64710
rect 629 64655 648 64689
rect 682 64655 701 64689
rect 629 64634 701 64655
rect 749 64689 821 64710
rect 749 64655 768 64689
rect 802 64655 821 64689
rect 749 64634 821 64655
rect 21068 64674 21140 64695
rect 21068 64640 21087 64674
rect 21121 64640 21140 64674
rect 21068 64619 21140 64640
rect 21194 64674 21266 64695
rect 21194 64640 21213 64674
rect 21247 64640 21266 64674
rect 21194 64619 21266 64640
rect 21314 64674 21386 64695
rect 21314 64640 21333 64674
rect 21367 64640 21386 64674
rect 21314 64619 21386 64640
rect 503 64571 575 64592
rect 503 64537 522 64571
rect 556 64537 575 64571
rect 503 64516 575 64537
rect 629 64571 701 64592
rect 629 64537 648 64571
rect 682 64537 701 64571
rect 629 64516 701 64537
rect 749 64571 821 64592
rect 749 64537 768 64571
rect 802 64537 821 64571
rect 749 64516 821 64537
rect 21068 64556 21140 64577
rect 21068 64522 21087 64556
rect 21121 64522 21140 64556
rect 21068 64501 21140 64522
rect 21194 64556 21266 64577
rect 21194 64522 21213 64556
rect 21247 64522 21266 64556
rect 21194 64501 21266 64522
rect 21314 64556 21386 64577
rect 21314 64522 21333 64556
rect 21367 64522 21386 64556
rect 21314 64501 21386 64522
rect 503 63511 575 63532
rect 503 63477 522 63511
rect 556 63477 575 63511
rect 503 63456 575 63477
rect 629 63511 701 63532
rect 629 63477 648 63511
rect 682 63477 701 63511
rect 629 63456 701 63477
rect 749 63511 821 63532
rect 749 63477 768 63511
rect 802 63477 821 63511
rect 749 63456 821 63477
rect 21068 63471 21140 63492
rect 21068 63437 21087 63471
rect 21121 63437 21140 63471
rect 21068 63416 21140 63437
rect 21194 63471 21266 63492
rect 21194 63437 21213 63471
rect 21247 63437 21266 63471
rect 21194 63416 21266 63437
rect 21314 63471 21386 63492
rect 21314 63437 21333 63471
rect 21367 63437 21386 63471
rect 21314 63416 21386 63437
rect 503 63393 575 63414
rect 503 63359 522 63393
rect 556 63359 575 63393
rect 503 63338 575 63359
rect 629 63393 701 63414
rect 629 63359 648 63393
rect 682 63359 701 63393
rect 629 63338 701 63359
rect 749 63393 821 63414
rect 749 63359 768 63393
rect 802 63359 821 63393
rect 749 63338 821 63359
rect 21068 63353 21140 63374
rect 21068 63319 21087 63353
rect 21121 63319 21140 63353
rect 21068 63298 21140 63319
rect 21194 63353 21266 63374
rect 21194 63319 21213 63353
rect 21247 63319 21266 63353
rect 21194 63298 21266 63319
rect 21314 63353 21386 63374
rect 21314 63319 21333 63353
rect 21367 63319 21386 63353
rect 21314 63298 21386 63319
rect 464 63068 947 63109
rect 463 63039 947 63068
rect 463 63005 523 63039
rect 557 63005 645 63039
rect 679 63005 771 63039
rect 805 63005 947 63039
rect 463 62892 947 63005
rect 463 62858 523 62892
rect 557 62858 645 62892
rect 679 62858 771 62892
rect 805 62858 947 62892
rect 463 62755 947 62858
rect 463 62721 523 62755
rect 557 62721 645 62755
rect 679 62721 771 62755
rect 805 62721 947 62755
rect 463 62650 947 62721
rect 22010 62036 22082 62057
rect 22010 62002 22029 62036
rect 22063 62002 22082 62036
rect 22010 61981 22082 62002
rect 22136 62036 22208 62057
rect 22136 62002 22155 62036
rect 22189 62002 22208 62036
rect 22136 61981 22208 62002
rect 22256 62036 22328 62057
rect 22256 62002 22275 62036
rect 22309 62002 22328 62036
rect 22256 61981 22328 62002
rect 22010 61918 22082 61939
rect 22010 61884 22029 61918
rect 22063 61884 22082 61918
rect 22010 61863 22082 61884
rect 22136 61918 22208 61939
rect 22136 61884 22155 61918
rect 22189 61884 22208 61918
rect 22136 61863 22208 61884
rect 22256 61918 22328 61939
rect 22256 61884 22275 61918
rect 22309 61884 22328 61918
rect 22256 61863 22328 61884
rect 463 61280 946 61350
rect 463 61246 523 61280
rect 557 61246 645 61280
rect 679 61246 771 61280
rect 805 61246 946 61280
rect 463 61133 946 61246
rect 463 61099 523 61133
rect 557 61099 645 61133
rect 679 61099 771 61133
rect 805 61099 946 61133
rect 463 60996 946 61099
rect 463 60962 523 60996
rect 557 60962 645 60996
rect 679 60962 771 60996
rect 805 60962 946 60996
rect 463 60891 946 60962
rect 503 60663 575 60684
rect 503 60629 522 60663
rect 556 60629 575 60663
rect 503 60608 575 60629
rect 629 60663 701 60684
rect 629 60629 648 60663
rect 682 60629 701 60663
rect 629 60608 701 60629
rect 749 60663 821 60684
rect 749 60629 768 60663
rect 802 60629 821 60663
rect 749 60608 821 60629
rect 21068 60674 21140 60695
rect 21068 60640 21087 60674
rect 21121 60640 21140 60674
rect 21068 60619 21140 60640
rect 21194 60674 21266 60695
rect 21194 60640 21213 60674
rect 21247 60640 21266 60674
rect 21194 60619 21266 60640
rect 21314 60674 21386 60695
rect 21314 60640 21333 60674
rect 21367 60640 21386 60674
rect 21314 60619 21386 60640
rect 503 60545 575 60566
rect 503 60511 522 60545
rect 556 60511 575 60545
rect 503 60490 575 60511
rect 629 60545 701 60566
rect 629 60511 648 60545
rect 682 60511 701 60545
rect 629 60490 701 60511
rect 749 60545 821 60566
rect 749 60511 768 60545
rect 802 60511 821 60545
rect 749 60490 821 60511
rect 21068 60556 21140 60577
rect 21068 60522 21087 60556
rect 21121 60522 21140 60556
rect 21068 60501 21140 60522
rect 21194 60556 21266 60577
rect 21194 60522 21213 60556
rect 21247 60522 21266 60556
rect 21194 60501 21266 60522
rect 21314 60556 21386 60577
rect 21314 60522 21333 60556
rect 21367 60522 21386 60556
rect 21314 60501 21386 60522
rect 21068 59525 21140 59546
rect 21068 59491 21087 59525
rect 21121 59491 21140 59525
rect 503 59460 575 59481
rect 503 59426 522 59460
rect 556 59426 575 59460
rect 503 59405 575 59426
rect 629 59460 701 59481
rect 629 59426 648 59460
rect 682 59426 701 59460
rect 629 59405 701 59426
rect 749 59460 821 59481
rect 21068 59470 21140 59491
rect 21194 59525 21266 59546
rect 21194 59491 21213 59525
rect 21247 59491 21266 59525
rect 21194 59470 21266 59491
rect 21314 59525 21386 59546
rect 21314 59491 21333 59525
rect 21367 59491 21386 59525
rect 21314 59470 21386 59491
rect 749 59426 768 59460
rect 802 59426 821 59460
rect 749 59405 821 59426
rect 21068 59407 21140 59428
rect 21068 59373 21087 59407
rect 21121 59373 21140 59407
rect 503 59342 575 59363
rect 503 59308 522 59342
rect 556 59308 575 59342
rect 503 59287 575 59308
rect 629 59342 701 59363
rect 629 59308 648 59342
rect 682 59308 701 59342
rect 629 59287 701 59308
rect 749 59342 821 59363
rect 21068 59352 21140 59373
rect 21194 59407 21266 59428
rect 21194 59373 21213 59407
rect 21247 59373 21266 59407
rect 21194 59352 21266 59373
rect 21314 59407 21386 59428
rect 21314 59373 21333 59407
rect 21367 59373 21386 59407
rect 21314 59352 21386 59373
rect 749 59308 768 59342
rect 802 59308 821 59342
rect 749 59287 821 59308
rect 464 59068 947 59109
rect 463 59039 947 59068
rect 463 59005 523 59039
rect 557 59005 645 59039
rect 679 59005 771 59039
rect 805 59005 947 59039
rect 463 58892 947 59005
rect 463 58858 523 58892
rect 557 58858 645 58892
rect 679 58858 771 58892
rect 805 58858 947 58892
rect 463 58755 947 58858
rect 463 58721 523 58755
rect 557 58721 645 58755
rect 679 58721 771 58755
rect 805 58721 947 58755
rect 463 58650 947 58721
rect 22010 58075 22082 58096
rect 22010 58041 22029 58075
rect 22063 58041 22082 58075
rect 22010 58020 22082 58041
rect 22136 58075 22208 58096
rect 22136 58041 22155 58075
rect 22189 58041 22208 58075
rect 22136 58020 22208 58041
rect 22256 58075 22328 58096
rect 22256 58041 22275 58075
rect 22309 58041 22328 58075
rect 22256 58020 22328 58041
rect 22010 57957 22082 57978
rect 22010 57923 22029 57957
rect 22063 57923 22082 57957
rect 22010 57902 22082 57923
rect 22136 57957 22208 57978
rect 22136 57923 22155 57957
rect 22189 57923 22208 57957
rect 22136 57902 22208 57923
rect 22256 57957 22328 57978
rect 22256 57923 22275 57957
rect 22309 57923 22328 57957
rect 22256 57902 22328 57923
rect 463 57278 946 57348
rect 463 57244 523 57278
rect 557 57244 645 57278
rect 679 57244 771 57278
rect 805 57244 946 57278
rect 463 57131 946 57244
rect 463 57097 523 57131
rect 557 57097 645 57131
rect 679 57097 771 57131
rect 805 57097 946 57131
rect 463 56994 946 57097
rect 463 56960 523 56994
rect 557 56960 645 56994
rect 679 56960 771 56994
rect 805 56960 946 56994
rect 463 56889 946 56960
rect 503 56683 575 56704
rect 503 56649 522 56683
rect 556 56649 575 56683
rect 503 56628 575 56649
rect 629 56683 701 56704
rect 629 56649 648 56683
rect 682 56649 701 56683
rect 629 56628 701 56649
rect 749 56683 821 56704
rect 749 56649 768 56683
rect 802 56649 821 56683
rect 749 56628 821 56649
rect 21068 56609 21140 56630
rect 503 56565 575 56586
rect 503 56531 522 56565
rect 556 56531 575 56565
rect 503 56510 575 56531
rect 629 56565 701 56586
rect 629 56531 648 56565
rect 682 56531 701 56565
rect 629 56510 701 56531
rect 749 56565 821 56586
rect 749 56531 768 56565
rect 802 56531 821 56565
rect 21068 56575 21087 56609
rect 21121 56575 21140 56609
rect 21068 56554 21140 56575
rect 21194 56609 21266 56630
rect 21194 56575 21213 56609
rect 21247 56575 21266 56609
rect 21194 56554 21266 56575
rect 21314 56609 21386 56630
rect 21314 56575 21333 56609
rect 21367 56575 21386 56609
rect 21314 56554 21386 56575
rect 749 56510 821 56531
rect 21068 56491 21140 56512
rect 21068 56457 21087 56491
rect 21121 56457 21140 56491
rect 21068 56436 21140 56457
rect 21194 56491 21266 56512
rect 21194 56457 21213 56491
rect 21247 56457 21266 56491
rect 21194 56436 21266 56457
rect 21314 56491 21386 56512
rect 21314 56457 21333 56491
rect 21367 56457 21386 56491
rect 21314 56436 21386 56457
rect 503 55476 575 55497
rect 503 55442 522 55476
rect 556 55442 575 55476
rect 503 55421 575 55442
rect 629 55476 701 55497
rect 629 55442 648 55476
rect 682 55442 701 55476
rect 629 55421 701 55442
rect 749 55476 821 55497
rect 749 55442 768 55476
rect 802 55442 821 55476
rect 749 55421 821 55442
rect 21068 55426 21140 55447
rect 21068 55392 21087 55426
rect 21121 55392 21140 55426
rect 503 55358 575 55379
rect 503 55324 522 55358
rect 556 55324 575 55358
rect 503 55303 575 55324
rect 629 55358 701 55379
rect 629 55324 648 55358
rect 682 55324 701 55358
rect 629 55303 701 55324
rect 749 55358 821 55379
rect 21068 55371 21140 55392
rect 21194 55426 21266 55447
rect 21194 55392 21213 55426
rect 21247 55392 21266 55426
rect 21194 55371 21266 55392
rect 21314 55426 21386 55447
rect 21314 55392 21333 55426
rect 21367 55392 21386 55426
rect 21314 55371 21386 55392
rect 749 55324 768 55358
rect 802 55324 821 55358
rect 749 55303 821 55324
rect 21068 55308 21140 55329
rect 21068 55274 21087 55308
rect 21121 55274 21140 55308
rect 21068 55253 21140 55274
rect 21194 55308 21266 55329
rect 21194 55274 21213 55308
rect 21247 55274 21266 55308
rect 21194 55253 21266 55274
rect 21314 55308 21386 55329
rect 21314 55274 21333 55308
rect 21367 55274 21386 55308
rect 21314 55253 21386 55274
rect 463 55039 946 55109
rect 463 55005 523 55039
rect 557 55005 645 55039
rect 679 55005 771 55039
rect 805 55005 946 55039
rect 463 54892 946 55005
rect 463 54858 523 54892
rect 557 54858 645 54892
rect 679 54858 771 54892
rect 805 54858 946 54892
rect 463 54755 946 54858
rect 463 54721 523 54755
rect 557 54721 645 54755
rect 679 54721 771 54755
rect 805 54721 946 54755
rect 463 54650 946 54721
rect 22010 54058 22082 54079
rect 22010 54024 22029 54058
rect 22063 54024 22082 54058
rect 22010 54003 22082 54024
rect 22136 54058 22208 54079
rect 22136 54024 22155 54058
rect 22189 54024 22208 54058
rect 22136 54003 22208 54024
rect 22256 54058 22328 54079
rect 22256 54024 22275 54058
rect 22309 54024 22328 54058
rect 22256 54003 22328 54024
rect 22010 53940 22082 53961
rect 22010 53906 22029 53940
rect 22063 53906 22082 53940
rect 22010 53885 22082 53906
rect 22136 53940 22208 53961
rect 22136 53906 22155 53940
rect 22189 53906 22208 53940
rect 22136 53885 22208 53906
rect 22256 53940 22328 53961
rect 22256 53906 22275 53940
rect 22309 53906 22328 53940
rect 22256 53885 22328 53906
rect 463 53280 946 53350
rect 463 53246 523 53280
rect 557 53246 645 53280
rect 679 53246 771 53280
rect 805 53246 946 53280
rect 463 53133 946 53246
rect 463 53099 523 53133
rect 557 53099 645 53133
rect 679 53099 771 53133
rect 805 53099 946 53133
rect 463 52996 946 53099
rect 463 52962 523 52996
rect 557 52962 645 52996
rect 679 52962 771 52996
rect 805 52962 946 52996
rect 463 52891 946 52962
rect 503 52710 575 52731
rect 503 52676 522 52710
rect 556 52676 575 52710
rect 503 52655 575 52676
rect 629 52710 701 52731
rect 629 52676 648 52710
rect 682 52676 701 52710
rect 629 52655 701 52676
rect 749 52710 821 52731
rect 749 52676 768 52710
rect 802 52676 821 52710
rect 749 52655 821 52676
rect 503 52592 575 52613
rect 503 52558 522 52592
rect 556 52558 575 52592
rect 503 52537 575 52558
rect 629 52592 701 52613
rect 629 52558 648 52592
rect 682 52558 701 52592
rect 629 52537 701 52558
rect 749 52592 821 52613
rect 749 52558 768 52592
rect 802 52558 821 52592
rect 749 52537 821 52558
rect 21068 52554 21140 52575
rect 21068 52520 21087 52554
rect 21121 52520 21140 52554
rect 21068 52499 21140 52520
rect 21194 52554 21266 52575
rect 21194 52520 21213 52554
rect 21247 52520 21266 52554
rect 21194 52499 21266 52520
rect 21314 52554 21386 52575
rect 21314 52520 21333 52554
rect 21367 52520 21386 52554
rect 21314 52499 21386 52520
rect 21068 52436 21140 52457
rect 21068 52402 21087 52436
rect 21121 52402 21140 52436
rect 21068 52381 21140 52402
rect 21194 52436 21266 52457
rect 21194 52402 21213 52436
rect 21247 52402 21266 52436
rect 21194 52381 21266 52402
rect 21314 52436 21386 52457
rect 21314 52402 21333 52436
rect 21367 52402 21386 52436
rect 21314 52381 21386 52402
rect 503 51523 575 51544
rect 503 51489 522 51523
rect 556 51489 575 51523
rect 503 51468 575 51489
rect 629 51523 701 51544
rect 629 51489 648 51523
rect 682 51489 701 51523
rect 629 51468 701 51489
rect 749 51523 821 51544
rect 749 51489 768 51523
rect 802 51489 821 51523
rect 749 51468 821 51489
rect 503 51405 575 51426
rect 503 51371 522 51405
rect 556 51371 575 51405
rect 503 51350 575 51371
rect 629 51405 701 51426
rect 629 51371 648 51405
rect 682 51371 701 51405
rect 629 51350 701 51371
rect 749 51405 821 51426
rect 749 51371 768 51405
rect 802 51371 821 51405
rect 749 51350 821 51371
rect 21068 51419 21140 51440
rect 21068 51385 21087 51419
rect 21121 51385 21140 51419
rect 21068 51364 21140 51385
rect 21194 51419 21266 51440
rect 21194 51385 21213 51419
rect 21247 51385 21266 51419
rect 21194 51364 21266 51385
rect 21314 51419 21386 51440
rect 21314 51385 21333 51419
rect 21367 51385 21386 51419
rect 21314 51364 21386 51385
rect 21068 51301 21140 51322
rect 21068 51267 21087 51301
rect 21121 51267 21140 51301
rect 21068 51246 21140 51267
rect 21194 51301 21266 51322
rect 21194 51267 21213 51301
rect 21247 51267 21266 51301
rect 21194 51246 21266 51267
rect 21314 51301 21386 51322
rect 21314 51267 21333 51301
rect 21367 51267 21386 51301
rect 21314 51246 21386 51267
rect 463 51039 946 51109
rect 463 51005 523 51039
rect 557 51005 645 51039
rect 679 51005 771 51039
rect 805 51005 946 51039
rect 463 50892 946 51005
rect 463 50858 523 50892
rect 557 50858 645 50892
rect 679 50858 771 50892
rect 805 50858 946 50892
rect 463 50755 946 50858
rect 463 50721 523 50755
rect 557 50721 645 50755
rect 679 50721 771 50755
rect 805 50721 946 50755
rect 463 50650 946 50721
rect 22010 50137 22082 50158
rect 22010 50103 22029 50137
rect 22063 50103 22082 50137
rect 22010 50082 22082 50103
rect 22136 50137 22208 50158
rect 22136 50103 22155 50137
rect 22189 50103 22208 50137
rect 22136 50082 22208 50103
rect 22256 50137 22328 50158
rect 22256 50103 22275 50137
rect 22309 50103 22328 50137
rect 22256 50082 22328 50103
rect 22010 50019 22082 50040
rect 22010 49985 22029 50019
rect 22063 49985 22082 50019
rect 22010 49964 22082 49985
rect 22136 50019 22208 50040
rect 22136 49985 22155 50019
rect 22189 49985 22208 50019
rect 22136 49964 22208 49985
rect 22256 50019 22328 50040
rect 22256 49985 22275 50019
rect 22309 49985 22328 50019
rect 22256 49964 22328 49985
rect 463 49280 946 49350
rect 463 49246 523 49280
rect 557 49246 645 49280
rect 679 49246 771 49280
rect 805 49246 946 49280
rect 463 49133 946 49246
rect 463 49099 523 49133
rect 557 49099 645 49133
rect 679 49099 771 49133
rect 805 49099 946 49133
rect 463 48996 946 49099
rect 463 48962 523 48996
rect 557 48962 645 48996
rect 679 48962 771 48996
rect 805 48962 946 48996
rect 463 48891 946 48962
rect 503 48701 575 48722
rect 503 48667 522 48701
rect 556 48667 575 48701
rect 503 48646 575 48667
rect 629 48701 701 48722
rect 629 48667 648 48701
rect 682 48667 701 48701
rect 629 48646 701 48667
rect 749 48701 821 48722
rect 749 48667 768 48701
rect 802 48667 821 48701
rect 749 48646 821 48667
rect 21068 48660 21140 48681
rect 21068 48626 21087 48660
rect 21121 48626 21140 48660
rect 21068 48605 21140 48626
rect 21194 48660 21266 48681
rect 21194 48626 21213 48660
rect 21247 48626 21266 48660
rect 21194 48605 21266 48626
rect 21314 48660 21386 48681
rect 21314 48626 21333 48660
rect 21367 48626 21386 48660
rect 21314 48605 21386 48626
rect 503 48583 575 48604
rect 503 48549 522 48583
rect 556 48549 575 48583
rect 503 48528 575 48549
rect 629 48583 701 48604
rect 629 48549 648 48583
rect 682 48549 701 48583
rect 629 48528 701 48549
rect 749 48583 821 48604
rect 749 48549 768 48583
rect 802 48549 821 48583
rect 749 48528 821 48549
rect 21068 48542 21140 48563
rect 21068 48508 21087 48542
rect 21121 48508 21140 48542
rect 21068 48487 21140 48508
rect 21194 48542 21266 48563
rect 21194 48508 21213 48542
rect 21247 48508 21266 48542
rect 21194 48487 21266 48508
rect 21314 48542 21386 48563
rect 21314 48508 21333 48542
rect 21367 48508 21386 48542
rect 21314 48487 21386 48508
rect 503 47548 575 47569
rect 503 47514 522 47548
rect 556 47514 575 47548
rect 503 47493 575 47514
rect 629 47548 701 47569
rect 629 47514 648 47548
rect 682 47514 701 47548
rect 629 47493 701 47514
rect 749 47548 821 47569
rect 749 47514 768 47548
rect 802 47514 821 47548
rect 749 47493 821 47514
rect 21068 47507 21140 47528
rect 21068 47473 21087 47507
rect 21121 47473 21140 47507
rect 21068 47452 21140 47473
rect 21194 47507 21266 47528
rect 21194 47473 21213 47507
rect 21247 47473 21266 47507
rect 21194 47452 21266 47473
rect 21314 47507 21386 47528
rect 21314 47473 21333 47507
rect 21367 47473 21386 47507
rect 21314 47452 21386 47473
rect 503 47430 575 47451
rect 503 47396 522 47430
rect 556 47396 575 47430
rect 503 47375 575 47396
rect 629 47430 701 47451
rect 629 47396 648 47430
rect 682 47396 701 47430
rect 629 47375 701 47396
rect 749 47430 821 47451
rect 749 47396 768 47430
rect 802 47396 821 47430
rect 749 47375 821 47396
rect 21068 47389 21140 47410
rect 21068 47355 21087 47389
rect 21121 47355 21140 47389
rect 21068 47334 21140 47355
rect 21194 47389 21266 47410
rect 21194 47355 21213 47389
rect 21247 47355 21266 47389
rect 21194 47334 21266 47355
rect 21314 47389 21386 47410
rect 21314 47355 21333 47389
rect 21367 47355 21386 47389
rect 21314 47334 21386 47355
rect 463 47039 946 47109
rect 463 47005 523 47039
rect 557 47005 645 47039
rect 679 47005 771 47039
rect 805 47005 946 47039
rect 463 46892 946 47005
rect 463 46858 523 46892
rect 557 46858 645 46892
rect 679 46858 771 46892
rect 805 46858 946 46892
rect 463 46755 946 46858
rect 463 46721 523 46755
rect 557 46721 645 46755
rect 679 46721 771 46755
rect 805 46721 946 46755
rect 463 46650 946 46721
rect 22010 45879 22082 45900
rect 22010 45845 22029 45879
rect 22063 45845 22082 45879
rect 22010 45824 22082 45845
rect 22136 45879 22208 45900
rect 22136 45845 22155 45879
rect 22189 45845 22208 45879
rect 22136 45824 22208 45845
rect 22256 45879 22328 45900
rect 22256 45845 22275 45879
rect 22309 45845 22328 45879
rect 22256 45824 22328 45845
rect 22010 45761 22082 45782
rect 22010 45727 22029 45761
rect 22063 45727 22082 45761
rect 22010 45706 22082 45727
rect 22136 45761 22208 45782
rect 22136 45727 22155 45761
rect 22189 45727 22208 45761
rect 22136 45706 22208 45727
rect 22256 45761 22328 45782
rect 22256 45727 22275 45761
rect 22309 45727 22328 45761
rect 22256 45706 22328 45727
rect 463 45279 946 45350
rect 463 45245 523 45279
rect 557 45245 645 45279
rect 679 45245 771 45279
rect 805 45245 946 45279
rect 463 45132 946 45245
rect 463 45098 523 45132
rect 557 45098 645 45132
rect 679 45098 771 45132
rect 805 45098 946 45132
rect 463 44995 946 45098
rect 463 44961 523 44995
rect 557 44961 645 44995
rect 679 44961 771 44995
rect 805 44961 946 44995
rect 463 44891 946 44961
rect 463 44890 836 44891
rect 503 44488 575 44509
rect 503 44454 522 44488
rect 556 44454 575 44488
rect 503 44433 575 44454
rect 629 44488 701 44509
rect 629 44454 648 44488
rect 682 44454 701 44488
rect 629 44433 701 44454
rect 749 44488 821 44509
rect 749 44454 768 44488
rect 802 44454 821 44488
rect 749 44433 821 44454
rect 21068 44391 21140 44412
rect 503 44370 575 44391
rect 503 44336 522 44370
rect 556 44336 575 44370
rect 503 44315 575 44336
rect 629 44370 701 44391
rect 629 44336 648 44370
rect 682 44336 701 44370
rect 629 44315 701 44336
rect 749 44370 821 44391
rect 749 44336 768 44370
rect 802 44336 821 44370
rect 21068 44357 21087 44391
rect 21121 44357 21140 44391
rect 21068 44336 21140 44357
rect 21194 44391 21266 44412
rect 21194 44357 21213 44391
rect 21247 44357 21266 44391
rect 21194 44336 21266 44357
rect 21314 44391 21386 44412
rect 21314 44357 21333 44391
rect 21367 44357 21386 44391
rect 21314 44336 21386 44357
rect 749 44315 821 44336
rect 21068 44273 21140 44294
rect 21068 44239 21087 44273
rect 21121 44239 21140 44273
rect 21068 44218 21140 44239
rect 21194 44273 21266 44294
rect 21194 44239 21213 44273
rect 21247 44239 21266 44273
rect 21194 44218 21266 44239
rect 21314 44273 21386 44294
rect 21314 44239 21333 44273
rect 21367 44239 21386 44273
rect 21314 44218 21386 44239
rect 924 39650 5204 39727
rect 924 39548 1335 39650
rect 1437 39548 1735 39650
rect 1837 39548 2135 39650
rect 2237 39548 2535 39650
rect 2637 39548 2935 39650
rect 3037 39548 3335 39650
rect 3437 39548 3735 39650
rect 3837 39548 4135 39650
rect 4237 39548 4535 39650
rect 4637 39548 5204 39650
rect 924 39476 5204 39548
rect 924 39467 1188 39476
rect 924 39365 1009 39467
rect 1111 39365 1188 39467
rect 4914 39467 5204 39476
rect 924 39117 1188 39365
rect 1868 39391 2503 39410
rect 1650 39317 1796 39329
rect 1650 39283 1666 39317
rect 1700 39283 1746 39317
rect 1780 39283 1796 39317
rect 1650 39237 1796 39283
rect 1868 39285 1891 39391
rect 1997 39285 2047 39391
rect 2153 39285 2203 39391
rect 2309 39285 2503 39391
rect 4914 39365 5012 39467
rect 5114 39365 5204 39467
rect 1868 39271 2503 39285
rect 1868 39270 2009 39271
rect 1650 39203 1666 39237
rect 1700 39203 1746 39237
rect 1780 39223 1796 39237
rect 2192 39227 2227 39237
rect 1780 39203 2192 39223
rect 1650 39193 2192 39203
rect 2226 39193 2227 39227
rect 1650 39189 2227 39193
rect 924 39116 1114 39117
rect 924 39082 960 39116
rect 994 39083 1114 39116
rect 1148 39083 1188 39117
rect 994 39082 1188 39083
rect 924 39067 1188 39082
rect 924 39000 1009 39067
rect 924 38966 963 39000
rect 997 38966 1009 39000
rect 924 38965 1009 38966
rect 1111 39003 1188 39067
rect 1604 39109 1638 39139
rect 1919 39113 1954 39139
rect 1604 39052 1638 39075
rect 1111 38969 1114 39003
rect 1148 38969 1188 39003
rect 1762 38999 1796 39090
rect 1919 39079 1920 39113
rect 1919 39069 1954 39079
rect 2192 39078 2227 39189
rect 2351 39085 2503 39271
rect 2539 39324 2685 39336
rect 2539 39290 2555 39324
rect 2589 39290 2635 39324
rect 2669 39290 2685 39324
rect 2539 39244 2685 39290
rect 2539 39210 2555 39244
rect 2589 39210 2635 39244
rect 2669 39210 2685 39244
rect 2539 39196 2685 39210
rect 2638 39085 2672 39196
rect 4914 39108 5204 39365
rect 1919 39058 1953 39069
rect 1111 38965 1188 38969
rect 924 38667 1188 38965
rect 1604 38933 1638 38989
rect 1604 38797 1638 38899
rect 1762 38798 1796 38977
rect 1920 38933 1954 38989
rect 1920 38797 1954 38899
rect 2035 38933 2069 38997
rect 2035 38796 2069 38899
rect 2193 38795 2227 38988
rect 2351 38977 2514 39085
rect 2793 38977 2831 39085
rect 4721 39074 5204 39108
rect 4914 39067 5204 39074
rect 2351 38933 2385 38977
rect 2351 38796 2385 38899
rect 2479 38936 2514 38977
rect 2513 38902 2514 38936
rect 2479 38851 2514 38902
rect 2480 38797 2514 38851
rect 2638 38797 2672 38977
rect 2796 38936 2831 38977
rect 2885 38981 2951 38982
rect 2885 38947 2901 38981
rect 2935 38947 2951 38981
rect 4914 38965 5012 39067
rect 5114 38965 5204 39067
rect 2885 38946 2951 38947
rect 2796 38902 2797 38936
rect 2796 38851 2831 38902
rect 4315 38870 4557 38876
rect 2796 38797 2830 38851
rect 2900 38836 2921 38870
rect 2955 38836 2973 38870
rect 3287 38836 3288 38870
rect 4315 38836 4339 38870
rect 4373 38836 4557 38870
rect 4315 38828 4557 38836
rect 4591 38870 4663 38876
rect 4591 38836 4615 38870
rect 4649 38836 4663 38870
rect 4591 38829 4663 38836
rect 4591 38828 4638 38829
rect 1762 38761 1796 38782
rect 3834 38779 3835 38813
rect 1762 38706 1796 38727
rect 924 38565 1009 38667
rect 1111 38565 1188 38667
rect 924 38267 1188 38565
rect 4914 38667 5204 38965
rect 4914 38565 5012 38667
rect 5114 38565 5204 38667
rect 924 38165 1009 38267
rect 1111 38165 1188 38267
rect 1339 38259 1523 38269
rect 1339 38225 1480 38259
rect 1514 38225 1523 38259
rect 1339 38217 1523 38225
rect 2818 38202 2942 38343
rect 3740 38202 3864 38343
rect 4914 38267 5204 38565
rect 4632 38258 4704 38262
rect 4632 38224 4662 38258
rect 4696 38224 4704 38258
rect 4632 38207 4704 38224
rect 924 37867 1188 38165
rect 4914 38165 5012 38267
rect 5114 38165 5204 38267
rect 4914 38020 5204 38165
rect 4812 37986 5204 38020
rect 924 37765 1009 37867
rect 1111 37765 1188 37867
rect 4914 37867 5204 37986
rect 924 37467 1188 37765
rect 1573 37745 1769 37788
rect 2818 37663 2942 37804
rect 3740 37663 3864 37804
rect 4696 37748 4704 37780
rect 4675 37745 4704 37748
rect 4914 37765 5012 37867
rect 5114 37765 5204 37867
rect 924 37365 1009 37467
rect 1111 37365 1188 37467
rect 4914 37467 5204 37765
rect 1963 37442 1997 37465
rect 924 37067 1188 37365
rect 1680 37351 1739 37375
rect 1680 37317 1692 37351
rect 1726 37317 1739 37351
rect 1680 37239 1739 37317
rect 2114 37312 2149 37451
rect 4914 37365 5012 37467
rect 5114 37365 5204 37467
rect 1680 37205 1692 37239
rect 1726 37205 1739 37239
rect 1680 37187 1739 37205
rect 924 37052 1009 37067
rect 1111 37052 1188 37067
rect 924 37018 977 37052
rect 1139 37018 1188 37052
rect 1957 37134 1991 37257
rect 1957 37029 1991 37100
rect 2115 37029 2149 37256
rect 2273 37133 2307 37257
rect 2273 37029 2307 37099
rect 2436 37137 2471 37255
rect 2470 37103 2471 37137
rect 2436 37029 2471 37103
rect 2595 37029 2629 37258
rect 2753 37134 2787 37267
rect 2884 37138 2902 37172
rect 2936 37138 2952 37172
rect 4315 37170 4557 37178
rect 4315 37136 4523 37170
rect 4315 37130 4557 37136
rect 4591 37170 4661 37178
rect 4591 37136 4615 37170
rect 4649 37136 4661 37170
rect 4591 37131 4661 37136
rect 4591 37130 4657 37131
rect 2753 37029 2787 37100
rect 2913 37037 2956 37058
rect 4914 37067 5204 37365
rect 924 36965 1009 37018
rect 1111 36965 1188 37018
rect 924 36922 1188 36965
rect 924 36888 977 36922
rect 1011 36888 1106 36922
rect 1140 36888 1188 36922
rect 1946 36921 1991 37029
rect 2273 36921 2318 37029
rect 2423 36921 2471 37029
rect 2753 36928 2800 37029
rect 2913 37003 2917 37037
rect 2951 37003 2956 37037
rect 2913 36987 2956 37003
rect 4914 36965 5012 37067
rect 5114 36965 5204 37067
rect 4914 36932 5204 36965
rect 924 36650 1188 36888
rect 2595 36838 2629 36921
rect 2753 36838 2879 36928
rect 4721 36898 5204 36932
rect 2538 36826 2685 36838
rect 2538 36792 2555 36826
rect 2589 36792 2635 36826
rect 2669 36792 2685 36826
rect 2538 36747 2685 36792
rect 2538 36713 2555 36747
rect 2589 36713 2635 36747
rect 2669 36713 2685 36747
rect 2538 36703 2685 36713
rect 2752 36826 2899 36838
rect 2752 36792 2769 36826
rect 2803 36792 2849 36826
rect 2883 36792 2899 36826
rect 2752 36747 2899 36792
rect 2752 36713 2769 36747
rect 2803 36713 2849 36747
rect 2883 36713 2899 36747
rect 2752 36707 2899 36713
rect 4914 36650 5204 36898
rect 924 36585 5204 36650
rect 924 36483 1009 36585
rect 1111 36483 1437 36585
rect 1539 36483 1837 36585
rect 1939 36483 2237 36585
rect 2339 36580 3437 36585
rect 2339 36483 2771 36580
rect 924 36478 2771 36483
rect 2873 36478 3098 36580
rect 3200 36483 3437 36580
rect 3539 36483 3837 36585
rect 3939 36483 4237 36585
rect 4339 36483 4637 36585
rect 4739 36483 5012 36585
rect 5114 36483 5204 36585
rect 3200 36478 5204 36483
rect 924 36449 5204 36478
rect 924 36411 5203 36449
rect 20526 35571 21428 35642
rect 20526 35537 21088 35571
rect 21122 35537 21210 35571
rect 21244 35537 21336 35571
rect 21370 35537 21428 35571
rect 20526 35424 21428 35537
rect 20526 35390 21088 35424
rect 21122 35390 21210 35424
rect 21244 35390 21336 35424
rect 21370 35390 21428 35424
rect 20526 35287 21428 35390
rect 20526 35253 21088 35287
rect 21122 35253 21210 35287
rect 21244 35253 21336 35287
rect 21370 35253 21428 35287
rect 20526 35183 21428 35253
rect 20526 35182 21401 35183
rect 20526 33811 21428 33882
rect 20526 33777 21088 33811
rect 21122 33777 21210 33811
rect 21244 33777 21336 33811
rect 21370 33777 21428 33811
rect 20526 33664 21428 33777
rect 20526 33630 21088 33664
rect 21122 33630 21210 33664
rect 21244 33630 21336 33664
rect 21370 33630 21428 33664
rect 20526 33527 21428 33630
rect 20526 33493 21088 33527
rect 21122 33493 21210 33527
rect 21244 33493 21336 33527
rect 21370 33493 21428 33527
rect 20526 33423 21428 33493
rect 20526 33422 21401 33423
rect 503 32281 575 32302
rect 503 32247 522 32281
rect 556 32247 575 32281
rect 503 32226 575 32247
rect 629 32281 701 32302
rect 629 32247 648 32281
rect 682 32247 701 32281
rect 629 32226 701 32247
rect 749 32281 821 32302
rect 749 32247 768 32281
rect 802 32247 821 32281
rect 749 32226 821 32247
rect 21068 32281 21140 32302
rect 21068 32247 21087 32281
rect 21121 32247 21140 32281
rect 21068 32226 21140 32247
rect 21194 32281 21266 32302
rect 21194 32247 21213 32281
rect 21247 32247 21266 32281
rect 21194 32226 21266 32247
rect 21314 32281 21386 32302
rect 21314 32247 21333 32281
rect 21367 32247 21386 32281
rect 21314 32226 21386 32247
rect 503 32163 575 32184
rect 503 32129 522 32163
rect 556 32129 575 32163
rect 503 32108 575 32129
rect 629 32163 701 32184
rect 629 32129 648 32163
rect 682 32129 701 32163
rect 629 32108 701 32129
rect 749 32163 821 32184
rect 749 32129 768 32163
rect 802 32129 821 32163
rect 749 32108 821 32129
rect 21068 32163 21140 32184
rect 21068 32129 21087 32163
rect 21121 32129 21140 32163
rect 21068 32108 21140 32129
rect 21194 32163 21266 32184
rect 21194 32129 21213 32163
rect 21247 32129 21266 32163
rect 21194 32108 21266 32129
rect 21314 32163 21386 32184
rect 21314 32129 21333 32163
rect 21367 32129 21386 32163
rect 21314 32108 21386 32129
rect 503 31499 575 31520
rect 503 31465 522 31499
rect 556 31465 575 31499
rect 503 31444 575 31465
rect 629 31499 701 31520
rect 629 31465 648 31499
rect 682 31465 701 31499
rect 629 31444 701 31465
rect 749 31499 821 31520
rect 749 31465 768 31499
rect 802 31465 821 31499
rect 749 31444 821 31465
rect 21068 31499 21140 31520
rect 21068 31465 21087 31499
rect 21121 31465 21140 31499
rect 21068 31444 21140 31465
rect 21194 31499 21266 31520
rect 21194 31465 21213 31499
rect 21247 31465 21266 31499
rect 21194 31444 21266 31465
rect 21314 31499 21386 31520
rect 21314 31465 21333 31499
rect 21367 31465 21386 31499
rect 21314 31444 21386 31465
rect 503 31381 575 31402
rect 503 31347 522 31381
rect 556 31347 575 31381
rect 503 31326 575 31347
rect 629 31381 701 31402
rect 629 31347 648 31381
rect 682 31347 701 31381
rect 629 31326 701 31347
rect 749 31381 821 31402
rect 749 31347 768 31381
rect 802 31347 821 31381
rect 749 31326 821 31347
rect 21068 31381 21140 31402
rect 21068 31347 21087 31381
rect 21121 31347 21140 31381
rect 21068 31326 21140 31347
rect 21194 31381 21266 31402
rect 21194 31347 21213 31381
rect 21247 31347 21266 31381
rect 21194 31326 21266 31347
rect 21314 31381 21386 31402
rect 21314 31347 21333 31381
rect 21367 31347 21386 31381
rect 21314 31326 21386 31347
rect 485 31110 847 31111
rect 463 31040 1116 31110
rect 463 31006 523 31040
rect 557 31006 645 31040
rect 679 31006 771 31040
rect 805 31006 1116 31040
rect 463 30893 1116 31006
rect 463 30859 523 30893
rect 557 30859 645 30893
rect 679 30859 771 30893
rect 805 30859 1116 30893
rect 463 30756 1116 30859
rect 463 30722 523 30756
rect 557 30722 645 30756
rect 679 30722 771 30756
rect 805 30722 1116 30756
rect 463 30652 1116 30722
rect 463 30651 946 30652
rect 22010 30109 22082 30130
rect 22010 30075 22029 30109
rect 22063 30075 22082 30109
rect 22010 30054 22082 30075
rect 22136 30109 22208 30130
rect 22136 30075 22155 30109
rect 22189 30075 22208 30109
rect 22136 30054 22208 30075
rect 22256 30109 22328 30130
rect 22256 30075 22275 30109
rect 22309 30075 22328 30109
rect 22256 30054 22328 30075
rect 22010 29991 22082 30012
rect 22010 29957 22029 29991
rect 22063 29957 22082 29991
rect 22010 29936 22082 29957
rect 22136 29991 22208 30012
rect 22136 29957 22155 29991
rect 22189 29957 22208 29991
rect 22136 29936 22208 29957
rect 22256 29991 22328 30012
rect 22256 29957 22275 29991
rect 22309 29957 22328 29991
rect 22256 29936 22328 29957
rect 463 29273 1026 29350
rect 463 29239 523 29273
rect 557 29239 645 29273
rect 679 29239 771 29273
rect 805 29239 1026 29273
rect 463 29126 1026 29239
rect 463 29092 523 29126
rect 557 29092 645 29126
rect 679 29092 771 29126
rect 805 29092 1026 29126
rect 463 28989 1026 29092
rect 463 28955 523 28989
rect 557 28955 645 28989
rect 679 28955 771 28989
rect 805 28955 1026 28989
rect 463 28890 1026 28955
rect 503 28587 575 28608
rect 503 28553 522 28587
rect 556 28553 575 28587
rect 503 28532 575 28553
rect 629 28587 701 28608
rect 629 28553 648 28587
rect 682 28553 701 28587
rect 629 28532 701 28553
rect 749 28587 821 28608
rect 749 28553 768 28587
rect 802 28553 821 28587
rect 749 28532 821 28553
rect 21068 28538 21140 28559
rect 21068 28504 21087 28538
rect 21121 28504 21140 28538
rect 503 28469 575 28490
rect 503 28435 522 28469
rect 556 28435 575 28469
rect 503 28414 575 28435
rect 629 28469 701 28490
rect 629 28435 648 28469
rect 682 28435 701 28469
rect 629 28414 701 28435
rect 749 28469 821 28490
rect 21068 28483 21140 28504
rect 21194 28538 21266 28559
rect 21194 28504 21213 28538
rect 21247 28504 21266 28538
rect 21194 28483 21266 28504
rect 21314 28538 21386 28559
rect 21314 28504 21333 28538
rect 21367 28504 21386 28538
rect 21314 28483 21386 28504
rect 749 28435 768 28469
rect 802 28435 821 28469
rect 749 28414 821 28435
rect 21068 28420 21140 28441
rect 21068 28386 21087 28420
rect 21121 28386 21140 28420
rect 21068 28365 21140 28386
rect 21194 28420 21266 28441
rect 21194 28386 21213 28420
rect 21247 28386 21266 28420
rect 21194 28365 21266 28386
rect 21314 28420 21386 28441
rect 21314 28386 21333 28420
rect 21367 28386 21386 28420
rect 21314 28365 21386 28386
rect 503 27583 575 27604
rect 503 27549 522 27583
rect 556 27549 575 27583
rect 503 27528 575 27549
rect 629 27583 701 27604
rect 629 27549 648 27583
rect 682 27549 701 27583
rect 629 27528 701 27549
rect 749 27583 821 27604
rect 749 27549 768 27583
rect 802 27549 821 27583
rect 749 27528 821 27549
rect 503 27465 575 27486
rect 503 27431 522 27465
rect 556 27431 575 27465
rect 503 27410 575 27431
rect 629 27465 701 27486
rect 629 27431 648 27465
rect 682 27431 701 27465
rect 629 27410 701 27431
rect 749 27465 821 27486
rect 749 27431 768 27465
rect 802 27431 821 27465
rect 749 27410 821 27431
rect 21068 27421 21140 27442
rect 21068 27387 21087 27421
rect 21121 27387 21140 27421
rect 21068 27366 21140 27387
rect 21194 27421 21266 27442
rect 21194 27387 21213 27421
rect 21247 27387 21266 27421
rect 21194 27366 21266 27387
rect 21314 27421 21386 27442
rect 21314 27387 21333 27421
rect 21367 27387 21386 27421
rect 21314 27366 21386 27387
rect 21068 27303 21140 27324
rect 21068 27269 21087 27303
rect 21121 27269 21140 27303
rect 21068 27248 21140 27269
rect 21194 27303 21266 27324
rect 21194 27269 21213 27303
rect 21247 27269 21266 27303
rect 21194 27248 21266 27269
rect 21314 27303 21386 27324
rect 21314 27269 21333 27303
rect 21367 27269 21386 27303
rect 21314 27248 21386 27269
rect 463 27039 946 27109
rect 463 27005 523 27039
rect 557 27005 645 27039
rect 679 27005 771 27039
rect 805 27005 946 27039
rect 463 26892 946 27005
rect 463 26858 523 26892
rect 557 26858 645 26892
rect 679 26858 771 26892
rect 805 26858 946 26892
rect 463 26755 946 26858
rect 463 26721 523 26755
rect 557 26721 645 26755
rect 679 26721 771 26755
rect 805 26721 946 26755
rect 463 26650 946 26721
rect 22010 25950 22082 25971
rect 22010 25916 22029 25950
rect 22063 25916 22082 25950
rect 22010 25895 22082 25916
rect 22136 25950 22208 25971
rect 22136 25916 22155 25950
rect 22189 25916 22208 25950
rect 22136 25895 22208 25916
rect 22256 25950 22328 25971
rect 22256 25916 22275 25950
rect 22309 25916 22328 25950
rect 22256 25895 22328 25916
rect 22010 25832 22082 25853
rect 22010 25798 22029 25832
rect 22063 25798 22082 25832
rect 22010 25777 22082 25798
rect 22136 25832 22208 25853
rect 22136 25798 22155 25832
rect 22189 25798 22208 25832
rect 22136 25777 22208 25798
rect 22256 25832 22328 25853
rect 22256 25798 22275 25832
rect 22309 25798 22328 25832
rect 22256 25777 22328 25798
rect 463 25279 946 25349
rect 463 25245 523 25279
rect 557 25245 645 25279
rect 679 25245 771 25279
rect 805 25245 946 25279
rect 463 25132 946 25245
rect 463 25098 523 25132
rect 557 25098 645 25132
rect 679 25098 771 25132
rect 805 25098 946 25132
rect 463 24995 946 25098
rect 463 24961 523 24995
rect 557 24961 645 24995
rect 679 24961 771 24995
rect 805 24961 946 24995
rect 463 24890 946 24961
rect 503 24605 575 24626
rect 503 24571 522 24605
rect 556 24571 575 24605
rect 503 24550 575 24571
rect 629 24605 701 24626
rect 629 24571 648 24605
rect 682 24571 701 24605
rect 629 24550 701 24571
rect 749 24605 821 24626
rect 749 24571 768 24605
rect 802 24571 821 24605
rect 749 24550 821 24571
rect 21068 24578 21140 24599
rect 21068 24544 21087 24578
rect 21121 24544 21140 24578
rect 21068 24523 21140 24544
rect 21194 24578 21266 24599
rect 21194 24544 21213 24578
rect 21247 24544 21266 24578
rect 21194 24523 21266 24544
rect 21314 24578 21386 24599
rect 21314 24544 21333 24578
rect 21367 24544 21386 24578
rect 21314 24523 21386 24544
rect 503 24487 575 24508
rect 503 24453 522 24487
rect 556 24453 575 24487
rect 503 24432 575 24453
rect 629 24487 701 24508
rect 629 24453 648 24487
rect 682 24453 701 24487
rect 629 24432 701 24453
rect 749 24487 821 24508
rect 749 24453 768 24487
rect 802 24453 821 24487
rect 749 24432 821 24453
rect 21068 24460 21140 24481
rect 21068 24426 21087 24460
rect 21121 24426 21140 24460
rect 21068 24405 21140 24426
rect 21194 24460 21266 24481
rect 21194 24426 21213 24460
rect 21247 24426 21266 24460
rect 21194 24405 21266 24426
rect 21314 24460 21386 24481
rect 21314 24426 21333 24460
rect 21367 24426 21386 24460
rect 21314 24405 21386 24426
rect 503 23523 575 23544
rect 503 23489 522 23523
rect 556 23489 575 23523
rect 503 23468 575 23489
rect 629 23523 701 23544
rect 629 23489 648 23523
rect 682 23489 701 23523
rect 629 23468 701 23489
rect 749 23523 821 23544
rect 749 23489 768 23523
rect 802 23489 821 23523
rect 749 23468 821 23489
rect 503 23405 575 23426
rect 503 23371 522 23405
rect 556 23371 575 23405
rect 503 23350 575 23371
rect 629 23405 701 23426
rect 629 23371 648 23405
rect 682 23371 701 23405
rect 629 23350 701 23371
rect 749 23405 821 23426
rect 749 23371 768 23405
rect 802 23371 821 23405
rect 749 23350 821 23371
rect 21068 23403 21140 23424
rect 21068 23369 21087 23403
rect 21121 23369 21140 23403
rect 21068 23348 21140 23369
rect 21194 23403 21266 23424
rect 21194 23369 21213 23403
rect 21247 23369 21266 23403
rect 21194 23348 21266 23369
rect 21314 23403 21386 23424
rect 21314 23369 21333 23403
rect 21367 23369 21386 23403
rect 21314 23348 21386 23369
rect 21068 23285 21140 23306
rect 21068 23251 21087 23285
rect 21121 23251 21140 23285
rect 21068 23230 21140 23251
rect 21194 23285 21266 23306
rect 21194 23251 21213 23285
rect 21247 23251 21266 23285
rect 21194 23230 21266 23251
rect 21314 23285 21386 23306
rect 21314 23251 21333 23285
rect 21367 23251 21386 23285
rect 21314 23230 21386 23251
rect 463 23039 946 23109
rect 463 23005 523 23039
rect 557 23005 645 23039
rect 679 23005 771 23039
rect 805 23005 946 23039
rect 463 22892 946 23005
rect 463 22858 523 22892
rect 557 22858 645 22892
rect 679 22858 771 22892
rect 805 22858 946 22892
rect 463 22755 946 22858
rect 463 22721 523 22755
rect 557 22721 645 22755
rect 679 22721 771 22755
rect 805 22721 946 22755
rect 463 22650 946 22721
rect 22010 22160 22082 22181
rect 22010 22126 22029 22160
rect 22063 22126 22082 22160
rect 22010 22105 22082 22126
rect 22136 22160 22208 22181
rect 22136 22126 22155 22160
rect 22189 22126 22208 22160
rect 22136 22105 22208 22126
rect 22256 22160 22328 22181
rect 22256 22126 22275 22160
rect 22309 22126 22328 22160
rect 22256 22105 22328 22126
rect 22010 22042 22082 22063
rect 22010 22008 22029 22042
rect 22063 22008 22082 22042
rect 22010 21987 22082 22008
rect 22136 22042 22208 22063
rect 22136 22008 22155 22042
rect 22189 22008 22208 22042
rect 22136 21987 22208 22008
rect 22256 22042 22328 22063
rect 22256 22008 22275 22042
rect 22309 22008 22328 22042
rect 22256 21987 22328 22008
rect 463 21280 946 21350
rect 463 21246 523 21280
rect 557 21246 645 21280
rect 679 21246 771 21280
rect 805 21246 946 21280
rect 463 21133 946 21246
rect 463 21099 523 21133
rect 557 21099 645 21133
rect 679 21099 771 21133
rect 805 21099 946 21133
rect 463 20996 946 21099
rect 463 20962 523 20996
rect 557 20962 645 20996
rect 679 20962 771 20996
rect 805 20962 946 20996
rect 463 20891 946 20962
rect 503 20648 575 20669
rect 503 20614 522 20648
rect 556 20614 575 20648
rect 503 20593 575 20614
rect 629 20648 701 20669
rect 629 20614 648 20648
rect 682 20614 701 20648
rect 629 20593 701 20614
rect 749 20648 821 20669
rect 749 20614 768 20648
rect 802 20614 821 20648
rect 749 20593 821 20614
rect 21068 20562 21140 20583
rect 503 20530 575 20551
rect 503 20496 522 20530
rect 556 20496 575 20530
rect 503 20475 575 20496
rect 629 20530 701 20551
rect 629 20496 648 20530
rect 682 20496 701 20530
rect 629 20475 701 20496
rect 749 20530 821 20551
rect 749 20496 768 20530
rect 802 20496 821 20530
rect 21068 20528 21087 20562
rect 21121 20528 21140 20562
rect 21068 20507 21140 20528
rect 21194 20562 21266 20583
rect 21194 20528 21213 20562
rect 21247 20528 21266 20562
rect 21194 20507 21266 20528
rect 21314 20562 21386 20583
rect 21314 20528 21333 20562
rect 21367 20528 21386 20562
rect 21314 20507 21386 20528
rect 749 20475 821 20496
rect 21068 20444 21140 20465
rect 21068 20410 21087 20444
rect 21121 20410 21140 20444
rect 21068 20389 21140 20410
rect 21194 20444 21266 20465
rect 21194 20410 21213 20444
rect 21247 20410 21266 20444
rect 21194 20389 21266 20410
rect 21314 20444 21386 20465
rect 21314 20410 21333 20444
rect 21367 20410 21386 20444
rect 21314 20389 21386 20410
rect 503 19547 575 19568
rect 503 19513 522 19547
rect 556 19513 575 19547
rect 503 19492 575 19513
rect 629 19547 701 19568
rect 629 19513 648 19547
rect 682 19513 701 19547
rect 629 19492 701 19513
rect 749 19547 821 19568
rect 749 19513 768 19547
rect 802 19513 821 19547
rect 749 19492 821 19513
rect 503 19429 575 19450
rect 503 19395 522 19429
rect 556 19395 575 19429
rect 503 19374 575 19395
rect 629 19429 701 19450
rect 629 19395 648 19429
rect 682 19395 701 19429
rect 629 19374 701 19395
rect 749 19429 821 19450
rect 749 19395 768 19429
rect 802 19395 821 19429
rect 749 19374 821 19395
rect 21068 19391 21140 19412
rect 21068 19357 21087 19391
rect 21121 19357 21140 19391
rect 21068 19336 21140 19357
rect 21194 19391 21266 19412
rect 21194 19357 21213 19391
rect 21247 19357 21266 19391
rect 21194 19336 21266 19357
rect 21314 19391 21386 19412
rect 21314 19357 21333 19391
rect 21367 19357 21386 19391
rect 21314 19336 21386 19357
rect 21068 19273 21140 19294
rect 21068 19239 21087 19273
rect 21121 19239 21140 19273
rect 21068 19218 21140 19239
rect 21194 19273 21266 19294
rect 21194 19239 21213 19273
rect 21247 19239 21266 19273
rect 21194 19218 21266 19239
rect 21314 19273 21386 19294
rect 21314 19239 21333 19273
rect 21367 19239 21386 19273
rect 21314 19218 21386 19239
rect 463 19039 946 19109
rect 463 19005 523 19039
rect 557 19005 645 19039
rect 679 19005 771 19039
rect 805 19005 946 19039
rect 463 18892 946 19005
rect 463 18858 523 18892
rect 557 18858 645 18892
rect 679 18858 771 18892
rect 805 18858 946 18892
rect 463 18755 946 18858
rect 463 18721 523 18755
rect 557 18721 645 18755
rect 679 18721 771 18755
rect 805 18721 946 18755
rect 463 18650 946 18721
rect 22010 18053 22082 18074
rect 22010 18019 22029 18053
rect 22063 18019 22082 18053
rect 22010 17998 22082 18019
rect 22136 18053 22208 18074
rect 22136 18019 22155 18053
rect 22189 18019 22208 18053
rect 22136 17998 22208 18019
rect 22256 18053 22328 18074
rect 22256 18019 22275 18053
rect 22309 18019 22328 18053
rect 22256 17998 22328 18019
rect 22010 17935 22082 17956
rect 22010 17901 22029 17935
rect 22063 17901 22082 17935
rect 22010 17880 22082 17901
rect 22136 17935 22208 17956
rect 22136 17901 22155 17935
rect 22189 17901 22208 17935
rect 22136 17880 22208 17901
rect 22256 17935 22328 17956
rect 22256 17901 22275 17935
rect 22309 17901 22328 17935
rect 22256 17880 22328 17901
rect 463 17279 946 17349
rect 463 17245 523 17279
rect 557 17245 645 17279
rect 679 17245 771 17279
rect 805 17245 946 17279
rect 463 17132 946 17245
rect 463 17098 523 17132
rect 557 17098 645 17132
rect 679 17098 771 17132
rect 805 17098 946 17132
rect 463 16995 946 17098
rect 463 16961 523 16995
rect 557 16961 645 16995
rect 679 16961 771 16995
rect 805 16961 946 16995
rect 463 16890 946 16961
rect 503 16681 575 16702
rect 503 16647 522 16681
rect 556 16647 575 16681
rect 503 16626 575 16647
rect 629 16681 701 16702
rect 629 16647 648 16681
rect 682 16647 701 16681
rect 629 16626 701 16647
rect 749 16681 821 16702
rect 749 16647 768 16681
rect 802 16647 821 16681
rect 749 16626 821 16647
rect 21068 16630 21140 16651
rect 21068 16596 21087 16630
rect 21121 16596 21140 16630
rect 503 16563 575 16584
rect 503 16529 522 16563
rect 556 16529 575 16563
rect 503 16508 575 16529
rect 629 16563 701 16584
rect 629 16529 648 16563
rect 682 16529 701 16563
rect 629 16508 701 16529
rect 749 16563 821 16584
rect 21068 16575 21140 16596
rect 21194 16630 21266 16651
rect 21194 16596 21213 16630
rect 21247 16596 21266 16630
rect 21194 16575 21266 16596
rect 21314 16630 21386 16651
rect 21314 16596 21333 16630
rect 21367 16596 21386 16630
rect 21314 16575 21386 16596
rect 749 16529 768 16563
rect 802 16529 821 16563
rect 749 16508 821 16529
rect 21068 16512 21140 16533
rect 21068 16478 21087 16512
rect 21121 16478 21140 16512
rect 21068 16457 21140 16478
rect 21194 16512 21266 16533
rect 21194 16478 21213 16512
rect 21247 16478 21266 16512
rect 21194 16457 21266 16478
rect 21314 16512 21386 16533
rect 21314 16478 21333 16512
rect 21367 16478 21386 16512
rect 21314 16457 21386 16478
rect 503 15465 575 15486
rect 503 15431 522 15465
rect 556 15431 575 15465
rect 503 15410 575 15431
rect 629 15465 701 15486
rect 629 15431 648 15465
rect 682 15431 701 15465
rect 629 15410 701 15431
rect 749 15465 821 15486
rect 749 15431 768 15465
rect 802 15431 821 15465
rect 749 15410 821 15431
rect 21068 15416 21140 15437
rect 21068 15382 21087 15416
rect 21121 15382 21140 15416
rect 503 15347 575 15368
rect 503 15313 522 15347
rect 556 15313 575 15347
rect 503 15292 575 15313
rect 629 15347 701 15368
rect 629 15313 648 15347
rect 682 15313 701 15347
rect 629 15292 701 15313
rect 749 15347 821 15368
rect 21068 15361 21140 15382
rect 21194 15416 21266 15437
rect 21194 15382 21213 15416
rect 21247 15382 21266 15416
rect 21194 15361 21266 15382
rect 21314 15416 21386 15437
rect 21314 15382 21333 15416
rect 21367 15382 21386 15416
rect 21314 15361 21386 15382
rect 749 15313 768 15347
rect 802 15313 821 15347
rect 749 15292 821 15313
rect 21068 15298 21140 15319
rect 21068 15264 21087 15298
rect 21121 15264 21140 15298
rect 21068 15243 21140 15264
rect 21194 15298 21266 15319
rect 21194 15264 21213 15298
rect 21247 15264 21266 15298
rect 21194 15243 21266 15264
rect 21314 15298 21386 15319
rect 21314 15264 21333 15298
rect 21367 15264 21386 15298
rect 21314 15243 21386 15264
rect 463 15039 946 15109
rect 463 15005 523 15039
rect 557 15005 645 15039
rect 679 15005 771 15039
rect 805 15005 946 15039
rect 463 14892 946 15005
rect 463 14858 523 14892
rect 557 14858 645 14892
rect 679 14858 771 14892
rect 805 14858 946 14892
rect 463 14755 946 14858
rect 463 14721 523 14755
rect 557 14721 645 14755
rect 679 14721 771 14755
rect 805 14721 946 14755
rect 463 14650 946 14721
rect 22010 14235 22082 14256
rect 22010 14201 22029 14235
rect 22063 14201 22082 14235
rect 22010 14180 22082 14201
rect 22136 14235 22208 14256
rect 22136 14201 22155 14235
rect 22189 14201 22208 14235
rect 22136 14180 22208 14201
rect 22256 14235 22328 14256
rect 22256 14201 22275 14235
rect 22309 14201 22328 14235
rect 22256 14180 22328 14201
rect 22010 14117 22082 14138
rect 22010 14083 22029 14117
rect 22063 14083 22082 14117
rect 22010 14062 22082 14083
rect 22136 14117 22208 14138
rect 22136 14083 22155 14117
rect 22189 14083 22208 14117
rect 22136 14062 22208 14083
rect 22256 14117 22328 14138
rect 22256 14083 22275 14117
rect 22309 14083 22328 14117
rect 22256 14062 22328 14083
rect 463 13279 946 13349
rect 463 13245 523 13279
rect 557 13245 645 13279
rect 679 13245 771 13279
rect 805 13245 946 13279
rect 463 13132 946 13245
rect 463 13098 523 13132
rect 557 13098 645 13132
rect 679 13098 771 13132
rect 805 13098 946 13132
rect 463 12995 946 13098
rect 463 12961 523 12995
rect 557 12961 645 12995
rect 679 12961 771 12995
rect 805 12961 946 12995
rect 463 12890 946 12961
rect 503 12600 575 12621
rect 503 12566 522 12600
rect 556 12566 575 12600
rect 503 12545 575 12566
rect 629 12600 701 12621
rect 629 12566 648 12600
rect 682 12566 701 12600
rect 629 12545 701 12566
rect 749 12600 821 12621
rect 749 12566 768 12600
rect 802 12566 821 12600
rect 749 12545 821 12566
rect 21068 12573 21140 12594
rect 21068 12539 21087 12573
rect 21121 12539 21140 12573
rect 21068 12518 21140 12539
rect 21194 12573 21266 12594
rect 21194 12539 21213 12573
rect 21247 12539 21266 12573
rect 21194 12518 21266 12539
rect 21314 12573 21386 12594
rect 21314 12539 21333 12573
rect 21367 12539 21386 12573
rect 21314 12518 21386 12539
rect 503 12482 575 12503
rect 503 12448 522 12482
rect 556 12448 575 12482
rect 503 12427 575 12448
rect 629 12482 701 12503
rect 629 12448 648 12482
rect 682 12448 701 12482
rect 629 12427 701 12448
rect 749 12482 821 12503
rect 749 12448 768 12482
rect 802 12448 821 12482
rect 749 12427 821 12448
rect 21068 12455 21140 12476
rect 21068 12421 21087 12455
rect 21121 12421 21140 12455
rect 21068 12400 21140 12421
rect 21194 12455 21266 12476
rect 21194 12421 21213 12455
rect 21247 12421 21266 12455
rect 21194 12400 21266 12421
rect 21314 12455 21386 12476
rect 21314 12421 21333 12455
rect 21367 12421 21386 12455
rect 21314 12400 21386 12421
rect 503 11478 575 11499
rect 503 11444 522 11478
rect 556 11444 575 11478
rect 503 11423 575 11444
rect 629 11478 701 11499
rect 629 11444 648 11478
rect 682 11444 701 11478
rect 629 11423 701 11444
rect 749 11478 821 11499
rect 749 11444 768 11478
rect 802 11444 821 11478
rect 749 11423 821 11444
rect 21068 11416 21140 11437
rect 21068 11382 21087 11416
rect 21121 11382 21140 11416
rect 503 11360 575 11381
rect 503 11326 522 11360
rect 556 11326 575 11360
rect 503 11305 575 11326
rect 629 11360 701 11381
rect 629 11326 648 11360
rect 682 11326 701 11360
rect 629 11305 701 11326
rect 749 11360 821 11381
rect 21068 11361 21140 11382
rect 21194 11416 21266 11437
rect 21194 11382 21213 11416
rect 21247 11382 21266 11416
rect 21194 11361 21266 11382
rect 21314 11416 21386 11437
rect 21314 11382 21333 11416
rect 21367 11382 21386 11416
rect 21314 11361 21386 11382
rect 749 11326 768 11360
rect 802 11326 821 11360
rect 749 11305 821 11326
rect 21068 11298 21140 11319
rect 21068 11264 21087 11298
rect 21121 11264 21140 11298
rect 21068 11243 21140 11264
rect 21194 11298 21266 11319
rect 21194 11264 21213 11298
rect 21247 11264 21266 11298
rect 21194 11243 21266 11264
rect 21314 11298 21386 11319
rect 21314 11264 21333 11298
rect 21367 11264 21386 11298
rect 21314 11243 21386 11264
rect 463 11040 946 11110
rect 463 11006 523 11040
rect 557 11006 645 11040
rect 679 11006 771 11040
rect 805 11006 946 11040
rect 463 10893 946 11006
rect 463 10859 523 10893
rect 557 10859 645 10893
rect 679 10859 771 10893
rect 805 10859 946 10893
rect 463 10756 946 10859
rect 463 10722 523 10756
rect 557 10722 645 10756
rect 679 10722 771 10756
rect 805 10722 946 10756
rect 463 10651 946 10722
rect 22010 10271 22082 10292
rect 22010 10237 22029 10271
rect 22063 10237 22082 10271
rect 22010 10216 22082 10237
rect 22136 10271 22208 10292
rect 22136 10237 22155 10271
rect 22189 10237 22208 10271
rect 22136 10216 22208 10237
rect 22256 10271 22328 10292
rect 22256 10237 22275 10271
rect 22309 10237 22328 10271
rect 22256 10216 22328 10237
rect 22010 10153 22082 10174
rect 22010 10119 22029 10153
rect 22063 10119 22082 10153
rect 22010 10098 22082 10119
rect 22136 10153 22208 10174
rect 22136 10119 22155 10153
rect 22189 10119 22208 10153
rect 22136 10098 22208 10119
rect 22256 10153 22328 10174
rect 22256 10119 22275 10153
rect 22309 10119 22328 10153
rect 22256 10098 22328 10119
rect 463 9278 946 9348
rect 463 9244 523 9278
rect 557 9244 645 9278
rect 679 9244 771 9278
rect 805 9244 946 9278
rect 463 9131 946 9244
rect 463 9097 523 9131
rect 557 9097 645 9131
rect 679 9097 771 9131
rect 805 9097 946 9131
rect 463 8994 946 9097
rect 463 8960 523 8994
rect 557 8960 645 8994
rect 679 8960 771 8994
rect 805 8960 946 8994
rect 463 8889 946 8960
rect 503 8618 575 8639
rect 503 8584 522 8618
rect 556 8584 575 8618
rect 503 8563 575 8584
rect 629 8618 701 8639
rect 629 8584 648 8618
rect 682 8584 701 8618
rect 629 8563 701 8584
rect 749 8618 821 8639
rect 749 8584 768 8618
rect 802 8584 821 8618
rect 749 8563 821 8584
rect 21068 8573 21140 8594
rect 21068 8539 21087 8573
rect 21121 8539 21140 8573
rect 503 8500 575 8521
rect 503 8466 522 8500
rect 556 8466 575 8500
rect 503 8445 575 8466
rect 629 8500 701 8521
rect 629 8466 648 8500
rect 682 8466 701 8500
rect 629 8445 701 8466
rect 749 8500 821 8521
rect 21068 8518 21140 8539
rect 21194 8573 21266 8594
rect 21194 8539 21213 8573
rect 21247 8539 21266 8573
rect 21194 8518 21266 8539
rect 21314 8573 21386 8594
rect 21314 8539 21333 8573
rect 21367 8539 21386 8573
rect 21314 8518 21386 8539
rect 749 8466 768 8500
rect 802 8466 821 8500
rect 749 8445 821 8466
rect 21068 8455 21140 8476
rect 21068 8421 21087 8455
rect 21121 8421 21140 8455
rect 21068 8400 21140 8421
rect 21194 8455 21266 8476
rect 21194 8421 21213 8455
rect 21247 8421 21266 8455
rect 21194 8400 21266 8421
rect 21314 8455 21386 8476
rect 21314 8421 21333 8455
rect 21367 8421 21386 8455
rect 21314 8400 21386 8421
rect 503 7507 575 7528
rect 503 7473 522 7507
rect 556 7473 575 7507
rect 503 7452 575 7473
rect 629 7507 701 7528
rect 629 7473 648 7507
rect 682 7473 701 7507
rect 629 7452 701 7473
rect 749 7507 821 7528
rect 749 7473 768 7507
rect 802 7473 821 7507
rect 749 7452 821 7473
rect 21068 7416 21140 7437
rect 503 7389 575 7410
rect 503 7355 522 7389
rect 556 7355 575 7389
rect 503 7334 575 7355
rect 629 7389 701 7410
rect 629 7355 648 7389
rect 682 7355 701 7389
rect 629 7334 701 7355
rect 749 7389 821 7410
rect 749 7355 768 7389
rect 802 7355 821 7389
rect 21068 7382 21087 7416
rect 21121 7382 21140 7416
rect 21068 7361 21140 7382
rect 21194 7416 21266 7437
rect 21194 7382 21213 7416
rect 21247 7382 21266 7416
rect 21194 7361 21266 7382
rect 21314 7416 21386 7437
rect 21314 7382 21333 7416
rect 21367 7382 21386 7416
rect 21314 7361 21386 7382
rect 749 7334 821 7355
rect 21068 7298 21140 7319
rect 21068 7264 21087 7298
rect 21121 7264 21140 7298
rect 21068 7243 21140 7264
rect 21194 7298 21266 7319
rect 21194 7264 21213 7298
rect 21247 7264 21266 7298
rect 21194 7243 21266 7264
rect 21314 7298 21386 7319
rect 21314 7264 21333 7298
rect 21367 7264 21386 7298
rect 21314 7243 21386 7264
rect 463 7040 946 7110
rect 463 7006 523 7040
rect 557 7006 645 7040
rect 679 7006 771 7040
rect 805 7006 946 7040
rect 463 6893 946 7006
rect 463 6859 523 6893
rect 557 6859 645 6893
rect 679 6859 771 6893
rect 805 6859 946 6893
rect 463 6756 946 6859
rect 463 6722 523 6756
rect 557 6722 645 6756
rect 679 6722 771 6756
rect 805 6722 946 6756
rect 463 6651 946 6722
rect 22010 6259 22082 6280
rect 22010 6225 22029 6259
rect 22063 6225 22082 6259
rect 22010 6204 22082 6225
rect 22136 6259 22208 6280
rect 22136 6225 22155 6259
rect 22189 6225 22208 6259
rect 22136 6204 22208 6225
rect 22256 6259 22328 6280
rect 22256 6225 22275 6259
rect 22309 6225 22328 6259
rect 22256 6204 22328 6225
rect 22010 6141 22082 6162
rect 22010 6107 22029 6141
rect 22063 6107 22082 6141
rect 22010 6086 22082 6107
rect 22136 6141 22208 6162
rect 22136 6107 22155 6141
rect 22189 6107 22208 6141
rect 22136 6086 22208 6107
rect 22256 6141 22328 6162
rect 22256 6107 22275 6141
rect 22309 6107 22328 6141
rect 22256 6086 22328 6107
rect 463 5279 946 5349
rect 463 5245 523 5279
rect 557 5245 645 5279
rect 679 5245 771 5279
rect 805 5245 946 5279
rect 463 5132 946 5245
rect 463 5098 523 5132
rect 557 5098 645 5132
rect 679 5098 771 5132
rect 805 5098 946 5132
rect 463 4995 946 5098
rect 463 4961 523 4995
rect 557 4961 645 4995
rect 679 4961 771 4995
rect 805 4961 946 4995
rect 463 4890 946 4961
rect 503 4684 575 4705
rect 503 4650 522 4684
rect 556 4650 575 4684
rect 503 4629 575 4650
rect 629 4684 701 4705
rect 629 4650 648 4684
rect 682 4650 701 4684
rect 629 4629 701 4650
rect 749 4684 821 4705
rect 749 4650 768 4684
rect 802 4650 821 4684
rect 749 4629 821 4650
rect 503 4566 575 4587
rect 503 4532 522 4566
rect 556 4532 575 4566
rect 503 4511 575 4532
rect 629 4566 701 4587
rect 629 4532 648 4566
rect 682 4532 701 4566
rect 629 4511 701 4532
rect 749 4566 821 4587
rect 749 4532 768 4566
rect 802 4532 821 4566
rect 749 4511 821 4532
rect 21068 4573 21140 4594
rect 21068 4539 21087 4573
rect 21121 4539 21140 4573
rect 21068 4518 21140 4539
rect 21194 4573 21266 4594
rect 21194 4539 21213 4573
rect 21247 4539 21266 4573
rect 21194 4518 21266 4539
rect 21314 4573 21386 4594
rect 21314 4539 21333 4573
rect 21367 4539 21386 4573
rect 21314 4518 21386 4539
rect 21068 4455 21140 4476
rect 21068 4421 21087 4455
rect 21121 4421 21140 4455
rect 21068 4400 21140 4421
rect 21194 4455 21266 4476
rect 21194 4421 21213 4455
rect 21247 4421 21266 4455
rect 21194 4400 21266 4421
rect 21314 4455 21386 4476
rect 21314 4421 21333 4455
rect 21367 4421 21386 4455
rect 21314 4400 21386 4421
rect 503 3507 575 3528
rect 503 3473 522 3507
rect 556 3473 575 3507
rect 503 3452 575 3473
rect 629 3507 701 3528
rect 629 3473 648 3507
rect 682 3473 701 3507
rect 629 3452 701 3473
rect 749 3507 821 3528
rect 749 3473 768 3507
rect 802 3473 821 3507
rect 749 3452 821 3473
rect 21068 3416 21140 3437
rect 503 3389 575 3410
rect 503 3355 522 3389
rect 556 3355 575 3389
rect 503 3334 575 3355
rect 629 3389 701 3410
rect 629 3355 648 3389
rect 682 3355 701 3389
rect 629 3334 701 3355
rect 749 3389 821 3410
rect 749 3355 768 3389
rect 802 3355 821 3389
rect 21068 3382 21087 3416
rect 21121 3382 21140 3416
rect 21068 3361 21140 3382
rect 21194 3416 21266 3437
rect 21194 3382 21213 3416
rect 21247 3382 21266 3416
rect 21194 3361 21266 3382
rect 21314 3416 21386 3437
rect 21314 3382 21333 3416
rect 21367 3382 21386 3416
rect 21314 3361 21386 3382
rect 749 3334 821 3355
rect 21068 3298 21140 3319
rect 21068 3264 21087 3298
rect 21121 3264 21140 3298
rect 21068 3243 21140 3264
rect 21194 3298 21266 3319
rect 21194 3264 21213 3298
rect 21247 3264 21266 3298
rect 21194 3243 21266 3264
rect 21314 3298 21386 3319
rect 21314 3264 21333 3298
rect 21367 3264 21386 3298
rect 21314 3243 21386 3264
rect 463 3040 946 3110
rect 463 3006 523 3040
rect 557 3006 645 3040
rect 679 3006 771 3040
rect 805 3006 946 3040
rect 463 2893 946 3006
rect 463 2859 523 2893
rect 557 2859 645 2893
rect 679 2859 771 2893
rect 805 2859 946 2893
rect 463 2756 946 2859
rect 463 2722 523 2756
rect 557 2722 645 2756
rect 679 2722 771 2756
rect 805 2722 946 2756
rect 463 2651 946 2722
rect 22010 2259 22082 2280
rect 22010 2225 22029 2259
rect 22063 2225 22082 2259
rect 22010 2204 22082 2225
rect 22136 2259 22208 2280
rect 22136 2225 22155 2259
rect 22189 2225 22208 2259
rect 22136 2204 22208 2225
rect 22256 2259 22328 2280
rect 22256 2225 22275 2259
rect 22309 2225 22328 2259
rect 22256 2204 22328 2225
rect 22010 2141 22082 2162
rect 22010 2107 22029 2141
rect 22063 2107 22082 2141
rect 22010 2086 22082 2107
rect 22136 2141 22208 2162
rect 22136 2107 22155 2141
rect 22189 2107 22208 2141
rect 22136 2086 22208 2107
rect 22256 2141 22328 2162
rect 22256 2107 22275 2141
rect 22309 2107 22328 2141
rect 22256 2086 22328 2107
rect 463 1279 946 1349
rect 463 1245 523 1279
rect 557 1245 645 1279
rect 679 1245 771 1279
rect 805 1245 946 1279
rect 463 1132 946 1245
rect 463 1098 523 1132
rect 557 1098 645 1132
rect 679 1098 771 1132
rect 805 1098 946 1132
rect 463 995 946 1098
rect 463 961 523 995
rect 557 961 645 995
rect 679 961 771 995
rect 805 961 946 995
rect 463 890 946 961
rect 503 684 575 705
rect 503 650 522 684
rect 556 650 575 684
rect 503 629 575 650
rect 629 684 701 705
rect 629 650 648 684
rect 682 650 701 684
rect 629 629 701 650
rect 749 684 821 705
rect 749 650 768 684
rect 802 650 821 684
rect 749 629 821 650
rect 503 566 575 587
rect 503 532 522 566
rect 556 532 575 566
rect 503 511 575 532
rect 629 566 701 587
rect 629 532 648 566
rect 682 532 701 566
rect 629 511 701 532
rect 749 566 821 587
rect 749 532 768 566
rect 802 532 821 566
rect 749 511 821 532
rect 21068 573 21140 594
rect 21068 539 21087 573
rect 21121 539 21140 573
rect 21068 518 21140 539
rect 21194 573 21266 594
rect 21194 539 21213 573
rect 21247 539 21266 573
rect 21194 518 21266 539
rect 21314 573 21386 594
rect 21314 539 21333 573
rect 21367 539 21386 573
rect 21314 518 21386 539
rect 21068 455 21140 476
rect 21068 421 21087 455
rect 21121 421 21140 455
rect 21068 400 21140 421
rect 21194 455 21266 476
rect 21194 421 21213 455
rect 21247 421 21266 455
rect 21194 400 21266 421
rect 21314 455 21386 476
rect 21314 421 21333 455
rect 21367 421 21386 455
rect 21314 400 21386 421
<< viali >>
rect 522 75397 556 75431
rect 648 75397 682 75431
rect 768 75397 802 75431
rect 21087 75437 21121 75471
rect 21213 75437 21247 75471
rect 21333 75437 21367 75471
rect 522 75279 556 75313
rect 648 75279 682 75313
rect 768 75279 802 75313
rect 21087 75319 21121 75353
rect 21213 75319 21247 75353
rect 21333 75319 21367 75353
rect 523 75005 557 75039
rect 645 75005 679 75039
rect 771 75005 805 75039
rect 523 74858 557 74892
rect 645 74858 679 74892
rect 771 74858 805 74892
rect 523 74721 557 74755
rect 645 74721 679 74755
rect 771 74721 805 74755
rect 22029 74016 22063 74050
rect 22155 74016 22189 74050
rect 22275 74016 22309 74050
rect 22029 73898 22063 73932
rect 22155 73898 22189 73932
rect 22275 73898 22309 73932
rect 523 73245 557 73279
rect 645 73245 679 73279
rect 771 73245 805 73279
rect 523 73098 557 73132
rect 645 73098 679 73132
rect 771 73098 805 73132
rect 523 72961 557 72995
rect 645 72961 679 72995
rect 771 72961 805 72995
rect 522 72724 556 72758
rect 648 72724 682 72758
rect 768 72724 802 72758
rect 522 72606 556 72640
rect 648 72606 682 72640
rect 768 72606 802 72640
rect 21087 72640 21121 72674
rect 21213 72640 21247 72674
rect 21333 72640 21367 72674
rect 21087 72522 21121 72556
rect 21213 72522 21247 72556
rect 21333 72522 21367 72556
rect 522 71397 556 71431
rect 648 71397 682 71431
rect 768 71397 802 71431
rect 21087 71437 21121 71471
rect 21213 71437 21247 71471
rect 21333 71437 21367 71471
rect 522 71279 556 71313
rect 648 71279 682 71313
rect 768 71279 802 71313
rect 21087 71319 21121 71353
rect 21213 71319 21247 71353
rect 21333 71319 21367 71353
rect 523 71005 557 71039
rect 645 71005 679 71039
rect 771 71005 805 71039
rect 523 70858 557 70892
rect 645 70858 679 70892
rect 771 70858 805 70892
rect 523 70721 557 70755
rect 645 70721 679 70755
rect 771 70721 805 70755
rect 22029 70016 22063 70050
rect 22155 70016 22189 70050
rect 22275 70016 22309 70050
rect 22029 69898 22063 69932
rect 22155 69898 22189 69932
rect 22275 69898 22309 69932
rect 523 69245 557 69279
rect 645 69245 679 69279
rect 771 69245 805 69279
rect 523 69098 557 69132
rect 645 69098 679 69132
rect 771 69098 805 69132
rect 523 68961 557 68995
rect 645 68961 679 68995
rect 771 68961 805 68995
rect 522 68724 556 68758
rect 648 68724 682 68758
rect 768 68724 802 68758
rect 522 68606 556 68640
rect 648 68606 682 68640
rect 768 68606 802 68640
rect 21087 68640 21121 68674
rect 21213 68640 21247 68674
rect 21333 68640 21367 68674
rect 21087 68522 21121 68556
rect 21213 68522 21247 68556
rect 21333 68522 21367 68556
rect 522 67395 556 67429
rect 648 67395 682 67429
rect 768 67395 802 67429
rect 21087 67437 21121 67471
rect 21213 67437 21247 67471
rect 21333 67437 21367 67471
rect 522 67277 556 67311
rect 648 67277 682 67311
rect 768 67277 802 67311
rect 21087 67319 21121 67353
rect 21213 67319 21247 67353
rect 21333 67319 21367 67353
rect 523 67005 557 67039
rect 645 67005 679 67039
rect 771 67005 805 67039
rect 523 66858 557 66892
rect 645 66858 679 66892
rect 771 66858 805 66892
rect 523 66721 557 66755
rect 645 66721 679 66755
rect 771 66721 805 66755
rect 22029 66003 22063 66037
rect 22155 66003 22189 66037
rect 22275 66003 22309 66037
rect 22029 65885 22063 65919
rect 22155 65885 22189 65919
rect 22275 65885 22309 65919
rect 523 65246 557 65280
rect 645 65246 679 65280
rect 771 65246 805 65280
rect 523 65099 557 65133
rect 645 65099 679 65133
rect 771 65099 805 65133
rect 523 64962 557 64996
rect 645 64962 679 64996
rect 771 64962 805 64996
rect 522 64655 556 64689
rect 648 64655 682 64689
rect 768 64655 802 64689
rect 21087 64640 21121 64674
rect 21213 64640 21247 64674
rect 21333 64640 21367 64674
rect 522 64537 556 64571
rect 648 64537 682 64571
rect 768 64537 802 64571
rect 21087 64522 21121 64556
rect 21213 64522 21247 64556
rect 21333 64522 21367 64556
rect 522 63477 556 63511
rect 648 63477 682 63511
rect 768 63477 802 63511
rect 21087 63437 21121 63471
rect 21213 63437 21247 63471
rect 21333 63437 21367 63471
rect 522 63359 556 63393
rect 648 63359 682 63393
rect 768 63359 802 63393
rect 21087 63319 21121 63353
rect 21213 63319 21247 63353
rect 21333 63319 21367 63353
rect 523 63005 557 63039
rect 645 63005 679 63039
rect 771 63005 805 63039
rect 523 62858 557 62892
rect 645 62858 679 62892
rect 771 62858 805 62892
rect 523 62721 557 62755
rect 645 62721 679 62755
rect 771 62721 805 62755
rect 22029 62002 22063 62036
rect 22155 62002 22189 62036
rect 22275 62002 22309 62036
rect 22029 61884 22063 61918
rect 22155 61884 22189 61918
rect 22275 61884 22309 61918
rect 523 61246 557 61280
rect 645 61246 679 61280
rect 771 61246 805 61280
rect 523 61099 557 61133
rect 645 61099 679 61133
rect 771 61099 805 61133
rect 523 60962 557 60996
rect 645 60962 679 60996
rect 771 60962 805 60996
rect 522 60629 556 60663
rect 648 60629 682 60663
rect 768 60629 802 60663
rect 21087 60640 21121 60674
rect 21213 60640 21247 60674
rect 21333 60640 21367 60674
rect 522 60511 556 60545
rect 648 60511 682 60545
rect 768 60511 802 60545
rect 21087 60522 21121 60556
rect 21213 60522 21247 60556
rect 21333 60522 21367 60556
rect 21087 59491 21121 59525
rect 522 59426 556 59460
rect 648 59426 682 59460
rect 21213 59491 21247 59525
rect 21333 59491 21367 59525
rect 768 59426 802 59460
rect 21087 59373 21121 59407
rect 522 59308 556 59342
rect 648 59308 682 59342
rect 21213 59373 21247 59407
rect 21333 59373 21367 59407
rect 768 59308 802 59342
rect 523 59005 557 59039
rect 645 59005 679 59039
rect 771 59005 805 59039
rect 523 58858 557 58892
rect 645 58858 679 58892
rect 771 58858 805 58892
rect 523 58721 557 58755
rect 645 58721 679 58755
rect 771 58721 805 58755
rect 22029 58041 22063 58075
rect 22155 58041 22189 58075
rect 22275 58041 22309 58075
rect 22029 57923 22063 57957
rect 22155 57923 22189 57957
rect 22275 57923 22309 57957
rect 523 57244 557 57278
rect 645 57244 679 57278
rect 771 57244 805 57278
rect 523 57097 557 57131
rect 645 57097 679 57131
rect 771 57097 805 57131
rect 523 56960 557 56994
rect 645 56960 679 56994
rect 771 56960 805 56994
rect 522 56649 556 56683
rect 648 56649 682 56683
rect 768 56649 802 56683
rect 522 56531 556 56565
rect 648 56531 682 56565
rect 768 56531 802 56565
rect 21087 56575 21121 56609
rect 21213 56575 21247 56609
rect 21333 56575 21367 56609
rect 21087 56457 21121 56491
rect 21213 56457 21247 56491
rect 21333 56457 21367 56491
rect 522 55442 556 55476
rect 648 55442 682 55476
rect 768 55442 802 55476
rect 21087 55392 21121 55426
rect 522 55324 556 55358
rect 648 55324 682 55358
rect 21213 55392 21247 55426
rect 21333 55392 21367 55426
rect 768 55324 802 55358
rect 21087 55274 21121 55308
rect 21213 55274 21247 55308
rect 21333 55274 21367 55308
rect 523 55005 557 55039
rect 645 55005 679 55039
rect 771 55005 805 55039
rect 523 54858 557 54892
rect 645 54858 679 54892
rect 771 54858 805 54892
rect 523 54721 557 54755
rect 645 54721 679 54755
rect 771 54721 805 54755
rect 22029 54024 22063 54058
rect 22155 54024 22189 54058
rect 22275 54024 22309 54058
rect 22029 53906 22063 53940
rect 22155 53906 22189 53940
rect 22275 53906 22309 53940
rect 523 53246 557 53280
rect 645 53246 679 53280
rect 771 53246 805 53280
rect 523 53099 557 53133
rect 645 53099 679 53133
rect 771 53099 805 53133
rect 523 52962 557 52996
rect 645 52962 679 52996
rect 771 52962 805 52996
rect 522 52676 556 52710
rect 648 52676 682 52710
rect 768 52676 802 52710
rect 522 52558 556 52592
rect 648 52558 682 52592
rect 768 52558 802 52592
rect 21087 52520 21121 52554
rect 21213 52520 21247 52554
rect 21333 52520 21367 52554
rect 21087 52402 21121 52436
rect 21213 52402 21247 52436
rect 21333 52402 21367 52436
rect 522 51489 556 51523
rect 648 51489 682 51523
rect 768 51489 802 51523
rect 522 51371 556 51405
rect 648 51371 682 51405
rect 768 51371 802 51405
rect 21087 51385 21121 51419
rect 21213 51385 21247 51419
rect 21333 51385 21367 51419
rect 21087 51267 21121 51301
rect 21213 51267 21247 51301
rect 21333 51267 21367 51301
rect 523 51005 557 51039
rect 645 51005 679 51039
rect 771 51005 805 51039
rect 523 50858 557 50892
rect 645 50858 679 50892
rect 771 50858 805 50892
rect 523 50721 557 50755
rect 645 50721 679 50755
rect 771 50721 805 50755
rect 22029 50103 22063 50137
rect 22155 50103 22189 50137
rect 22275 50103 22309 50137
rect 22029 49985 22063 50019
rect 22155 49985 22189 50019
rect 22275 49985 22309 50019
rect 523 49246 557 49280
rect 645 49246 679 49280
rect 771 49246 805 49280
rect 523 49099 557 49133
rect 645 49099 679 49133
rect 771 49099 805 49133
rect 523 48962 557 48996
rect 645 48962 679 48996
rect 771 48962 805 48996
rect 522 48667 556 48701
rect 648 48667 682 48701
rect 768 48667 802 48701
rect 21087 48626 21121 48660
rect 21213 48626 21247 48660
rect 21333 48626 21367 48660
rect 522 48549 556 48583
rect 648 48549 682 48583
rect 768 48549 802 48583
rect 21087 48508 21121 48542
rect 21213 48508 21247 48542
rect 21333 48508 21367 48542
rect 522 47514 556 47548
rect 648 47514 682 47548
rect 768 47514 802 47548
rect 21087 47473 21121 47507
rect 21213 47473 21247 47507
rect 21333 47473 21367 47507
rect 522 47396 556 47430
rect 648 47396 682 47430
rect 768 47396 802 47430
rect 21087 47355 21121 47389
rect 21213 47355 21247 47389
rect 21333 47355 21367 47389
rect 523 47005 557 47039
rect 645 47005 679 47039
rect 771 47005 805 47039
rect 523 46858 557 46892
rect 645 46858 679 46892
rect 771 46858 805 46892
rect 523 46721 557 46755
rect 645 46721 679 46755
rect 771 46721 805 46755
rect 22029 45845 22063 45879
rect 22155 45845 22189 45879
rect 22275 45845 22309 45879
rect 22029 45727 22063 45761
rect 22155 45727 22189 45761
rect 22275 45727 22309 45761
rect 523 45245 557 45279
rect 645 45245 679 45279
rect 771 45245 805 45279
rect 523 45098 557 45132
rect 645 45098 679 45132
rect 771 45098 805 45132
rect 523 44961 557 44995
rect 645 44961 679 44995
rect 771 44961 805 44995
rect 522 44454 556 44488
rect 648 44454 682 44488
rect 768 44454 802 44488
rect 522 44336 556 44370
rect 648 44336 682 44370
rect 768 44336 802 44370
rect 21087 44357 21121 44391
rect 21213 44357 21247 44391
rect 21333 44357 21367 44391
rect 21087 44239 21121 44273
rect 21213 44239 21247 44273
rect 21333 44239 21367 44273
rect 1666 39283 1700 39317
rect 1746 39283 1780 39317
rect 1891 39285 1997 39391
rect 2047 39285 2153 39391
rect 2203 39285 2309 39391
rect 1666 39203 1700 39237
rect 1746 39203 1780 39237
rect 2192 39193 2226 39227
rect 960 39082 994 39116
rect 1114 39083 1148 39117
rect 963 38966 997 39000
rect 1604 39075 1638 39109
rect 1114 38969 1148 39003
rect 1920 39079 1954 39113
rect 2555 39290 2589 39324
rect 2635 39290 2669 39324
rect 2555 39210 2589 39244
rect 2635 39210 2669 39244
rect 1604 38899 1638 38933
rect 1920 38899 1954 38933
rect 2035 38899 2069 38933
rect 2351 38899 2385 38933
rect 2479 38902 2513 38936
rect 2901 38947 2935 38981
rect 2797 38902 2831 38936
rect 4251 38926 4285 38960
rect 2921 38836 2955 38870
rect 3253 38836 3287 38870
rect 3553 38836 3587 38870
rect 4105 38836 4139 38870
rect 4339 38836 4373 38870
rect 4615 38836 4649 38870
rect 3800 38779 3834 38813
rect 1762 38727 1796 38761
rect 1480 38225 1514 38259
rect 1715 38224 1749 38258
rect 1807 38227 1841 38261
rect 1899 38224 1933 38258
rect 2029 38218 2063 38252
rect 4662 38224 4696 38258
rect 1481 37748 1515 37782
rect 1805 37753 1839 37787
rect 1889 37754 1923 37788
rect 1986 37748 2020 37782
rect 4662 37748 4696 37782
rect 1692 37317 1726 37351
rect 1692 37205 1726 37239
rect 977 37018 1009 37052
rect 1009 37018 1011 37052
rect 1105 37018 1111 37052
rect 1111 37018 1139 37052
rect 1957 37100 1991 37134
rect 2273 37099 2307 37133
rect 2436 37103 2470 37137
rect 3807 37193 3841 37227
rect 2902 37138 2936 37172
rect 3237 37137 3271 37171
rect 3553 37136 3587 37170
rect 4105 37136 4139 37170
rect 4523 37136 4557 37170
rect 2753 37100 2787 37134
rect 4615 37136 4649 37170
rect 4251 37046 4285 37080
rect 977 36888 1011 36922
rect 1106 36888 1140 36922
rect 2917 37003 2951 37037
rect 2555 36792 2589 36826
rect 2635 36792 2669 36826
rect 2555 36713 2589 36747
rect 2635 36713 2669 36747
rect 2769 36792 2803 36826
rect 2849 36792 2883 36826
rect 2769 36713 2803 36747
rect 2849 36713 2883 36747
rect 21088 35537 21122 35571
rect 21210 35537 21244 35571
rect 21336 35537 21370 35571
rect 21088 35390 21122 35424
rect 21210 35390 21244 35424
rect 21336 35390 21370 35424
rect 21088 35253 21122 35287
rect 21210 35253 21244 35287
rect 21336 35253 21370 35287
rect 21088 33777 21122 33811
rect 21210 33777 21244 33811
rect 21336 33777 21370 33811
rect 21088 33630 21122 33664
rect 21210 33630 21244 33664
rect 21336 33630 21370 33664
rect 21088 33493 21122 33527
rect 21210 33493 21244 33527
rect 21336 33493 21370 33527
rect 522 32247 556 32281
rect 648 32247 682 32281
rect 768 32247 802 32281
rect 21087 32247 21121 32281
rect 21213 32247 21247 32281
rect 21333 32247 21367 32281
rect 522 32129 556 32163
rect 648 32129 682 32163
rect 768 32129 802 32163
rect 21087 32129 21121 32163
rect 21213 32129 21247 32163
rect 21333 32129 21367 32163
rect 522 31465 556 31499
rect 648 31465 682 31499
rect 768 31465 802 31499
rect 21087 31465 21121 31499
rect 21213 31465 21247 31499
rect 21333 31465 21367 31499
rect 522 31347 556 31381
rect 648 31347 682 31381
rect 768 31347 802 31381
rect 21087 31347 21121 31381
rect 21213 31347 21247 31381
rect 21333 31347 21367 31381
rect 523 31006 557 31040
rect 645 31006 679 31040
rect 771 31006 805 31040
rect 523 30859 557 30893
rect 645 30859 679 30893
rect 771 30859 805 30893
rect 523 30722 557 30756
rect 645 30722 679 30756
rect 771 30722 805 30756
rect 22029 30075 22063 30109
rect 22155 30075 22189 30109
rect 22275 30075 22309 30109
rect 22029 29957 22063 29991
rect 22155 29957 22189 29991
rect 22275 29957 22309 29991
rect 523 29239 557 29273
rect 645 29239 679 29273
rect 771 29239 805 29273
rect 523 29092 557 29126
rect 645 29092 679 29126
rect 771 29092 805 29126
rect 523 28955 557 28989
rect 645 28955 679 28989
rect 771 28955 805 28989
rect 522 28553 556 28587
rect 648 28553 682 28587
rect 768 28553 802 28587
rect 21087 28504 21121 28538
rect 522 28435 556 28469
rect 648 28435 682 28469
rect 21213 28504 21247 28538
rect 21333 28504 21367 28538
rect 768 28435 802 28469
rect 21087 28386 21121 28420
rect 21213 28386 21247 28420
rect 21333 28386 21367 28420
rect 522 27549 556 27583
rect 648 27549 682 27583
rect 768 27549 802 27583
rect 522 27431 556 27465
rect 648 27431 682 27465
rect 768 27431 802 27465
rect 21087 27387 21121 27421
rect 21213 27387 21247 27421
rect 21333 27387 21367 27421
rect 21087 27269 21121 27303
rect 21213 27269 21247 27303
rect 21333 27269 21367 27303
rect 523 27005 557 27039
rect 645 27005 679 27039
rect 771 27005 805 27039
rect 523 26858 557 26892
rect 645 26858 679 26892
rect 771 26858 805 26892
rect 523 26721 557 26755
rect 645 26721 679 26755
rect 771 26721 805 26755
rect 22029 25916 22063 25950
rect 22155 25916 22189 25950
rect 22275 25916 22309 25950
rect 22029 25798 22063 25832
rect 22155 25798 22189 25832
rect 22275 25798 22309 25832
rect 523 25245 557 25279
rect 645 25245 679 25279
rect 771 25245 805 25279
rect 523 25098 557 25132
rect 645 25098 679 25132
rect 771 25098 805 25132
rect 523 24961 557 24995
rect 645 24961 679 24995
rect 771 24961 805 24995
rect 522 24571 556 24605
rect 648 24571 682 24605
rect 768 24571 802 24605
rect 21087 24544 21121 24578
rect 21213 24544 21247 24578
rect 21333 24544 21367 24578
rect 522 24453 556 24487
rect 648 24453 682 24487
rect 768 24453 802 24487
rect 21087 24426 21121 24460
rect 21213 24426 21247 24460
rect 21333 24426 21367 24460
rect 522 23489 556 23523
rect 648 23489 682 23523
rect 768 23489 802 23523
rect 522 23371 556 23405
rect 648 23371 682 23405
rect 768 23371 802 23405
rect 21087 23369 21121 23403
rect 21213 23369 21247 23403
rect 21333 23369 21367 23403
rect 21087 23251 21121 23285
rect 21213 23251 21247 23285
rect 21333 23251 21367 23285
rect 523 23005 557 23039
rect 645 23005 679 23039
rect 771 23005 805 23039
rect 523 22858 557 22892
rect 645 22858 679 22892
rect 771 22858 805 22892
rect 523 22721 557 22755
rect 645 22721 679 22755
rect 771 22721 805 22755
rect 22029 22126 22063 22160
rect 22155 22126 22189 22160
rect 22275 22126 22309 22160
rect 22029 22008 22063 22042
rect 22155 22008 22189 22042
rect 22275 22008 22309 22042
rect 523 21246 557 21280
rect 645 21246 679 21280
rect 771 21246 805 21280
rect 523 21099 557 21133
rect 645 21099 679 21133
rect 771 21099 805 21133
rect 523 20962 557 20996
rect 645 20962 679 20996
rect 771 20962 805 20996
rect 522 20614 556 20648
rect 648 20614 682 20648
rect 768 20614 802 20648
rect 522 20496 556 20530
rect 648 20496 682 20530
rect 768 20496 802 20530
rect 21087 20528 21121 20562
rect 21213 20528 21247 20562
rect 21333 20528 21367 20562
rect 21087 20410 21121 20444
rect 21213 20410 21247 20444
rect 21333 20410 21367 20444
rect 522 19513 556 19547
rect 648 19513 682 19547
rect 768 19513 802 19547
rect 522 19395 556 19429
rect 648 19395 682 19429
rect 768 19395 802 19429
rect 21087 19357 21121 19391
rect 21213 19357 21247 19391
rect 21333 19357 21367 19391
rect 21087 19239 21121 19273
rect 21213 19239 21247 19273
rect 21333 19239 21367 19273
rect 523 19005 557 19039
rect 645 19005 679 19039
rect 771 19005 805 19039
rect 523 18858 557 18892
rect 645 18858 679 18892
rect 771 18858 805 18892
rect 523 18721 557 18755
rect 645 18721 679 18755
rect 771 18721 805 18755
rect 22029 18019 22063 18053
rect 22155 18019 22189 18053
rect 22275 18019 22309 18053
rect 22029 17901 22063 17935
rect 22155 17901 22189 17935
rect 22275 17901 22309 17935
rect 523 17245 557 17279
rect 645 17245 679 17279
rect 771 17245 805 17279
rect 523 17098 557 17132
rect 645 17098 679 17132
rect 771 17098 805 17132
rect 523 16961 557 16995
rect 645 16961 679 16995
rect 771 16961 805 16995
rect 522 16647 556 16681
rect 648 16647 682 16681
rect 768 16647 802 16681
rect 21087 16596 21121 16630
rect 522 16529 556 16563
rect 648 16529 682 16563
rect 21213 16596 21247 16630
rect 21333 16596 21367 16630
rect 768 16529 802 16563
rect 21087 16478 21121 16512
rect 21213 16478 21247 16512
rect 21333 16478 21367 16512
rect 522 15431 556 15465
rect 648 15431 682 15465
rect 768 15431 802 15465
rect 21087 15382 21121 15416
rect 522 15313 556 15347
rect 648 15313 682 15347
rect 21213 15382 21247 15416
rect 21333 15382 21367 15416
rect 768 15313 802 15347
rect 21087 15264 21121 15298
rect 21213 15264 21247 15298
rect 21333 15264 21367 15298
rect 523 15005 557 15039
rect 645 15005 679 15039
rect 771 15005 805 15039
rect 523 14858 557 14892
rect 645 14858 679 14892
rect 771 14858 805 14892
rect 523 14721 557 14755
rect 645 14721 679 14755
rect 771 14721 805 14755
rect 22029 14201 22063 14235
rect 22155 14201 22189 14235
rect 22275 14201 22309 14235
rect 22029 14083 22063 14117
rect 22155 14083 22189 14117
rect 22275 14083 22309 14117
rect 523 13245 557 13279
rect 645 13245 679 13279
rect 771 13245 805 13279
rect 523 13098 557 13132
rect 645 13098 679 13132
rect 771 13098 805 13132
rect 523 12961 557 12995
rect 645 12961 679 12995
rect 771 12961 805 12995
rect 522 12566 556 12600
rect 648 12566 682 12600
rect 768 12566 802 12600
rect 21087 12539 21121 12573
rect 21213 12539 21247 12573
rect 21333 12539 21367 12573
rect 522 12448 556 12482
rect 648 12448 682 12482
rect 768 12448 802 12482
rect 21087 12421 21121 12455
rect 21213 12421 21247 12455
rect 21333 12421 21367 12455
rect 522 11444 556 11478
rect 648 11444 682 11478
rect 768 11444 802 11478
rect 21087 11382 21121 11416
rect 522 11326 556 11360
rect 648 11326 682 11360
rect 21213 11382 21247 11416
rect 21333 11382 21367 11416
rect 768 11326 802 11360
rect 21087 11264 21121 11298
rect 21213 11264 21247 11298
rect 21333 11264 21367 11298
rect 523 11006 557 11040
rect 645 11006 679 11040
rect 771 11006 805 11040
rect 523 10859 557 10893
rect 645 10859 679 10893
rect 771 10859 805 10893
rect 523 10722 557 10756
rect 645 10722 679 10756
rect 771 10722 805 10756
rect 22029 10237 22063 10271
rect 22155 10237 22189 10271
rect 22275 10237 22309 10271
rect 22029 10119 22063 10153
rect 22155 10119 22189 10153
rect 22275 10119 22309 10153
rect 523 9244 557 9278
rect 645 9244 679 9278
rect 771 9244 805 9278
rect 523 9097 557 9131
rect 645 9097 679 9131
rect 771 9097 805 9131
rect 523 8960 557 8994
rect 645 8960 679 8994
rect 771 8960 805 8994
rect 522 8584 556 8618
rect 648 8584 682 8618
rect 768 8584 802 8618
rect 21087 8539 21121 8573
rect 522 8466 556 8500
rect 648 8466 682 8500
rect 21213 8539 21247 8573
rect 21333 8539 21367 8573
rect 768 8466 802 8500
rect 21087 8421 21121 8455
rect 21213 8421 21247 8455
rect 21333 8421 21367 8455
rect 522 7473 556 7507
rect 648 7473 682 7507
rect 768 7473 802 7507
rect 522 7355 556 7389
rect 648 7355 682 7389
rect 768 7355 802 7389
rect 21087 7382 21121 7416
rect 21213 7382 21247 7416
rect 21333 7382 21367 7416
rect 21087 7264 21121 7298
rect 21213 7264 21247 7298
rect 21333 7264 21367 7298
rect 523 7006 557 7040
rect 645 7006 679 7040
rect 771 7006 805 7040
rect 523 6859 557 6893
rect 645 6859 679 6893
rect 771 6859 805 6893
rect 523 6722 557 6756
rect 645 6722 679 6756
rect 771 6722 805 6756
rect 22029 6225 22063 6259
rect 22155 6225 22189 6259
rect 22275 6225 22309 6259
rect 22029 6107 22063 6141
rect 22155 6107 22189 6141
rect 22275 6107 22309 6141
rect 523 5245 557 5279
rect 645 5245 679 5279
rect 771 5245 805 5279
rect 523 5098 557 5132
rect 645 5098 679 5132
rect 771 5098 805 5132
rect 523 4961 557 4995
rect 645 4961 679 4995
rect 771 4961 805 4995
rect 522 4650 556 4684
rect 648 4650 682 4684
rect 768 4650 802 4684
rect 522 4532 556 4566
rect 648 4532 682 4566
rect 768 4532 802 4566
rect 21087 4539 21121 4573
rect 21213 4539 21247 4573
rect 21333 4539 21367 4573
rect 21087 4421 21121 4455
rect 21213 4421 21247 4455
rect 21333 4421 21367 4455
rect 522 3473 556 3507
rect 648 3473 682 3507
rect 768 3473 802 3507
rect 522 3355 556 3389
rect 648 3355 682 3389
rect 768 3355 802 3389
rect 21087 3382 21121 3416
rect 21213 3382 21247 3416
rect 21333 3382 21367 3416
rect 21087 3264 21121 3298
rect 21213 3264 21247 3298
rect 21333 3264 21367 3298
rect 523 3006 557 3040
rect 645 3006 679 3040
rect 771 3006 805 3040
rect 523 2859 557 2893
rect 645 2859 679 2893
rect 771 2859 805 2893
rect 523 2722 557 2756
rect 645 2722 679 2756
rect 771 2722 805 2756
rect 22029 2225 22063 2259
rect 22155 2225 22189 2259
rect 22275 2225 22309 2259
rect 22029 2107 22063 2141
rect 22155 2107 22189 2141
rect 22275 2107 22309 2141
rect 523 1245 557 1279
rect 645 1245 679 1279
rect 771 1245 805 1279
rect 523 1098 557 1132
rect 645 1098 679 1132
rect 771 1098 805 1132
rect 523 961 557 995
rect 645 961 679 995
rect 771 961 805 995
rect 522 650 556 684
rect 648 650 682 684
rect 768 650 802 684
rect 522 532 556 566
rect 648 532 682 566
rect 768 532 802 566
rect 21087 539 21121 573
rect 21213 539 21247 573
rect 21333 539 21367 573
rect 21087 421 21121 455
rect 21213 421 21247 455
rect 21333 421 21367 455
<< metal1 >>
rect 20946 75480 21426 75517
rect 463 75440 946 75477
rect 463 75388 513 75440
rect 565 75388 639 75440
rect 691 75388 759 75440
rect 811 75388 946 75440
rect 463 75322 946 75388
rect 463 75270 513 75322
rect 565 75270 639 75322
rect 691 75270 759 75322
rect 811 75270 946 75322
rect 463 75222 946 75270
rect 20946 75428 21078 75480
rect 21130 75428 21204 75480
rect 21256 75428 21324 75480
rect 21376 75428 21426 75480
rect 20946 75362 21426 75428
rect 20946 75310 21078 75362
rect 21130 75310 21204 75362
rect 21256 75310 21324 75362
rect 21376 75310 21426 75362
rect 20946 75262 21426 75310
rect 463 75048 863 75109
rect 463 74996 514 75048
rect 566 74996 636 75048
rect 688 74996 762 75048
rect 814 74996 863 75048
rect 463 74901 863 74996
rect 463 74849 514 74901
rect 566 74849 636 74901
rect 688 74849 762 74901
rect 814 74849 863 74901
rect 463 74764 863 74849
rect 463 74712 514 74764
rect 566 74712 636 74764
rect 688 74712 762 74764
rect 814 74712 863 74764
rect 463 74650 863 74712
rect 20946 74059 22370 74096
rect 20946 74007 22020 74059
rect 22072 74007 22146 74059
rect 22198 74007 22266 74059
rect 22318 74007 22370 74059
rect 20946 73941 22370 74007
rect 20946 73889 22020 73941
rect 22072 73889 22146 73941
rect 22198 73889 22266 73941
rect 22318 73889 22370 73941
rect 20946 73841 22370 73889
rect 463 73288 863 73349
rect 463 73236 514 73288
rect 566 73236 636 73288
rect 688 73236 762 73288
rect 814 73236 863 73288
rect 463 73141 863 73236
rect 463 73089 514 73141
rect 566 73089 636 73141
rect 688 73089 762 73141
rect 814 73089 863 73141
rect 463 73004 863 73089
rect 463 72952 514 73004
rect 566 72952 636 73004
rect 688 72952 762 73004
rect 814 72952 863 73004
rect 463 72890 863 72952
rect 463 72767 946 72804
rect 463 72715 513 72767
rect 565 72715 639 72767
rect 691 72715 759 72767
rect 811 72715 946 72767
rect 463 72649 946 72715
rect 463 72597 513 72649
rect 565 72597 639 72649
rect 691 72597 759 72649
rect 811 72597 946 72649
rect 463 72549 946 72597
rect 20946 72683 21428 72720
rect 20946 72631 21078 72683
rect 21130 72631 21204 72683
rect 21256 72631 21324 72683
rect 21376 72631 21428 72683
rect 20946 72565 21428 72631
rect 20946 72513 21078 72565
rect 21130 72513 21204 72565
rect 21256 72513 21324 72565
rect 21376 72513 21428 72565
rect 20946 72465 21428 72513
rect 20946 71480 21426 71517
rect 463 71440 947 71477
rect 463 71388 513 71440
rect 565 71388 639 71440
rect 691 71388 759 71440
rect 811 71388 947 71440
rect 463 71322 947 71388
rect 463 71270 513 71322
rect 565 71270 639 71322
rect 691 71270 759 71322
rect 811 71270 947 71322
rect 463 71222 947 71270
rect 20946 71428 21078 71480
rect 21130 71428 21204 71480
rect 21256 71428 21324 71480
rect 21376 71428 21426 71480
rect 20946 71362 21426 71428
rect 20946 71310 21078 71362
rect 21130 71310 21204 71362
rect 21256 71310 21324 71362
rect 21376 71310 21426 71362
rect 20946 71262 21426 71310
rect 463 71048 863 71109
rect 463 70996 514 71048
rect 566 70996 636 71048
rect 688 70996 762 71048
rect 814 70996 863 71048
rect 463 70901 863 70996
rect 463 70849 514 70901
rect 566 70849 636 70901
rect 688 70849 762 70901
rect 814 70849 863 70901
rect 463 70764 863 70849
rect 463 70712 514 70764
rect 566 70712 636 70764
rect 688 70712 762 70764
rect 814 70712 863 70764
rect 463 70650 863 70712
rect 20946 70059 22370 70096
rect 20946 70007 22020 70059
rect 22072 70007 22146 70059
rect 22198 70007 22266 70059
rect 22318 70007 22370 70059
rect 20946 69941 22370 70007
rect 20946 69889 22020 69941
rect 22072 69889 22146 69941
rect 22198 69889 22266 69941
rect 22318 69889 22370 69941
rect 20946 69841 22370 69889
rect 463 69288 863 69349
rect 463 69236 514 69288
rect 566 69236 636 69288
rect 688 69236 762 69288
rect 814 69236 863 69288
rect 463 69141 863 69236
rect 463 69089 514 69141
rect 566 69089 636 69141
rect 688 69089 762 69141
rect 814 69089 863 69141
rect 463 69004 863 69089
rect 463 68952 514 69004
rect 566 68952 636 69004
rect 688 68952 762 69004
rect 814 68952 863 69004
rect 463 68890 863 68952
rect 463 68767 947 68804
rect 463 68715 513 68767
rect 565 68715 639 68767
rect 691 68715 759 68767
rect 811 68715 947 68767
rect 463 68649 947 68715
rect 463 68597 513 68649
rect 565 68597 639 68649
rect 691 68597 759 68649
rect 811 68597 947 68649
rect 463 68549 947 68597
rect 20946 68683 21428 68720
rect 20946 68631 21078 68683
rect 21130 68631 21204 68683
rect 21256 68631 21324 68683
rect 21376 68631 21428 68683
rect 20946 68565 21428 68631
rect 20946 68513 21078 68565
rect 21130 68513 21204 68565
rect 21256 68513 21324 68565
rect 21376 68513 21428 68565
rect 20946 68465 21428 68513
rect 20945 67517 20946 67530
rect 20945 67480 21426 67517
rect 463 67438 947 67475
rect 463 67386 513 67438
rect 565 67386 639 67438
rect 691 67386 759 67438
rect 811 67386 947 67438
rect 463 67320 947 67386
rect 463 67268 513 67320
rect 565 67268 639 67320
rect 691 67268 759 67320
rect 811 67268 947 67320
rect 20945 67428 21078 67480
rect 21130 67428 21204 67480
rect 21256 67428 21324 67480
rect 21376 67428 21426 67480
rect 20945 67362 21426 67428
rect 20945 67310 21078 67362
rect 21130 67310 21204 67362
rect 21256 67310 21324 67362
rect 21376 67310 21426 67362
rect 20945 67275 21426 67310
rect 463 67220 947 67268
rect 20946 67262 21426 67275
rect 463 67048 863 67109
rect 463 66996 514 67048
rect 566 66996 636 67048
rect 688 66996 762 67048
rect 814 66996 863 67048
rect 463 66901 863 66996
rect 463 66849 514 66901
rect 566 66849 636 66901
rect 688 66849 762 66901
rect 814 66849 863 66901
rect 463 66764 863 66849
rect 463 66712 514 66764
rect 566 66712 636 66764
rect 688 66712 762 66764
rect 814 66712 863 66764
rect 463 66650 863 66712
rect 20946 66046 22370 66083
rect 20946 65994 22020 66046
rect 22072 65994 22146 66046
rect 22198 65994 22266 66046
rect 22318 65994 22370 66046
rect 20946 65928 22370 65994
rect 20946 65876 22020 65928
rect 22072 65876 22146 65928
rect 22198 65876 22266 65928
rect 22318 65876 22370 65928
rect 20946 65828 22370 65876
rect 463 65289 863 65350
rect 463 65237 514 65289
rect 566 65237 636 65289
rect 688 65237 762 65289
rect 814 65237 863 65289
rect 463 65142 863 65237
rect 463 65090 514 65142
rect 566 65090 636 65142
rect 688 65090 762 65142
rect 814 65090 863 65142
rect 463 65005 863 65090
rect 463 64953 514 65005
rect 566 64953 636 65005
rect 688 64953 762 65005
rect 814 64953 863 65005
rect 463 64891 863 64953
rect 463 64698 947 64735
rect 463 64646 513 64698
rect 565 64646 639 64698
rect 691 64646 759 64698
rect 811 64646 947 64698
rect 463 64580 947 64646
rect 463 64528 513 64580
rect 565 64528 639 64580
rect 691 64528 759 64580
rect 811 64528 947 64580
rect 463 64480 947 64528
rect 20945 64720 20946 64760
rect 20945 64683 21428 64720
rect 20945 64631 21078 64683
rect 21130 64631 21204 64683
rect 21256 64631 21324 64683
rect 21376 64631 21428 64683
rect 20945 64565 21428 64631
rect 20945 64513 21078 64565
rect 21130 64513 21204 64565
rect 21256 64513 21324 64565
rect 21376 64513 21428 64565
rect 20945 64505 21428 64513
rect 20946 64465 21428 64505
rect 463 63520 947 63557
rect 463 63468 513 63520
rect 565 63468 639 63520
rect 691 63468 759 63520
rect 811 63468 947 63520
rect 463 63402 947 63468
rect 463 63350 513 63402
rect 565 63350 639 63402
rect 691 63350 759 63402
rect 811 63350 947 63402
rect 463 63302 947 63350
rect 20944 63480 21426 63517
rect 20944 63428 21078 63480
rect 21130 63428 21204 63480
rect 21256 63428 21324 63480
rect 21376 63428 21426 63480
rect 20944 63362 21426 63428
rect 20944 63310 21078 63362
rect 21130 63310 21204 63362
rect 21256 63310 21324 63362
rect 21376 63310 21426 63362
rect 20944 63262 21426 63310
rect 464 63068 864 63109
rect 463 63048 864 63068
rect 463 62996 514 63048
rect 566 62996 636 63048
rect 688 62996 762 63048
rect 814 62996 864 63048
rect 463 62901 864 62996
rect 463 62849 514 62901
rect 566 62849 636 62901
rect 688 62849 762 62901
rect 814 62849 864 62901
rect 463 62764 864 62849
rect 463 62712 514 62764
rect 566 62712 636 62764
rect 688 62712 762 62764
rect 814 62712 864 62764
rect 463 62650 864 62712
rect 20946 62045 22370 62082
rect 20946 61993 22020 62045
rect 22072 61993 22146 62045
rect 22198 61993 22266 62045
rect 22318 61993 22370 62045
rect 20946 61927 22370 61993
rect 20946 61875 22020 61927
rect 22072 61875 22146 61927
rect 22198 61875 22266 61927
rect 22318 61875 22370 61927
rect 20946 61827 22370 61875
rect 463 61289 863 61350
rect 463 61237 514 61289
rect 566 61237 636 61289
rect 688 61237 762 61289
rect 814 61237 863 61289
rect 463 61142 863 61237
rect 463 61090 514 61142
rect 566 61090 636 61142
rect 688 61090 762 61142
rect 814 61090 863 61142
rect 463 61005 863 61090
rect 463 60953 514 61005
rect 566 60953 636 61005
rect 688 60953 762 61005
rect 814 60953 863 61005
rect 463 60891 863 60953
rect 463 60672 949 60709
rect 463 60620 513 60672
rect 565 60620 639 60672
rect 691 60620 759 60672
rect 811 60620 949 60672
rect 463 60554 949 60620
rect 463 60502 513 60554
rect 565 60502 639 60554
rect 691 60502 759 60554
rect 811 60502 949 60554
rect 463 60454 949 60502
rect 20946 60683 21428 60720
rect 20946 60631 21078 60683
rect 21130 60631 21204 60683
rect 21256 60631 21324 60683
rect 21376 60631 21428 60683
rect 20946 60565 21428 60631
rect 20946 60513 21078 60565
rect 21130 60513 21204 60565
rect 21256 60513 21324 60565
rect 21376 60513 21428 60565
rect 20946 60465 21428 60513
rect 20945 59534 21427 59571
rect 463 59469 947 59506
rect 463 59417 513 59469
rect 565 59417 639 59469
rect 691 59417 759 59469
rect 811 59417 947 59469
rect 463 59351 947 59417
rect 463 59299 513 59351
rect 565 59299 639 59351
rect 691 59299 759 59351
rect 811 59299 947 59351
rect 20945 59482 21078 59534
rect 21130 59482 21204 59534
rect 21256 59482 21324 59534
rect 21376 59482 21427 59534
rect 20945 59416 21427 59482
rect 20945 59364 21078 59416
rect 21130 59364 21204 59416
rect 21256 59364 21324 59416
rect 21376 59364 21427 59416
rect 20945 59316 21427 59364
rect 463 59251 947 59299
rect 464 59068 864 59109
rect 463 59048 864 59068
rect 463 58996 514 59048
rect 566 58996 636 59048
rect 688 58996 762 59048
rect 814 58996 864 59048
rect 463 58901 864 58996
rect 463 58849 514 58901
rect 566 58849 636 58901
rect 688 58849 762 58901
rect 814 58849 864 58901
rect 463 58764 864 58849
rect 463 58712 514 58764
rect 566 58712 636 58764
rect 688 58712 762 58764
rect 814 58712 864 58764
rect 463 58650 864 58712
rect 20946 58084 22370 58121
rect 20946 58032 22020 58084
rect 22072 58032 22146 58084
rect 22198 58032 22266 58084
rect 22318 58032 22370 58084
rect 20946 57966 22370 58032
rect 20946 57914 22020 57966
rect 22072 57914 22146 57966
rect 22198 57914 22266 57966
rect 22318 57914 22370 57966
rect 20946 57866 22370 57914
rect 463 57287 863 57348
rect 463 57235 514 57287
rect 566 57235 636 57287
rect 688 57235 762 57287
rect 814 57235 863 57287
rect 463 57140 863 57235
rect 463 57088 514 57140
rect 566 57088 636 57140
rect 688 57088 762 57140
rect 814 57088 863 57140
rect 463 57003 863 57088
rect 463 56951 514 57003
rect 566 56951 636 57003
rect 688 56951 762 57003
rect 814 56951 863 57003
rect 463 56889 863 56951
rect 463 56692 947 56729
rect 463 56640 513 56692
rect 565 56640 639 56692
rect 691 56640 759 56692
rect 811 56640 947 56692
rect 463 56574 947 56640
rect 463 56522 513 56574
rect 565 56522 639 56574
rect 691 56522 759 56574
rect 811 56522 947 56574
rect 463 56474 947 56522
rect 20946 56618 21428 56655
rect 20946 56566 21078 56618
rect 21130 56566 21204 56618
rect 21256 56566 21324 56618
rect 21376 56566 21428 56618
rect 20946 56500 21428 56566
rect 20946 56448 21078 56500
rect 21130 56448 21204 56500
rect 21256 56448 21324 56500
rect 21376 56448 21428 56500
rect 20946 56400 21428 56448
rect 463 55485 949 55522
rect 463 55433 513 55485
rect 565 55433 639 55485
rect 691 55433 759 55485
rect 811 55433 949 55485
rect 463 55367 949 55433
rect 463 55315 513 55367
rect 565 55315 639 55367
rect 691 55315 759 55367
rect 811 55315 949 55367
rect 463 55267 949 55315
rect 20945 55435 21427 55472
rect 20945 55383 21078 55435
rect 21130 55383 21204 55435
rect 21256 55383 21324 55435
rect 21376 55383 21427 55435
rect 20945 55317 21427 55383
rect 20945 55265 21078 55317
rect 21130 55265 21204 55317
rect 21256 55265 21324 55317
rect 21376 55265 21427 55317
rect 20945 55217 21427 55265
rect 463 55048 863 55109
rect 463 54996 514 55048
rect 566 54996 636 55048
rect 688 54996 762 55048
rect 814 54996 863 55048
rect 463 54901 863 54996
rect 463 54849 514 54901
rect 566 54849 636 54901
rect 688 54849 762 54901
rect 814 54849 863 54901
rect 463 54764 863 54849
rect 463 54712 514 54764
rect 566 54712 636 54764
rect 688 54712 762 54764
rect 814 54712 863 54764
rect 463 54650 863 54712
rect 20946 54067 22370 54104
rect 20946 54015 22020 54067
rect 22072 54015 22146 54067
rect 22198 54015 22266 54067
rect 22318 54015 22370 54067
rect 20946 53949 22370 54015
rect 20946 53897 22020 53949
rect 22072 53897 22146 53949
rect 22198 53897 22266 53949
rect 22318 53897 22370 53949
rect 20946 53849 22370 53897
rect 463 53289 863 53350
rect 463 53237 514 53289
rect 566 53237 636 53289
rect 688 53237 762 53289
rect 814 53237 863 53289
rect 463 53142 863 53237
rect 463 53090 514 53142
rect 566 53090 636 53142
rect 688 53090 762 53142
rect 814 53090 863 53142
rect 463 53005 863 53090
rect 463 52953 514 53005
rect 566 52953 636 53005
rect 688 52953 762 53005
rect 814 52953 863 53005
rect 463 52891 863 52953
rect 463 52719 947 52756
rect 463 52667 513 52719
rect 565 52667 639 52719
rect 691 52667 759 52719
rect 811 52667 947 52719
rect 463 52601 947 52667
rect 463 52549 513 52601
rect 565 52549 639 52601
rect 691 52549 759 52601
rect 811 52549 947 52601
rect 463 52501 947 52549
rect 20946 52563 21428 52600
rect 20946 52511 21078 52563
rect 21130 52511 21204 52563
rect 21256 52511 21324 52563
rect 21376 52511 21428 52563
rect 20946 52445 21428 52511
rect 20946 52393 21078 52445
rect 21130 52393 21204 52445
rect 21256 52393 21324 52445
rect 21376 52393 21428 52445
rect 20946 52345 21428 52393
rect 463 51532 947 51569
rect 463 51480 513 51532
rect 565 51480 639 51532
rect 691 51480 759 51532
rect 811 51480 947 51532
rect 463 51414 947 51480
rect 463 51362 513 51414
rect 565 51362 639 51414
rect 691 51362 759 51414
rect 811 51362 947 51414
rect 463 51314 947 51362
rect 20946 51428 21428 51465
rect 20946 51376 21078 51428
rect 21130 51376 21204 51428
rect 21256 51376 21324 51428
rect 21376 51376 21428 51428
rect 20946 51310 21428 51376
rect 20946 51258 21078 51310
rect 21130 51258 21204 51310
rect 21256 51258 21324 51310
rect 21376 51258 21428 51310
rect 20946 51210 21428 51258
rect 463 51048 863 51109
rect 463 50996 514 51048
rect 566 50996 636 51048
rect 688 50996 762 51048
rect 814 50996 863 51048
rect 463 50901 863 50996
rect 463 50849 514 50901
rect 566 50849 636 50901
rect 688 50849 762 50901
rect 814 50849 863 50901
rect 463 50764 863 50849
rect 463 50712 514 50764
rect 566 50712 636 50764
rect 688 50712 762 50764
rect 814 50712 863 50764
rect 463 50650 863 50712
rect 20946 50146 22370 50183
rect 20946 50094 22020 50146
rect 22072 50094 22146 50146
rect 22198 50094 22266 50146
rect 22318 50094 22370 50146
rect 20946 50028 22370 50094
rect 20946 49976 22020 50028
rect 22072 49976 22146 50028
rect 22198 49976 22266 50028
rect 22318 49976 22370 50028
rect 20946 49928 22370 49976
rect 463 49289 863 49350
rect 463 49237 514 49289
rect 566 49237 636 49289
rect 688 49237 762 49289
rect 814 49237 863 49289
rect 463 49142 863 49237
rect 463 49090 514 49142
rect 566 49090 636 49142
rect 688 49090 762 49142
rect 814 49090 863 49142
rect 463 49005 863 49090
rect 463 48953 514 49005
rect 566 48953 636 49005
rect 688 48953 762 49005
rect 814 48953 863 49005
rect 463 48891 863 48953
rect 463 48710 947 48747
rect 463 48658 513 48710
rect 565 48658 639 48710
rect 691 48658 759 48710
rect 811 48658 947 48710
rect 463 48592 947 48658
rect 463 48540 513 48592
rect 565 48540 639 48592
rect 691 48540 759 48592
rect 811 48540 947 48592
rect 463 48492 947 48540
rect 20946 48669 21428 48706
rect 20946 48617 21078 48669
rect 21130 48617 21204 48669
rect 21256 48617 21324 48669
rect 21376 48617 21428 48669
rect 20946 48551 21428 48617
rect 20946 48499 21078 48551
rect 21130 48499 21204 48551
rect 21256 48499 21324 48551
rect 21376 48499 21428 48551
rect 20946 48451 21428 48499
rect 463 47557 947 47594
rect 463 47505 513 47557
rect 565 47505 639 47557
rect 691 47505 759 47557
rect 811 47505 947 47557
rect 463 47439 947 47505
rect 463 47387 513 47439
rect 565 47387 639 47439
rect 691 47387 759 47439
rect 811 47387 947 47439
rect 463 47339 947 47387
rect 20946 47516 21428 47553
rect 20946 47464 21078 47516
rect 21130 47464 21204 47516
rect 21256 47464 21324 47516
rect 21376 47464 21428 47516
rect 20946 47398 21428 47464
rect 20946 47346 21078 47398
rect 21130 47346 21204 47398
rect 21256 47346 21324 47398
rect 21376 47346 21428 47398
rect 20946 47298 21428 47346
rect 463 47048 863 47109
rect 463 46996 514 47048
rect 566 46996 636 47048
rect 688 46996 762 47048
rect 814 46996 863 47048
rect 463 46901 863 46996
rect 463 46849 514 46901
rect 566 46849 636 46901
rect 688 46849 762 46901
rect 814 46849 863 46901
rect 463 46764 863 46849
rect 463 46712 514 46764
rect 566 46712 636 46764
rect 688 46712 762 46764
rect 814 46712 863 46764
rect 463 46650 863 46712
rect 20946 45888 22370 45925
rect 20946 45836 22020 45888
rect 22072 45836 22146 45888
rect 22198 45836 22266 45888
rect 22318 45836 22370 45888
rect 20946 45770 22370 45836
rect 20946 45718 22020 45770
rect 22072 45718 22146 45770
rect 22198 45718 22266 45770
rect 22318 45718 22370 45770
rect 20946 45670 22370 45718
rect 463 45288 863 45350
rect 463 45236 514 45288
rect 566 45236 636 45288
rect 688 45236 762 45288
rect 814 45236 863 45288
rect 463 45141 863 45236
rect 463 45089 514 45141
rect 566 45089 636 45141
rect 688 45089 762 45141
rect 814 45089 863 45141
rect 463 45004 863 45089
rect 463 44952 514 45004
rect 566 44952 636 45004
rect 688 44952 762 45004
rect 814 44952 863 45004
rect 463 44891 863 44952
rect 463 44890 836 44891
rect 463 44497 946 44534
rect 463 44445 513 44497
rect 565 44445 639 44497
rect 691 44445 759 44497
rect 811 44445 946 44497
rect 463 44379 946 44445
rect 463 44327 513 44379
rect 565 44327 639 44379
rect 691 44327 759 44379
rect 811 44327 946 44379
rect 463 44279 946 44327
rect 20946 44400 21428 44437
rect 20946 44348 21078 44400
rect 21130 44348 21204 44400
rect 21256 44348 21324 44400
rect 21376 44348 21428 44400
rect 20946 44282 21428 44348
rect 20946 44230 21078 44282
rect 21130 44230 21204 44282
rect 21256 44230 21324 44282
rect 21376 44230 21428 44282
rect 20946 44182 21428 44230
rect 3287 39752 4421 39753
rect 0 39727 21902 39752
rect 0 39675 46 39727
rect 98 39675 171 39727
rect 223 39675 296 39727
rect 348 39712 21902 39727
rect 348 39675 21549 39712
rect 0 39660 21549 39675
rect 21601 39660 21674 39712
rect 21726 39660 21799 39712
rect 21851 39660 21902 39712
rect 0 39621 21902 39660
rect 0 39569 46 39621
rect 98 39569 171 39621
rect 223 39569 296 39621
rect 348 39592 21902 39621
rect 348 39569 21548 39592
rect 0 39540 21548 39569
rect 21600 39540 21673 39592
rect 21725 39540 21798 39592
rect 21850 39540 21902 39592
rect 0 39497 21902 39540
rect 1868 39391 2335 39410
rect 1868 39364 1891 39391
rect 1997 39364 2047 39391
rect 2153 39364 2203 39391
rect 2309 39364 2335 39391
rect 1650 39321 1796 39329
rect 1650 39269 1662 39321
rect 1714 39269 1732 39321
rect 1784 39269 1796 39321
rect 1868 39312 1886 39364
rect 2002 39312 2042 39364
rect 2158 39312 2198 39364
rect 2314 39312 2335 39364
rect 1868 39285 1891 39312
rect 1997 39285 2047 39312
rect 2153 39285 2203 39312
rect 2309 39285 2335 39312
rect 1868 39270 2335 39285
rect 2539 39328 2685 39336
rect 2539 39276 2551 39328
rect 2603 39276 2621 39328
rect 2673 39276 2685 39328
rect 1650 39251 1796 39269
rect 1650 39199 1662 39251
rect 1714 39199 1732 39251
rect 1784 39233 1796 39251
rect 2539 39258 2685 39276
rect 2167 39233 2239 39236
rect 1784 39227 2239 39233
rect 1784 39199 2192 39227
rect 1650 39193 2192 39199
rect 2226 39193 2239 39227
rect 2539 39206 2551 39258
rect 2603 39206 2621 39258
rect 2673 39206 2685 39258
rect 2539 39196 2685 39206
rect 1650 39189 2239 39193
rect 2167 39185 2239 39189
rect 924 39139 1188 39173
rect 463 39117 2973 39139
rect 463 39065 494 39117
rect 546 39065 608 39117
rect 660 39065 722 39117
rect 774 39116 1114 39117
rect 774 39082 960 39116
rect 994 39083 1114 39116
rect 1148 39113 2973 39117
rect 1148 39109 1920 39113
rect 1148 39083 1604 39109
rect 994 39082 1604 39083
rect 774 39075 1604 39082
rect 1638 39079 1920 39109
rect 1954 39079 2973 39113
rect 1638 39075 2973 39079
rect 774 39065 2973 39075
rect 463 39043 2973 39065
rect 924 39003 1188 39043
rect 924 39000 1114 39003
rect 924 38966 963 39000
rect 997 38969 1114 39000
rect 1148 38969 1188 39003
rect 997 38966 1188 38969
rect 924 38923 1188 38966
rect 2889 38982 2950 38987
rect 2889 38981 3370 38982
rect 1592 38933 1966 38954
rect 1592 38899 1604 38933
rect 1638 38899 1920 38933
rect 1954 38899 1966 38933
rect 1592 38882 1966 38899
rect 2022 38933 2397 38954
rect 2022 38899 2035 38933
rect 2069 38899 2351 38933
rect 2385 38899 2397 38933
rect 2022 38882 2397 38899
rect 2467 38936 2843 38955
rect 2889 38947 2901 38981
rect 2935 38947 3370 38981
rect 2889 38946 3370 38947
rect 2889 38941 2950 38946
rect 2467 38902 2479 38936
rect 2513 38902 2797 38936
rect 2831 38902 2843 38936
rect 2467 38883 2843 38902
rect 2900 38870 3301 38876
rect 2900 38836 2921 38870
rect 2955 38836 3253 38870
rect 3287 38836 3301 38870
rect 2900 38829 3301 38836
rect 1495 38774 1569 38781
rect 1495 38722 1507 38774
rect 1559 38770 1569 38774
rect 1755 38770 1802 38794
rect 3342 38772 3370 38946
rect 3615 38960 4297 38966
rect 3615 38926 4251 38960
rect 4285 38926 4297 38960
rect 3615 38920 4297 38926
rect 3523 38828 3529 38880
rect 3581 38876 3587 38880
rect 3615 38876 3650 38920
rect 4610 38879 4662 38885
rect 4092 38876 4156 38878
rect 3581 38870 3650 38876
rect 3587 38836 3650 38870
rect 3581 38830 3650 38836
rect 4075 38870 4385 38876
rect 4075 38836 4105 38870
rect 4139 38836 4339 38870
rect 4373 38836 4385 38870
rect 4075 38830 4385 38836
rect 3581 38828 3587 38830
rect 4092 38826 4156 38830
rect 4608 38829 4610 38877
rect 3792 38813 3841 38825
rect 4610 38821 4662 38827
rect 3792 38779 3800 38813
rect 3834 38779 3841 38813
rect 3792 38772 3841 38779
rect 1559 38761 1802 38770
rect 1559 38727 1762 38761
rect 1796 38727 1802 38761
rect 3341 38737 3841 38772
rect 1559 38722 1802 38727
rect 1495 38717 1802 38722
rect 1755 38694 1802 38717
rect 0 38573 1593 38595
rect 0 38521 31 38573
rect 83 38521 145 38573
rect 197 38521 259 38573
rect 311 38521 1593 38573
rect 0 38499 1593 38521
rect 3608 38348 3660 38354
rect 1893 38305 3608 38334
rect 1465 38217 1471 38269
rect 1523 38268 1529 38269
rect 1523 38258 1773 38268
rect 1523 38224 1715 38258
rect 1749 38224 1773 38258
rect 1523 38218 1773 38224
rect 1801 38261 1847 38275
rect 1801 38227 1807 38261
rect 1841 38227 1847 38261
rect 1523 38217 1529 38218
rect 1801 38210 1847 38227
rect 1893 38258 1941 38305
rect 3608 38290 3660 38296
rect 1893 38224 1899 38258
rect 1933 38224 1941 38258
rect 1893 38212 1941 38224
rect 2019 38252 2076 38275
rect 2019 38218 2029 38252
rect 2063 38218 2076 38252
rect 1805 38184 1847 38210
rect 2019 38202 2076 38218
rect 4652 38267 4704 38273
rect 4652 38209 4704 38215
rect 2019 38184 2063 38202
rect 1805 38155 2063 38184
rect 463 38029 2056 38051
rect 463 37977 494 38029
rect 546 37977 608 38029
rect 660 37977 722 38029
rect 774 37977 2056 38029
rect 463 37955 2056 37977
rect 3517 37889 3523 37897
rect 1874 37854 3523 37889
rect 1457 37738 1463 37790
rect 1515 37738 1539 37790
rect 1799 37787 1845 37851
rect 1799 37753 1805 37787
rect 1839 37753 1845 37787
rect 1799 37708 1845 37753
rect 1874 37788 1940 37854
rect 3517 37845 3523 37854
rect 3575 37845 3581 37897
rect 1874 37754 1889 37788
rect 1923 37754 1940 37788
rect 1874 37738 1940 37754
rect 1980 37782 2032 37795
rect 1980 37748 1986 37782
rect 2020 37748 2032 37782
rect 1980 37708 2032 37748
rect 4652 37791 4704 37797
rect 4652 37733 4704 37739
rect 1799 37680 2032 37708
rect 0 37485 1317 37507
rect 0 37433 31 37485
rect 83 37433 145 37485
rect 197 37433 259 37485
rect 311 37433 1317 37485
rect 0 37411 1317 37433
rect 1680 37358 1739 37375
rect 1680 37306 1683 37358
rect 1735 37306 1739 37358
rect 1680 37252 1739 37306
rect 1680 37200 1683 37252
rect 1735 37200 1739 37252
rect 1680 37150 1739 37200
rect 3332 37265 3841 37300
rect 2867 37172 3295 37178
rect 1680 37134 2320 37150
rect 924 37052 1188 37111
rect 1680 37100 1957 37134
rect 1991 37133 2320 37134
rect 1991 37100 2273 37133
rect 1680 37099 2273 37100
rect 2307 37099 2320 37133
rect 1680 37084 2320 37099
rect 2416 37137 2804 37152
rect 2416 37103 2436 37137
rect 2470 37134 2804 37137
rect 2470 37103 2753 37134
rect 2416 37100 2753 37103
rect 2787 37100 2804 37134
rect 2867 37138 2902 37172
rect 2936 37171 3295 37172
rect 2936 37138 3237 37171
rect 2867 37137 3237 37138
rect 3271 37137 3295 37171
rect 2867 37131 3295 37137
rect 2416 37085 2804 37100
rect 1680 37083 1739 37084
rect 1945 37083 2320 37084
rect 3332 37069 3375 37265
rect 3806 37233 3841 37265
rect 3801 37227 3848 37233
rect 3801 37193 3807 37227
rect 3841 37193 3848 37227
rect 3547 37176 3553 37182
rect 3523 37130 3553 37176
rect 3605 37130 3646 37182
rect 3801 37181 3848 37193
rect 4609 37181 4661 37187
rect 2969 37058 3375 37069
rect 924 37018 977 37052
rect 1011 37018 1105 37052
rect 1139 37018 1188 37052
rect 924 36963 1188 37018
rect 2910 37037 3375 37058
rect 3610 37086 3646 37130
rect 4075 37178 4156 37180
rect 4075 37170 4569 37178
rect 4075 37136 4105 37170
rect 4139 37136 4523 37170
rect 4557 37136 4569 37170
rect 4075 37130 4569 37136
rect 4075 37128 4156 37130
rect 4609 37123 4661 37129
rect 3610 37080 4297 37086
rect 3610 37046 4251 37080
rect 4285 37046 4297 37080
rect 3610 37038 4297 37046
rect 2910 37003 2917 37037
rect 2951 37034 3375 37037
rect 2951 37023 2987 37034
rect 2951 37003 2959 37023
rect 2910 36991 2959 37003
rect 463 36941 2973 36963
rect 463 36889 494 36941
rect 546 36889 608 36941
rect 660 36889 722 36941
rect 774 36922 2973 36941
rect 774 36889 977 36922
rect 463 36888 977 36889
rect 1011 36888 1106 36922
rect 1140 36888 2973 36922
rect 463 36867 2973 36888
rect 924 36835 1188 36867
rect 2538 36830 2685 36838
rect 2538 36778 2551 36830
rect 2603 36778 2621 36830
rect 2673 36778 2685 36830
rect 2538 36763 2685 36778
rect 2538 36711 2551 36763
rect 2603 36711 2621 36763
rect 2673 36711 2685 36763
rect 2538 36649 2685 36711
rect 2752 36830 2899 36838
rect 2752 36778 2765 36830
rect 2817 36778 2835 36830
rect 2887 36778 2899 36830
rect 2752 36765 2899 36778
rect 2752 36713 2765 36765
rect 2817 36713 2835 36765
rect 2887 36713 2899 36765
rect 2752 36707 2899 36713
rect 20527 36158 21428 36198
rect 20527 36106 21075 36158
rect 21127 36106 21200 36158
rect 21252 36106 21325 36158
rect 21377 36106 21428 36158
rect 20527 36038 21428 36106
rect 20527 35986 21074 36038
rect 21126 35986 21199 36038
rect 21251 35986 21324 36038
rect 21376 35986 21428 36038
rect 20527 35943 21428 35986
rect 21028 35580 21428 35642
rect 21028 35528 21079 35580
rect 21131 35528 21201 35580
rect 21253 35528 21327 35580
rect 21379 35528 21428 35580
rect 21028 35433 21428 35528
rect 21028 35381 21079 35433
rect 21131 35381 21201 35433
rect 21253 35381 21327 35433
rect 21379 35381 21428 35433
rect 21028 35296 21428 35381
rect 21028 35244 21079 35296
rect 21131 35244 21201 35296
rect 21253 35244 21327 35296
rect 21379 35244 21428 35296
rect 21028 35183 21428 35244
rect 21028 35182 21401 35183
rect 20526 34662 21902 34702
rect 20526 34610 20574 34662
rect 20626 34610 20699 34662
rect 20751 34610 20824 34662
rect 20876 34610 21549 34662
rect 21601 34610 21674 34662
rect 21726 34610 21799 34662
rect 21851 34610 21902 34662
rect 20526 34542 21902 34610
rect 20526 34490 20573 34542
rect 20625 34490 20698 34542
rect 20750 34490 20823 34542
rect 20875 34490 21548 34542
rect 21600 34490 21673 34542
rect 21725 34490 21798 34542
rect 21850 34490 21902 34542
rect 20526 34447 21902 34490
rect 21028 33820 21428 33882
rect 21028 33768 21079 33820
rect 21131 33768 21201 33820
rect 21253 33768 21327 33820
rect 21379 33768 21428 33820
rect 21028 33673 21428 33768
rect 21028 33621 21079 33673
rect 21131 33621 21201 33673
rect 21253 33621 21327 33673
rect 21379 33621 21428 33673
rect 21028 33536 21428 33621
rect 21028 33484 21079 33536
rect 21131 33484 21201 33536
rect 21253 33484 21327 33536
rect 21379 33484 21428 33536
rect 21028 33423 21428 33484
rect 21028 33422 21401 33423
rect 20514 33103 21427 33143
rect 20514 33051 21074 33103
rect 21126 33051 21199 33103
rect 21251 33051 21324 33103
rect 21376 33051 21427 33103
rect 20514 32983 21427 33051
rect 20514 32931 21073 32983
rect 21125 32931 21198 32983
rect 21250 32931 21323 32983
rect 21375 32931 21427 32983
rect 20514 32888 21427 32931
rect 463 32290 21428 32360
rect 463 32238 513 32290
rect 565 32238 639 32290
rect 691 32238 759 32290
rect 811 32238 21078 32290
rect 21130 32238 21204 32290
rect 21256 32238 21324 32290
rect 21376 32238 21428 32290
rect 463 32172 21428 32238
rect 463 32120 513 32172
rect 565 32120 639 32172
rect 691 32120 759 32172
rect 811 32120 21078 32172
rect 21130 32120 21204 32172
rect 21256 32120 21324 32172
rect 21376 32120 21428 32172
rect 463 32073 21428 32120
rect 463 32072 1825 32073
rect 2313 32072 21428 32073
rect 463 31508 946 31545
rect 463 31456 513 31508
rect 565 31456 639 31508
rect 691 31456 759 31508
rect 811 31456 946 31508
rect 463 31390 946 31456
rect 463 31338 513 31390
rect 565 31338 639 31390
rect 691 31338 759 31390
rect 811 31338 946 31390
rect 463 31290 946 31338
rect 20946 31508 21428 31545
rect 20946 31456 21078 31508
rect 21130 31456 21204 31508
rect 21256 31456 21324 31508
rect 21376 31456 21428 31508
rect 20946 31390 21428 31456
rect 20946 31338 21078 31390
rect 21130 31338 21204 31390
rect 21256 31338 21324 31390
rect 21376 31338 21428 31390
rect 20946 31290 21428 31338
rect 463 31049 863 31111
rect 463 30997 514 31049
rect 566 30997 636 31049
rect 688 30997 762 31049
rect 814 30997 863 31049
rect 463 30902 863 30997
rect 463 30850 514 30902
rect 566 30850 636 30902
rect 688 30850 762 30902
rect 814 30850 863 30902
rect 463 30765 863 30850
rect 463 30713 514 30765
rect 566 30713 636 30765
rect 688 30713 762 30765
rect 814 30713 863 30765
rect 463 30651 863 30713
rect 20946 30118 22370 30155
rect 20946 30066 22020 30118
rect 22072 30066 22146 30118
rect 22198 30066 22266 30118
rect 22318 30066 22370 30118
rect 20946 30000 22370 30066
rect 20946 29948 22020 30000
rect 22072 29948 22146 30000
rect 22198 29948 22266 30000
rect 22318 29948 22370 30000
rect 20946 29900 22370 29948
rect 463 29282 863 29350
rect 463 29230 514 29282
rect 566 29230 636 29282
rect 688 29230 762 29282
rect 814 29230 863 29282
rect 463 29135 863 29230
rect 463 29083 514 29135
rect 566 29083 636 29135
rect 688 29083 762 29135
rect 814 29083 863 29135
rect 463 28998 863 29083
rect 463 28946 514 28998
rect 566 28946 636 28998
rect 688 28946 762 28998
rect 814 28946 863 28998
rect 463 28890 863 28946
rect 463 28596 946 28633
rect 463 28544 513 28596
rect 565 28544 639 28596
rect 691 28544 759 28596
rect 811 28544 946 28596
rect 463 28478 946 28544
rect 463 28426 513 28478
rect 565 28426 639 28478
rect 691 28426 759 28478
rect 811 28426 946 28478
rect 463 28378 946 28426
rect 20946 28547 21428 28584
rect 20946 28495 21078 28547
rect 21130 28495 21204 28547
rect 21256 28495 21324 28547
rect 21376 28495 21428 28547
rect 20946 28429 21428 28495
rect 20946 28377 21078 28429
rect 21130 28377 21204 28429
rect 21256 28377 21324 28429
rect 21376 28377 21428 28429
rect 20946 28329 21428 28377
rect 463 27592 946 27629
rect 463 27540 513 27592
rect 565 27540 639 27592
rect 691 27540 759 27592
rect 811 27540 946 27592
rect 463 27474 946 27540
rect 463 27422 513 27474
rect 565 27422 639 27474
rect 691 27422 759 27474
rect 811 27422 946 27474
rect 463 27374 946 27422
rect 20945 27430 21427 27467
rect 20945 27378 21078 27430
rect 21130 27378 21204 27430
rect 21256 27378 21324 27430
rect 21376 27378 21427 27430
rect 20945 27312 21427 27378
rect 20945 27260 21078 27312
rect 21130 27260 21204 27312
rect 21256 27260 21324 27312
rect 21376 27260 21427 27312
rect 20945 27212 21427 27260
rect 463 27048 863 27109
rect 463 26996 514 27048
rect 566 26996 636 27048
rect 688 26996 762 27048
rect 814 26996 863 27048
rect 463 26901 863 26996
rect 463 26849 514 26901
rect 566 26849 636 26901
rect 688 26849 762 26901
rect 814 26849 863 26901
rect 463 26764 863 26849
rect 463 26712 514 26764
rect 566 26712 636 26764
rect 688 26712 762 26764
rect 814 26712 863 26764
rect 463 26650 863 26712
rect 20946 25959 22370 25996
rect 20946 25907 22020 25959
rect 22072 25907 22146 25959
rect 22198 25907 22266 25959
rect 22318 25907 22370 25959
rect 20946 25841 22370 25907
rect 20946 25789 22020 25841
rect 22072 25789 22146 25841
rect 22198 25789 22266 25841
rect 22318 25789 22370 25841
rect 20946 25741 22370 25789
rect 463 25288 863 25349
rect 463 25236 514 25288
rect 566 25236 636 25288
rect 688 25236 762 25288
rect 814 25236 863 25288
rect 463 25141 863 25236
rect 463 25089 514 25141
rect 566 25089 636 25141
rect 688 25089 762 25141
rect 814 25089 863 25141
rect 463 25004 863 25089
rect 463 24952 514 25004
rect 566 24952 636 25004
rect 688 24952 762 25004
rect 814 24952 863 25004
rect 463 24890 863 24952
rect 463 24614 947 24651
rect 463 24562 513 24614
rect 565 24562 639 24614
rect 691 24562 759 24614
rect 811 24562 947 24614
rect 463 24496 947 24562
rect 463 24444 513 24496
rect 565 24444 639 24496
rect 691 24444 759 24496
rect 811 24444 947 24496
rect 463 24396 947 24444
rect 20946 24587 21428 24624
rect 20946 24535 21078 24587
rect 21130 24535 21204 24587
rect 21256 24535 21324 24587
rect 21376 24535 21428 24587
rect 20946 24469 21428 24535
rect 20946 24417 21078 24469
rect 21130 24417 21204 24469
rect 21256 24417 21324 24469
rect 21376 24417 21428 24469
rect 20946 24369 21428 24417
rect 463 23532 947 23569
rect 463 23480 513 23532
rect 565 23480 639 23532
rect 691 23480 759 23532
rect 811 23480 947 23532
rect 463 23414 947 23480
rect 463 23362 513 23414
rect 565 23362 639 23414
rect 691 23362 759 23414
rect 811 23362 947 23414
rect 463 23314 947 23362
rect 20946 23412 21428 23449
rect 20946 23360 21078 23412
rect 21130 23360 21204 23412
rect 21256 23360 21324 23412
rect 21376 23360 21428 23412
rect 20946 23294 21428 23360
rect 20946 23242 21078 23294
rect 21130 23242 21204 23294
rect 21256 23242 21324 23294
rect 21376 23242 21428 23294
rect 20946 23194 21428 23242
rect 463 23048 863 23109
rect 463 22996 514 23048
rect 566 22996 636 23048
rect 688 22996 762 23048
rect 814 22996 863 23048
rect 463 22901 863 22996
rect 463 22849 514 22901
rect 566 22849 636 22901
rect 688 22849 762 22901
rect 814 22849 863 22901
rect 463 22764 863 22849
rect 463 22712 514 22764
rect 566 22712 636 22764
rect 688 22712 762 22764
rect 814 22712 863 22764
rect 463 22650 863 22712
rect 20946 22169 22370 22206
rect 20946 22117 22020 22169
rect 22072 22117 22146 22169
rect 22198 22117 22266 22169
rect 22318 22117 22370 22169
rect 20946 22051 22370 22117
rect 20946 21999 22020 22051
rect 22072 21999 22146 22051
rect 22198 21999 22266 22051
rect 22318 21999 22370 22051
rect 20946 21951 22370 21999
rect 463 21289 863 21350
rect 463 21237 514 21289
rect 566 21237 636 21289
rect 688 21237 762 21289
rect 814 21237 863 21289
rect 463 21142 863 21237
rect 463 21090 514 21142
rect 566 21090 636 21142
rect 688 21090 762 21142
rect 814 21090 863 21142
rect 463 21005 863 21090
rect 463 20953 514 21005
rect 566 20953 636 21005
rect 688 20953 762 21005
rect 814 20953 863 21005
rect 463 20891 863 20953
rect 463 20657 947 20694
rect 463 20605 513 20657
rect 565 20605 639 20657
rect 691 20605 759 20657
rect 811 20605 947 20657
rect 463 20539 947 20605
rect 463 20487 513 20539
rect 565 20487 639 20539
rect 691 20487 759 20539
rect 811 20487 947 20539
rect 463 20439 947 20487
rect 20945 20571 21427 20608
rect 20945 20519 21078 20571
rect 21130 20519 21204 20571
rect 21256 20519 21324 20571
rect 21376 20519 21427 20571
rect 20945 20453 21427 20519
rect 20945 20401 21078 20453
rect 21130 20401 21204 20453
rect 21256 20401 21324 20453
rect 21376 20401 21427 20453
rect 20945 20353 21427 20401
rect 463 19556 947 19593
rect 463 19504 513 19556
rect 565 19504 639 19556
rect 691 19504 759 19556
rect 811 19504 947 19556
rect 463 19438 947 19504
rect 463 19386 513 19438
rect 565 19386 639 19438
rect 691 19386 759 19438
rect 811 19386 947 19438
rect 463 19338 947 19386
rect 20945 19400 21427 19437
rect 20945 19348 21078 19400
rect 21130 19348 21204 19400
rect 21256 19348 21324 19400
rect 21376 19348 21427 19400
rect 20945 19282 21427 19348
rect 20945 19230 21078 19282
rect 21130 19230 21204 19282
rect 21256 19230 21324 19282
rect 21376 19230 21427 19282
rect 20945 19182 21427 19230
rect 463 19048 863 19109
rect 463 18996 514 19048
rect 566 18996 636 19048
rect 688 18996 762 19048
rect 814 18996 863 19048
rect 463 18901 863 18996
rect 463 18849 514 18901
rect 566 18849 636 18901
rect 688 18849 762 18901
rect 814 18849 863 18901
rect 463 18764 863 18849
rect 463 18712 514 18764
rect 566 18712 636 18764
rect 688 18712 762 18764
rect 814 18712 863 18764
rect 463 18650 863 18712
rect 20946 18062 22370 18099
rect 20946 18010 22020 18062
rect 22072 18010 22146 18062
rect 22198 18010 22266 18062
rect 22318 18010 22370 18062
rect 20946 17944 22370 18010
rect 20946 17892 22020 17944
rect 22072 17892 22146 17944
rect 22198 17892 22266 17944
rect 22318 17892 22370 17944
rect 20946 17844 22370 17892
rect 463 17288 863 17349
rect 463 17236 514 17288
rect 566 17236 636 17288
rect 688 17236 762 17288
rect 814 17236 863 17288
rect 463 17141 863 17236
rect 463 17089 514 17141
rect 566 17089 636 17141
rect 688 17089 762 17141
rect 814 17089 863 17141
rect 463 17004 863 17089
rect 463 16952 514 17004
rect 566 16952 636 17004
rect 688 16952 762 17004
rect 814 16952 863 17004
rect 463 16890 863 16952
rect 463 16690 948 16727
rect 463 16638 513 16690
rect 565 16638 639 16690
rect 691 16638 759 16690
rect 811 16638 948 16690
rect 463 16572 948 16638
rect 463 16520 513 16572
rect 565 16520 639 16572
rect 691 16520 759 16572
rect 811 16520 948 16572
rect 463 16472 948 16520
rect 20945 16639 21427 16676
rect 20945 16587 21078 16639
rect 21130 16587 21204 16639
rect 21256 16587 21324 16639
rect 21376 16587 21427 16639
rect 20945 16521 21427 16587
rect 20945 16469 21078 16521
rect 21130 16469 21204 16521
rect 21256 16469 21324 16521
rect 21376 16469 21427 16521
rect 20945 16421 21427 16469
rect 463 15474 949 15511
rect 463 15422 513 15474
rect 565 15422 639 15474
rect 691 15422 759 15474
rect 811 15422 949 15474
rect 463 15356 949 15422
rect 463 15304 513 15356
rect 565 15304 639 15356
rect 691 15304 759 15356
rect 811 15304 949 15356
rect 463 15256 949 15304
rect 20945 15425 21427 15462
rect 20945 15373 21078 15425
rect 21130 15373 21204 15425
rect 21256 15373 21324 15425
rect 21376 15373 21427 15425
rect 20945 15307 21427 15373
rect 20945 15255 21078 15307
rect 21130 15255 21204 15307
rect 21256 15255 21324 15307
rect 21376 15255 21427 15307
rect 20945 15207 21427 15255
rect 463 15048 863 15109
rect 463 14996 514 15048
rect 566 14996 636 15048
rect 688 14996 762 15048
rect 814 14996 863 15048
rect 463 14901 863 14996
rect 463 14849 514 14901
rect 566 14849 636 14901
rect 688 14849 762 14901
rect 814 14849 863 14901
rect 463 14764 863 14849
rect 463 14712 514 14764
rect 566 14712 636 14764
rect 688 14712 762 14764
rect 814 14712 863 14764
rect 463 14650 863 14712
rect 20946 14244 22370 14281
rect 20946 14192 22020 14244
rect 22072 14192 22146 14244
rect 22198 14192 22266 14244
rect 22318 14192 22370 14244
rect 20946 14126 22370 14192
rect 20946 14074 22020 14126
rect 22072 14074 22146 14126
rect 22198 14074 22266 14126
rect 22318 14074 22370 14126
rect 20946 14026 22370 14074
rect 463 13288 863 13349
rect 463 13236 514 13288
rect 566 13236 636 13288
rect 688 13236 762 13288
rect 814 13236 863 13288
rect 463 13141 863 13236
rect 463 13089 514 13141
rect 566 13089 636 13141
rect 688 13089 762 13141
rect 814 13089 863 13141
rect 463 13004 863 13089
rect 463 12952 514 13004
rect 566 12952 636 13004
rect 688 12952 762 13004
rect 814 12952 863 13004
rect 463 12890 863 12952
rect 463 12609 947 12646
rect 463 12557 513 12609
rect 565 12557 639 12609
rect 691 12557 759 12609
rect 811 12557 947 12609
rect 463 12491 947 12557
rect 463 12439 513 12491
rect 565 12439 639 12491
rect 691 12439 759 12491
rect 811 12439 947 12491
rect 463 12391 947 12439
rect 20946 12582 21428 12619
rect 20946 12530 21078 12582
rect 21130 12530 21204 12582
rect 21256 12530 21324 12582
rect 21376 12530 21428 12582
rect 20946 12464 21428 12530
rect 20946 12412 21078 12464
rect 21130 12412 21204 12464
rect 21256 12412 21324 12464
rect 21376 12412 21428 12464
rect 20946 12364 21428 12412
rect 463 11487 947 11524
rect 463 11435 513 11487
rect 565 11435 639 11487
rect 691 11435 759 11487
rect 811 11435 947 11487
rect 463 11369 947 11435
rect 463 11317 513 11369
rect 565 11317 639 11369
rect 691 11317 759 11369
rect 811 11317 947 11369
rect 463 11269 947 11317
rect 20946 11425 21427 11462
rect 20946 11373 21078 11425
rect 21130 11373 21204 11425
rect 21256 11373 21324 11425
rect 21376 11373 21427 11425
rect 20946 11307 21427 11373
rect 20946 11255 21078 11307
rect 21130 11255 21204 11307
rect 21256 11255 21324 11307
rect 21376 11255 21427 11307
rect 20946 11207 21427 11255
rect 463 11049 863 11110
rect 463 10997 514 11049
rect 566 10997 636 11049
rect 688 10997 762 11049
rect 814 10997 863 11049
rect 463 10902 863 10997
rect 463 10850 514 10902
rect 566 10850 636 10902
rect 688 10850 762 10902
rect 814 10850 863 10902
rect 463 10765 863 10850
rect 463 10713 514 10765
rect 566 10713 636 10765
rect 688 10713 762 10765
rect 814 10713 863 10765
rect 463 10651 863 10713
rect 20946 10280 22370 10317
rect 20946 10228 22020 10280
rect 22072 10228 22146 10280
rect 22198 10228 22266 10280
rect 22318 10228 22370 10280
rect 20946 10162 22370 10228
rect 20946 10110 22020 10162
rect 22072 10110 22146 10162
rect 22198 10110 22266 10162
rect 22318 10110 22370 10162
rect 20946 10062 22370 10110
rect 463 9287 863 9348
rect 463 9235 514 9287
rect 566 9235 636 9287
rect 688 9235 762 9287
rect 814 9235 863 9287
rect 463 9140 863 9235
rect 463 9088 514 9140
rect 566 9088 636 9140
rect 688 9088 762 9140
rect 814 9088 863 9140
rect 463 9003 863 9088
rect 463 8951 514 9003
rect 566 8951 636 9003
rect 688 8951 762 9003
rect 814 8951 863 9003
rect 463 8889 863 8951
rect 463 8627 946 8664
rect 463 8575 513 8627
rect 565 8575 639 8627
rect 691 8575 759 8627
rect 811 8575 946 8627
rect 463 8509 946 8575
rect 463 8457 513 8509
rect 565 8457 639 8509
rect 691 8457 759 8509
rect 811 8457 946 8509
rect 463 8409 946 8457
rect 20946 8582 21428 8619
rect 20946 8530 21078 8582
rect 21130 8530 21204 8582
rect 21256 8530 21324 8582
rect 21376 8530 21428 8582
rect 20946 8464 21428 8530
rect 20946 8412 21078 8464
rect 21130 8412 21204 8464
rect 21256 8412 21324 8464
rect 21376 8412 21428 8464
rect 20946 8364 21428 8412
rect 463 7516 946 7553
rect 463 7464 513 7516
rect 565 7464 639 7516
rect 691 7464 759 7516
rect 811 7464 946 7516
rect 463 7398 946 7464
rect 463 7346 513 7398
rect 565 7346 639 7398
rect 691 7346 759 7398
rect 811 7346 946 7398
rect 463 7298 946 7346
rect 20946 7425 21427 7462
rect 20946 7373 21078 7425
rect 21130 7373 21204 7425
rect 21256 7373 21324 7425
rect 21376 7373 21427 7425
rect 20946 7307 21427 7373
rect 20946 7255 21078 7307
rect 21130 7255 21204 7307
rect 21256 7255 21324 7307
rect 21376 7255 21427 7307
rect 20946 7207 21427 7255
rect 463 7049 863 7110
rect 463 6997 514 7049
rect 566 6997 636 7049
rect 688 6997 762 7049
rect 814 6997 863 7049
rect 463 6902 863 6997
rect 463 6850 514 6902
rect 566 6850 636 6902
rect 688 6850 762 6902
rect 814 6850 863 6902
rect 463 6765 863 6850
rect 463 6713 514 6765
rect 566 6713 636 6765
rect 688 6713 762 6765
rect 814 6713 863 6765
rect 463 6651 863 6713
rect 20946 6268 22370 6305
rect 20946 6216 22020 6268
rect 22072 6216 22146 6268
rect 22198 6216 22266 6268
rect 22318 6216 22370 6268
rect 20946 6150 22370 6216
rect 20946 6098 22020 6150
rect 22072 6098 22146 6150
rect 22198 6098 22266 6150
rect 22318 6098 22370 6150
rect 20946 6050 22370 6098
rect 463 5288 863 5349
rect 463 5236 514 5288
rect 566 5236 636 5288
rect 688 5236 762 5288
rect 814 5236 863 5288
rect 463 5141 863 5236
rect 463 5089 514 5141
rect 566 5089 636 5141
rect 688 5089 762 5141
rect 814 5089 863 5141
rect 463 5004 863 5089
rect 463 4952 514 5004
rect 566 4952 636 5004
rect 688 4952 762 5004
rect 814 4952 863 5004
rect 463 4890 863 4952
rect 463 4693 948 4730
rect 463 4641 513 4693
rect 565 4641 639 4693
rect 691 4641 759 4693
rect 811 4641 948 4693
rect 463 4575 948 4641
rect 463 4523 513 4575
rect 565 4523 639 4575
rect 691 4523 759 4575
rect 811 4523 948 4575
rect 463 4475 948 4523
rect 20946 4582 21428 4619
rect 20946 4530 21078 4582
rect 21130 4530 21204 4582
rect 21256 4530 21324 4582
rect 21376 4530 21428 4582
rect 20946 4464 21428 4530
rect 20946 4412 21078 4464
rect 21130 4412 21204 4464
rect 21256 4412 21324 4464
rect 21376 4412 21428 4464
rect 20946 4364 21428 4412
rect 463 3516 946 3553
rect 463 3464 513 3516
rect 565 3464 639 3516
rect 691 3464 759 3516
rect 811 3464 946 3516
rect 463 3398 946 3464
rect 463 3346 513 3398
rect 565 3346 639 3398
rect 691 3346 759 3398
rect 811 3346 946 3398
rect 463 3298 946 3346
rect 20946 3425 21427 3462
rect 20946 3373 21078 3425
rect 21130 3373 21204 3425
rect 21256 3373 21324 3425
rect 21376 3373 21427 3425
rect 20946 3307 21427 3373
rect 20946 3255 21078 3307
rect 21130 3255 21204 3307
rect 21256 3255 21324 3307
rect 21376 3255 21427 3307
rect 20946 3207 21427 3255
rect 463 3049 863 3110
rect 463 2997 514 3049
rect 566 2997 636 3049
rect 688 2997 762 3049
rect 814 2997 863 3049
rect 463 2902 863 2997
rect 463 2850 514 2902
rect 566 2850 636 2902
rect 688 2850 762 2902
rect 814 2850 863 2902
rect 463 2765 863 2850
rect 463 2713 514 2765
rect 566 2713 636 2765
rect 688 2713 762 2765
rect 814 2713 863 2765
rect 463 2651 863 2713
rect 20946 2268 22370 2305
rect 20946 2216 22020 2268
rect 22072 2216 22146 2268
rect 22198 2216 22266 2268
rect 22318 2216 22370 2268
rect 20946 2150 22370 2216
rect 20946 2098 22020 2150
rect 22072 2098 22146 2150
rect 22198 2098 22266 2150
rect 22318 2098 22370 2150
rect 20946 2050 22370 2098
rect 463 1288 863 1349
rect 463 1236 514 1288
rect 566 1236 636 1288
rect 688 1236 762 1288
rect 814 1236 863 1288
rect 463 1141 863 1236
rect 463 1089 514 1141
rect 566 1089 636 1141
rect 688 1089 762 1141
rect 814 1089 863 1141
rect 463 1004 863 1089
rect 463 952 514 1004
rect 566 952 636 1004
rect 688 952 762 1004
rect 814 952 863 1004
rect 463 890 863 952
rect 463 693 946 730
rect 463 641 513 693
rect 565 641 639 693
rect 691 641 759 693
rect 811 641 946 693
rect 463 575 946 641
rect 463 523 513 575
rect 565 523 639 575
rect 691 523 759 575
rect 811 523 946 575
rect 463 475 946 523
rect 20946 582 21428 619
rect 20946 530 21078 582
rect 21130 530 21204 582
rect 21256 530 21324 582
rect 21376 530 21428 582
rect 20946 464 21428 530
rect 20946 412 21078 464
rect 21130 412 21204 464
rect 21256 412 21324 464
rect 21376 412 21428 464
rect 20946 364 21428 412
<< via1 >>
rect 513 75431 565 75440
rect 513 75397 522 75431
rect 522 75397 556 75431
rect 556 75397 565 75431
rect 513 75388 565 75397
rect 639 75431 691 75440
rect 639 75397 648 75431
rect 648 75397 682 75431
rect 682 75397 691 75431
rect 639 75388 691 75397
rect 759 75431 811 75440
rect 759 75397 768 75431
rect 768 75397 802 75431
rect 802 75397 811 75431
rect 759 75388 811 75397
rect 513 75313 565 75322
rect 513 75279 522 75313
rect 522 75279 556 75313
rect 556 75279 565 75313
rect 513 75270 565 75279
rect 639 75313 691 75322
rect 639 75279 648 75313
rect 648 75279 682 75313
rect 682 75279 691 75313
rect 639 75270 691 75279
rect 759 75313 811 75322
rect 759 75279 768 75313
rect 768 75279 802 75313
rect 802 75279 811 75313
rect 759 75270 811 75279
rect 21078 75471 21130 75480
rect 21078 75437 21087 75471
rect 21087 75437 21121 75471
rect 21121 75437 21130 75471
rect 21078 75428 21130 75437
rect 21204 75471 21256 75480
rect 21204 75437 21213 75471
rect 21213 75437 21247 75471
rect 21247 75437 21256 75471
rect 21204 75428 21256 75437
rect 21324 75471 21376 75480
rect 21324 75437 21333 75471
rect 21333 75437 21367 75471
rect 21367 75437 21376 75471
rect 21324 75428 21376 75437
rect 21078 75353 21130 75362
rect 21078 75319 21087 75353
rect 21087 75319 21121 75353
rect 21121 75319 21130 75353
rect 21078 75310 21130 75319
rect 21204 75353 21256 75362
rect 21204 75319 21213 75353
rect 21213 75319 21247 75353
rect 21247 75319 21256 75353
rect 21204 75310 21256 75319
rect 21324 75353 21376 75362
rect 21324 75319 21333 75353
rect 21333 75319 21367 75353
rect 21367 75319 21376 75353
rect 21324 75310 21376 75319
rect 514 75039 566 75048
rect 514 75005 523 75039
rect 523 75005 557 75039
rect 557 75005 566 75039
rect 514 74996 566 75005
rect 636 75039 688 75048
rect 636 75005 645 75039
rect 645 75005 679 75039
rect 679 75005 688 75039
rect 636 74996 688 75005
rect 762 75039 814 75048
rect 762 75005 771 75039
rect 771 75005 805 75039
rect 805 75005 814 75039
rect 762 74996 814 75005
rect 514 74892 566 74901
rect 514 74858 523 74892
rect 523 74858 557 74892
rect 557 74858 566 74892
rect 514 74849 566 74858
rect 636 74892 688 74901
rect 636 74858 645 74892
rect 645 74858 679 74892
rect 679 74858 688 74892
rect 636 74849 688 74858
rect 762 74892 814 74901
rect 762 74858 771 74892
rect 771 74858 805 74892
rect 805 74858 814 74892
rect 762 74849 814 74858
rect 514 74755 566 74764
rect 514 74721 523 74755
rect 523 74721 557 74755
rect 557 74721 566 74755
rect 514 74712 566 74721
rect 636 74755 688 74764
rect 636 74721 645 74755
rect 645 74721 679 74755
rect 679 74721 688 74755
rect 636 74712 688 74721
rect 762 74755 814 74764
rect 762 74721 771 74755
rect 771 74721 805 74755
rect 805 74721 814 74755
rect 762 74712 814 74721
rect 22020 74050 22072 74059
rect 22020 74016 22029 74050
rect 22029 74016 22063 74050
rect 22063 74016 22072 74050
rect 22020 74007 22072 74016
rect 22146 74050 22198 74059
rect 22146 74016 22155 74050
rect 22155 74016 22189 74050
rect 22189 74016 22198 74050
rect 22146 74007 22198 74016
rect 22266 74050 22318 74059
rect 22266 74016 22275 74050
rect 22275 74016 22309 74050
rect 22309 74016 22318 74050
rect 22266 74007 22318 74016
rect 22020 73932 22072 73941
rect 22020 73898 22029 73932
rect 22029 73898 22063 73932
rect 22063 73898 22072 73932
rect 22020 73889 22072 73898
rect 22146 73932 22198 73941
rect 22146 73898 22155 73932
rect 22155 73898 22189 73932
rect 22189 73898 22198 73932
rect 22146 73889 22198 73898
rect 22266 73932 22318 73941
rect 22266 73898 22275 73932
rect 22275 73898 22309 73932
rect 22309 73898 22318 73932
rect 22266 73889 22318 73898
rect 514 73279 566 73288
rect 514 73245 523 73279
rect 523 73245 557 73279
rect 557 73245 566 73279
rect 514 73236 566 73245
rect 636 73279 688 73288
rect 636 73245 645 73279
rect 645 73245 679 73279
rect 679 73245 688 73279
rect 636 73236 688 73245
rect 762 73279 814 73288
rect 762 73245 771 73279
rect 771 73245 805 73279
rect 805 73245 814 73279
rect 762 73236 814 73245
rect 514 73132 566 73141
rect 514 73098 523 73132
rect 523 73098 557 73132
rect 557 73098 566 73132
rect 514 73089 566 73098
rect 636 73132 688 73141
rect 636 73098 645 73132
rect 645 73098 679 73132
rect 679 73098 688 73132
rect 636 73089 688 73098
rect 762 73132 814 73141
rect 762 73098 771 73132
rect 771 73098 805 73132
rect 805 73098 814 73132
rect 762 73089 814 73098
rect 514 72995 566 73004
rect 514 72961 523 72995
rect 523 72961 557 72995
rect 557 72961 566 72995
rect 514 72952 566 72961
rect 636 72995 688 73004
rect 636 72961 645 72995
rect 645 72961 679 72995
rect 679 72961 688 72995
rect 636 72952 688 72961
rect 762 72995 814 73004
rect 762 72961 771 72995
rect 771 72961 805 72995
rect 805 72961 814 72995
rect 762 72952 814 72961
rect 513 72758 565 72767
rect 513 72724 522 72758
rect 522 72724 556 72758
rect 556 72724 565 72758
rect 513 72715 565 72724
rect 639 72758 691 72767
rect 639 72724 648 72758
rect 648 72724 682 72758
rect 682 72724 691 72758
rect 639 72715 691 72724
rect 759 72758 811 72767
rect 759 72724 768 72758
rect 768 72724 802 72758
rect 802 72724 811 72758
rect 759 72715 811 72724
rect 513 72640 565 72649
rect 513 72606 522 72640
rect 522 72606 556 72640
rect 556 72606 565 72640
rect 513 72597 565 72606
rect 639 72640 691 72649
rect 639 72606 648 72640
rect 648 72606 682 72640
rect 682 72606 691 72640
rect 639 72597 691 72606
rect 759 72640 811 72649
rect 759 72606 768 72640
rect 768 72606 802 72640
rect 802 72606 811 72640
rect 759 72597 811 72606
rect 21078 72674 21130 72683
rect 21078 72640 21087 72674
rect 21087 72640 21121 72674
rect 21121 72640 21130 72674
rect 21078 72631 21130 72640
rect 21204 72674 21256 72683
rect 21204 72640 21213 72674
rect 21213 72640 21247 72674
rect 21247 72640 21256 72674
rect 21204 72631 21256 72640
rect 21324 72674 21376 72683
rect 21324 72640 21333 72674
rect 21333 72640 21367 72674
rect 21367 72640 21376 72674
rect 21324 72631 21376 72640
rect 21078 72556 21130 72565
rect 21078 72522 21087 72556
rect 21087 72522 21121 72556
rect 21121 72522 21130 72556
rect 21078 72513 21130 72522
rect 21204 72556 21256 72565
rect 21204 72522 21213 72556
rect 21213 72522 21247 72556
rect 21247 72522 21256 72556
rect 21204 72513 21256 72522
rect 21324 72556 21376 72565
rect 21324 72522 21333 72556
rect 21333 72522 21367 72556
rect 21367 72522 21376 72556
rect 21324 72513 21376 72522
rect 513 71431 565 71440
rect 513 71397 522 71431
rect 522 71397 556 71431
rect 556 71397 565 71431
rect 513 71388 565 71397
rect 639 71431 691 71440
rect 639 71397 648 71431
rect 648 71397 682 71431
rect 682 71397 691 71431
rect 639 71388 691 71397
rect 759 71431 811 71440
rect 759 71397 768 71431
rect 768 71397 802 71431
rect 802 71397 811 71431
rect 759 71388 811 71397
rect 513 71313 565 71322
rect 513 71279 522 71313
rect 522 71279 556 71313
rect 556 71279 565 71313
rect 513 71270 565 71279
rect 639 71313 691 71322
rect 639 71279 648 71313
rect 648 71279 682 71313
rect 682 71279 691 71313
rect 639 71270 691 71279
rect 759 71313 811 71322
rect 759 71279 768 71313
rect 768 71279 802 71313
rect 802 71279 811 71313
rect 759 71270 811 71279
rect 21078 71471 21130 71480
rect 21078 71437 21087 71471
rect 21087 71437 21121 71471
rect 21121 71437 21130 71471
rect 21078 71428 21130 71437
rect 21204 71471 21256 71480
rect 21204 71437 21213 71471
rect 21213 71437 21247 71471
rect 21247 71437 21256 71471
rect 21204 71428 21256 71437
rect 21324 71471 21376 71480
rect 21324 71437 21333 71471
rect 21333 71437 21367 71471
rect 21367 71437 21376 71471
rect 21324 71428 21376 71437
rect 21078 71353 21130 71362
rect 21078 71319 21087 71353
rect 21087 71319 21121 71353
rect 21121 71319 21130 71353
rect 21078 71310 21130 71319
rect 21204 71353 21256 71362
rect 21204 71319 21213 71353
rect 21213 71319 21247 71353
rect 21247 71319 21256 71353
rect 21204 71310 21256 71319
rect 21324 71353 21376 71362
rect 21324 71319 21333 71353
rect 21333 71319 21367 71353
rect 21367 71319 21376 71353
rect 21324 71310 21376 71319
rect 514 71039 566 71048
rect 514 71005 523 71039
rect 523 71005 557 71039
rect 557 71005 566 71039
rect 514 70996 566 71005
rect 636 71039 688 71048
rect 636 71005 645 71039
rect 645 71005 679 71039
rect 679 71005 688 71039
rect 636 70996 688 71005
rect 762 71039 814 71048
rect 762 71005 771 71039
rect 771 71005 805 71039
rect 805 71005 814 71039
rect 762 70996 814 71005
rect 514 70892 566 70901
rect 514 70858 523 70892
rect 523 70858 557 70892
rect 557 70858 566 70892
rect 514 70849 566 70858
rect 636 70892 688 70901
rect 636 70858 645 70892
rect 645 70858 679 70892
rect 679 70858 688 70892
rect 636 70849 688 70858
rect 762 70892 814 70901
rect 762 70858 771 70892
rect 771 70858 805 70892
rect 805 70858 814 70892
rect 762 70849 814 70858
rect 514 70755 566 70764
rect 514 70721 523 70755
rect 523 70721 557 70755
rect 557 70721 566 70755
rect 514 70712 566 70721
rect 636 70755 688 70764
rect 636 70721 645 70755
rect 645 70721 679 70755
rect 679 70721 688 70755
rect 636 70712 688 70721
rect 762 70755 814 70764
rect 762 70721 771 70755
rect 771 70721 805 70755
rect 805 70721 814 70755
rect 762 70712 814 70721
rect 22020 70050 22072 70059
rect 22020 70016 22029 70050
rect 22029 70016 22063 70050
rect 22063 70016 22072 70050
rect 22020 70007 22072 70016
rect 22146 70050 22198 70059
rect 22146 70016 22155 70050
rect 22155 70016 22189 70050
rect 22189 70016 22198 70050
rect 22146 70007 22198 70016
rect 22266 70050 22318 70059
rect 22266 70016 22275 70050
rect 22275 70016 22309 70050
rect 22309 70016 22318 70050
rect 22266 70007 22318 70016
rect 22020 69932 22072 69941
rect 22020 69898 22029 69932
rect 22029 69898 22063 69932
rect 22063 69898 22072 69932
rect 22020 69889 22072 69898
rect 22146 69932 22198 69941
rect 22146 69898 22155 69932
rect 22155 69898 22189 69932
rect 22189 69898 22198 69932
rect 22146 69889 22198 69898
rect 22266 69932 22318 69941
rect 22266 69898 22275 69932
rect 22275 69898 22309 69932
rect 22309 69898 22318 69932
rect 22266 69889 22318 69898
rect 514 69279 566 69288
rect 514 69245 523 69279
rect 523 69245 557 69279
rect 557 69245 566 69279
rect 514 69236 566 69245
rect 636 69279 688 69288
rect 636 69245 645 69279
rect 645 69245 679 69279
rect 679 69245 688 69279
rect 636 69236 688 69245
rect 762 69279 814 69288
rect 762 69245 771 69279
rect 771 69245 805 69279
rect 805 69245 814 69279
rect 762 69236 814 69245
rect 514 69132 566 69141
rect 514 69098 523 69132
rect 523 69098 557 69132
rect 557 69098 566 69132
rect 514 69089 566 69098
rect 636 69132 688 69141
rect 636 69098 645 69132
rect 645 69098 679 69132
rect 679 69098 688 69132
rect 636 69089 688 69098
rect 762 69132 814 69141
rect 762 69098 771 69132
rect 771 69098 805 69132
rect 805 69098 814 69132
rect 762 69089 814 69098
rect 514 68995 566 69004
rect 514 68961 523 68995
rect 523 68961 557 68995
rect 557 68961 566 68995
rect 514 68952 566 68961
rect 636 68995 688 69004
rect 636 68961 645 68995
rect 645 68961 679 68995
rect 679 68961 688 68995
rect 636 68952 688 68961
rect 762 68995 814 69004
rect 762 68961 771 68995
rect 771 68961 805 68995
rect 805 68961 814 68995
rect 762 68952 814 68961
rect 513 68758 565 68767
rect 513 68724 522 68758
rect 522 68724 556 68758
rect 556 68724 565 68758
rect 513 68715 565 68724
rect 639 68758 691 68767
rect 639 68724 648 68758
rect 648 68724 682 68758
rect 682 68724 691 68758
rect 639 68715 691 68724
rect 759 68758 811 68767
rect 759 68724 768 68758
rect 768 68724 802 68758
rect 802 68724 811 68758
rect 759 68715 811 68724
rect 513 68640 565 68649
rect 513 68606 522 68640
rect 522 68606 556 68640
rect 556 68606 565 68640
rect 513 68597 565 68606
rect 639 68640 691 68649
rect 639 68606 648 68640
rect 648 68606 682 68640
rect 682 68606 691 68640
rect 639 68597 691 68606
rect 759 68640 811 68649
rect 759 68606 768 68640
rect 768 68606 802 68640
rect 802 68606 811 68640
rect 759 68597 811 68606
rect 21078 68674 21130 68683
rect 21078 68640 21087 68674
rect 21087 68640 21121 68674
rect 21121 68640 21130 68674
rect 21078 68631 21130 68640
rect 21204 68674 21256 68683
rect 21204 68640 21213 68674
rect 21213 68640 21247 68674
rect 21247 68640 21256 68674
rect 21204 68631 21256 68640
rect 21324 68674 21376 68683
rect 21324 68640 21333 68674
rect 21333 68640 21367 68674
rect 21367 68640 21376 68674
rect 21324 68631 21376 68640
rect 21078 68556 21130 68565
rect 21078 68522 21087 68556
rect 21087 68522 21121 68556
rect 21121 68522 21130 68556
rect 21078 68513 21130 68522
rect 21204 68556 21256 68565
rect 21204 68522 21213 68556
rect 21213 68522 21247 68556
rect 21247 68522 21256 68556
rect 21204 68513 21256 68522
rect 21324 68556 21376 68565
rect 21324 68522 21333 68556
rect 21333 68522 21367 68556
rect 21367 68522 21376 68556
rect 21324 68513 21376 68522
rect 513 67429 565 67438
rect 513 67395 522 67429
rect 522 67395 556 67429
rect 556 67395 565 67429
rect 513 67386 565 67395
rect 639 67429 691 67438
rect 639 67395 648 67429
rect 648 67395 682 67429
rect 682 67395 691 67429
rect 639 67386 691 67395
rect 759 67429 811 67438
rect 759 67395 768 67429
rect 768 67395 802 67429
rect 802 67395 811 67429
rect 759 67386 811 67395
rect 513 67311 565 67320
rect 513 67277 522 67311
rect 522 67277 556 67311
rect 556 67277 565 67311
rect 513 67268 565 67277
rect 639 67311 691 67320
rect 639 67277 648 67311
rect 648 67277 682 67311
rect 682 67277 691 67311
rect 639 67268 691 67277
rect 759 67311 811 67320
rect 759 67277 768 67311
rect 768 67277 802 67311
rect 802 67277 811 67311
rect 759 67268 811 67277
rect 21078 67471 21130 67480
rect 21078 67437 21087 67471
rect 21087 67437 21121 67471
rect 21121 67437 21130 67471
rect 21078 67428 21130 67437
rect 21204 67471 21256 67480
rect 21204 67437 21213 67471
rect 21213 67437 21247 67471
rect 21247 67437 21256 67471
rect 21204 67428 21256 67437
rect 21324 67471 21376 67480
rect 21324 67437 21333 67471
rect 21333 67437 21367 67471
rect 21367 67437 21376 67471
rect 21324 67428 21376 67437
rect 21078 67353 21130 67362
rect 21078 67319 21087 67353
rect 21087 67319 21121 67353
rect 21121 67319 21130 67353
rect 21078 67310 21130 67319
rect 21204 67353 21256 67362
rect 21204 67319 21213 67353
rect 21213 67319 21247 67353
rect 21247 67319 21256 67353
rect 21204 67310 21256 67319
rect 21324 67353 21376 67362
rect 21324 67319 21333 67353
rect 21333 67319 21367 67353
rect 21367 67319 21376 67353
rect 21324 67310 21376 67319
rect 514 67039 566 67048
rect 514 67005 523 67039
rect 523 67005 557 67039
rect 557 67005 566 67039
rect 514 66996 566 67005
rect 636 67039 688 67048
rect 636 67005 645 67039
rect 645 67005 679 67039
rect 679 67005 688 67039
rect 636 66996 688 67005
rect 762 67039 814 67048
rect 762 67005 771 67039
rect 771 67005 805 67039
rect 805 67005 814 67039
rect 762 66996 814 67005
rect 514 66892 566 66901
rect 514 66858 523 66892
rect 523 66858 557 66892
rect 557 66858 566 66892
rect 514 66849 566 66858
rect 636 66892 688 66901
rect 636 66858 645 66892
rect 645 66858 679 66892
rect 679 66858 688 66892
rect 636 66849 688 66858
rect 762 66892 814 66901
rect 762 66858 771 66892
rect 771 66858 805 66892
rect 805 66858 814 66892
rect 762 66849 814 66858
rect 514 66755 566 66764
rect 514 66721 523 66755
rect 523 66721 557 66755
rect 557 66721 566 66755
rect 514 66712 566 66721
rect 636 66755 688 66764
rect 636 66721 645 66755
rect 645 66721 679 66755
rect 679 66721 688 66755
rect 636 66712 688 66721
rect 762 66755 814 66764
rect 762 66721 771 66755
rect 771 66721 805 66755
rect 805 66721 814 66755
rect 762 66712 814 66721
rect 22020 66037 22072 66046
rect 22020 66003 22029 66037
rect 22029 66003 22063 66037
rect 22063 66003 22072 66037
rect 22020 65994 22072 66003
rect 22146 66037 22198 66046
rect 22146 66003 22155 66037
rect 22155 66003 22189 66037
rect 22189 66003 22198 66037
rect 22146 65994 22198 66003
rect 22266 66037 22318 66046
rect 22266 66003 22275 66037
rect 22275 66003 22309 66037
rect 22309 66003 22318 66037
rect 22266 65994 22318 66003
rect 22020 65919 22072 65928
rect 22020 65885 22029 65919
rect 22029 65885 22063 65919
rect 22063 65885 22072 65919
rect 22020 65876 22072 65885
rect 22146 65919 22198 65928
rect 22146 65885 22155 65919
rect 22155 65885 22189 65919
rect 22189 65885 22198 65919
rect 22146 65876 22198 65885
rect 22266 65919 22318 65928
rect 22266 65885 22275 65919
rect 22275 65885 22309 65919
rect 22309 65885 22318 65919
rect 22266 65876 22318 65885
rect 514 65280 566 65289
rect 514 65246 523 65280
rect 523 65246 557 65280
rect 557 65246 566 65280
rect 514 65237 566 65246
rect 636 65280 688 65289
rect 636 65246 645 65280
rect 645 65246 679 65280
rect 679 65246 688 65280
rect 636 65237 688 65246
rect 762 65280 814 65289
rect 762 65246 771 65280
rect 771 65246 805 65280
rect 805 65246 814 65280
rect 762 65237 814 65246
rect 514 65133 566 65142
rect 514 65099 523 65133
rect 523 65099 557 65133
rect 557 65099 566 65133
rect 514 65090 566 65099
rect 636 65133 688 65142
rect 636 65099 645 65133
rect 645 65099 679 65133
rect 679 65099 688 65133
rect 636 65090 688 65099
rect 762 65133 814 65142
rect 762 65099 771 65133
rect 771 65099 805 65133
rect 805 65099 814 65133
rect 762 65090 814 65099
rect 514 64996 566 65005
rect 514 64962 523 64996
rect 523 64962 557 64996
rect 557 64962 566 64996
rect 514 64953 566 64962
rect 636 64996 688 65005
rect 636 64962 645 64996
rect 645 64962 679 64996
rect 679 64962 688 64996
rect 636 64953 688 64962
rect 762 64996 814 65005
rect 762 64962 771 64996
rect 771 64962 805 64996
rect 805 64962 814 64996
rect 762 64953 814 64962
rect 513 64689 565 64698
rect 513 64655 522 64689
rect 522 64655 556 64689
rect 556 64655 565 64689
rect 513 64646 565 64655
rect 639 64689 691 64698
rect 639 64655 648 64689
rect 648 64655 682 64689
rect 682 64655 691 64689
rect 639 64646 691 64655
rect 759 64689 811 64698
rect 759 64655 768 64689
rect 768 64655 802 64689
rect 802 64655 811 64689
rect 759 64646 811 64655
rect 513 64571 565 64580
rect 513 64537 522 64571
rect 522 64537 556 64571
rect 556 64537 565 64571
rect 513 64528 565 64537
rect 639 64571 691 64580
rect 639 64537 648 64571
rect 648 64537 682 64571
rect 682 64537 691 64571
rect 639 64528 691 64537
rect 759 64571 811 64580
rect 759 64537 768 64571
rect 768 64537 802 64571
rect 802 64537 811 64571
rect 759 64528 811 64537
rect 21078 64674 21130 64683
rect 21078 64640 21087 64674
rect 21087 64640 21121 64674
rect 21121 64640 21130 64674
rect 21078 64631 21130 64640
rect 21204 64674 21256 64683
rect 21204 64640 21213 64674
rect 21213 64640 21247 64674
rect 21247 64640 21256 64674
rect 21204 64631 21256 64640
rect 21324 64674 21376 64683
rect 21324 64640 21333 64674
rect 21333 64640 21367 64674
rect 21367 64640 21376 64674
rect 21324 64631 21376 64640
rect 21078 64556 21130 64565
rect 21078 64522 21087 64556
rect 21087 64522 21121 64556
rect 21121 64522 21130 64556
rect 21078 64513 21130 64522
rect 21204 64556 21256 64565
rect 21204 64522 21213 64556
rect 21213 64522 21247 64556
rect 21247 64522 21256 64556
rect 21204 64513 21256 64522
rect 21324 64556 21376 64565
rect 21324 64522 21333 64556
rect 21333 64522 21367 64556
rect 21367 64522 21376 64556
rect 21324 64513 21376 64522
rect 513 63511 565 63520
rect 513 63477 522 63511
rect 522 63477 556 63511
rect 556 63477 565 63511
rect 513 63468 565 63477
rect 639 63511 691 63520
rect 639 63477 648 63511
rect 648 63477 682 63511
rect 682 63477 691 63511
rect 639 63468 691 63477
rect 759 63511 811 63520
rect 759 63477 768 63511
rect 768 63477 802 63511
rect 802 63477 811 63511
rect 759 63468 811 63477
rect 513 63393 565 63402
rect 513 63359 522 63393
rect 522 63359 556 63393
rect 556 63359 565 63393
rect 513 63350 565 63359
rect 639 63393 691 63402
rect 639 63359 648 63393
rect 648 63359 682 63393
rect 682 63359 691 63393
rect 639 63350 691 63359
rect 759 63393 811 63402
rect 759 63359 768 63393
rect 768 63359 802 63393
rect 802 63359 811 63393
rect 759 63350 811 63359
rect 21078 63471 21130 63480
rect 21078 63437 21087 63471
rect 21087 63437 21121 63471
rect 21121 63437 21130 63471
rect 21078 63428 21130 63437
rect 21204 63471 21256 63480
rect 21204 63437 21213 63471
rect 21213 63437 21247 63471
rect 21247 63437 21256 63471
rect 21204 63428 21256 63437
rect 21324 63471 21376 63480
rect 21324 63437 21333 63471
rect 21333 63437 21367 63471
rect 21367 63437 21376 63471
rect 21324 63428 21376 63437
rect 21078 63353 21130 63362
rect 21078 63319 21087 63353
rect 21087 63319 21121 63353
rect 21121 63319 21130 63353
rect 21078 63310 21130 63319
rect 21204 63353 21256 63362
rect 21204 63319 21213 63353
rect 21213 63319 21247 63353
rect 21247 63319 21256 63353
rect 21204 63310 21256 63319
rect 21324 63353 21376 63362
rect 21324 63319 21333 63353
rect 21333 63319 21367 63353
rect 21367 63319 21376 63353
rect 21324 63310 21376 63319
rect 514 63039 566 63048
rect 514 63005 523 63039
rect 523 63005 557 63039
rect 557 63005 566 63039
rect 514 62996 566 63005
rect 636 63039 688 63048
rect 636 63005 645 63039
rect 645 63005 679 63039
rect 679 63005 688 63039
rect 636 62996 688 63005
rect 762 63039 814 63048
rect 762 63005 771 63039
rect 771 63005 805 63039
rect 805 63005 814 63039
rect 762 62996 814 63005
rect 514 62892 566 62901
rect 514 62858 523 62892
rect 523 62858 557 62892
rect 557 62858 566 62892
rect 514 62849 566 62858
rect 636 62892 688 62901
rect 636 62858 645 62892
rect 645 62858 679 62892
rect 679 62858 688 62892
rect 636 62849 688 62858
rect 762 62892 814 62901
rect 762 62858 771 62892
rect 771 62858 805 62892
rect 805 62858 814 62892
rect 762 62849 814 62858
rect 514 62755 566 62764
rect 514 62721 523 62755
rect 523 62721 557 62755
rect 557 62721 566 62755
rect 514 62712 566 62721
rect 636 62755 688 62764
rect 636 62721 645 62755
rect 645 62721 679 62755
rect 679 62721 688 62755
rect 636 62712 688 62721
rect 762 62755 814 62764
rect 762 62721 771 62755
rect 771 62721 805 62755
rect 805 62721 814 62755
rect 762 62712 814 62721
rect 22020 62036 22072 62045
rect 22020 62002 22029 62036
rect 22029 62002 22063 62036
rect 22063 62002 22072 62036
rect 22020 61993 22072 62002
rect 22146 62036 22198 62045
rect 22146 62002 22155 62036
rect 22155 62002 22189 62036
rect 22189 62002 22198 62036
rect 22146 61993 22198 62002
rect 22266 62036 22318 62045
rect 22266 62002 22275 62036
rect 22275 62002 22309 62036
rect 22309 62002 22318 62036
rect 22266 61993 22318 62002
rect 22020 61918 22072 61927
rect 22020 61884 22029 61918
rect 22029 61884 22063 61918
rect 22063 61884 22072 61918
rect 22020 61875 22072 61884
rect 22146 61918 22198 61927
rect 22146 61884 22155 61918
rect 22155 61884 22189 61918
rect 22189 61884 22198 61918
rect 22146 61875 22198 61884
rect 22266 61918 22318 61927
rect 22266 61884 22275 61918
rect 22275 61884 22309 61918
rect 22309 61884 22318 61918
rect 22266 61875 22318 61884
rect 514 61280 566 61289
rect 514 61246 523 61280
rect 523 61246 557 61280
rect 557 61246 566 61280
rect 514 61237 566 61246
rect 636 61280 688 61289
rect 636 61246 645 61280
rect 645 61246 679 61280
rect 679 61246 688 61280
rect 636 61237 688 61246
rect 762 61280 814 61289
rect 762 61246 771 61280
rect 771 61246 805 61280
rect 805 61246 814 61280
rect 762 61237 814 61246
rect 514 61133 566 61142
rect 514 61099 523 61133
rect 523 61099 557 61133
rect 557 61099 566 61133
rect 514 61090 566 61099
rect 636 61133 688 61142
rect 636 61099 645 61133
rect 645 61099 679 61133
rect 679 61099 688 61133
rect 636 61090 688 61099
rect 762 61133 814 61142
rect 762 61099 771 61133
rect 771 61099 805 61133
rect 805 61099 814 61133
rect 762 61090 814 61099
rect 514 60996 566 61005
rect 514 60962 523 60996
rect 523 60962 557 60996
rect 557 60962 566 60996
rect 514 60953 566 60962
rect 636 60996 688 61005
rect 636 60962 645 60996
rect 645 60962 679 60996
rect 679 60962 688 60996
rect 636 60953 688 60962
rect 762 60996 814 61005
rect 762 60962 771 60996
rect 771 60962 805 60996
rect 805 60962 814 60996
rect 762 60953 814 60962
rect 513 60663 565 60672
rect 513 60629 522 60663
rect 522 60629 556 60663
rect 556 60629 565 60663
rect 513 60620 565 60629
rect 639 60663 691 60672
rect 639 60629 648 60663
rect 648 60629 682 60663
rect 682 60629 691 60663
rect 639 60620 691 60629
rect 759 60663 811 60672
rect 759 60629 768 60663
rect 768 60629 802 60663
rect 802 60629 811 60663
rect 759 60620 811 60629
rect 513 60545 565 60554
rect 513 60511 522 60545
rect 522 60511 556 60545
rect 556 60511 565 60545
rect 513 60502 565 60511
rect 639 60545 691 60554
rect 639 60511 648 60545
rect 648 60511 682 60545
rect 682 60511 691 60545
rect 639 60502 691 60511
rect 759 60545 811 60554
rect 759 60511 768 60545
rect 768 60511 802 60545
rect 802 60511 811 60545
rect 759 60502 811 60511
rect 21078 60674 21130 60683
rect 21078 60640 21087 60674
rect 21087 60640 21121 60674
rect 21121 60640 21130 60674
rect 21078 60631 21130 60640
rect 21204 60674 21256 60683
rect 21204 60640 21213 60674
rect 21213 60640 21247 60674
rect 21247 60640 21256 60674
rect 21204 60631 21256 60640
rect 21324 60674 21376 60683
rect 21324 60640 21333 60674
rect 21333 60640 21367 60674
rect 21367 60640 21376 60674
rect 21324 60631 21376 60640
rect 21078 60556 21130 60565
rect 21078 60522 21087 60556
rect 21087 60522 21121 60556
rect 21121 60522 21130 60556
rect 21078 60513 21130 60522
rect 21204 60556 21256 60565
rect 21204 60522 21213 60556
rect 21213 60522 21247 60556
rect 21247 60522 21256 60556
rect 21204 60513 21256 60522
rect 21324 60556 21376 60565
rect 21324 60522 21333 60556
rect 21333 60522 21367 60556
rect 21367 60522 21376 60556
rect 21324 60513 21376 60522
rect 513 59460 565 59469
rect 513 59426 522 59460
rect 522 59426 556 59460
rect 556 59426 565 59460
rect 513 59417 565 59426
rect 639 59460 691 59469
rect 639 59426 648 59460
rect 648 59426 682 59460
rect 682 59426 691 59460
rect 639 59417 691 59426
rect 759 59460 811 59469
rect 759 59426 768 59460
rect 768 59426 802 59460
rect 802 59426 811 59460
rect 759 59417 811 59426
rect 513 59342 565 59351
rect 513 59308 522 59342
rect 522 59308 556 59342
rect 556 59308 565 59342
rect 513 59299 565 59308
rect 639 59342 691 59351
rect 639 59308 648 59342
rect 648 59308 682 59342
rect 682 59308 691 59342
rect 639 59299 691 59308
rect 759 59342 811 59351
rect 759 59308 768 59342
rect 768 59308 802 59342
rect 802 59308 811 59342
rect 759 59299 811 59308
rect 21078 59525 21130 59534
rect 21078 59491 21087 59525
rect 21087 59491 21121 59525
rect 21121 59491 21130 59525
rect 21078 59482 21130 59491
rect 21204 59525 21256 59534
rect 21204 59491 21213 59525
rect 21213 59491 21247 59525
rect 21247 59491 21256 59525
rect 21204 59482 21256 59491
rect 21324 59525 21376 59534
rect 21324 59491 21333 59525
rect 21333 59491 21367 59525
rect 21367 59491 21376 59525
rect 21324 59482 21376 59491
rect 21078 59407 21130 59416
rect 21078 59373 21087 59407
rect 21087 59373 21121 59407
rect 21121 59373 21130 59407
rect 21078 59364 21130 59373
rect 21204 59407 21256 59416
rect 21204 59373 21213 59407
rect 21213 59373 21247 59407
rect 21247 59373 21256 59407
rect 21204 59364 21256 59373
rect 21324 59407 21376 59416
rect 21324 59373 21333 59407
rect 21333 59373 21367 59407
rect 21367 59373 21376 59407
rect 21324 59364 21376 59373
rect 514 59039 566 59048
rect 514 59005 523 59039
rect 523 59005 557 59039
rect 557 59005 566 59039
rect 514 58996 566 59005
rect 636 59039 688 59048
rect 636 59005 645 59039
rect 645 59005 679 59039
rect 679 59005 688 59039
rect 636 58996 688 59005
rect 762 59039 814 59048
rect 762 59005 771 59039
rect 771 59005 805 59039
rect 805 59005 814 59039
rect 762 58996 814 59005
rect 514 58892 566 58901
rect 514 58858 523 58892
rect 523 58858 557 58892
rect 557 58858 566 58892
rect 514 58849 566 58858
rect 636 58892 688 58901
rect 636 58858 645 58892
rect 645 58858 679 58892
rect 679 58858 688 58892
rect 636 58849 688 58858
rect 762 58892 814 58901
rect 762 58858 771 58892
rect 771 58858 805 58892
rect 805 58858 814 58892
rect 762 58849 814 58858
rect 514 58755 566 58764
rect 514 58721 523 58755
rect 523 58721 557 58755
rect 557 58721 566 58755
rect 514 58712 566 58721
rect 636 58755 688 58764
rect 636 58721 645 58755
rect 645 58721 679 58755
rect 679 58721 688 58755
rect 636 58712 688 58721
rect 762 58755 814 58764
rect 762 58721 771 58755
rect 771 58721 805 58755
rect 805 58721 814 58755
rect 762 58712 814 58721
rect 22020 58075 22072 58084
rect 22020 58041 22029 58075
rect 22029 58041 22063 58075
rect 22063 58041 22072 58075
rect 22020 58032 22072 58041
rect 22146 58075 22198 58084
rect 22146 58041 22155 58075
rect 22155 58041 22189 58075
rect 22189 58041 22198 58075
rect 22146 58032 22198 58041
rect 22266 58075 22318 58084
rect 22266 58041 22275 58075
rect 22275 58041 22309 58075
rect 22309 58041 22318 58075
rect 22266 58032 22318 58041
rect 22020 57957 22072 57966
rect 22020 57923 22029 57957
rect 22029 57923 22063 57957
rect 22063 57923 22072 57957
rect 22020 57914 22072 57923
rect 22146 57957 22198 57966
rect 22146 57923 22155 57957
rect 22155 57923 22189 57957
rect 22189 57923 22198 57957
rect 22146 57914 22198 57923
rect 22266 57957 22318 57966
rect 22266 57923 22275 57957
rect 22275 57923 22309 57957
rect 22309 57923 22318 57957
rect 22266 57914 22318 57923
rect 514 57278 566 57287
rect 514 57244 523 57278
rect 523 57244 557 57278
rect 557 57244 566 57278
rect 514 57235 566 57244
rect 636 57278 688 57287
rect 636 57244 645 57278
rect 645 57244 679 57278
rect 679 57244 688 57278
rect 636 57235 688 57244
rect 762 57278 814 57287
rect 762 57244 771 57278
rect 771 57244 805 57278
rect 805 57244 814 57278
rect 762 57235 814 57244
rect 514 57131 566 57140
rect 514 57097 523 57131
rect 523 57097 557 57131
rect 557 57097 566 57131
rect 514 57088 566 57097
rect 636 57131 688 57140
rect 636 57097 645 57131
rect 645 57097 679 57131
rect 679 57097 688 57131
rect 636 57088 688 57097
rect 762 57131 814 57140
rect 762 57097 771 57131
rect 771 57097 805 57131
rect 805 57097 814 57131
rect 762 57088 814 57097
rect 514 56994 566 57003
rect 514 56960 523 56994
rect 523 56960 557 56994
rect 557 56960 566 56994
rect 514 56951 566 56960
rect 636 56994 688 57003
rect 636 56960 645 56994
rect 645 56960 679 56994
rect 679 56960 688 56994
rect 636 56951 688 56960
rect 762 56994 814 57003
rect 762 56960 771 56994
rect 771 56960 805 56994
rect 805 56960 814 56994
rect 762 56951 814 56960
rect 513 56683 565 56692
rect 513 56649 522 56683
rect 522 56649 556 56683
rect 556 56649 565 56683
rect 513 56640 565 56649
rect 639 56683 691 56692
rect 639 56649 648 56683
rect 648 56649 682 56683
rect 682 56649 691 56683
rect 639 56640 691 56649
rect 759 56683 811 56692
rect 759 56649 768 56683
rect 768 56649 802 56683
rect 802 56649 811 56683
rect 759 56640 811 56649
rect 513 56565 565 56574
rect 513 56531 522 56565
rect 522 56531 556 56565
rect 556 56531 565 56565
rect 513 56522 565 56531
rect 639 56565 691 56574
rect 639 56531 648 56565
rect 648 56531 682 56565
rect 682 56531 691 56565
rect 639 56522 691 56531
rect 759 56565 811 56574
rect 759 56531 768 56565
rect 768 56531 802 56565
rect 802 56531 811 56565
rect 759 56522 811 56531
rect 21078 56609 21130 56618
rect 21078 56575 21087 56609
rect 21087 56575 21121 56609
rect 21121 56575 21130 56609
rect 21078 56566 21130 56575
rect 21204 56609 21256 56618
rect 21204 56575 21213 56609
rect 21213 56575 21247 56609
rect 21247 56575 21256 56609
rect 21204 56566 21256 56575
rect 21324 56609 21376 56618
rect 21324 56575 21333 56609
rect 21333 56575 21367 56609
rect 21367 56575 21376 56609
rect 21324 56566 21376 56575
rect 21078 56491 21130 56500
rect 21078 56457 21087 56491
rect 21087 56457 21121 56491
rect 21121 56457 21130 56491
rect 21078 56448 21130 56457
rect 21204 56491 21256 56500
rect 21204 56457 21213 56491
rect 21213 56457 21247 56491
rect 21247 56457 21256 56491
rect 21204 56448 21256 56457
rect 21324 56491 21376 56500
rect 21324 56457 21333 56491
rect 21333 56457 21367 56491
rect 21367 56457 21376 56491
rect 21324 56448 21376 56457
rect 513 55476 565 55485
rect 513 55442 522 55476
rect 522 55442 556 55476
rect 556 55442 565 55476
rect 513 55433 565 55442
rect 639 55476 691 55485
rect 639 55442 648 55476
rect 648 55442 682 55476
rect 682 55442 691 55476
rect 639 55433 691 55442
rect 759 55476 811 55485
rect 759 55442 768 55476
rect 768 55442 802 55476
rect 802 55442 811 55476
rect 759 55433 811 55442
rect 513 55358 565 55367
rect 513 55324 522 55358
rect 522 55324 556 55358
rect 556 55324 565 55358
rect 513 55315 565 55324
rect 639 55358 691 55367
rect 639 55324 648 55358
rect 648 55324 682 55358
rect 682 55324 691 55358
rect 639 55315 691 55324
rect 759 55358 811 55367
rect 759 55324 768 55358
rect 768 55324 802 55358
rect 802 55324 811 55358
rect 759 55315 811 55324
rect 21078 55426 21130 55435
rect 21078 55392 21087 55426
rect 21087 55392 21121 55426
rect 21121 55392 21130 55426
rect 21078 55383 21130 55392
rect 21204 55426 21256 55435
rect 21204 55392 21213 55426
rect 21213 55392 21247 55426
rect 21247 55392 21256 55426
rect 21204 55383 21256 55392
rect 21324 55426 21376 55435
rect 21324 55392 21333 55426
rect 21333 55392 21367 55426
rect 21367 55392 21376 55426
rect 21324 55383 21376 55392
rect 21078 55308 21130 55317
rect 21078 55274 21087 55308
rect 21087 55274 21121 55308
rect 21121 55274 21130 55308
rect 21078 55265 21130 55274
rect 21204 55308 21256 55317
rect 21204 55274 21213 55308
rect 21213 55274 21247 55308
rect 21247 55274 21256 55308
rect 21204 55265 21256 55274
rect 21324 55308 21376 55317
rect 21324 55274 21333 55308
rect 21333 55274 21367 55308
rect 21367 55274 21376 55308
rect 21324 55265 21376 55274
rect 514 55039 566 55048
rect 514 55005 523 55039
rect 523 55005 557 55039
rect 557 55005 566 55039
rect 514 54996 566 55005
rect 636 55039 688 55048
rect 636 55005 645 55039
rect 645 55005 679 55039
rect 679 55005 688 55039
rect 636 54996 688 55005
rect 762 55039 814 55048
rect 762 55005 771 55039
rect 771 55005 805 55039
rect 805 55005 814 55039
rect 762 54996 814 55005
rect 514 54892 566 54901
rect 514 54858 523 54892
rect 523 54858 557 54892
rect 557 54858 566 54892
rect 514 54849 566 54858
rect 636 54892 688 54901
rect 636 54858 645 54892
rect 645 54858 679 54892
rect 679 54858 688 54892
rect 636 54849 688 54858
rect 762 54892 814 54901
rect 762 54858 771 54892
rect 771 54858 805 54892
rect 805 54858 814 54892
rect 762 54849 814 54858
rect 514 54755 566 54764
rect 514 54721 523 54755
rect 523 54721 557 54755
rect 557 54721 566 54755
rect 514 54712 566 54721
rect 636 54755 688 54764
rect 636 54721 645 54755
rect 645 54721 679 54755
rect 679 54721 688 54755
rect 636 54712 688 54721
rect 762 54755 814 54764
rect 762 54721 771 54755
rect 771 54721 805 54755
rect 805 54721 814 54755
rect 762 54712 814 54721
rect 22020 54058 22072 54067
rect 22020 54024 22029 54058
rect 22029 54024 22063 54058
rect 22063 54024 22072 54058
rect 22020 54015 22072 54024
rect 22146 54058 22198 54067
rect 22146 54024 22155 54058
rect 22155 54024 22189 54058
rect 22189 54024 22198 54058
rect 22146 54015 22198 54024
rect 22266 54058 22318 54067
rect 22266 54024 22275 54058
rect 22275 54024 22309 54058
rect 22309 54024 22318 54058
rect 22266 54015 22318 54024
rect 22020 53940 22072 53949
rect 22020 53906 22029 53940
rect 22029 53906 22063 53940
rect 22063 53906 22072 53940
rect 22020 53897 22072 53906
rect 22146 53940 22198 53949
rect 22146 53906 22155 53940
rect 22155 53906 22189 53940
rect 22189 53906 22198 53940
rect 22146 53897 22198 53906
rect 22266 53940 22318 53949
rect 22266 53906 22275 53940
rect 22275 53906 22309 53940
rect 22309 53906 22318 53940
rect 22266 53897 22318 53906
rect 514 53280 566 53289
rect 514 53246 523 53280
rect 523 53246 557 53280
rect 557 53246 566 53280
rect 514 53237 566 53246
rect 636 53280 688 53289
rect 636 53246 645 53280
rect 645 53246 679 53280
rect 679 53246 688 53280
rect 636 53237 688 53246
rect 762 53280 814 53289
rect 762 53246 771 53280
rect 771 53246 805 53280
rect 805 53246 814 53280
rect 762 53237 814 53246
rect 514 53133 566 53142
rect 514 53099 523 53133
rect 523 53099 557 53133
rect 557 53099 566 53133
rect 514 53090 566 53099
rect 636 53133 688 53142
rect 636 53099 645 53133
rect 645 53099 679 53133
rect 679 53099 688 53133
rect 636 53090 688 53099
rect 762 53133 814 53142
rect 762 53099 771 53133
rect 771 53099 805 53133
rect 805 53099 814 53133
rect 762 53090 814 53099
rect 514 52996 566 53005
rect 514 52962 523 52996
rect 523 52962 557 52996
rect 557 52962 566 52996
rect 514 52953 566 52962
rect 636 52996 688 53005
rect 636 52962 645 52996
rect 645 52962 679 52996
rect 679 52962 688 52996
rect 636 52953 688 52962
rect 762 52996 814 53005
rect 762 52962 771 52996
rect 771 52962 805 52996
rect 805 52962 814 52996
rect 762 52953 814 52962
rect 513 52710 565 52719
rect 513 52676 522 52710
rect 522 52676 556 52710
rect 556 52676 565 52710
rect 513 52667 565 52676
rect 639 52710 691 52719
rect 639 52676 648 52710
rect 648 52676 682 52710
rect 682 52676 691 52710
rect 639 52667 691 52676
rect 759 52710 811 52719
rect 759 52676 768 52710
rect 768 52676 802 52710
rect 802 52676 811 52710
rect 759 52667 811 52676
rect 513 52592 565 52601
rect 513 52558 522 52592
rect 522 52558 556 52592
rect 556 52558 565 52592
rect 513 52549 565 52558
rect 639 52592 691 52601
rect 639 52558 648 52592
rect 648 52558 682 52592
rect 682 52558 691 52592
rect 639 52549 691 52558
rect 759 52592 811 52601
rect 759 52558 768 52592
rect 768 52558 802 52592
rect 802 52558 811 52592
rect 759 52549 811 52558
rect 21078 52554 21130 52563
rect 21078 52520 21087 52554
rect 21087 52520 21121 52554
rect 21121 52520 21130 52554
rect 21078 52511 21130 52520
rect 21204 52554 21256 52563
rect 21204 52520 21213 52554
rect 21213 52520 21247 52554
rect 21247 52520 21256 52554
rect 21204 52511 21256 52520
rect 21324 52554 21376 52563
rect 21324 52520 21333 52554
rect 21333 52520 21367 52554
rect 21367 52520 21376 52554
rect 21324 52511 21376 52520
rect 21078 52436 21130 52445
rect 21078 52402 21087 52436
rect 21087 52402 21121 52436
rect 21121 52402 21130 52436
rect 21078 52393 21130 52402
rect 21204 52436 21256 52445
rect 21204 52402 21213 52436
rect 21213 52402 21247 52436
rect 21247 52402 21256 52436
rect 21204 52393 21256 52402
rect 21324 52436 21376 52445
rect 21324 52402 21333 52436
rect 21333 52402 21367 52436
rect 21367 52402 21376 52436
rect 21324 52393 21376 52402
rect 513 51523 565 51532
rect 513 51489 522 51523
rect 522 51489 556 51523
rect 556 51489 565 51523
rect 513 51480 565 51489
rect 639 51523 691 51532
rect 639 51489 648 51523
rect 648 51489 682 51523
rect 682 51489 691 51523
rect 639 51480 691 51489
rect 759 51523 811 51532
rect 759 51489 768 51523
rect 768 51489 802 51523
rect 802 51489 811 51523
rect 759 51480 811 51489
rect 513 51405 565 51414
rect 513 51371 522 51405
rect 522 51371 556 51405
rect 556 51371 565 51405
rect 513 51362 565 51371
rect 639 51405 691 51414
rect 639 51371 648 51405
rect 648 51371 682 51405
rect 682 51371 691 51405
rect 639 51362 691 51371
rect 759 51405 811 51414
rect 759 51371 768 51405
rect 768 51371 802 51405
rect 802 51371 811 51405
rect 759 51362 811 51371
rect 21078 51419 21130 51428
rect 21078 51385 21087 51419
rect 21087 51385 21121 51419
rect 21121 51385 21130 51419
rect 21078 51376 21130 51385
rect 21204 51419 21256 51428
rect 21204 51385 21213 51419
rect 21213 51385 21247 51419
rect 21247 51385 21256 51419
rect 21204 51376 21256 51385
rect 21324 51419 21376 51428
rect 21324 51385 21333 51419
rect 21333 51385 21367 51419
rect 21367 51385 21376 51419
rect 21324 51376 21376 51385
rect 21078 51301 21130 51310
rect 21078 51267 21087 51301
rect 21087 51267 21121 51301
rect 21121 51267 21130 51301
rect 21078 51258 21130 51267
rect 21204 51301 21256 51310
rect 21204 51267 21213 51301
rect 21213 51267 21247 51301
rect 21247 51267 21256 51301
rect 21204 51258 21256 51267
rect 21324 51301 21376 51310
rect 21324 51267 21333 51301
rect 21333 51267 21367 51301
rect 21367 51267 21376 51301
rect 21324 51258 21376 51267
rect 514 51039 566 51048
rect 514 51005 523 51039
rect 523 51005 557 51039
rect 557 51005 566 51039
rect 514 50996 566 51005
rect 636 51039 688 51048
rect 636 51005 645 51039
rect 645 51005 679 51039
rect 679 51005 688 51039
rect 636 50996 688 51005
rect 762 51039 814 51048
rect 762 51005 771 51039
rect 771 51005 805 51039
rect 805 51005 814 51039
rect 762 50996 814 51005
rect 514 50892 566 50901
rect 514 50858 523 50892
rect 523 50858 557 50892
rect 557 50858 566 50892
rect 514 50849 566 50858
rect 636 50892 688 50901
rect 636 50858 645 50892
rect 645 50858 679 50892
rect 679 50858 688 50892
rect 636 50849 688 50858
rect 762 50892 814 50901
rect 762 50858 771 50892
rect 771 50858 805 50892
rect 805 50858 814 50892
rect 762 50849 814 50858
rect 514 50755 566 50764
rect 514 50721 523 50755
rect 523 50721 557 50755
rect 557 50721 566 50755
rect 514 50712 566 50721
rect 636 50755 688 50764
rect 636 50721 645 50755
rect 645 50721 679 50755
rect 679 50721 688 50755
rect 636 50712 688 50721
rect 762 50755 814 50764
rect 762 50721 771 50755
rect 771 50721 805 50755
rect 805 50721 814 50755
rect 762 50712 814 50721
rect 22020 50137 22072 50146
rect 22020 50103 22029 50137
rect 22029 50103 22063 50137
rect 22063 50103 22072 50137
rect 22020 50094 22072 50103
rect 22146 50137 22198 50146
rect 22146 50103 22155 50137
rect 22155 50103 22189 50137
rect 22189 50103 22198 50137
rect 22146 50094 22198 50103
rect 22266 50137 22318 50146
rect 22266 50103 22275 50137
rect 22275 50103 22309 50137
rect 22309 50103 22318 50137
rect 22266 50094 22318 50103
rect 22020 50019 22072 50028
rect 22020 49985 22029 50019
rect 22029 49985 22063 50019
rect 22063 49985 22072 50019
rect 22020 49976 22072 49985
rect 22146 50019 22198 50028
rect 22146 49985 22155 50019
rect 22155 49985 22189 50019
rect 22189 49985 22198 50019
rect 22146 49976 22198 49985
rect 22266 50019 22318 50028
rect 22266 49985 22275 50019
rect 22275 49985 22309 50019
rect 22309 49985 22318 50019
rect 22266 49976 22318 49985
rect 514 49280 566 49289
rect 514 49246 523 49280
rect 523 49246 557 49280
rect 557 49246 566 49280
rect 514 49237 566 49246
rect 636 49280 688 49289
rect 636 49246 645 49280
rect 645 49246 679 49280
rect 679 49246 688 49280
rect 636 49237 688 49246
rect 762 49280 814 49289
rect 762 49246 771 49280
rect 771 49246 805 49280
rect 805 49246 814 49280
rect 762 49237 814 49246
rect 514 49133 566 49142
rect 514 49099 523 49133
rect 523 49099 557 49133
rect 557 49099 566 49133
rect 514 49090 566 49099
rect 636 49133 688 49142
rect 636 49099 645 49133
rect 645 49099 679 49133
rect 679 49099 688 49133
rect 636 49090 688 49099
rect 762 49133 814 49142
rect 762 49099 771 49133
rect 771 49099 805 49133
rect 805 49099 814 49133
rect 762 49090 814 49099
rect 514 48996 566 49005
rect 514 48962 523 48996
rect 523 48962 557 48996
rect 557 48962 566 48996
rect 514 48953 566 48962
rect 636 48996 688 49005
rect 636 48962 645 48996
rect 645 48962 679 48996
rect 679 48962 688 48996
rect 636 48953 688 48962
rect 762 48996 814 49005
rect 762 48962 771 48996
rect 771 48962 805 48996
rect 805 48962 814 48996
rect 762 48953 814 48962
rect 513 48701 565 48710
rect 513 48667 522 48701
rect 522 48667 556 48701
rect 556 48667 565 48701
rect 513 48658 565 48667
rect 639 48701 691 48710
rect 639 48667 648 48701
rect 648 48667 682 48701
rect 682 48667 691 48701
rect 639 48658 691 48667
rect 759 48701 811 48710
rect 759 48667 768 48701
rect 768 48667 802 48701
rect 802 48667 811 48701
rect 759 48658 811 48667
rect 513 48583 565 48592
rect 513 48549 522 48583
rect 522 48549 556 48583
rect 556 48549 565 48583
rect 513 48540 565 48549
rect 639 48583 691 48592
rect 639 48549 648 48583
rect 648 48549 682 48583
rect 682 48549 691 48583
rect 639 48540 691 48549
rect 759 48583 811 48592
rect 759 48549 768 48583
rect 768 48549 802 48583
rect 802 48549 811 48583
rect 759 48540 811 48549
rect 21078 48660 21130 48669
rect 21078 48626 21087 48660
rect 21087 48626 21121 48660
rect 21121 48626 21130 48660
rect 21078 48617 21130 48626
rect 21204 48660 21256 48669
rect 21204 48626 21213 48660
rect 21213 48626 21247 48660
rect 21247 48626 21256 48660
rect 21204 48617 21256 48626
rect 21324 48660 21376 48669
rect 21324 48626 21333 48660
rect 21333 48626 21367 48660
rect 21367 48626 21376 48660
rect 21324 48617 21376 48626
rect 21078 48542 21130 48551
rect 21078 48508 21087 48542
rect 21087 48508 21121 48542
rect 21121 48508 21130 48542
rect 21078 48499 21130 48508
rect 21204 48542 21256 48551
rect 21204 48508 21213 48542
rect 21213 48508 21247 48542
rect 21247 48508 21256 48542
rect 21204 48499 21256 48508
rect 21324 48542 21376 48551
rect 21324 48508 21333 48542
rect 21333 48508 21367 48542
rect 21367 48508 21376 48542
rect 21324 48499 21376 48508
rect 513 47548 565 47557
rect 513 47514 522 47548
rect 522 47514 556 47548
rect 556 47514 565 47548
rect 513 47505 565 47514
rect 639 47548 691 47557
rect 639 47514 648 47548
rect 648 47514 682 47548
rect 682 47514 691 47548
rect 639 47505 691 47514
rect 759 47548 811 47557
rect 759 47514 768 47548
rect 768 47514 802 47548
rect 802 47514 811 47548
rect 759 47505 811 47514
rect 513 47430 565 47439
rect 513 47396 522 47430
rect 522 47396 556 47430
rect 556 47396 565 47430
rect 513 47387 565 47396
rect 639 47430 691 47439
rect 639 47396 648 47430
rect 648 47396 682 47430
rect 682 47396 691 47430
rect 639 47387 691 47396
rect 759 47430 811 47439
rect 759 47396 768 47430
rect 768 47396 802 47430
rect 802 47396 811 47430
rect 759 47387 811 47396
rect 21078 47507 21130 47516
rect 21078 47473 21087 47507
rect 21087 47473 21121 47507
rect 21121 47473 21130 47507
rect 21078 47464 21130 47473
rect 21204 47507 21256 47516
rect 21204 47473 21213 47507
rect 21213 47473 21247 47507
rect 21247 47473 21256 47507
rect 21204 47464 21256 47473
rect 21324 47507 21376 47516
rect 21324 47473 21333 47507
rect 21333 47473 21367 47507
rect 21367 47473 21376 47507
rect 21324 47464 21376 47473
rect 21078 47389 21130 47398
rect 21078 47355 21087 47389
rect 21087 47355 21121 47389
rect 21121 47355 21130 47389
rect 21078 47346 21130 47355
rect 21204 47389 21256 47398
rect 21204 47355 21213 47389
rect 21213 47355 21247 47389
rect 21247 47355 21256 47389
rect 21204 47346 21256 47355
rect 21324 47389 21376 47398
rect 21324 47355 21333 47389
rect 21333 47355 21367 47389
rect 21367 47355 21376 47389
rect 21324 47346 21376 47355
rect 514 47039 566 47048
rect 514 47005 523 47039
rect 523 47005 557 47039
rect 557 47005 566 47039
rect 514 46996 566 47005
rect 636 47039 688 47048
rect 636 47005 645 47039
rect 645 47005 679 47039
rect 679 47005 688 47039
rect 636 46996 688 47005
rect 762 47039 814 47048
rect 762 47005 771 47039
rect 771 47005 805 47039
rect 805 47005 814 47039
rect 762 46996 814 47005
rect 514 46892 566 46901
rect 514 46858 523 46892
rect 523 46858 557 46892
rect 557 46858 566 46892
rect 514 46849 566 46858
rect 636 46892 688 46901
rect 636 46858 645 46892
rect 645 46858 679 46892
rect 679 46858 688 46892
rect 636 46849 688 46858
rect 762 46892 814 46901
rect 762 46858 771 46892
rect 771 46858 805 46892
rect 805 46858 814 46892
rect 762 46849 814 46858
rect 514 46755 566 46764
rect 514 46721 523 46755
rect 523 46721 557 46755
rect 557 46721 566 46755
rect 514 46712 566 46721
rect 636 46755 688 46764
rect 636 46721 645 46755
rect 645 46721 679 46755
rect 679 46721 688 46755
rect 636 46712 688 46721
rect 762 46755 814 46764
rect 762 46721 771 46755
rect 771 46721 805 46755
rect 805 46721 814 46755
rect 762 46712 814 46721
rect 22020 45879 22072 45888
rect 22020 45845 22029 45879
rect 22029 45845 22063 45879
rect 22063 45845 22072 45879
rect 22020 45836 22072 45845
rect 22146 45879 22198 45888
rect 22146 45845 22155 45879
rect 22155 45845 22189 45879
rect 22189 45845 22198 45879
rect 22146 45836 22198 45845
rect 22266 45879 22318 45888
rect 22266 45845 22275 45879
rect 22275 45845 22309 45879
rect 22309 45845 22318 45879
rect 22266 45836 22318 45845
rect 22020 45761 22072 45770
rect 22020 45727 22029 45761
rect 22029 45727 22063 45761
rect 22063 45727 22072 45761
rect 22020 45718 22072 45727
rect 22146 45761 22198 45770
rect 22146 45727 22155 45761
rect 22155 45727 22189 45761
rect 22189 45727 22198 45761
rect 22146 45718 22198 45727
rect 22266 45761 22318 45770
rect 22266 45727 22275 45761
rect 22275 45727 22309 45761
rect 22309 45727 22318 45761
rect 22266 45718 22318 45727
rect 514 45279 566 45288
rect 514 45245 523 45279
rect 523 45245 557 45279
rect 557 45245 566 45279
rect 514 45236 566 45245
rect 636 45279 688 45288
rect 636 45245 645 45279
rect 645 45245 679 45279
rect 679 45245 688 45279
rect 636 45236 688 45245
rect 762 45279 814 45288
rect 762 45245 771 45279
rect 771 45245 805 45279
rect 805 45245 814 45279
rect 762 45236 814 45245
rect 514 45132 566 45141
rect 514 45098 523 45132
rect 523 45098 557 45132
rect 557 45098 566 45132
rect 514 45089 566 45098
rect 636 45132 688 45141
rect 636 45098 645 45132
rect 645 45098 679 45132
rect 679 45098 688 45132
rect 636 45089 688 45098
rect 762 45132 814 45141
rect 762 45098 771 45132
rect 771 45098 805 45132
rect 805 45098 814 45132
rect 762 45089 814 45098
rect 514 44995 566 45004
rect 514 44961 523 44995
rect 523 44961 557 44995
rect 557 44961 566 44995
rect 514 44952 566 44961
rect 636 44995 688 45004
rect 636 44961 645 44995
rect 645 44961 679 44995
rect 679 44961 688 44995
rect 636 44952 688 44961
rect 762 44995 814 45004
rect 762 44961 771 44995
rect 771 44961 805 44995
rect 805 44961 814 44995
rect 762 44952 814 44961
rect 513 44488 565 44497
rect 513 44454 522 44488
rect 522 44454 556 44488
rect 556 44454 565 44488
rect 513 44445 565 44454
rect 639 44488 691 44497
rect 639 44454 648 44488
rect 648 44454 682 44488
rect 682 44454 691 44488
rect 639 44445 691 44454
rect 759 44488 811 44497
rect 759 44454 768 44488
rect 768 44454 802 44488
rect 802 44454 811 44488
rect 759 44445 811 44454
rect 513 44370 565 44379
rect 513 44336 522 44370
rect 522 44336 556 44370
rect 556 44336 565 44370
rect 513 44327 565 44336
rect 639 44370 691 44379
rect 639 44336 648 44370
rect 648 44336 682 44370
rect 682 44336 691 44370
rect 639 44327 691 44336
rect 759 44370 811 44379
rect 759 44336 768 44370
rect 768 44336 802 44370
rect 802 44336 811 44370
rect 759 44327 811 44336
rect 21078 44391 21130 44400
rect 21078 44357 21087 44391
rect 21087 44357 21121 44391
rect 21121 44357 21130 44391
rect 21078 44348 21130 44357
rect 21204 44391 21256 44400
rect 21204 44357 21213 44391
rect 21213 44357 21247 44391
rect 21247 44357 21256 44391
rect 21204 44348 21256 44357
rect 21324 44391 21376 44400
rect 21324 44357 21333 44391
rect 21333 44357 21367 44391
rect 21367 44357 21376 44391
rect 21324 44348 21376 44357
rect 21078 44273 21130 44282
rect 21078 44239 21087 44273
rect 21087 44239 21121 44273
rect 21121 44239 21130 44273
rect 21078 44230 21130 44239
rect 21204 44273 21256 44282
rect 21204 44239 21213 44273
rect 21213 44239 21247 44273
rect 21247 44239 21256 44273
rect 21204 44230 21256 44239
rect 21324 44273 21376 44282
rect 21324 44239 21333 44273
rect 21333 44239 21367 44273
rect 21367 44239 21376 44273
rect 21324 44230 21376 44239
rect 46 39675 98 39727
rect 171 39675 223 39727
rect 296 39675 348 39727
rect 21549 39660 21601 39712
rect 21674 39660 21726 39712
rect 21799 39660 21851 39712
rect 46 39569 98 39621
rect 171 39569 223 39621
rect 296 39569 348 39621
rect 21548 39540 21600 39592
rect 21673 39540 21725 39592
rect 21798 39540 21850 39592
rect 1662 39317 1714 39321
rect 1662 39283 1666 39317
rect 1666 39283 1700 39317
rect 1700 39283 1714 39317
rect 1662 39269 1714 39283
rect 1732 39317 1784 39321
rect 1732 39283 1746 39317
rect 1746 39283 1780 39317
rect 1780 39283 1784 39317
rect 1732 39269 1784 39283
rect 1886 39312 1891 39364
rect 1891 39312 1938 39364
rect 1950 39312 1997 39364
rect 1997 39312 2002 39364
rect 2042 39312 2047 39364
rect 2047 39312 2094 39364
rect 2106 39312 2153 39364
rect 2153 39312 2158 39364
rect 2198 39312 2203 39364
rect 2203 39312 2250 39364
rect 2262 39312 2309 39364
rect 2309 39312 2314 39364
rect 2551 39324 2603 39328
rect 2551 39290 2555 39324
rect 2555 39290 2589 39324
rect 2589 39290 2603 39324
rect 2551 39276 2603 39290
rect 2621 39324 2673 39328
rect 2621 39290 2635 39324
rect 2635 39290 2669 39324
rect 2669 39290 2673 39324
rect 2621 39276 2673 39290
rect 1662 39237 1714 39251
rect 1662 39203 1666 39237
rect 1666 39203 1700 39237
rect 1700 39203 1714 39237
rect 1662 39199 1714 39203
rect 1732 39237 1784 39251
rect 1732 39203 1746 39237
rect 1746 39203 1780 39237
rect 1780 39203 1784 39237
rect 1732 39199 1784 39203
rect 2551 39244 2603 39258
rect 2551 39210 2555 39244
rect 2555 39210 2589 39244
rect 2589 39210 2603 39244
rect 2551 39206 2603 39210
rect 2621 39244 2673 39258
rect 2621 39210 2635 39244
rect 2635 39210 2669 39244
rect 2669 39210 2673 39244
rect 2621 39206 2673 39210
rect 494 39065 546 39117
rect 608 39065 660 39117
rect 722 39065 774 39117
rect 1507 38722 1559 38774
rect 3529 38870 3581 38880
rect 3529 38836 3553 38870
rect 3553 38836 3581 38870
rect 3529 38828 3581 38836
rect 4610 38870 4662 38879
rect 4610 38836 4615 38870
rect 4615 38836 4649 38870
rect 4649 38836 4662 38870
rect 4610 38827 4662 38836
rect 31 38521 83 38573
rect 145 38521 197 38573
rect 259 38521 311 38573
rect 1471 38259 1523 38269
rect 1471 38225 1480 38259
rect 1480 38225 1514 38259
rect 1514 38225 1523 38259
rect 1471 38217 1523 38225
rect 3608 38296 3660 38348
rect 4652 38258 4704 38267
rect 4652 38224 4662 38258
rect 4662 38224 4696 38258
rect 4696 38224 4704 38258
rect 4652 38215 4704 38224
rect 494 37977 546 38029
rect 608 37977 660 38029
rect 722 37977 774 38029
rect 1463 37782 1515 37790
rect 1463 37748 1481 37782
rect 1481 37748 1515 37782
rect 1463 37738 1515 37748
rect 3523 37845 3575 37897
rect 4652 37782 4704 37791
rect 4652 37748 4662 37782
rect 4662 37748 4696 37782
rect 4696 37748 4704 37782
rect 4652 37739 4704 37748
rect 31 37433 83 37485
rect 145 37433 197 37485
rect 259 37433 311 37485
rect 1683 37351 1735 37358
rect 1683 37317 1692 37351
rect 1692 37317 1726 37351
rect 1726 37317 1735 37351
rect 1683 37306 1735 37317
rect 1683 37239 1735 37252
rect 1683 37205 1692 37239
rect 1692 37205 1726 37239
rect 1726 37205 1735 37239
rect 1683 37200 1735 37205
rect 3553 37170 3605 37182
rect 3553 37136 3587 37170
rect 3587 37136 3605 37170
rect 3553 37130 3605 37136
rect 4609 37170 4661 37181
rect 4609 37136 4615 37170
rect 4615 37136 4649 37170
rect 4649 37136 4661 37170
rect 4609 37129 4661 37136
rect 494 36889 546 36941
rect 608 36889 660 36941
rect 722 36889 774 36941
rect 2551 36826 2603 36830
rect 2551 36792 2555 36826
rect 2555 36792 2589 36826
rect 2589 36792 2603 36826
rect 2551 36778 2603 36792
rect 2621 36826 2673 36830
rect 2621 36792 2635 36826
rect 2635 36792 2669 36826
rect 2669 36792 2673 36826
rect 2621 36778 2673 36792
rect 2551 36747 2603 36763
rect 2551 36713 2555 36747
rect 2555 36713 2589 36747
rect 2589 36713 2603 36747
rect 2551 36711 2603 36713
rect 2621 36747 2673 36763
rect 2621 36713 2635 36747
rect 2635 36713 2669 36747
rect 2669 36713 2673 36747
rect 2621 36711 2673 36713
rect 2765 36826 2817 36830
rect 2765 36792 2769 36826
rect 2769 36792 2803 36826
rect 2803 36792 2817 36826
rect 2765 36778 2817 36792
rect 2835 36826 2887 36830
rect 2835 36792 2849 36826
rect 2849 36792 2883 36826
rect 2883 36792 2887 36826
rect 2835 36778 2887 36792
rect 2765 36747 2817 36765
rect 2765 36713 2769 36747
rect 2769 36713 2803 36747
rect 2803 36713 2817 36747
rect 2835 36747 2887 36765
rect 2835 36713 2849 36747
rect 2849 36713 2883 36747
rect 2883 36713 2887 36747
rect 21075 36106 21127 36158
rect 21200 36106 21252 36158
rect 21325 36106 21377 36158
rect 21074 35986 21126 36038
rect 21199 35986 21251 36038
rect 21324 35986 21376 36038
rect 21079 35571 21131 35580
rect 21079 35537 21088 35571
rect 21088 35537 21122 35571
rect 21122 35537 21131 35571
rect 21079 35528 21131 35537
rect 21201 35571 21253 35580
rect 21201 35537 21210 35571
rect 21210 35537 21244 35571
rect 21244 35537 21253 35571
rect 21201 35528 21253 35537
rect 21327 35571 21379 35580
rect 21327 35537 21336 35571
rect 21336 35537 21370 35571
rect 21370 35537 21379 35571
rect 21327 35528 21379 35537
rect 21079 35424 21131 35433
rect 21079 35390 21088 35424
rect 21088 35390 21122 35424
rect 21122 35390 21131 35424
rect 21079 35381 21131 35390
rect 21201 35424 21253 35433
rect 21201 35390 21210 35424
rect 21210 35390 21244 35424
rect 21244 35390 21253 35424
rect 21201 35381 21253 35390
rect 21327 35424 21379 35433
rect 21327 35390 21336 35424
rect 21336 35390 21370 35424
rect 21370 35390 21379 35424
rect 21327 35381 21379 35390
rect 21079 35287 21131 35296
rect 21079 35253 21088 35287
rect 21088 35253 21122 35287
rect 21122 35253 21131 35287
rect 21079 35244 21131 35253
rect 21201 35287 21253 35296
rect 21201 35253 21210 35287
rect 21210 35253 21244 35287
rect 21244 35253 21253 35287
rect 21201 35244 21253 35253
rect 21327 35287 21379 35296
rect 21327 35253 21336 35287
rect 21336 35253 21370 35287
rect 21370 35253 21379 35287
rect 21327 35244 21379 35253
rect 20574 34610 20626 34662
rect 20699 34610 20751 34662
rect 20824 34610 20876 34662
rect 21549 34610 21601 34662
rect 21674 34610 21726 34662
rect 21799 34610 21851 34662
rect 20573 34490 20625 34542
rect 20698 34490 20750 34542
rect 20823 34490 20875 34542
rect 21548 34490 21600 34542
rect 21673 34490 21725 34542
rect 21798 34490 21850 34542
rect 21079 33811 21131 33820
rect 21079 33777 21088 33811
rect 21088 33777 21122 33811
rect 21122 33777 21131 33811
rect 21079 33768 21131 33777
rect 21201 33811 21253 33820
rect 21201 33777 21210 33811
rect 21210 33777 21244 33811
rect 21244 33777 21253 33811
rect 21201 33768 21253 33777
rect 21327 33811 21379 33820
rect 21327 33777 21336 33811
rect 21336 33777 21370 33811
rect 21370 33777 21379 33811
rect 21327 33768 21379 33777
rect 21079 33664 21131 33673
rect 21079 33630 21088 33664
rect 21088 33630 21122 33664
rect 21122 33630 21131 33664
rect 21079 33621 21131 33630
rect 21201 33664 21253 33673
rect 21201 33630 21210 33664
rect 21210 33630 21244 33664
rect 21244 33630 21253 33664
rect 21201 33621 21253 33630
rect 21327 33664 21379 33673
rect 21327 33630 21336 33664
rect 21336 33630 21370 33664
rect 21370 33630 21379 33664
rect 21327 33621 21379 33630
rect 21079 33527 21131 33536
rect 21079 33493 21088 33527
rect 21088 33493 21122 33527
rect 21122 33493 21131 33527
rect 21079 33484 21131 33493
rect 21201 33527 21253 33536
rect 21201 33493 21210 33527
rect 21210 33493 21244 33527
rect 21244 33493 21253 33527
rect 21201 33484 21253 33493
rect 21327 33527 21379 33536
rect 21327 33493 21336 33527
rect 21336 33493 21370 33527
rect 21370 33493 21379 33527
rect 21327 33484 21379 33493
rect 21074 33051 21126 33103
rect 21199 33051 21251 33103
rect 21324 33051 21376 33103
rect 21073 32931 21125 32983
rect 21198 32931 21250 32983
rect 21323 32931 21375 32983
rect 513 32281 565 32290
rect 513 32247 522 32281
rect 522 32247 556 32281
rect 556 32247 565 32281
rect 513 32238 565 32247
rect 639 32281 691 32290
rect 639 32247 648 32281
rect 648 32247 682 32281
rect 682 32247 691 32281
rect 639 32238 691 32247
rect 759 32281 811 32290
rect 759 32247 768 32281
rect 768 32247 802 32281
rect 802 32247 811 32281
rect 759 32238 811 32247
rect 21078 32281 21130 32290
rect 21078 32247 21087 32281
rect 21087 32247 21121 32281
rect 21121 32247 21130 32281
rect 21078 32238 21130 32247
rect 21204 32281 21256 32290
rect 21204 32247 21213 32281
rect 21213 32247 21247 32281
rect 21247 32247 21256 32281
rect 21204 32238 21256 32247
rect 21324 32281 21376 32290
rect 21324 32247 21333 32281
rect 21333 32247 21367 32281
rect 21367 32247 21376 32281
rect 21324 32238 21376 32247
rect 513 32163 565 32172
rect 513 32129 522 32163
rect 522 32129 556 32163
rect 556 32129 565 32163
rect 513 32120 565 32129
rect 639 32163 691 32172
rect 639 32129 648 32163
rect 648 32129 682 32163
rect 682 32129 691 32163
rect 639 32120 691 32129
rect 759 32163 811 32172
rect 759 32129 768 32163
rect 768 32129 802 32163
rect 802 32129 811 32163
rect 759 32120 811 32129
rect 21078 32163 21130 32172
rect 21078 32129 21087 32163
rect 21087 32129 21121 32163
rect 21121 32129 21130 32163
rect 21078 32120 21130 32129
rect 21204 32163 21256 32172
rect 21204 32129 21213 32163
rect 21213 32129 21247 32163
rect 21247 32129 21256 32163
rect 21204 32120 21256 32129
rect 21324 32163 21376 32172
rect 21324 32129 21333 32163
rect 21333 32129 21367 32163
rect 21367 32129 21376 32163
rect 21324 32120 21376 32129
rect 513 31499 565 31508
rect 513 31465 522 31499
rect 522 31465 556 31499
rect 556 31465 565 31499
rect 513 31456 565 31465
rect 639 31499 691 31508
rect 639 31465 648 31499
rect 648 31465 682 31499
rect 682 31465 691 31499
rect 639 31456 691 31465
rect 759 31499 811 31508
rect 759 31465 768 31499
rect 768 31465 802 31499
rect 802 31465 811 31499
rect 759 31456 811 31465
rect 513 31381 565 31390
rect 513 31347 522 31381
rect 522 31347 556 31381
rect 556 31347 565 31381
rect 513 31338 565 31347
rect 639 31381 691 31390
rect 639 31347 648 31381
rect 648 31347 682 31381
rect 682 31347 691 31381
rect 639 31338 691 31347
rect 759 31381 811 31390
rect 759 31347 768 31381
rect 768 31347 802 31381
rect 802 31347 811 31381
rect 759 31338 811 31347
rect 21078 31499 21130 31508
rect 21078 31465 21087 31499
rect 21087 31465 21121 31499
rect 21121 31465 21130 31499
rect 21078 31456 21130 31465
rect 21204 31499 21256 31508
rect 21204 31465 21213 31499
rect 21213 31465 21247 31499
rect 21247 31465 21256 31499
rect 21204 31456 21256 31465
rect 21324 31499 21376 31508
rect 21324 31465 21333 31499
rect 21333 31465 21367 31499
rect 21367 31465 21376 31499
rect 21324 31456 21376 31465
rect 21078 31381 21130 31390
rect 21078 31347 21087 31381
rect 21087 31347 21121 31381
rect 21121 31347 21130 31381
rect 21078 31338 21130 31347
rect 21204 31381 21256 31390
rect 21204 31347 21213 31381
rect 21213 31347 21247 31381
rect 21247 31347 21256 31381
rect 21204 31338 21256 31347
rect 21324 31381 21376 31390
rect 21324 31347 21333 31381
rect 21333 31347 21367 31381
rect 21367 31347 21376 31381
rect 21324 31338 21376 31347
rect 514 31040 566 31049
rect 514 31006 523 31040
rect 523 31006 557 31040
rect 557 31006 566 31040
rect 514 30997 566 31006
rect 636 31040 688 31049
rect 636 31006 645 31040
rect 645 31006 679 31040
rect 679 31006 688 31040
rect 636 30997 688 31006
rect 762 31040 814 31049
rect 762 31006 771 31040
rect 771 31006 805 31040
rect 805 31006 814 31040
rect 762 30997 814 31006
rect 514 30893 566 30902
rect 514 30859 523 30893
rect 523 30859 557 30893
rect 557 30859 566 30893
rect 514 30850 566 30859
rect 636 30893 688 30902
rect 636 30859 645 30893
rect 645 30859 679 30893
rect 679 30859 688 30893
rect 636 30850 688 30859
rect 762 30893 814 30902
rect 762 30859 771 30893
rect 771 30859 805 30893
rect 805 30859 814 30893
rect 762 30850 814 30859
rect 514 30756 566 30765
rect 514 30722 523 30756
rect 523 30722 557 30756
rect 557 30722 566 30756
rect 514 30713 566 30722
rect 636 30756 688 30765
rect 636 30722 645 30756
rect 645 30722 679 30756
rect 679 30722 688 30756
rect 636 30713 688 30722
rect 762 30756 814 30765
rect 762 30722 771 30756
rect 771 30722 805 30756
rect 805 30722 814 30756
rect 762 30713 814 30722
rect 22020 30109 22072 30118
rect 22020 30075 22029 30109
rect 22029 30075 22063 30109
rect 22063 30075 22072 30109
rect 22020 30066 22072 30075
rect 22146 30109 22198 30118
rect 22146 30075 22155 30109
rect 22155 30075 22189 30109
rect 22189 30075 22198 30109
rect 22146 30066 22198 30075
rect 22266 30109 22318 30118
rect 22266 30075 22275 30109
rect 22275 30075 22309 30109
rect 22309 30075 22318 30109
rect 22266 30066 22318 30075
rect 22020 29991 22072 30000
rect 22020 29957 22029 29991
rect 22029 29957 22063 29991
rect 22063 29957 22072 29991
rect 22020 29948 22072 29957
rect 22146 29991 22198 30000
rect 22146 29957 22155 29991
rect 22155 29957 22189 29991
rect 22189 29957 22198 29991
rect 22146 29948 22198 29957
rect 22266 29991 22318 30000
rect 22266 29957 22275 29991
rect 22275 29957 22309 29991
rect 22309 29957 22318 29991
rect 22266 29948 22318 29957
rect 514 29273 566 29282
rect 514 29239 523 29273
rect 523 29239 557 29273
rect 557 29239 566 29273
rect 514 29230 566 29239
rect 636 29273 688 29282
rect 636 29239 645 29273
rect 645 29239 679 29273
rect 679 29239 688 29273
rect 636 29230 688 29239
rect 762 29273 814 29282
rect 762 29239 771 29273
rect 771 29239 805 29273
rect 805 29239 814 29273
rect 762 29230 814 29239
rect 514 29126 566 29135
rect 514 29092 523 29126
rect 523 29092 557 29126
rect 557 29092 566 29126
rect 514 29083 566 29092
rect 636 29126 688 29135
rect 636 29092 645 29126
rect 645 29092 679 29126
rect 679 29092 688 29126
rect 636 29083 688 29092
rect 762 29126 814 29135
rect 762 29092 771 29126
rect 771 29092 805 29126
rect 805 29092 814 29126
rect 762 29083 814 29092
rect 514 28989 566 28998
rect 514 28955 523 28989
rect 523 28955 557 28989
rect 557 28955 566 28989
rect 514 28946 566 28955
rect 636 28989 688 28998
rect 636 28955 645 28989
rect 645 28955 679 28989
rect 679 28955 688 28989
rect 636 28946 688 28955
rect 762 28989 814 28998
rect 762 28955 771 28989
rect 771 28955 805 28989
rect 805 28955 814 28989
rect 762 28946 814 28955
rect 513 28587 565 28596
rect 513 28553 522 28587
rect 522 28553 556 28587
rect 556 28553 565 28587
rect 513 28544 565 28553
rect 639 28587 691 28596
rect 639 28553 648 28587
rect 648 28553 682 28587
rect 682 28553 691 28587
rect 639 28544 691 28553
rect 759 28587 811 28596
rect 759 28553 768 28587
rect 768 28553 802 28587
rect 802 28553 811 28587
rect 759 28544 811 28553
rect 513 28469 565 28478
rect 513 28435 522 28469
rect 522 28435 556 28469
rect 556 28435 565 28469
rect 513 28426 565 28435
rect 639 28469 691 28478
rect 639 28435 648 28469
rect 648 28435 682 28469
rect 682 28435 691 28469
rect 639 28426 691 28435
rect 759 28469 811 28478
rect 759 28435 768 28469
rect 768 28435 802 28469
rect 802 28435 811 28469
rect 759 28426 811 28435
rect 21078 28538 21130 28547
rect 21078 28504 21087 28538
rect 21087 28504 21121 28538
rect 21121 28504 21130 28538
rect 21078 28495 21130 28504
rect 21204 28538 21256 28547
rect 21204 28504 21213 28538
rect 21213 28504 21247 28538
rect 21247 28504 21256 28538
rect 21204 28495 21256 28504
rect 21324 28538 21376 28547
rect 21324 28504 21333 28538
rect 21333 28504 21367 28538
rect 21367 28504 21376 28538
rect 21324 28495 21376 28504
rect 21078 28420 21130 28429
rect 21078 28386 21087 28420
rect 21087 28386 21121 28420
rect 21121 28386 21130 28420
rect 21078 28377 21130 28386
rect 21204 28420 21256 28429
rect 21204 28386 21213 28420
rect 21213 28386 21247 28420
rect 21247 28386 21256 28420
rect 21204 28377 21256 28386
rect 21324 28420 21376 28429
rect 21324 28386 21333 28420
rect 21333 28386 21367 28420
rect 21367 28386 21376 28420
rect 21324 28377 21376 28386
rect 513 27583 565 27592
rect 513 27549 522 27583
rect 522 27549 556 27583
rect 556 27549 565 27583
rect 513 27540 565 27549
rect 639 27583 691 27592
rect 639 27549 648 27583
rect 648 27549 682 27583
rect 682 27549 691 27583
rect 639 27540 691 27549
rect 759 27583 811 27592
rect 759 27549 768 27583
rect 768 27549 802 27583
rect 802 27549 811 27583
rect 759 27540 811 27549
rect 513 27465 565 27474
rect 513 27431 522 27465
rect 522 27431 556 27465
rect 556 27431 565 27465
rect 513 27422 565 27431
rect 639 27465 691 27474
rect 639 27431 648 27465
rect 648 27431 682 27465
rect 682 27431 691 27465
rect 639 27422 691 27431
rect 759 27465 811 27474
rect 759 27431 768 27465
rect 768 27431 802 27465
rect 802 27431 811 27465
rect 759 27422 811 27431
rect 21078 27421 21130 27430
rect 21078 27387 21087 27421
rect 21087 27387 21121 27421
rect 21121 27387 21130 27421
rect 21078 27378 21130 27387
rect 21204 27421 21256 27430
rect 21204 27387 21213 27421
rect 21213 27387 21247 27421
rect 21247 27387 21256 27421
rect 21204 27378 21256 27387
rect 21324 27421 21376 27430
rect 21324 27387 21333 27421
rect 21333 27387 21367 27421
rect 21367 27387 21376 27421
rect 21324 27378 21376 27387
rect 21078 27303 21130 27312
rect 21078 27269 21087 27303
rect 21087 27269 21121 27303
rect 21121 27269 21130 27303
rect 21078 27260 21130 27269
rect 21204 27303 21256 27312
rect 21204 27269 21213 27303
rect 21213 27269 21247 27303
rect 21247 27269 21256 27303
rect 21204 27260 21256 27269
rect 21324 27303 21376 27312
rect 21324 27269 21333 27303
rect 21333 27269 21367 27303
rect 21367 27269 21376 27303
rect 21324 27260 21376 27269
rect 514 27039 566 27048
rect 514 27005 523 27039
rect 523 27005 557 27039
rect 557 27005 566 27039
rect 514 26996 566 27005
rect 636 27039 688 27048
rect 636 27005 645 27039
rect 645 27005 679 27039
rect 679 27005 688 27039
rect 636 26996 688 27005
rect 762 27039 814 27048
rect 762 27005 771 27039
rect 771 27005 805 27039
rect 805 27005 814 27039
rect 762 26996 814 27005
rect 514 26892 566 26901
rect 514 26858 523 26892
rect 523 26858 557 26892
rect 557 26858 566 26892
rect 514 26849 566 26858
rect 636 26892 688 26901
rect 636 26858 645 26892
rect 645 26858 679 26892
rect 679 26858 688 26892
rect 636 26849 688 26858
rect 762 26892 814 26901
rect 762 26858 771 26892
rect 771 26858 805 26892
rect 805 26858 814 26892
rect 762 26849 814 26858
rect 514 26755 566 26764
rect 514 26721 523 26755
rect 523 26721 557 26755
rect 557 26721 566 26755
rect 514 26712 566 26721
rect 636 26755 688 26764
rect 636 26721 645 26755
rect 645 26721 679 26755
rect 679 26721 688 26755
rect 636 26712 688 26721
rect 762 26755 814 26764
rect 762 26721 771 26755
rect 771 26721 805 26755
rect 805 26721 814 26755
rect 762 26712 814 26721
rect 22020 25950 22072 25959
rect 22020 25916 22029 25950
rect 22029 25916 22063 25950
rect 22063 25916 22072 25950
rect 22020 25907 22072 25916
rect 22146 25950 22198 25959
rect 22146 25916 22155 25950
rect 22155 25916 22189 25950
rect 22189 25916 22198 25950
rect 22146 25907 22198 25916
rect 22266 25950 22318 25959
rect 22266 25916 22275 25950
rect 22275 25916 22309 25950
rect 22309 25916 22318 25950
rect 22266 25907 22318 25916
rect 22020 25832 22072 25841
rect 22020 25798 22029 25832
rect 22029 25798 22063 25832
rect 22063 25798 22072 25832
rect 22020 25789 22072 25798
rect 22146 25832 22198 25841
rect 22146 25798 22155 25832
rect 22155 25798 22189 25832
rect 22189 25798 22198 25832
rect 22146 25789 22198 25798
rect 22266 25832 22318 25841
rect 22266 25798 22275 25832
rect 22275 25798 22309 25832
rect 22309 25798 22318 25832
rect 22266 25789 22318 25798
rect 514 25279 566 25288
rect 514 25245 523 25279
rect 523 25245 557 25279
rect 557 25245 566 25279
rect 514 25236 566 25245
rect 636 25279 688 25288
rect 636 25245 645 25279
rect 645 25245 679 25279
rect 679 25245 688 25279
rect 636 25236 688 25245
rect 762 25279 814 25288
rect 762 25245 771 25279
rect 771 25245 805 25279
rect 805 25245 814 25279
rect 762 25236 814 25245
rect 514 25132 566 25141
rect 514 25098 523 25132
rect 523 25098 557 25132
rect 557 25098 566 25132
rect 514 25089 566 25098
rect 636 25132 688 25141
rect 636 25098 645 25132
rect 645 25098 679 25132
rect 679 25098 688 25132
rect 636 25089 688 25098
rect 762 25132 814 25141
rect 762 25098 771 25132
rect 771 25098 805 25132
rect 805 25098 814 25132
rect 762 25089 814 25098
rect 514 24995 566 25004
rect 514 24961 523 24995
rect 523 24961 557 24995
rect 557 24961 566 24995
rect 514 24952 566 24961
rect 636 24995 688 25004
rect 636 24961 645 24995
rect 645 24961 679 24995
rect 679 24961 688 24995
rect 636 24952 688 24961
rect 762 24995 814 25004
rect 762 24961 771 24995
rect 771 24961 805 24995
rect 805 24961 814 24995
rect 762 24952 814 24961
rect 513 24605 565 24614
rect 513 24571 522 24605
rect 522 24571 556 24605
rect 556 24571 565 24605
rect 513 24562 565 24571
rect 639 24605 691 24614
rect 639 24571 648 24605
rect 648 24571 682 24605
rect 682 24571 691 24605
rect 639 24562 691 24571
rect 759 24605 811 24614
rect 759 24571 768 24605
rect 768 24571 802 24605
rect 802 24571 811 24605
rect 759 24562 811 24571
rect 513 24487 565 24496
rect 513 24453 522 24487
rect 522 24453 556 24487
rect 556 24453 565 24487
rect 513 24444 565 24453
rect 639 24487 691 24496
rect 639 24453 648 24487
rect 648 24453 682 24487
rect 682 24453 691 24487
rect 639 24444 691 24453
rect 759 24487 811 24496
rect 759 24453 768 24487
rect 768 24453 802 24487
rect 802 24453 811 24487
rect 759 24444 811 24453
rect 21078 24578 21130 24587
rect 21078 24544 21087 24578
rect 21087 24544 21121 24578
rect 21121 24544 21130 24578
rect 21078 24535 21130 24544
rect 21204 24578 21256 24587
rect 21204 24544 21213 24578
rect 21213 24544 21247 24578
rect 21247 24544 21256 24578
rect 21204 24535 21256 24544
rect 21324 24578 21376 24587
rect 21324 24544 21333 24578
rect 21333 24544 21367 24578
rect 21367 24544 21376 24578
rect 21324 24535 21376 24544
rect 21078 24460 21130 24469
rect 21078 24426 21087 24460
rect 21087 24426 21121 24460
rect 21121 24426 21130 24460
rect 21078 24417 21130 24426
rect 21204 24460 21256 24469
rect 21204 24426 21213 24460
rect 21213 24426 21247 24460
rect 21247 24426 21256 24460
rect 21204 24417 21256 24426
rect 21324 24460 21376 24469
rect 21324 24426 21333 24460
rect 21333 24426 21367 24460
rect 21367 24426 21376 24460
rect 21324 24417 21376 24426
rect 513 23523 565 23532
rect 513 23489 522 23523
rect 522 23489 556 23523
rect 556 23489 565 23523
rect 513 23480 565 23489
rect 639 23523 691 23532
rect 639 23489 648 23523
rect 648 23489 682 23523
rect 682 23489 691 23523
rect 639 23480 691 23489
rect 759 23523 811 23532
rect 759 23489 768 23523
rect 768 23489 802 23523
rect 802 23489 811 23523
rect 759 23480 811 23489
rect 513 23405 565 23414
rect 513 23371 522 23405
rect 522 23371 556 23405
rect 556 23371 565 23405
rect 513 23362 565 23371
rect 639 23405 691 23414
rect 639 23371 648 23405
rect 648 23371 682 23405
rect 682 23371 691 23405
rect 639 23362 691 23371
rect 759 23405 811 23414
rect 759 23371 768 23405
rect 768 23371 802 23405
rect 802 23371 811 23405
rect 759 23362 811 23371
rect 21078 23403 21130 23412
rect 21078 23369 21087 23403
rect 21087 23369 21121 23403
rect 21121 23369 21130 23403
rect 21078 23360 21130 23369
rect 21204 23403 21256 23412
rect 21204 23369 21213 23403
rect 21213 23369 21247 23403
rect 21247 23369 21256 23403
rect 21204 23360 21256 23369
rect 21324 23403 21376 23412
rect 21324 23369 21333 23403
rect 21333 23369 21367 23403
rect 21367 23369 21376 23403
rect 21324 23360 21376 23369
rect 21078 23285 21130 23294
rect 21078 23251 21087 23285
rect 21087 23251 21121 23285
rect 21121 23251 21130 23285
rect 21078 23242 21130 23251
rect 21204 23285 21256 23294
rect 21204 23251 21213 23285
rect 21213 23251 21247 23285
rect 21247 23251 21256 23285
rect 21204 23242 21256 23251
rect 21324 23285 21376 23294
rect 21324 23251 21333 23285
rect 21333 23251 21367 23285
rect 21367 23251 21376 23285
rect 21324 23242 21376 23251
rect 514 23039 566 23048
rect 514 23005 523 23039
rect 523 23005 557 23039
rect 557 23005 566 23039
rect 514 22996 566 23005
rect 636 23039 688 23048
rect 636 23005 645 23039
rect 645 23005 679 23039
rect 679 23005 688 23039
rect 636 22996 688 23005
rect 762 23039 814 23048
rect 762 23005 771 23039
rect 771 23005 805 23039
rect 805 23005 814 23039
rect 762 22996 814 23005
rect 514 22892 566 22901
rect 514 22858 523 22892
rect 523 22858 557 22892
rect 557 22858 566 22892
rect 514 22849 566 22858
rect 636 22892 688 22901
rect 636 22858 645 22892
rect 645 22858 679 22892
rect 679 22858 688 22892
rect 636 22849 688 22858
rect 762 22892 814 22901
rect 762 22858 771 22892
rect 771 22858 805 22892
rect 805 22858 814 22892
rect 762 22849 814 22858
rect 514 22755 566 22764
rect 514 22721 523 22755
rect 523 22721 557 22755
rect 557 22721 566 22755
rect 514 22712 566 22721
rect 636 22755 688 22764
rect 636 22721 645 22755
rect 645 22721 679 22755
rect 679 22721 688 22755
rect 636 22712 688 22721
rect 762 22755 814 22764
rect 762 22721 771 22755
rect 771 22721 805 22755
rect 805 22721 814 22755
rect 762 22712 814 22721
rect 22020 22160 22072 22169
rect 22020 22126 22029 22160
rect 22029 22126 22063 22160
rect 22063 22126 22072 22160
rect 22020 22117 22072 22126
rect 22146 22160 22198 22169
rect 22146 22126 22155 22160
rect 22155 22126 22189 22160
rect 22189 22126 22198 22160
rect 22146 22117 22198 22126
rect 22266 22160 22318 22169
rect 22266 22126 22275 22160
rect 22275 22126 22309 22160
rect 22309 22126 22318 22160
rect 22266 22117 22318 22126
rect 22020 22042 22072 22051
rect 22020 22008 22029 22042
rect 22029 22008 22063 22042
rect 22063 22008 22072 22042
rect 22020 21999 22072 22008
rect 22146 22042 22198 22051
rect 22146 22008 22155 22042
rect 22155 22008 22189 22042
rect 22189 22008 22198 22042
rect 22146 21999 22198 22008
rect 22266 22042 22318 22051
rect 22266 22008 22275 22042
rect 22275 22008 22309 22042
rect 22309 22008 22318 22042
rect 22266 21999 22318 22008
rect 514 21280 566 21289
rect 514 21246 523 21280
rect 523 21246 557 21280
rect 557 21246 566 21280
rect 514 21237 566 21246
rect 636 21280 688 21289
rect 636 21246 645 21280
rect 645 21246 679 21280
rect 679 21246 688 21280
rect 636 21237 688 21246
rect 762 21280 814 21289
rect 762 21246 771 21280
rect 771 21246 805 21280
rect 805 21246 814 21280
rect 762 21237 814 21246
rect 514 21133 566 21142
rect 514 21099 523 21133
rect 523 21099 557 21133
rect 557 21099 566 21133
rect 514 21090 566 21099
rect 636 21133 688 21142
rect 636 21099 645 21133
rect 645 21099 679 21133
rect 679 21099 688 21133
rect 636 21090 688 21099
rect 762 21133 814 21142
rect 762 21099 771 21133
rect 771 21099 805 21133
rect 805 21099 814 21133
rect 762 21090 814 21099
rect 514 20996 566 21005
rect 514 20962 523 20996
rect 523 20962 557 20996
rect 557 20962 566 20996
rect 514 20953 566 20962
rect 636 20996 688 21005
rect 636 20962 645 20996
rect 645 20962 679 20996
rect 679 20962 688 20996
rect 636 20953 688 20962
rect 762 20996 814 21005
rect 762 20962 771 20996
rect 771 20962 805 20996
rect 805 20962 814 20996
rect 762 20953 814 20962
rect 513 20648 565 20657
rect 513 20614 522 20648
rect 522 20614 556 20648
rect 556 20614 565 20648
rect 513 20605 565 20614
rect 639 20648 691 20657
rect 639 20614 648 20648
rect 648 20614 682 20648
rect 682 20614 691 20648
rect 639 20605 691 20614
rect 759 20648 811 20657
rect 759 20614 768 20648
rect 768 20614 802 20648
rect 802 20614 811 20648
rect 759 20605 811 20614
rect 513 20530 565 20539
rect 513 20496 522 20530
rect 522 20496 556 20530
rect 556 20496 565 20530
rect 513 20487 565 20496
rect 639 20530 691 20539
rect 639 20496 648 20530
rect 648 20496 682 20530
rect 682 20496 691 20530
rect 639 20487 691 20496
rect 759 20530 811 20539
rect 759 20496 768 20530
rect 768 20496 802 20530
rect 802 20496 811 20530
rect 759 20487 811 20496
rect 21078 20562 21130 20571
rect 21078 20528 21087 20562
rect 21087 20528 21121 20562
rect 21121 20528 21130 20562
rect 21078 20519 21130 20528
rect 21204 20562 21256 20571
rect 21204 20528 21213 20562
rect 21213 20528 21247 20562
rect 21247 20528 21256 20562
rect 21204 20519 21256 20528
rect 21324 20562 21376 20571
rect 21324 20528 21333 20562
rect 21333 20528 21367 20562
rect 21367 20528 21376 20562
rect 21324 20519 21376 20528
rect 21078 20444 21130 20453
rect 21078 20410 21087 20444
rect 21087 20410 21121 20444
rect 21121 20410 21130 20444
rect 21078 20401 21130 20410
rect 21204 20444 21256 20453
rect 21204 20410 21213 20444
rect 21213 20410 21247 20444
rect 21247 20410 21256 20444
rect 21204 20401 21256 20410
rect 21324 20444 21376 20453
rect 21324 20410 21333 20444
rect 21333 20410 21367 20444
rect 21367 20410 21376 20444
rect 21324 20401 21376 20410
rect 513 19547 565 19556
rect 513 19513 522 19547
rect 522 19513 556 19547
rect 556 19513 565 19547
rect 513 19504 565 19513
rect 639 19547 691 19556
rect 639 19513 648 19547
rect 648 19513 682 19547
rect 682 19513 691 19547
rect 639 19504 691 19513
rect 759 19547 811 19556
rect 759 19513 768 19547
rect 768 19513 802 19547
rect 802 19513 811 19547
rect 759 19504 811 19513
rect 513 19429 565 19438
rect 513 19395 522 19429
rect 522 19395 556 19429
rect 556 19395 565 19429
rect 513 19386 565 19395
rect 639 19429 691 19438
rect 639 19395 648 19429
rect 648 19395 682 19429
rect 682 19395 691 19429
rect 639 19386 691 19395
rect 759 19429 811 19438
rect 759 19395 768 19429
rect 768 19395 802 19429
rect 802 19395 811 19429
rect 759 19386 811 19395
rect 21078 19391 21130 19400
rect 21078 19357 21087 19391
rect 21087 19357 21121 19391
rect 21121 19357 21130 19391
rect 21078 19348 21130 19357
rect 21204 19391 21256 19400
rect 21204 19357 21213 19391
rect 21213 19357 21247 19391
rect 21247 19357 21256 19391
rect 21204 19348 21256 19357
rect 21324 19391 21376 19400
rect 21324 19357 21333 19391
rect 21333 19357 21367 19391
rect 21367 19357 21376 19391
rect 21324 19348 21376 19357
rect 21078 19273 21130 19282
rect 21078 19239 21087 19273
rect 21087 19239 21121 19273
rect 21121 19239 21130 19273
rect 21078 19230 21130 19239
rect 21204 19273 21256 19282
rect 21204 19239 21213 19273
rect 21213 19239 21247 19273
rect 21247 19239 21256 19273
rect 21204 19230 21256 19239
rect 21324 19273 21376 19282
rect 21324 19239 21333 19273
rect 21333 19239 21367 19273
rect 21367 19239 21376 19273
rect 21324 19230 21376 19239
rect 514 19039 566 19048
rect 514 19005 523 19039
rect 523 19005 557 19039
rect 557 19005 566 19039
rect 514 18996 566 19005
rect 636 19039 688 19048
rect 636 19005 645 19039
rect 645 19005 679 19039
rect 679 19005 688 19039
rect 636 18996 688 19005
rect 762 19039 814 19048
rect 762 19005 771 19039
rect 771 19005 805 19039
rect 805 19005 814 19039
rect 762 18996 814 19005
rect 514 18892 566 18901
rect 514 18858 523 18892
rect 523 18858 557 18892
rect 557 18858 566 18892
rect 514 18849 566 18858
rect 636 18892 688 18901
rect 636 18858 645 18892
rect 645 18858 679 18892
rect 679 18858 688 18892
rect 636 18849 688 18858
rect 762 18892 814 18901
rect 762 18858 771 18892
rect 771 18858 805 18892
rect 805 18858 814 18892
rect 762 18849 814 18858
rect 514 18755 566 18764
rect 514 18721 523 18755
rect 523 18721 557 18755
rect 557 18721 566 18755
rect 514 18712 566 18721
rect 636 18755 688 18764
rect 636 18721 645 18755
rect 645 18721 679 18755
rect 679 18721 688 18755
rect 636 18712 688 18721
rect 762 18755 814 18764
rect 762 18721 771 18755
rect 771 18721 805 18755
rect 805 18721 814 18755
rect 762 18712 814 18721
rect 22020 18053 22072 18062
rect 22020 18019 22029 18053
rect 22029 18019 22063 18053
rect 22063 18019 22072 18053
rect 22020 18010 22072 18019
rect 22146 18053 22198 18062
rect 22146 18019 22155 18053
rect 22155 18019 22189 18053
rect 22189 18019 22198 18053
rect 22146 18010 22198 18019
rect 22266 18053 22318 18062
rect 22266 18019 22275 18053
rect 22275 18019 22309 18053
rect 22309 18019 22318 18053
rect 22266 18010 22318 18019
rect 22020 17935 22072 17944
rect 22020 17901 22029 17935
rect 22029 17901 22063 17935
rect 22063 17901 22072 17935
rect 22020 17892 22072 17901
rect 22146 17935 22198 17944
rect 22146 17901 22155 17935
rect 22155 17901 22189 17935
rect 22189 17901 22198 17935
rect 22146 17892 22198 17901
rect 22266 17935 22318 17944
rect 22266 17901 22275 17935
rect 22275 17901 22309 17935
rect 22309 17901 22318 17935
rect 22266 17892 22318 17901
rect 514 17279 566 17288
rect 514 17245 523 17279
rect 523 17245 557 17279
rect 557 17245 566 17279
rect 514 17236 566 17245
rect 636 17279 688 17288
rect 636 17245 645 17279
rect 645 17245 679 17279
rect 679 17245 688 17279
rect 636 17236 688 17245
rect 762 17279 814 17288
rect 762 17245 771 17279
rect 771 17245 805 17279
rect 805 17245 814 17279
rect 762 17236 814 17245
rect 514 17132 566 17141
rect 514 17098 523 17132
rect 523 17098 557 17132
rect 557 17098 566 17132
rect 514 17089 566 17098
rect 636 17132 688 17141
rect 636 17098 645 17132
rect 645 17098 679 17132
rect 679 17098 688 17132
rect 636 17089 688 17098
rect 762 17132 814 17141
rect 762 17098 771 17132
rect 771 17098 805 17132
rect 805 17098 814 17132
rect 762 17089 814 17098
rect 514 16995 566 17004
rect 514 16961 523 16995
rect 523 16961 557 16995
rect 557 16961 566 16995
rect 514 16952 566 16961
rect 636 16995 688 17004
rect 636 16961 645 16995
rect 645 16961 679 16995
rect 679 16961 688 16995
rect 636 16952 688 16961
rect 762 16995 814 17004
rect 762 16961 771 16995
rect 771 16961 805 16995
rect 805 16961 814 16995
rect 762 16952 814 16961
rect 513 16681 565 16690
rect 513 16647 522 16681
rect 522 16647 556 16681
rect 556 16647 565 16681
rect 513 16638 565 16647
rect 639 16681 691 16690
rect 639 16647 648 16681
rect 648 16647 682 16681
rect 682 16647 691 16681
rect 639 16638 691 16647
rect 759 16681 811 16690
rect 759 16647 768 16681
rect 768 16647 802 16681
rect 802 16647 811 16681
rect 759 16638 811 16647
rect 513 16563 565 16572
rect 513 16529 522 16563
rect 522 16529 556 16563
rect 556 16529 565 16563
rect 513 16520 565 16529
rect 639 16563 691 16572
rect 639 16529 648 16563
rect 648 16529 682 16563
rect 682 16529 691 16563
rect 639 16520 691 16529
rect 759 16563 811 16572
rect 759 16529 768 16563
rect 768 16529 802 16563
rect 802 16529 811 16563
rect 759 16520 811 16529
rect 21078 16630 21130 16639
rect 21078 16596 21087 16630
rect 21087 16596 21121 16630
rect 21121 16596 21130 16630
rect 21078 16587 21130 16596
rect 21204 16630 21256 16639
rect 21204 16596 21213 16630
rect 21213 16596 21247 16630
rect 21247 16596 21256 16630
rect 21204 16587 21256 16596
rect 21324 16630 21376 16639
rect 21324 16596 21333 16630
rect 21333 16596 21367 16630
rect 21367 16596 21376 16630
rect 21324 16587 21376 16596
rect 21078 16512 21130 16521
rect 21078 16478 21087 16512
rect 21087 16478 21121 16512
rect 21121 16478 21130 16512
rect 21078 16469 21130 16478
rect 21204 16512 21256 16521
rect 21204 16478 21213 16512
rect 21213 16478 21247 16512
rect 21247 16478 21256 16512
rect 21204 16469 21256 16478
rect 21324 16512 21376 16521
rect 21324 16478 21333 16512
rect 21333 16478 21367 16512
rect 21367 16478 21376 16512
rect 21324 16469 21376 16478
rect 513 15465 565 15474
rect 513 15431 522 15465
rect 522 15431 556 15465
rect 556 15431 565 15465
rect 513 15422 565 15431
rect 639 15465 691 15474
rect 639 15431 648 15465
rect 648 15431 682 15465
rect 682 15431 691 15465
rect 639 15422 691 15431
rect 759 15465 811 15474
rect 759 15431 768 15465
rect 768 15431 802 15465
rect 802 15431 811 15465
rect 759 15422 811 15431
rect 513 15347 565 15356
rect 513 15313 522 15347
rect 522 15313 556 15347
rect 556 15313 565 15347
rect 513 15304 565 15313
rect 639 15347 691 15356
rect 639 15313 648 15347
rect 648 15313 682 15347
rect 682 15313 691 15347
rect 639 15304 691 15313
rect 759 15347 811 15356
rect 759 15313 768 15347
rect 768 15313 802 15347
rect 802 15313 811 15347
rect 759 15304 811 15313
rect 21078 15416 21130 15425
rect 21078 15382 21087 15416
rect 21087 15382 21121 15416
rect 21121 15382 21130 15416
rect 21078 15373 21130 15382
rect 21204 15416 21256 15425
rect 21204 15382 21213 15416
rect 21213 15382 21247 15416
rect 21247 15382 21256 15416
rect 21204 15373 21256 15382
rect 21324 15416 21376 15425
rect 21324 15382 21333 15416
rect 21333 15382 21367 15416
rect 21367 15382 21376 15416
rect 21324 15373 21376 15382
rect 21078 15298 21130 15307
rect 21078 15264 21087 15298
rect 21087 15264 21121 15298
rect 21121 15264 21130 15298
rect 21078 15255 21130 15264
rect 21204 15298 21256 15307
rect 21204 15264 21213 15298
rect 21213 15264 21247 15298
rect 21247 15264 21256 15298
rect 21204 15255 21256 15264
rect 21324 15298 21376 15307
rect 21324 15264 21333 15298
rect 21333 15264 21367 15298
rect 21367 15264 21376 15298
rect 21324 15255 21376 15264
rect 514 15039 566 15048
rect 514 15005 523 15039
rect 523 15005 557 15039
rect 557 15005 566 15039
rect 514 14996 566 15005
rect 636 15039 688 15048
rect 636 15005 645 15039
rect 645 15005 679 15039
rect 679 15005 688 15039
rect 636 14996 688 15005
rect 762 15039 814 15048
rect 762 15005 771 15039
rect 771 15005 805 15039
rect 805 15005 814 15039
rect 762 14996 814 15005
rect 514 14892 566 14901
rect 514 14858 523 14892
rect 523 14858 557 14892
rect 557 14858 566 14892
rect 514 14849 566 14858
rect 636 14892 688 14901
rect 636 14858 645 14892
rect 645 14858 679 14892
rect 679 14858 688 14892
rect 636 14849 688 14858
rect 762 14892 814 14901
rect 762 14858 771 14892
rect 771 14858 805 14892
rect 805 14858 814 14892
rect 762 14849 814 14858
rect 514 14755 566 14764
rect 514 14721 523 14755
rect 523 14721 557 14755
rect 557 14721 566 14755
rect 514 14712 566 14721
rect 636 14755 688 14764
rect 636 14721 645 14755
rect 645 14721 679 14755
rect 679 14721 688 14755
rect 636 14712 688 14721
rect 762 14755 814 14764
rect 762 14721 771 14755
rect 771 14721 805 14755
rect 805 14721 814 14755
rect 762 14712 814 14721
rect 22020 14235 22072 14244
rect 22020 14201 22029 14235
rect 22029 14201 22063 14235
rect 22063 14201 22072 14235
rect 22020 14192 22072 14201
rect 22146 14235 22198 14244
rect 22146 14201 22155 14235
rect 22155 14201 22189 14235
rect 22189 14201 22198 14235
rect 22146 14192 22198 14201
rect 22266 14235 22318 14244
rect 22266 14201 22275 14235
rect 22275 14201 22309 14235
rect 22309 14201 22318 14235
rect 22266 14192 22318 14201
rect 22020 14117 22072 14126
rect 22020 14083 22029 14117
rect 22029 14083 22063 14117
rect 22063 14083 22072 14117
rect 22020 14074 22072 14083
rect 22146 14117 22198 14126
rect 22146 14083 22155 14117
rect 22155 14083 22189 14117
rect 22189 14083 22198 14117
rect 22146 14074 22198 14083
rect 22266 14117 22318 14126
rect 22266 14083 22275 14117
rect 22275 14083 22309 14117
rect 22309 14083 22318 14117
rect 22266 14074 22318 14083
rect 514 13279 566 13288
rect 514 13245 523 13279
rect 523 13245 557 13279
rect 557 13245 566 13279
rect 514 13236 566 13245
rect 636 13279 688 13288
rect 636 13245 645 13279
rect 645 13245 679 13279
rect 679 13245 688 13279
rect 636 13236 688 13245
rect 762 13279 814 13288
rect 762 13245 771 13279
rect 771 13245 805 13279
rect 805 13245 814 13279
rect 762 13236 814 13245
rect 514 13132 566 13141
rect 514 13098 523 13132
rect 523 13098 557 13132
rect 557 13098 566 13132
rect 514 13089 566 13098
rect 636 13132 688 13141
rect 636 13098 645 13132
rect 645 13098 679 13132
rect 679 13098 688 13132
rect 636 13089 688 13098
rect 762 13132 814 13141
rect 762 13098 771 13132
rect 771 13098 805 13132
rect 805 13098 814 13132
rect 762 13089 814 13098
rect 514 12995 566 13004
rect 514 12961 523 12995
rect 523 12961 557 12995
rect 557 12961 566 12995
rect 514 12952 566 12961
rect 636 12995 688 13004
rect 636 12961 645 12995
rect 645 12961 679 12995
rect 679 12961 688 12995
rect 636 12952 688 12961
rect 762 12995 814 13004
rect 762 12961 771 12995
rect 771 12961 805 12995
rect 805 12961 814 12995
rect 762 12952 814 12961
rect 513 12600 565 12609
rect 513 12566 522 12600
rect 522 12566 556 12600
rect 556 12566 565 12600
rect 513 12557 565 12566
rect 639 12600 691 12609
rect 639 12566 648 12600
rect 648 12566 682 12600
rect 682 12566 691 12600
rect 639 12557 691 12566
rect 759 12600 811 12609
rect 759 12566 768 12600
rect 768 12566 802 12600
rect 802 12566 811 12600
rect 759 12557 811 12566
rect 513 12482 565 12491
rect 513 12448 522 12482
rect 522 12448 556 12482
rect 556 12448 565 12482
rect 513 12439 565 12448
rect 639 12482 691 12491
rect 639 12448 648 12482
rect 648 12448 682 12482
rect 682 12448 691 12482
rect 639 12439 691 12448
rect 759 12482 811 12491
rect 759 12448 768 12482
rect 768 12448 802 12482
rect 802 12448 811 12482
rect 759 12439 811 12448
rect 21078 12573 21130 12582
rect 21078 12539 21087 12573
rect 21087 12539 21121 12573
rect 21121 12539 21130 12573
rect 21078 12530 21130 12539
rect 21204 12573 21256 12582
rect 21204 12539 21213 12573
rect 21213 12539 21247 12573
rect 21247 12539 21256 12573
rect 21204 12530 21256 12539
rect 21324 12573 21376 12582
rect 21324 12539 21333 12573
rect 21333 12539 21367 12573
rect 21367 12539 21376 12573
rect 21324 12530 21376 12539
rect 21078 12455 21130 12464
rect 21078 12421 21087 12455
rect 21087 12421 21121 12455
rect 21121 12421 21130 12455
rect 21078 12412 21130 12421
rect 21204 12455 21256 12464
rect 21204 12421 21213 12455
rect 21213 12421 21247 12455
rect 21247 12421 21256 12455
rect 21204 12412 21256 12421
rect 21324 12455 21376 12464
rect 21324 12421 21333 12455
rect 21333 12421 21367 12455
rect 21367 12421 21376 12455
rect 21324 12412 21376 12421
rect 513 11478 565 11487
rect 513 11444 522 11478
rect 522 11444 556 11478
rect 556 11444 565 11478
rect 513 11435 565 11444
rect 639 11478 691 11487
rect 639 11444 648 11478
rect 648 11444 682 11478
rect 682 11444 691 11478
rect 639 11435 691 11444
rect 759 11478 811 11487
rect 759 11444 768 11478
rect 768 11444 802 11478
rect 802 11444 811 11478
rect 759 11435 811 11444
rect 513 11360 565 11369
rect 513 11326 522 11360
rect 522 11326 556 11360
rect 556 11326 565 11360
rect 513 11317 565 11326
rect 639 11360 691 11369
rect 639 11326 648 11360
rect 648 11326 682 11360
rect 682 11326 691 11360
rect 639 11317 691 11326
rect 759 11360 811 11369
rect 759 11326 768 11360
rect 768 11326 802 11360
rect 802 11326 811 11360
rect 759 11317 811 11326
rect 21078 11416 21130 11425
rect 21078 11382 21087 11416
rect 21087 11382 21121 11416
rect 21121 11382 21130 11416
rect 21078 11373 21130 11382
rect 21204 11416 21256 11425
rect 21204 11382 21213 11416
rect 21213 11382 21247 11416
rect 21247 11382 21256 11416
rect 21204 11373 21256 11382
rect 21324 11416 21376 11425
rect 21324 11382 21333 11416
rect 21333 11382 21367 11416
rect 21367 11382 21376 11416
rect 21324 11373 21376 11382
rect 21078 11298 21130 11307
rect 21078 11264 21087 11298
rect 21087 11264 21121 11298
rect 21121 11264 21130 11298
rect 21078 11255 21130 11264
rect 21204 11298 21256 11307
rect 21204 11264 21213 11298
rect 21213 11264 21247 11298
rect 21247 11264 21256 11298
rect 21204 11255 21256 11264
rect 21324 11298 21376 11307
rect 21324 11264 21333 11298
rect 21333 11264 21367 11298
rect 21367 11264 21376 11298
rect 21324 11255 21376 11264
rect 514 11040 566 11049
rect 514 11006 523 11040
rect 523 11006 557 11040
rect 557 11006 566 11040
rect 514 10997 566 11006
rect 636 11040 688 11049
rect 636 11006 645 11040
rect 645 11006 679 11040
rect 679 11006 688 11040
rect 636 10997 688 11006
rect 762 11040 814 11049
rect 762 11006 771 11040
rect 771 11006 805 11040
rect 805 11006 814 11040
rect 762 10997 814 11006
rect 514 10893 566 10902
rect 514 10859 523 10893
rect 523 10859 557 10893
rect 557 10859 566 10893
rect 514 10850 566 10859
rect 636 10893 688 10902
rect 636 10859 645 10893
rect 645 10859 679 10893
rect 679 10859 688 10893
rect 636 10850 688 10859
rect 762 10893 814 10902
rect 762 10859 771 10893
rect 771 10859 805 10893
rect 805 10859 814 10893
rect 762 10850 814 10859
rect 514 10756 566 10765
rect 514 10722 523 10756
rect 523 10722 557 10756
rect 557 10722 566 10756
rect 514 10713 566 10722
rect 636 10756 688 10765
rect 636 10722 645 10756
rect 645 10722 679 10756
rect 679 10722 688 10756
rect 636 10713 688 10722
rect 762 10756 814 10765
rect 762 10722 771 10756
rect 771 10722 805 10756
rect 805 10722 814 10756
rect 762 10713 814 10722
rect 22020 10271 22072 10280
rect 22020 10237 22029 10271
rect 22029 10237 22063 10271
rect 22063 10237 22072 10271
rect 22020 10228 22072 10237
rect 22146 10271 22198 10280
rect 22146 10237 22155 10271
rect 22155 10237 22189 10271
rect 22189 10237 22198 10271
rect 22146 10228 22198 10237
rect 22266 10271 22318 10280
rect 22266 10237 22275 10271
rect 22275 10237 22309 10271
rect 22309 10237 22318 10271
rect 22266 10228 22318 10237
rect 22020 10153 22072 10162
rect 22020 10119 22029 10153
rect 22029 10119 22063 10153
rect 22063 10119 22072 10153
rect 22020 10110 22072 10119
rect 22146 10153 22198 10162
rect 22146 10119 22155 10153
rect 22155 10119 22189 10153
rect 22189 10119 22198 10153
rect 22146 10110 22198 10119
rect 22266 10153 22318 10162
rect 22266 10119 22275 10153
rect 22275 10119 22309 10153
rect 22309 10119 22318 10153
rect 22266 10110 22318 10119
rect 514 9278 566 9287
rect 514 9244 523 9278
rect 523 9244 557 9278
rect 557 9244 566 9278
rect 514 9235 566 9244
rect 636 9278 688 9287
rect 636 9244 645 9278
rect 645 9244 679 9278
rect 679 9244 688 9278
rect 636 9235 688 9244
rect 762 9278 814 9287
rect 762 9244 771 9278
rect 771 9244 805 9278
rect 805 9244 814 9278
rect 762 9235 814 9244
rect 514 9131 566 9140
rect 514 9097 523 9131
rect 523 9097 557 9131
rect 557 9097 566 9131
rect 514 9088 566 9097
rect 636 9131 688 9140
rect 636 9097 645 9131
rect 645 9097 679 9131
rect 679 9097 688 9131
rect 636 9088 688 9097
rect 762 9131 814 9140
rect 762 9097 771 9131
rect 771 9097 805 9131
rect 805 9097 814 9131
rect 762 9088 814 9097
rect 514 8994 566 9003
rect 514 8960 523 8994
rect 523 8960 557 8994
rect 557 8960 566 8994
rect 514 8951 566 8960
rect 636 8994 688 9003
rect 636 8960 645 8994
rect 645 8960 679 8994
rect 679 8960 688 8994
rect 636 8951 688 8960
rect 762 8994 814 9003
rect 762 8960 771 8994
rect 771 8960 805 8994
rect 805 8960 814 8994
rect 762 8951 814 8960
rect 513 8618 565 8627
rect 513 8584 522 8618
rect 522 8584 556 8618
rect 556 8584 565 8618
rect 513 8575 565 8584
rect 639 8618 691 8627
rect 639 8584 648 8618
rect 648 8584 682 8618
rect 682 8584 691 8618
rect 639 8575 691 8584
rect 759 8618 811 8627
rect 759 8584 768 8618
rect 768 8584 802 8618
rect 802 8584 811 8618
rect 759 8575 811 8584
rect 513 8500 565 8509
rect 513 8466 522 8500
rect 522 8466 556 8500
rect 556 8466 565 8500
rect 513 8457 565 8466
rect 639 8500 691 8509
rect 639 8466 648 8500
rect 648 8466 682 8500
rect 682 8466 691 8500
rect 639 8457 691 8466
rect 759 8500 811 8509
rect 759 8466 768 8500
rect 768 8466 802 8500
rect 802 8466 811 8500
rect 759 8457 811 8466
rect 21078 8573 21130 8582
rect 21078 8539 21087 8573
rect 21087 8539 21121 8573
rect 21121 8539 21130 8573
rect 21078 8530 21130 8539
rect 21204 8573 21256 8582
rect 21204 8539 21213 8573
rect 21213 8539 21247 8573
rect 21247 8539 21256 8573
rect 21204 8530 21256 8539
rect 21324 8573 21376 8582
rect 21324 8539 21333 8573
rect 21333 8539 21367 8573
rect 21367 8539 21376 8573
rect 21324 8530 21376 8539
rect 21078 8455 21130 8464
rect 21078 8421 21087 8455
rect 21087 8421 21121 8455
rect 21121 8421 21130 8455
rect 21078 8412 21130 8421
rect 21204 8455 21256 8464
rect 21204 8421 21213 8455
rect 21213 8421 21247 8455
rect 21247 8421 21256 8455
rect 21204 8412 21256 8421
rect 21324 8455 21376 8464
rect 21324 8421 21333 8455
rect 21333 8421 21367 8455
rect 21367 8421 21376 8455
rect 21324 8412 21376 8421
rect 513 7507 565 7516
rect 513 7473 522 7507
rect 522 7473 556 7507
rect 556 7473 565 7507
rect 513 7464 565 7473
rect 639 7507 691 7516
rect 639 7473 648 7507
rect 648 7473 682 7507
rect 682 7473 691 7507
rect 639 7464 691 7473
rect 759 7507 811 7516
rect 759 7473 768 7507
rect 768 7473 802 7507
rect 802 7473 811 7507
rect 759 7464 811 7473
rect 513 7389 565 7398
rect 513 7355 522 7389
rect 522 7355 556 7389
rect 556 7355 565 7389
rect 513 7346 565 7355
rect 639 7389 691 7398
rect 639 7355 648 7389
rect 648 7355 682 7389
rect 682 7355 691 7389
rect 639 7346 691 7355
rect 759 7389 811 7398
rect 759 7355 768 7389
rect 768 7355 802 7389
rect 802 7355 811 7389
rect 759 7346 811 7355
rect 21078 7416 21130 7425
rect 21078 7382 21087 7416
rect 21087 7382 21121 7416
rect 21121 7382 21130 7416
rect 21078 7373 21130 7382
rect 21204 7416 21256 7425
rect 21204 7382 21213 7416
rect 21213 7382 21247 7416
rect 21247 7382 21256 7416
rect 21204 7373 21256 7382
rect 21324 7416 21376 7425
rect 21324 7382 21333 7416
rect 21333 7382 21367 7416
rect 21367 7382 21376 7416
rect 21324 7373 21376 7382
rect 21078 7298 21130 7307
rect 21078 7264 21087 7298
rect 21087 7264 21121 7298
rect 21121 7264 21130 7298
rect 21078 7255 21130 7264
rect 21204 7298 21256 7307
rect 21204 7264 21213 7298
rect 21213 7264 21247 7298
rect 21247 7264 21256 7298
rect 21204 7255 21256 7264
rect 21324 7298 21376 7307
rect 21324 7264 21333 7298
rect 21333 7264 21367 7298
rect 21367 7264 21376 7298
rect 21324 7255 21376 7264
rect 514 7040 566 7049
rect 514 7006 523 7040
rect 523 7006 557 7040
rect 557 7006 566 7040
rect 514 6997 566 7006
rect 636 7040 688 7049
rect 636 7006 645 7040
rect 645 7006 679 7040
rect 679 7006 688 7040
rect 636 6997 688 7006
rect 762 7040 814 7049
rect 762 7006 771 7040
rect 771 7006 805 7040
rect 805 7006 814 7040
rect 762 6997 814 7006
rect 514 6893 566 6902
rect 514 6859 523 6893
rect 523 6859 557 6893
rect 557 6859 566 6893
rect 514 6850 566 6859
rect 636 6893 688 6902
rect 636 6859 645 6893
rect 645 6859 679 6893
rect 679 6859 688 6893
rect 636 6850 688 6859
rect 762 6893 814 6902
rect 762 6859 771 6893
rect 771 6859 805 6893
rect 805 6859 814 6893
rect 762 6850 814 6859
rect 514 6756 566 6765
rect 514 6722 523 6756
rect 523 6722 557 6756
rect 557 6722 566 6756
rect 514 6713 566 6722
rect 636 6756 688 6765
rect 636 6722 645 6756
rect 645 6722 679 6756
rect 679 6722 688 6756
rect 636 6713 688 6722
rect 762 6756 814 6765
rect 762 6722 771 6756
rect 771 6722 805 6756
rect 805 6722 814 6756
rect 762 6713 814 6722
rect 22020 6259 22072 6268
rect 22020 6225 22029 6259
rect 22029 6225 22063 6259
rect 22063 6225 22072 6259
rect 22020 6216 22072 6225
rect 22146 6259 22198 6268
rect 22146 6225 22155 6259
rect 22155 6225 22189 6259
rect 22189 6225 22198 6259
rect 22146 6216 22198 6225
rect 22266 6259 22318 6268
rect 22266 6225 22275 6259
rect 22275 6225 22309 6259
rect 22309 6225 22318 6259
rect 22266 6216 22318 6225
rect 22020 6141 22072 6150
rect 22020 6107 22029 6141
rect 22029 6107 22063 6141
rect 22063 6107 22072 6141
rect 22020 6098 22072 6107
rect 22146 6141 22198 6150
rect 22146 6107 22155 6141
rect 22155 6107 22189 6141
rect 22189 6107 22198 6141
rect 22146 6098 22198 6107
rect 22266 6141 22318 6150
rect 22266 6107 22275 6141
rect 22275 6107 22309 6141
rect 22309 6107 22318 6141
rect 22266 6098 22318 6107
rect 514 5279 566 5288
rect 514 5245 523 5279
rect 523 5245 557 5279
rect 557 5245 566 5279
rect 514 5236 566 5245
rect 636 5279 688 5288
rect 636 5245 645 5279
rect 645 5245 679 5279
rect 679 5245 688 5279
rect 636 5236 688 5245
rect 762 5279 814 5288
rect 762 5245 771 5279
rect 771 5245 805 5279
rect 805 5245 814 5279
rect 762 5236 814 5245
rect 514 5132 566 5141
rect 514 5098 523 5132
rect 523 5098 557 5132
rect 557 5098 566 5132
rect 514 5089 566 5098
rect 636 5132 688 5141
rect 636 5098 645 5132
rect 645 5098 679 5132
rect 679 5098 688 5132
rect 636 5089 688 5098
rect 762 5132 814 5141
rect 762 5098 771 5132
rect 771 5098 805 5132
rect 805 5098 814 5132
rect 762 5089 814 5098
rect 514 4995 566 5004
rect 514 4961 523 4995
rect 523 4961 557 4995
rect 557 4961 566 4995
rect 514 4952 566 4961
rect 636 4995 688 5004
rect 636 4961 645 4995
rect 645 4961 679 4995
rect 679 4961 688 4995
rect 636 4952 688 4961
rect 762 4995 814 5004
rect 762 4961 771 4995
rect 771 4961 805 4995
rect 805 4961 814 4995
rect 762 4952 814 4961
rect 513 4684 565 4693
rect 513 4650 522 4684
rect 522 4650 556 4684
rect 556 4650 565 4684
rect 513 4641 565 4650
rect 639 4684 691 4693
rect 639 4650 648 4684
rect 648 4650 682 4684
rect 682 4650 691 4684
rect 639 4641 691 4650
rect 759 4684 811 4693
rect 759 4650 768 4684
rect 768 4650 802 4684
rect 802 4650 811 4684
rect 759 4641 811 4650
rect 513 4566 565 4575
rect 513 4532 522 4566
rect 522 4532 556 4566
rect 556 4532 565 4566
rect 513 4523 565 4532
rect 639 4566 691 4575
rect 639 4532 648 4566
rect 648 4532 682 4566
rect 682 4532 691 4566
rect 639 4523 691 4532
rect 759 4566 811 4575
rect 759 4532 768 4566
rect 768 4532 802 4566
rect 802 4532 811 4566
rect 759 4523 811 4532
rect 21078 4573 21130 4582
rect 21078 4539 21087 4573
rect 21087 4539 21121 4573
rect 21121 4539 21130 4573
rect 21078 4530 21130 4539
rect 21204 4573 21256 4582
rect 21204 4539 21213 4573
rect 21213 4539 21247 4573
rect 21247 4539 21256 4573
rect 21204 4530 21256 4539
rect 21324 4573 21376 4582
rect 21324 4539 21333 4573
rect 21333 4539 21367 4573
rect 21367 4539 21376 4573
rect 21324 4530 21376 4539
rect 21078 4455 21130 4464
rect 21078 4421 21087 4455
rect 21087 4421 21121 4455
rect 21121 4421 21130 4455
rect 21078 4412 21130 4421
rect 21204 4455 21256 4464
rect 21204 4421 21213 4455
rect 21213 4421 21247 4455
rect 21247 4421 21256 4455
rect 21204 4412 21256 4421
rect 21324 4455 21376 4464
rect 21324 4421 21333 4455
rect 21333 4421 21367 4455
rect 21367 4421 21376 4455
rect 21324 4412 21376 4421
rect 513 3507 565 3516
rect 513 3473 522 3507
rect 522 3473 556 3507
rect 556 3473 565 3507
rect 513 3464 565 3473
rect 639 3507 691 3516
rect 639 3473 648 3507
rect 648 3473 682 3507
rect 682 3473 691 3507
rect 639 3464 691 3473
rect 759 3507 811 3516
rect 759 3473 768 3507
rect 768 3473 802 3507
rect 802 3473 811 3507
rect 759 3464 811 3473
rect 513 3389 565 3398
rect 513 3355 522 3389
rect 522 3355 556 3389
rect 556 3355 565 3389
rect 513 3346 565 3355
rect 639 3389 691 3398
rect 639 3355 648 3389
rect 648 3355 682 3389
rect 682 3355 691 3389
rect 639 3346 691 3355
rect 759 3389 811 3398
rect 759 3355 768 3389
rect 768 3355 802 3389
rect 802 3355 811 3389
rect 759 3346 811 3355
rect 21078 3416 21130 3425
rect 21078 3382 21087 3416
rect 21087 3382 21121 3416
rect 21121 3382 21130 3416
rect 21078 3373 21130 3382
rect 21204 3416 21256 3425
rect 21204 3382 21213 3416
rect 21213 3382 21247 3416
rect 21247 3382 21256 3416
rect 21204 3373 21256 3382
rect 21324 3416 21376 3425
rect 21324 3382 21333 3416
rect 21333 3382 21367 3416
rect 21367 3382 21376 3416
rect 21324 3373 21376 3382
rect 21078 3298 21130 3307
rect 21078 3264 21087 3298
rect 21087 3264 21121 3298
rect 21121 3264 21130 3298
rect 21078 3255 21130 3264
rect 21204 3298 21256 3307
rect 21204 3264 21213 3298
rect 21213 3264 21247 3298
rect 21247 3264 21256 3298
rect 21204 3255 21256 3264
rect 21324 3298 21376 3307
rect 21324 3264 21333 3298
rect 21333 3264 21367 3298
rect 21367 3264 21376 3298
rect 21324 3255 21376 3264
rect 514 3040 566 3049
rect 514 3006 523 3040
rect 523 3006 557 3040
rect 557 3006 566 3040
rect 514 2997 566 3006
rect 636 3040 688 3049
rect 636 3006 645 3040
rect 645 3006 679 3040
rect 679 3006 688 3040
rect 636 2997 688 3006
rect 762 3040 814 3049
rect 762 3006 771 3040
rect 771 3006 805 3040
rect 805 3006 814 3040
rect 762 2997 814 3006
rect 514 2893 566 2902
rect 514 2859 523 2893
rect 523 2859 557 2893
rect 557 2859 566 2893
rect 514 2850 566 2859
rect 636 2893 688 2902
rect 636 2859 645 2893
rect 645 2859 679 2893
rect 679 2859 688 2893
rect 636 2850 688 2859
rect 762 2893 814 2902
rect 762 2859 771 2893
rect 771 2859 805 2893
rect 805 2859 814 2893
rect 762 2850 814 2859
rect 514 2756 566 2765
rect 514 2722 523 2756
rect 523 2722 557 2756
rect 557 2722 566 2756
rect 514 2713 566 2722
rect 636 2756 688 2765
rect 636 2722 645 2756
rect 645 2722 679 2756
rect 679 2722 688 2756
rect 636 2713 688 2722
rect 762 2756 814 2765
rect 762 2722 771 2756
rect 771 2722 805 2756
rect 805 2722 814 2756
rect 762 2713 814 2722
rect 22020 2259 22072 2268
rect 22020 2225 22029 2259
rect 22029 2225 22063 2259
rect 22063 2225 22072 2259
rect 22020 2216 22072 2225
rect 22146 2259 22198 2268
rect 22146 2225 22155 2259
rect 22155 2225 22189 2259
rect 22189 2225 22198 2259
rect 22146 2216 22198 2225
rect 22266 2259 22318 2268
rect 22266 2225 22275 2259
rect 22275 2225 22309 2259
rect 22309 2225 22318 2259
rect 22266 2216 22318 2225
rect 22020 2141 22072 2150
rect 22020 2107 22029 2141
rect 22029 2107 22063 2141
rect 22063 2107 22072 2141
rect 22020 2098 22072 2107
rect 22146 2141 22198 2150
rect 22146 2107 22155 2141
rect 22155 2107 22189 2141
rect 22189 2107 22198 2141
rect 22146 2098 22198 2107
rect 22266 2141 22318 2150
rect 22266 2107 22275 2141
rect 22275 2107 22309 2141
rect 22309 2107 22318 2141
rect 22266 2098 22318 2107
rect 514 1279 566 1288
rect 514 1245 523 1279
rect 523 1245 557 1279
rect 557 1245 566 1279
rect 514 1236 566 1245
rect 636 1279 688 1288
rect 636 1245 645 1279
rect 645 1245 679 1279
rect 679 1245 688 1279
rect 636 1236 688 1245
rect 762 1279 814 1288
rect 762 1245 771 1279
rect 771 1245 805 1279
rect 805 1245 814 1279
rect 762 1236 814 1245
rect 514 1132 566 1141
rect 514 1098 523 1132
rect 523 1098 557 1132
rect 557 1098 566 1132
rect 514 1089 566 1098
rect 636 1132 688 1141
rect 636 1098 645 1132
rect 645 1098 679 1132
rect 679 1098 688 1132
rect 636 1089 688 1098
rect 762 1132 814 1141
rect 762 1098 771 1132
rect 771 1098 805 1132
rect 805 1098 814 1132
rect 762 1089 814 1098
rect 514 995 566 1004
rect 514 961 523 995
rect 523 961 557 995
rect 557 961 566 995
rect 514 952 566 961
rect 636 995 688 1004
rect 636 961 645 995
rect 645 961 679 995
rect 679 961 688 995
rect 636 952 688 961
rect 762 995 814 1004
rect 762 961 771 995
rect 771 961 805 995
rect 805 961 814 995
rect 762 952 814 961
rect 513 684 565 693
rect 513 650 522 684
rect 522 650 556 684
rect 556 650 565 684
rect 513 641 565 650
rect 639 684 691 693
rect 639 650 648 684
rect 648 650 682 684
rect 682 650 691 684
rect 639 641 691 650
rect 759 684 811 693
rect 759 650 768 684
rect 768 650 802 684
rect 802 650 811 684
rect 759 641 811 650
rect 513 566 565 575
rect 513 532 522 566
rect 522 532 556 566
rect 556 532 565 566
rect 513 523 565 532
rect 639 566 691 575
rect 639 532 648 566
rect 648 532 682 566
rect 682 532 691 566
rect 639 523 691 532
rect 759 566 811 575
rect 759 532 768 566
rect 768 532 802 566
rect 802 532 811 566
rect 759 523 811 532
rect 21078 573 21130 582
rect 21078 539 21087 573
rect 21087 539 21121 573
rect 21121 539 21130 573
rect 21078 530 21130 539
rect 21204 573 21256 582
rect 21204 539 21213 573
rect 21213 539 21247 573
rect 21247 539 21256 573
rect 21204 530 21256 539
rect 21324 573 21376 582
rect 21324 539 21333 573
rect 21333 539 21367 573
rect 21367 539 21376 573
rect 21324 530 21376 539
rect 21078 455 21130 464
rect 21078 421 21087 455
rect 21087 421 21121 455
rect 21121 421 21130 455
rect 21078 412 21130 421
rect 21204 455 21256 464
rect 21204 421 21213 455
rect 21213 421 21247 455
rect 21247 421 21256 455
rect 21204 412 21256 421
rect 21324 455 21376 464
rect 21324 421 21333 455
rect 21333 421 21367 455
rect 21367 421 21376 455
rect 21324 412 21376 421
<< metal2 >>
rect 21026 75482 21426 75517
rect 463 75442 864 75477
rect 463 75386 511 75442
rect 567 75386 637 75442
rect 693 75386 757 75442
rect 813 75386 864 75442
rect 463 75324 864 75386
rect 463 75268 511 75324
rect 567 75268 637 75324
rect 693 75268 757 75324
rect 813 75268 864 75324
rect 463 75222 864 75268
rect 21026 75426 21076 75482
rect 21132 75426 21202 75482
rect 21258 75426 21322 75482
rect 21378 75426 21426 75482
rect 21026 75364 21426 75426
rect 21026 75308 21076 75364
rect 21132 75308 21202 75364
rect 21258 75308 21322 75364
rect 21378 75308 21426 75364
rect 21026 75262 21426 75308
rect 463 75050 863 75109
rect 463 74994 512 75050
rect 568 74994 634 75050
rect 690 74994 760 75050
rect 816 74994 863 75050
rect 463 74903 863 74994
rect 463 74847 512 74903
rect 568 74847 634 74903
rect 690 74847 760 74903
rect 816 74847 863 74903
rect 463 74766 863 74847
rect 463 74710 512 74766
rect 568 74710 634 74766
rect 690 74710 760 74766
rect 816 74710 863 74766
rect 463 74650 863 74710
rect 21970 74061 22370 74096
rect 21970 74005 22018 74061
rect 22074 74005 22144 74061
rect 22200 74005 22264 74061
rect 22320 74005 22370 74061
rect 21970 73943 22370 74005
rect 21970 73887 22018 73943
rect 22074 73887 22144 73943
rect 22200 73887 22264 73943
rect 22320 73887 22370 73943
rect 21970 73841 22370 73887
rect 463 73290 863 73349
rect 463 73234 512 73290
rect 568 73234 634 73290
rect 690 73234 760 73290
rect 816 73234 863 73290
rect 463 73143 863 73234
rect 463 73087 512 73143
rect 568 73087 634 73143
rect 690 73087 760 73143
rect 816 73087 863 73143
rect 463 73006 863 73087
rect 463 72950 512 73006
rect 568 72950 634 73006
rect 690 72950 760 73006
rect 816 72950 863 73006
rect 463 72890 863 72950
rect 463 72769 864 72804
rect 463 72713 511 72769
rect 567 72713 637 72769
rect 693 72713 757 72769
rect 813 72713 864 72769
rect 463 72651 864 72713
rect 463 72595 511 72651
rect 567 72595 637 72651
rect 693 72595 757 72651
rect 813 72595 864 72651
rect 463 72549 864 72595
rect 21028 72685 21428 72720
rect 21028 72629 21076 72685
rect 21132 72629 21202 72685
rect 21258 72629 21322 72685
rect 21378 72629 21428 72685
rect 21028 72567 21428 72629
rect 21028 72511 21076 72567
rect 21132 72511 21202 72567
rect 21258 72511 21322 72567
rect 21378 72511 21428 72567
rect 21028 72465 21428 72511
rect 21026 71482 21426 71517
rect 463 71442 864 71477
rect 463 71386 511 71442
rect 567 71386 637 71442
rect 693 71386 757 71442
rect 813 71386 864 71442
rect 463 71324 864 71386
rect 463 71268 511 71324
rect 567 71268 637 71324
rect 693 71268 757 71324
rect 813 71268 864 71324
rect 463 71222 864 71268
rect 21026 71426 21076 71482
rect 21132 71426 21202 71482
rect 21258 71426 21322 71482
rect 21378 71426 21426 71482
rect 21026 71364 21426 71426
rect 21026 71308 21076 71364
rect 21132 71308 21202 71364
rect 21258 71308 21322 71364
rect 21378 71308 21426 71364
rect 21026 71262 21426 71308
rect 463 71050 863 71109
rect 463 70994 512 71050
rect 568 70994 634 71050
rect 690 70994 760 71050
rect 816 70994 863 71050
rect 463 70903 863 70994
rect 463 70847 512 70903
rect 568 70847 634 70903
rect 690 70847 760 70903
rect 816 70847 863 70903
rect 463 70766 863 70847
rect 463 70710 512 70766
rect 568 70710 634 70766
rect 690 70710 760 70766
rect 816 70710 863 70766
rect 463 70650 863 70710
rect 21970 70061 22370 70096
rect 21970 70005 22018 70061
rect 22074 70005 22144 70061
rect 22200 70005 22264 70061
rect 22320 70005 22370 70061
rect 21970 69943 22370 70005
rect 21970 69887 22018 69943
rect 22074 69887 22144 69943
rect 22200 69887 22264 69943
rect 22320 69887 22370 69943
rect 21970 69841 22370 69887
rect 463 69290 863 69349
rect 463 69234 512 69290
rect 568 69234 634 69290
rect 690 69234 760 69290
rect 816 69234 863 69290
rect 463 69143 863 69234
rect 463 69087 512 69143
rect 568 69087 634 69143
rect 690 69087 760 69143
rect 816 69087 863 69143
rect 463 69006 863 69087
rect 463 68950 512 69006
rect 568 68950 634 69006
rect 690 68950 760 69006
rect 816 68950 863 69006
rect 463 68890 863 68950
rect 463 68769 864 68804
rect 463 68713 511 68769
rect 567 68713 637 68769
rect 693 68713 757 68769
rect 813 68713 864 68769
rect 463 68651 864 68713
rect 463 68595 511 68651
rect 567 68595 637 68651
rect 693 68595 757 68651
rect 813 68595 864 68651
rect 463 68549 864 68595
rect 21028 68685 21428 68720
rect 21028 68629 21076 68685
rect 21132 68629 21202 68685
rect 21258 68629 21322 68685
rect 21378 68629 21428 68685
rect 21028 68567 21428 68629
rect 21028 68511 21076 68567
rect 21132 68511 21202 68567
rect 21258 68511 21322 68567
rect 21378 68511 21428 68567
rect 21028 68465 21428 68511
rect 21026 67482 21426 67517
rect 463 67440 864 67475
rect 463 67384 511 67440
rect 567 67384 637 67440
rect 693 67384 757 67440
rect 813 67384 864 67440
rect 463 67322 864 67384
rect 463 67266 511 67322
rect 567 67266 637 67322
rect 693 67266 757 67322
rect 813 67266 864 67322
rect 463 67220 864 67266
rect 21026 67426 21076 67482
rect 21132 67426 21202 67482
rect 21258 67426 21322 67482
rect 21378 67426 21426 67482
rect 21026 67364 21426 67426
rect 21026 67308 21076 67364
rect 21132 67308 21202 67364
rect 21258 67308 21322 67364
rect 21378 67308 21426 67364
rect 21026 67262 21426 67308
rect 463 67050 863 67109
rect 463 66994 512 67050
rect 568 66994 634 67050
rect 690 66994 760 67050
rect 816 66994 863 67050
rect 463 66903 863 66994
rect 463 66847 512 66903
rect 568 66847 634 66903
rect 690 66847 760 66903
rect 816 66847 863 66903
rect 463 66766 863 66847
rect 463 66710 512 66766
rect 568 66710 634 66766
rect 690 66710 760 66766
rect 816 66710 863 66766
rect 463 66650 863 66710
rect 21970 66048 22370 66083
rect 21970 65992 22018 66048
rect 22074 65992 22144 66048
rect 22200 65992 22264 66048
rect 22320 65992 22370 66048
rect 21970 65930 22370 65992
rect 21970 65874 22018 65930
rect 22074 65874 22144 65930
rect 22200 65874 22264 65930
rect 22320 65874 22370 65930
rect 21970 65828 22370 65874
rect 463 65291 863 65350
rect 463 65235 512 65291
rect 568 65235 634 65291
rect 690 65235 760 65291
rect 816 65235 863 65291
rect 463 65144 863 65235
rect 463 65088 512 65144
rect 568 65088 634 65144
rect 690 65088 760 65144
rect 816 65088 863 65144
rect 463 65007 863 65088
rect 463 64951 512 65007
rect 568 64951 634 65007
rect 690 64951 760 65007
rect 816 64951 863 65007
rect 463 64891 863 64951
rect 463 64700 864 64735
rect 463 64644 511 64700
rect 567 64644 637 64700
rect 693 64644 757 64700
rect 813 64644 864 64700
rect 463 64582 864 64644
rect 463 64526 511 64582
rect 567 64526 637 64582
rect 693 64526 757 64582
rect 813 64526 864 64582
rect 463 64480 864 64526
rect 21028 64685 21428 64720
rect 21028 64629 21076 64685
rect 21132 64629 21202 64685
rect 21258 64629 21322 64685
rect 21378 64629 21428 64685
rect 21028 64567 21428 64629
rect 21028 64511 21076 64567
rect 21132 64511 21202 64567
rect 21258 64511 21322 64567
rect 21378 64511 21428 64567
rect 21028 64465 21428 64511
rect 463 63522 864 63557
rect 463 63466 511 63522
rect 567 63466 637 63522
rect 693 63466 757 63522
rect 813 63466 864 63522
rect 463 63404 864 63466
rect 463 63348 511 63404
rect 567 63348 637 63404
rect 693 63348 757 63404
rect 813 63348 864 63404
rect 463 63302 864 63348
rect 21026 63482 21426 63517
rect 21026 63426 21076 63482
rect 21132 63426 21202 63482
rect 21258 63426 21322 63482
rect 21378 63426 21426 63482
rect 21026 63364 21426 63426
rect 21026 63308 21076 63364
rect 21132 63308 21202 63364
rect 21258 63308 21322 63364
rect 21378 63308 21426 63364
rect 21026 63262 21426 63308
rect 464 63068 864 63109
rect 463 63050 864 63068
rect 463 62994 512 63050
rect 568 62994 634 63050
rect 690 62994 760 63050
rect 816 62994 864 63050
rect 463 62903 864 62994
rect 463 62847 512 62903
rect 568 62847 634 62903
rect 690 62847 760 62903
rect 816 62847 864 62903
rect 463 62766 864 62847
rect 463 62710 512 62766
rect 568 62710 634 62766
rect 690 62710 760 62766
rect 816 62710 864 62766
rect 463 62650 864 62710
rect 21970 62047 22370 62082
rect 21970 61991 22018 62047
rect 22074 61991 22144 62047
rect 22200 61991 22264 62047
rect 22320 61991 22370 62047
rect 21970 61929 22370 61991
rect 21970 61873 22018 61929
rect 22074 61873 22144 61929
rect 22200 61873 22264 61929
rect 22320 61873 22370 61929
rect 21970 61827 22370 61873
rect 463 61291 863 61350
rect 463 61235 512 61291
rect 568 61235 634 61291
rect 690 61235 760 61291
rect 816 61235 863 61291
rect 463 61144 863 61235
rect 463 61088 512 61144
rect 568 61088 634 61144
rect 690 61088 760 61144
rect 816 61088 863 61144
rect 463 61007 863 61088
rect 463 60951 512 61007
rect 568 60951 634 61007
rect 690 60951 760 61007
rect 816 60951 863 61007
rect 463 60891 863 60951
rect 463 60674 866 60709
rect 463 60618 511 60674
rect 567 60618 637 60674
rect 693 60618 757 60674
rect 813 60618 866 60674
rect 463 60556 866 60618
rect 463 60500 511 60556
rect 567 60500 637 60556
rect 693 60500 757 60556
rect 813 60500 866 60556
rect 463 60454 866 60500
rect 21028 60685 21428 60720
rect 21028 60629 21076 60685
rect 21132 60629 21202 60685
rect 21258 60629 21322 60685
rect 21378 60629 21428 60685
rect 21028 60567 21428 60629
rect 21028 60511 21076 60567
rect 21132 60511 21202 60567
rect 21258 60511 21322 60567
rect 21378 60511 21428 60567
rect 21028 60465 21428 60511
rect 21027 59536 21427 59571
rect 463 59471 864 59506
rect 463 59415 511 59471
rect 567 59415 637 59471
rect 693 59415 757 59471
rect 813 59415 864 59471
rect 463 59353 864 59415
rect 463 59297 511 59353
rect 567 59297 637 59353
rect 693 59297 757 59353
rect 813 59297 864 59353
rect 21027 59480 21076 59536
rect 21132 59480 21202 59536
rect 21258 59480 21322 59536
rect 21378 59480 21427 59536
rect 21027 59418 21427 59480
rect 21027 59362 21076 59418
rect 21132 59362 21202 59418
rect 21258 59362 21322 59418
rect 21378 59362 21427 59418
rect 21027 59316 21427 59362
rect 463 59251 864 59297
rect 464 59068 864 59109
rect 463 59050 864 59068
rect 463 58994 512 59050
rect 568 58994 634 59050
rect 690 58994 760 59050
rect 816 58994 864 59050
rect 463 58903 864 58994
rect 463 58847 512 58903
rect 568 58847 634 58903
rect 690 58847 760 58903
rect 816 58847 864 58903
rect 463 58766 864 58847
rect 463 58710 512 58766
rect 568 58710 634 58766
rect 690 58710 760 58766
rect 816 58710 864 58766
rect 463 58650 864 58710
rect 21970 58086 22370 58121
rect 21970 58030 22018 58086
rect 22074 58030 22144 58086
rect 22200 58030 22264 58086
rect 22320 58030 22370 58086
rect 21970 57968 22370 58030
rect 21970 57912 22018 57968
rect 22074 57912 22144 57968
rect 22200 57912 22264 57968
rect 22320 57912 22370 57968
rect 21970 57866 22370 57912
rect 463 57289 863 57348
rect 463 57233 512 57289
rect 568 57233 634 57289
rect 690 57233 760 57289
rect 816 57233 863 57289
rect 463 57142 863 57233
rect 463 57086 512 57142
rect 568 57086 634 57142
rect 690 57086 760 57142
rect 816 57086 863 57142
rect 463 57005 863 57086
rect 463 56949 512 57005
rect 568 56949 634 57005
rect 690 56949 760 57005
rect 816 56949 863 57005
rect 463 56889 863 56949
rect 463 56694 864 56729
rect 463 56638 511 56694
rect 567 56638 637 56694
rect 693 56638 757 56694
rect 813 56638 864 56694
rect 463 56576 864 56638
rect 463 56520 511 56576
rect 567 56520 637 56576
rect 693 56520 757 56576
rect 813 56520 864 56576
rect 463 56474 864 56520
rect 21028 56620 21428 56655
rect 21028 56564 21076 56620
rect 21132 56564 21202 56620
rect 21258 56564 21322 56620
rect 21378 56564 21428 56620
rect 21028 56502 21428 56564
rect 21028 56446 21076 56502
rect 21132 56446 21202 56502
rect 21258 56446 21322 56502
rect 21378 56446 21428 56502
rect 21028 56400 21428 56446
rect 463 55487 866 55522
rect 463 55431 511 55487
rect 567 55431 637 55487
rect 693 55431 757 55487
rect 813 55431 866 55487
rect 463 55369 866 55431
rect 463 55313 511 55369
rect 567 55313 637 55369
rect 693 55313 757 55369
rect 813 55313 866 55369
rect 463 55267 866 55313
rect 21027 55437 21427 55472
rect 21027 55381 21076 55437
rect 21132 55381 21202 55437
rect 21258 55381 21322 55437
rect 21378 55381 21427 55437
rect 21027 55319 21427 55381
rect 21027 55263 21076 55319
rect 21132 55263 21202 55319
rect 21258 55263 21322 55319
rect 21378 55263 21427 55319
rect 21027 55217 21427 55263
rect 463 55050 863 55109
rect 463 54994 512 55050
rect 568 54994 634 55050
rect 690 54994 760 55050
rect 816 54994 863 55050
rect 463 54903 863 54994
rect 463 54847 512 54903
rect 568 54847 634 54903
rect 690 54847 760 54903
rect 816 54847 863 54903
rect 463 54766 863 54847
rect 463 54710 512 54766
rect 568 54710 634 54766
rect 690 54710 760 54766
rect 816 54710 863 54766
rect 463 54650 863 54710
rect 21970 54069 22370 54104
rect 21970 54013 22018 54069
rect 22074 54013 22144 54069
rect 22200 54013 22264 54069
rect 22320 54013 22370 54069
rect 21970 53951 22370 54013
rect 21970 53895 22018 53951
rect 22074 53895 22144 53951
rect 22200 53895 22264 53951
rect 22320 53895 22370 53951
rect 21970 53849 22370 53895
rect 463 53291 863 53350
rect 463 53235 512 53291
rect 568 53235 634 53291
rect 690 53235 760 53291
rect 816 53235 863 53291
rect 463 53144 863 53235
rect 463 53088 512 53144
rect 568 53088 634 53144
rect 690 53088 760 53144
rect 816 53088 863 53144
rect 463 53007 863 53088
rect 463 52951 512 53007
rect 568 52951 634 53007
rect 690 52951 760 53007
rect 816 52951 863 53007
rect 463 52891 863 52951
rect 463 52721 864 52756
rect 463 52665 511 52721
rect 567 52665 637 52721
rect 693 52665 757 52721
rect 813 52665 864 52721
rect 463 52603 864 52665
rect 463 52547 511 52603
rect 567 52547 637 52603
rect 693 52547 757 52603
rect 813 52547 864 52603
rect 463 52501 864 52547
rect 21028 52565 21428 52600
rect 21028 52509 21076 52565
rect 21132 52509 21202 52565
rect 21258 52509 21322 52565
rect 21378 52509 21428 52565
rect 21028 52447 21428 52509
rect 21028 52391 21076 52447
rect 21132 52391 21202 52447
rect 21258 52391 21322 52447
rect 21378 52391 21428 52447
rect 21028 52345 21428 52391
rect 463 51534 864 51569
rect 463 51478 511 51534
rect 567 51478 637 51534
rect 693 51478 757 51534
rect 813 51478 864 51534
rect 463 51416 864 51478
rect 463 51360 511 51416
rect 567 51360 637 51416
rect 693 51360 757 51416
rect 813 51360 864 51416
rect 463 51314 864 51360
rect 21028 51430 21428 51465
rect 21028 51374 21076 51430
rect 21132 51374 21202 51430
rect 21258 51374 21322 51430
rect 21378 51374 21428 51430
rect 21028 51312 21428 51374
rect 21028 51256 21076 51312
rect 21132 51256 21202 51312
rect 21258 51256 21322 51312
rect 21378 51256 21428 51312
rect 21028 51210 21428 51256
rect 463 51050 863 51109
rect 463 50994 512 51050
rect 568 50994 634 51050
rect 690 50994 760 51050
rect 816 50994 863 51050
rect 463 50903 863 50994
rect 463 50847 512 50903
rect 568 50847 634 50903
rect 690 50847 760 50903
rect 816 50847 863 50903
rect 463 50766 863 50847
rect 463 50710 512 50766
rect 568 50710 634 50766
rect 690 50710 760 50766
rect 816 50710 863 50766
rect 463 50650 863 50710
rect 21970 50148 22370 50183
rect 21970 50092 22018 50148
rect 22074 50092 22144 50148
rect 22200 50092 22264 50148
rect 22320 50092 22370 50148
rect 21970 50030 22370 50092
rect 21970 49974 22018 50030
rect 22074 49974 22144 50030
rect 22200 49974 22264 50030
rect 22320 49974 22370 50030
rect 21970 49928 22370 49974
rect 463 49291 863 49350
rect 463 49235 512 49291
rect 568 49235 634 49291
rect 690 49235 760 49291
rect 816 49235 863 49291
rect 463 49144 863 49235
rect 463 49088 512 49144
rect 568 49088 634 49144
rect 690 49088 760 49144
rect 816 49088 863 49144
rect 463 49007 863 49088
rect 463 48951 512 49007
rect 568 48951 634 49007
rect 690 48951 760 49007
rect 816 48951 863 49007
rect 463 48891 863 48951
rect 463 48712 864 48747
rect 463 48656 511 48712
rect 567 48656 637 48712
rect 693 48656 757 48712
rect 813 48656 864 48712
rect 463 48594 864 48656
rect 463 48538 511 48594
rect 567 48538 637 48594
rect 693 48538 757 48594
rect 813 48538 864 48594
rect 463 48492 864 48538
rect 21028 48671 21428 48706
rect 21028 48615 21076 48671
rect 21132 48615 21202 48671
rect 21258 48615 21322 48671
rect 21378 48615 21428 48671
rect 21028 48553 21428 48615
rect 21028 48497 21076 48553
rect 21132 48497 21202 48553
rect 21258 48497 21322 48553
rect 21378 48497 21428 48553
rect 21028 48451 21428 48497
rect 463 47559 864 47594
rect 463 47503 511 47559
rect 567 47503 637 47559
rect 693 47503 757 47559
rect 813 47503 864 47559
rect 463 47441 864 47503
rect 463 47385 511 47441
rect 567 47385 637 47441
rect 693 47385 757 47441
rect 813 47385 864 47441
rect 463 47339 864 47385
rect 21028 47518 21428 47553
rect 21028 47462 21076 47518
rect 21132 47462 21202 47518
rect 21258 47462 21322 47518
rect 21378 47462 21428 47518
rect 21028 47400 21428 47462
rect 21028 47344 21076 47400
rect 21132 47344 21202 47400
rect 21258 47344 21322 47400
rect 21378 47344 21428 47400
rect 21028 47298 21428 47344
rect 463 47050 863 47109
rect 463 46994 512 47050
rect 568 46994 634 47050
rect 690 46994 760 47050
rect 816 46994 863 47050
rect 463 46903 863 46994
rect 463 46847 512 46903
rect 568 46847 634 46903
rect 690 46847 760 46903
rect 816 46847 863 46903
rect 463 46766 863 46847
rect 463 46710 512 46766
rect 568 46710 634 46766
rect 690 46710 760 46766
rect 816 46710 863 46766
rect 463 46650 863 46710
rect 21970 45890 22370 45925
rect 21970 45834 22018 45890
rect 22074 45834 22144 45890
rect 22200 45834 22264 45890
rect 22320 45834 22370 45890
rect 21970 45772 22370 45834
rect 21970 45716 22018 45772
rect 22074 45716 22144 45772
rect 22200 45716 22264 45772
rect 22320 45716 22370 45772
rect 21970 45670 22370 45716
rect 463 45290 863 45350
rect 463 45234 512 45290
rect 568 45234 634 45290
rect 690 45234 760 45290
rect 816 45234 863 45290
rect 463 45143 863 45234
rect 463 45087 512 45143
rect 568 45087 634 45143
rect 690 45087 760 45143
rect 816 45087 863 45143
rect 463 45006 863 45087
rect 463 44950 512 45006
rect 568 44950 634 45006
rect 690 44950 760 45006
rect 816 44950 863 45006
rect 463 44891 863 44950
rect 463 44890 836 44891
rect 463 44499 863 44534
rect 463 44443 511 44499
rect 567 44443 637 44499
rect 693 44443 757 44499
rect 813 44443 863 44499
rect 463 44381 863 44443
rect 463 44325 511 44381
rect 567 44325 637 44381
rect 693 44325 757 44381
rect 813 44325 863 44381
rect 463 44279 863 44325
rect 21028 44402 21428 44437
rect 21028 44346 21076 44402
rect 21132 44346 21202 44402
rect 21258 44346 21322 44402
rect 21378 44346 21428 44402
rect 21028 44284 21428 44346
rect 21028 44228 21076 44284
rect 21132 44228 21202 44284
rect 21258 44228 21322 44284
rect 21378 44228 21428 44284
rect 21028 44182 21428 44228
rect 1650 39925 2398 39940
rect 1650 39789 2257 39925
rect 2393 39789 2398 39925
rect 1650 39776 2398 39789
rect 1650 39774 2396 39776
rect 0 39729 400 39752
rect 0 39673 44 39729
rect 100 39673 169 39729
rect 225 39673 294 39729
rect 350 39673 400 39729
rect 0 39623 400 39673
rect 0 39567 44 39623
rect 100 39567 169 39623
rect 225 39567 294 39623
rect 350 39567 400 39623
rect 0 39528 400 39567
rect 1411 39320 1569 39333
rect 1411 39319 1498 39320
rect 1411 39263 1416 39319
rect 1472 39264 1498 39319
rect 1554 39264 1569 39320
rect 1472 39263 1569 39264
rect 1411 39240 1569 39263
rect 1411 39239 1499 39240
rect 1411 39183 1417 39239
rect 1473 39184 1499 39239
rect 1555 39184 1569 39240
rect 1650 39321 1796 39774
rect 2468 39711 2867 44000
rect 21970 43824 22370 43870
rect 21970 43528 22044 43824
rect 22260 43528 22370 43824
rect 21970 43480 22370 43528
rect 3352 39904 3502 39919
rect 3352 39768 3361 39904
rect 3497 39768 3502 39904
rect 3352 39755 3502 39768
rect 3352 39754 3500 39755
rect 1867 39438 2868 39711
rect 1650 39269 1662 39321
rect 1714 39269 1732 39321
rect 1784 39269 1796 39321
rect 1650 39251 1796 39269
rect 1650 39199 1662 39251
rect 1714 39199 1732 39251
rect 1784 39199 1796 39251
rect 1650 39189 1796 39199
rect 1868 39410 2267 39438
rect 1868 39364 2335 39410
rect 1868 39312 1886 39364
rect 1938 39312 1950 39364
rect 2002 39312 2042 39364
rect 2094 39312 2106 39364
rect 2158 39312 2198 39364
rect 2250 39312 2262 39364
rect 2314 39312 2335 39364
rect 1868 39270 2335 39312
rect 2538 39328 2685 39336
rect 2538 39276 2551 39328
rect 2603 39276 2621 39328
rect 2673 39276 2685 39328
rect 1473 39183 1569 39184
rect 1411 39169 1569 39183
rect 463 39119 805 39139
rect 463 39063 492 39119
rect 548 39063 606 39119
rect 662 39063 720 39119
rect 776 39063 805 39119
rect 463 39043 805 39063
rect 1495 38774 1569 39169
rect 1495 38722 1507 38774
rect 1559 38722 1569 38774
rect 1495 38717 1569 38722
rect 0 38575 342 38595
rect 0 38519 29 38575
rect 85 38519 143 38575
rect 199 38519 257 38575
rect 313 38519 342 38575
rect 0 38499 342 38519
rect 1471 38269 1523 38275
rect 1471 38211 1523 38217
rect 463 38031 805 38051
rect 463 37975 492 38031
rect 548 37975 606 38031
rect 662 37975 720 38031
rect 776 37975 805 38031
rect 463 37955 805 37975
rect 1471 37797 1504 38211
rect 1463 37790 1515 37797
rect 1463 37732 1515 37738
rect 0 37487 342 37507
rect 0 37431 29 37487
rect 85 37431 143 37487
rect 199 37431 257 37487
rect 313 37431 342 37487
rect 0 37411 342 37431
rect 1680 37358 1739 39189
rect 1680 37306 1683 37358
rect 1735 37306 1739 37358
rect 1680 37252 1739 37306
rect 1680 37200 1683 37252
rect 1735 37200 1739 37252
rect 1680 37187 1739 37200
rect 463 36943 805 36963
rect 463 36887 492 36943
rect 548 36887 606 36943
rect 662 36887 720 36943
rect 776 36887 805 36943
rect 463 36867 805 36887
rect 1868 32936 2267 39270
rect 2538 39258 2685 39276
rect 2538 39206 2551 39258
rect 2603 39206 2621 39258
rect 2673 39206 2685 39258
rect 2751 39318 2899 39332
rect 2751 39262 2760 39318
rect 2816 39317 2899 39318
rect 2816 39262 2840 39317
rect 2751 39261 2840 39262
rect 2896 39261 2899 39317
rect 2751 39253 2899 39261
rect 2538 36830 2685 39206
rect 2538 36778 2551 36830
rect 2603 36778 2621 36830
rect 2673 36778 2685 36830
rect 2538 36763 2685 36778
rect 2538 36711 2551 36763
rect 2603 36711 2621 36763
rect 2673 36711 2685 36763
rect 2538 36476 2685 36711
rect 2752 39237 2899 39253
rect 2752 39181 2761 39237
rect 2817 39181 2841 39237
rect 2897 39181 2899 39237
rect 2752 36830 2899 39181
rect 3352 39317 3499 39754
rect 21502 39714 21902 39752
rect 21502 39658 21547 39714
rect 21603 39658 21672 39714
rect 21728 39658 21797 39714
rect 21853 39658 21902 39714
rect 21502 39594 21902 39658
rect 21502 39538 21546 39594
rect 21602 39538 21671 39594
rect 21727 39538 21796 39594
rect 21852 39538 21902 39594
rect 21502 39497 21902 39538
rect 3352 39261 3360 39317
rect 3416 39316 3499 39317
rect 3416 39261 3440 39316
rect 3352 39260 3440 39261
rect 3496 39260 3499 39316
rect 3352 39236 3499 39260
rect 3352 39180 3361 39236
rect 3417 39180 3441 39236
rect 3497 39180 3499 39236
rect 3352 39169 3499 39180
rect 3523 38828 3529 38880
rect 3581 38828 3587 38880
rect 4610 38879 4704 38885
rect 3537 37897 3568 38828
rect 4662 38827 4704 38879
rect 4610 38821 4704 38827
rect 3608 38348 3660 38354
rect 3608 38290 3660 38296
rect 3517 37845 3523 37897
rect 3575 37845 3581 37897
rect 3620 37185 3649 38290
rect 4652 38267 4704 38821
rect 4652 38209 4704 38215
rect 4652 37791 4704 37797
rect 4652 37187 4704 37739
rect 3536 37182 3649 37185
rect 3536 37130 3553 37182
rect 3605 37130 3649 37182
rect 3536 37126 3649 37130
rect 4609 37181 4704 37187
rect 4661 37129 4704 37181
rect 4609 37123 4704 37129
rect 2752 36778 2765 36830
rect 2817 36778 2835 36830
rect 2887 36778 2899 36830
rect 2752 36765 2899 36778
rect 2752 36713 2765 36765
rect 2817 36713 2835 36765
rect 2887 36713 2899 36765
rect 2752 36707 2899 36713
rect 21970 36940 22370 36986
rect 21970 36644 22044 36940
rect 22260 36644 22370 36940
rect 21970 36596 22370 36644
rect 2535 36475 2685 36476
rect 2535 36460 2689 36475
rect 2535 36404 2544 36460
rect 2600 36404 2624 36460
rect 2680 36404 2689 36460
rect 2535 36391 2689 36404
rect 21028 36160 21428 36198
rect 21028 36104 21073 36160
rect 21129 36104 21198 36160
rect 21254 36104 21323 36160
rect 21379 36104 21428 36160
rect 21028 36040 21428 36104
rect 21028 35984 21072 36040
rect 21128 35984 21197 36040
rect 21253 35984 21322 36040
rect 21378 35984 21428 36040
rect 21028 35943 21428 35984
rect 21028 35582 21428 35642
rect 21028 35526 21077 35582
rect 21133 35526 21199 35582
rect 21255 35526 21325 35582
rect 21381 35526 21428 35582
rect 21028 35435 21428 35526
rect 21028 35379 21077 35435
rect 21133 35379 21199 35435
rect 21255 35379 21325 35435
rect 21381 35379 21428 35435
rect 21028 35298 21428 35379
rect 21028 35242 21077 35298
rect 21133 35242 21199 35298
rect 21255 35242 21325 35298
rect 21381 35242 21428 35298
rect 21028 35183 21428 35242
rect 21028 35182 21401 35183
rect 20527 34664 20927 34702
rect 20527 34608 20572 34664
rect 20628 34608 20697 34664
rect 20753 34608 20822 34664
rect 20878 34608 20927 34664
rect 20527 34544 20927 34608
rect 20527 34488 20571 34544
rect 20627 34488 20696 34544
rect 20752 34488 20821 34544
rect 20877 34488 20927 34544
rect 20527 34447 20927 34488
rect 21502 34664 21902 34702
rect 21502 34608 21547 34664
rect 21603 34608 21672 34664
rect 21728 34608 21797 34664
rect 21853 34608 21902 34664
rect 21502 34544 21902 34608
rect 21502 34488 21546 34544
rect 21602 34488 21671 34544
rect 21727 34488 21796 34544
rect 21852 34488 21902 34544
rect 21502 34447 21902 34488
rect 21028 33822 21428 33882
rect 21028 33766 21077 33822
rect 21133 33766 21199 33822
rect 21255 33766 21325 33822
rect 21381 33766 21428 33822
rect 21028 33675 21428 33766
rect 21028 33619 21077 33675
rect 21133 33619 21199 33675
rect 21255 33619 21325 33675
rect 21381 33619 21428 33675
rect 21028 33538 21428 33619
rect 21028 33482 21077 33538
rect 21133 33482 21199 33538
rect 21255 33482 21325 33538
rect 21381 33482 21428 33538
rect 21028 33423 21428 33482
rect 21028 33422 21401 33423
rect 21027 33105 21427 33143
rect 21027 33049 21072 33105
rect 21128 33049 21197 33105
rect 21253 33049 21322 33105
rect 21378 33049 21427 33105
rect 21027 32985 21427 33049
rect 1868 32710 2742 32936
rect 21027 32929 21071 32985
rect 21127 32929 21196 32985
rect 21252 32929 21321 32985
rect 21377 32929 21427 32985
rect 21027 32888 21427 32929
rect 1866 32485 2742 32710
rect 463 32292 866 32360
rect 463 32236 511 32292
rect 567 32236 637 32292
rect 693 32236 757 32292
rect 813 32236 866 32292
rect 463 32174 866 32236
rect 463 32118 511 32174
rect 567 32118 637 32174
rect 693 32118 757 32174
rect 813 32118 866 32174
rect 463 32072 866 32118
rect 2306 31967 2742 32485
rect 21025 32292 21428 32360
rect 21025 32236 21076 32292
rect 21132 32236 21202 32292
rect 21258 32236 21322 32292
rect 21378 32236 21428 32292
rect 21025 32174 21428 32236
rect 21025 32118 21076 32174
rect 21132 32118 21202 32174
rect 21258 32118 21322 32174
rect 21378 32118 21428 32174
rect 21025 32072 21428 32118
rect 463 31510 863 31545
rect 463 31454 511 31510
rect 567 31454 637 31510
rect 693 31454 757 31510
rect 813 31454 863 31510
rect 463 31392 863 31454
rect 463 31336 511 31392
rect 567 31336 637 31392
rect 693 31336 757 31392
rect 813 31336 863 31392
rect 463 31290 863 31336
rect 21028 31510 21428 31545
rect 21028 31454 21076 31510
rect 21132 31454 21202 31510
rect 21258 31454 21322 31510
rect 21378 31454 21428 31510
rect 21028 31392 21428 31454
rect 21028 31336 21076 31392
rect 21132 31336 21202 31392
rect 21258 31336 21322 31392
rect 21378 31336 21428 31392
rect 21028 31290 21428 31336
rect 463 31051 863 31111
rect 463 30995 512 31051
rect 568 30995 634 31051
rect 690 30995 760 31051
rect 816 30995 863 31051
rect 463 30904 863 30995
rect 463 30848 512 30904
rect 568 30848 634 30904
rect 690 30848 760 30904
rect 816 30848 863 30904
rect 463 30767 863 30848
rect 463 30711 512 30767
rect 568 30711 634 30767
rect 690 30711 760 30767
rect 816 30711 863 30767
rect 463 30651 863 30711
rect 21970 30120 22370 30155
rect 21970 30064 22018 30120
rect 22074 30064 22144 30120
rect 22200 30064 22264 30120
rect 22320 30064 22370 30120
rect 21970 30002 22370 30064
rect 21970 29946 22018 30002
rect 22074 29946 22144 30002
rect 22200 29946 22264 30002
rect 22320 29946 22370 30002
rect 21970 29900 22370 29946
rect 463 29284 863 29349
rect 463 29228 512 29284
rect 568 29228 634 29284
rect 690 29228 760 29284
rect 816 29228 863 29284
rect 463 29137 863 29228
rect 463 29081 512 29137
rect 568 29081 634 29137
rect 690 29081 760 29137
rect 816 29081 863 29137
rect 463 29000 863 29081
rect 463 28944 512 29000
rect 568 28944 634 29000
rect 690 28944 760 29000
rect 816 28944 863 29000
rect 463 28890 863 28944
rect 463 28598 863 28633
rect 463 28542 511 28598
rect 567 28542 637 28598
rect 693 28542 757 28598
rect 813 28542 863 28598
rect 463 28480 863 28542
rect 463 28424 511 28480
rect 567 28424 637 28480
rect 693 28424 757 28480
rect 813 28424 863 28480
rect 463 28378 863 28424
rect 21028 28549 21428 28584
rect 21028 28493 21076 28549
rect 21132 28493 21202 28549
rect 21258 28493 21322 28549
rect 21378 28493 21428 28549
rect 21028 28431 21428 28493
rect 21028 28375 21076 28431
rect 21132 28375 21202 28431
rect 21258 28375 21322 28431
rect 21378 28375 21428 28431
rect 21028 28329 21428 28375
rect 463 27594 863 27629
rect 463 27538 511 27594
rect 567 27538 637 27594
rect 693 27538 757 27594
rect 813 27538 863 27594
rect 463 27476 863 27538
rect 463 27420 511 27476
rect 567 27420 637 27476
rect 693 27420 757 27476
rect 813 27420 863 27476
rect 463 27374 863 27420
rect 21027 27432 21427 27467
rect 21027 27376 21076 27432
rect 21132 27376 21202 27432
rect 21258 27376 21322 27432
rect 21378 27376 21427 27432
rect 21027 27314 21427 27376
rect 21027 27258 21076 27314
rect 21132 27258 21202 27314
rect 21258 27258 21322 27314
rect 21378 27258 21427 27314
rect 21027 27212 21427 27258
rect 463 27050 863 27109
rect 463 26994 512 27050
rect 568 26994 634 27050
rect 690 26994 760 27050
rect 816 26994 863 27050
rect 463 26903 863 26994
rect 463 26847 512 26903
rect 568 26847 634 26903
rect 690 26847 760 26903
rect 816 26847 863 26903
rect 463 26766 863 26847
rect 463 26710 512 26766
rect 568 26710 634 26766
rect 690 26710 760 26766
rect 816 26710 863 26766
rect 463 26650 863 26710
rect 21970 25961 22370 25996
rect 21970 25905 22018 25961
rect 22074 25905 22144 25961
rect 22200 25905 22264 25961
rect 22320 25905 22370 25961
rect 21970 25843 22370 25905
rect 21970 25787 22018 25843
rect 22074 25787 22144 25843
rect 22200 25787 22264 25843
rect 22320 25787 22370 25843
rect 21970 25741 22370 25787
rect 463 25290 863 25349
rect 463 25234 512 25290
rect 568 25234 634 25290
rect 690 25234 760 25290
rect 816 25234 863 25290
rect 463 25143 863 25234
rect 463 25087 512 25143
rect 568 25087 634 25143
rect 690 25087 760 25143
rect 816 25087 863 25143
rect 463 25006 863 25087
rect 463 24950 512 25006
rect 568 24950 634 25006
rect 690 24950 760 25006
rect 816 24950 863 25006
rect 463 24890 863 24950
rect 463 24616 864 24651
rect 463 24560 511 24616
rect 567 24560 637 24616
rect 693 24560 757 24616
rect 813 24560 864 24616
rect 463 24498 864 24560
rect 463 24442 511 24498
rect 567 24442 637 24498
rect 693 24442 757 24498
rect 813 24442 864 24498
rect 463 24396 864 24442
rect 21028 24589 21428 24624
rect 21028 24533 21076 24589
rect 21132 24533 21202 24589
rect 21258 24533 21322 24589
rect 21378 24533 21428 24589
rect 21028 24471 21428 24533
rect 21028 24415 21076 24471
rect 21132 24415 21202 24471
rect 21258 24415 21322 24471
rect 21378 24415 21428 24471
rect 21028 24369 21428 24415
rect 463 23534 864 23569
rect 463 23478 511 23534
rect 567 23478 637 23534
rect 693 23478 757 23534
rect 813 23478 864 23534
rect 463 23416 864 23478
rect 463 23360 511 23416
rect 567 23360 637 23416
rect 693 23360 757 23416
rect 813 23360 864 23416
rect 463 23314 864 23360
rect 21028 23414 21428 23449
rect 21028 23358 21076 23414
rect 21132 23358 21202 23414
rect 21258 23358 21322 23414
rect 21378 23358 21428 23414
rect 21028 23296 21428 23358
rect 21028 23240 21076 23296
rect 21132 23240 21202 23296
rect 21258 23240 21322 23296
rect 21378 23240 21428 23296
rect 21028 23194 21428 23240
rect 463 23050 863 23109
rect 463 22994 512 23050
rect 568 22994 634 23050
rect 690 22994 760 23050
rect 816 22994 863 23050
rect 463 22903 863 22994
rect 463 22847 512 22903
rect 568 22847 634 22903
rect 690 22847 760 22903
rect 816 22847 863 22903
rect 463 22766 863 22847
rect 463 22710 512 22766
rect 568 22710 634 22766
rect 690 22710 760 22766
rect 816 22710 863 22766
rect 463 22650 863 22710
rect 21970 22171 22370 22206
rect 21970 22115 22018 22171
rect 22074 22115 22144 22171
rect 22200 22115 22264 22171
rect 22320 22115 22370 22171
rect 21970 22053 22370 22115
rect 21970 21997 22018 22053
rect 22074 21997 22144 22053
rect 22200 21997 22264 22053
rect 22320 21997 22370 22053
rect 21970 21951 22370 21997
rect 463 21291 863 21350
rect 463 21235 512 21291
rect 568 21235 634 21291
rect 690 21235 760 21291
rect 816 21235 863 21291
rect 463 21144 863 21235
rect 463 21088 512 21144
rect 568 21088 634 21144
rect 690 21088 760 21144
rect 816 21088 863 21144
rect 463 21007 863 21088
rect 463 20951 512 21007
rect 568 20951 634 21007
rect 690 20951 760 21007
rect 816 20951 863 21007
rect 463 20891 863 20951
rect 463 20659 864 20694
rect 463 20603 511 20659
rect 567 20603 637 20659
rect 693 20603 757 20659
rect 813 20603 864 20659
rect 463 20541 864 20603
rect 463 20485 511 20541
rect 567 20485 637 20541
rect 693 20485 757 20541
rect 813 20485 864 20541
rect 463 20439 864 20485
rect 21027 20573 21427 20608
rect 21027 20517 21076 20573
rect 21132 20517 21202 20573
rect 21258 20517 21322 20573
rect 21378 20517 21427 20573
rect 21027 20455 21427 20517
rect 21027 20399 21076 20455
rect 21132 20399 21202 20455
rect 21258 20399 21322 20455
rect 21378 20399 21427 20455
rect 21027 20353 21427 20399
rect 463 19558 864 19593
rect 463 19502 511 19558
rect 567 19502 637 19558
rect 693 19502 757 19558
rect 813 19502 864 19558
rect 463 19440 864 19502
rect 463 19384 511 19440
rect 567 19384 637 19440
rect 693 19384 757 19440
rect 813 19384 864 19440
rect 463 19338 864 19384
rect 21027 19402 21427 19437
rect 21027 19346 21076 19402
rect 21132 19346 21202 19402
rect 21258 19346 21322 19402
rect 21378 19346 21427 19402
rect 21027 19284 21427 19346
rect 21027 19228 21076 19284
rect 21132 19228 21202 19284
rect 21258 19228 21322 19284
rect 21378 19228 21427 19284
rect 21027 19182 21427 19228
rect 463 19050 863 19109
rect 463 18994 512 19050
rect 568 18994 634 19050
rect 690 18994 760 19050
rect 816 18994 863 19050
rect 463 18903 863 18994
rect 463 18847 512 18903
rect 568 18847 634 18903
rect 690 18847 760 18903
rect 816 18847 863 18903
rect 463 18766 863 18847
rect 463 18710 512 18766
rect 568 18710 634 18766
rect 690 18710 760 18766
rect 816 18710 863 18766
rect 463 18650 863 18710
rect 21970 18064 22370 18099
rect 21970 18008 22018 18064
rect 22074 18008 22144 18064
rect 22200 18008 22264 18064
rect 22320 18008 22370 18064
rect 21970 17946 22370 18008
rect 21970 17890 22018 17946
rect 22074 17890 22144 17946
rect 22200 17890 22264 17946
rect 22320 17890 22370 17946
rect 21970 17844 22370 17890
rect 463 17290 863 17349
rect 463 17234 512 17290
rect 568 17234 634 17290
rect 690 17234 760 17290
rect 816 17234 863 17290
rect 463 17143 863 17234
rect 463 17087 512 17143
rect 568 17087 634 17143
rect 690 17087 760 17143
rect 816 17087 863 17143
rect 463 17006 863 17087
rect 463 16950 512 17006
rect 568 16950 634 17006
rect 690 16950 760 17006
rect 816 16950 863 17006
rect 463 16890 863 16950
rect 463 16692 865 16727
rect 463 16636 511 16692
rect 567 16636 637 16692
rect 693 16636 757 16692
rect 813 16636 865 16692
rect 463 16574 865 16636
rect 463 16518 511 16574
rect 567 16518 637 16574
rect 693 16518 757 16574
rect 813 16518 865 16574
rect 463 16472 865 16518
rect 21027 16641 21427 16676
rect 21027 16585 21076 16641
rect 21132 16585 21202 16641
rect 21258 16585 21322 16641
rect 21378 16585 21427 16641
rect 21027 16523 21427 16585
rect 21027 16467 21076 16523
rect 21132 16467 21202 16523
rect 21258 16467 21322 16523
rect 21378 16467 21427 16523
rect 21027 16421 21427 16467
rect 463 15476 866 15511
rect 463 15420 511 15476
rect 567 15420 637 15476
rect 693 15420 757 15476
rect 813 15420 866 15476
rect 463 15358 866 15420
rect 463 15302 511 15358
rect 567 15302 637 15358
rect 693 15302 757 15358
rect 813 15302 866 15358
rect 463 15256 866 15302
rect 21027 15427 21427 15462
rect 21027 15371 21076 15427
rect 21132 15371 21202 15427
rect 21258 15371 21322 15427
rect 21378 15371 21427 15427
rect 21027 15309 21427 15371
rect 21027 15253 21076 15309
rect 21132 15253 21202 15309
rect 21258 15253 21322 15309
rect 21378 15253 21427 15309
rect 21027 15207 21427 15253
rect 463 15050 863 15109
rect 463 14994 512 15050
rect 568 14994 634 15050
rect 690 14994 760 15050
rect 816 14994 863 15050
rect 463 14903 863 14994
rect 463 14847 512 14903
rect 568 14847 634 14903
rect 690 14847 760 14903
rect 816 14847 863 14903
rect 463 14766 863 14847
rect 463 14710 512 14766
rect 568 14710 634 14766
rect 690 14710 760 14766
rect 816 14710 863 14766
rect 463 14650 863 14710
rect 21970 14246 22370 14281
rect 21970 14190 22018 14246
rect 22074 14190 22144 14246
rect 22200 14190 22264 14246
rect 22320 14190 22370 14246
rect 21970 14128 22370 14190
rect 21970 14072 22018 14128
rect 22074 14072 22144 14128
rect 22200 14072 22264 14128
rect 22320 14072 22370 14128
rect 21970 14026 22370 14072
rect 463 13290 863 13349
rect 463 13234 512 13290
rect 568 13234 634 13290
rect 690 13234 760 13290
rect 816 13234 863 13290
rect 463 13143 863 13234
rect 463 13087 512 13143
rect 568 13087 634 13143
rect 690 13087 760 13143
rect 816 13087 863 13143
rect 463 13006 863 13087
rect 463 12950 512 13006
rect 568 12950 634 13006
rect 690 12950 760 13006
rect 816 12950 863 13006
rect 463 12890 863 12950
rect 463 12611 864 12646
rect 463 12555 511 12611
rect 567 12555 637 12611
rect 693 12555 757 12611
rect 813 12555 864 12611
rect 463 12493 864 12555
rect 463 12437 511 12493
rect 567 12437 637 12493
rect 693 12437 757 12493
rect 813 12437 864 12493
rect 463 12391 864 12437
rect 21028 12584 21428 12619
rect 21028 12528 21076 12584
rect 21132 12528 21202 12584
rect 21258 12528 21322 12584
rect 21378 12528 21428 12584
rect 21028 12466 21428 12528
rect 21028 12410 21076 12466
rect 21132 12410 21202 12466
rect 21258 12410 21322 12466
rect 21378 12410 21428 12466
rect 21028 12364 21428 12410
rect 463 11489 864 11524
rect 463 11433 511 11489
rect 567 11433 637 11489
rect 693 11433 757 11489
rect 813 11433 864 11489
rect 463 11371 864 11433
rect 463 11315 511 11371
rect 567 11315 637 11371
rect 693 11315 757 11371
rect 813 11315 864 11371
rect 463 11269 864 11315
rect 21027 11427 21427 11462
rect 21027 11371 21076 11427
rect 21132 11371 21202 11427
rect 21258 11371 21322 11427
rect 21378 11371 21427 11427
rect 21027 11309 21427 11371
rect 21027 11253 21076 11309
rect 21132 11253 21202 11309
rect 21258 11253 21322 11309
rect 21378 11253 21427 11309
rect 21027 11207 21427 11253
rect 463 11051 863 11110
rect 463 10995 512 11051
rect 568 10995 634 11051
rect 690 10995 760 11051
rect 816 10995 863 11051
rect 463 10904 863 10995
rect 463 10848 512 10904
rect 568 10848 634 10904
rect 690 10848 760 10904
rect 816 10848 863 10904
rect 463 10767 863 10848
rect 463 10711 512 10767
rect 568 10711 634 10767
rect 690 10711 760 10767
rect 816 10711 863 10767
rect 463 10651 863 10711
rect 21970 10282 22370 10317
rect 21970 10226 22018 10282
rect 22074 10226 22144 10282
rect 22200 10226 22264 10282
rect 22320 10226 22370 10282
rect 21970 10164 22370 10226
rect 21970 10108 22018 10164
rect 22074 10108 22144 10164
rect 22200 10108 22264 10164
rect 22320 10108 22370 10164
rect 21970 10062 22370 10108
rect 463 9289 863 9348
rect 463 9233 512 9289
rect 568 9233 634 9289
rect 690 9233 760 9289
rect 816 9233 863 9289
rect 463 9142 863 9233
rect 463 9086 512 9142
rect 568 9086 634 9142
rect 690 9086 760 9142
rect 816 9086 863 9142
rect 463 9005 863 9086
rect 463 8949 512 9005
rect 568 8949 634 9005
rect 690 8949 760 9005
rect 816 8949 863 9005
rect 463 8889 863 8949
rect 463 8629 863 8664
rect 463 8573 511 8629
rect 567 8573 637 8629
rect 693 8573 757 8629
rect 813 8573 863 8629
rect 463 8511 863 8573
rect 463 8455 511 8511
rect 567 8455 637 8511
rect 693 8455 757 8511
rect 813 8455 863 8511
rect 463 8409 863 8455
rect 21028 8584 21428 8619
rect 21028 8528 21076 8584
rect 21132 8528 21202 8584
rect 21258 8528 21322 8584
rect 21378 8528 21428 8584
rect 21028 8466 21428 8528
rect 21028 8410 21076 8466
rect 21132 8410 21202 8466
rect 21258 8410 21322 8466
rect 21378 8410 21428 8466
rect 21028 8364 21428 8410
rect 463 7518 863 7553
rect 463 7462 511 7518
rect 567 7462 637 7518
rect 693 7462 757 7518
rect 813 7462 863 7518
rect 463 7400 863 7462
rect 463 7344 511 7400
rect 567 7344 637 7400
rect 693 7344 757 7400
rect 813 7344 863 7400
rect 463 7298 863 7344
rect 21027 7427 21427 7462
rect 21027 7371 21076 7427
rect 21132 7371 21202 7427
rect 21258 7371 21322 7427
rect 21378 7371 21427 7427
rect 21027 7309 21427 7371
rect 21027 7253 21076 7309
rect 21132 7253 21202 7309
rect 21258 7253 21322 7309
rect 21378 7253 21427 7309
rect 21027 7207 21427 7253
rect 463 7051 863 7110
rect 463 6995 512 7051
rect 568 6995 634 7051
rect 690 6995 760 7051
rect 816 6995 863 7051
rect 463 6904 863 6995
rect 463 6848 512 6904
rect 568 6848 634 6904
rect 690 6848 760 6904
rect 816 6848 863 6904
rect 463 6767 863 6848
rect 463 6711 512 6767
rect 568 6711 634 6767
rect 690 6711 760 6767
rect 816 6711 863 6767
rect 463 6651 863 6711
rect 21970 6270 22370 6305
rect 21970 6214 22018 6270
rect 22074 6214 22144 6270
rect 22200 6214 22264 6270
rect 22320 6214 22370 6270
rect 21970 6152 22370 6214
rect 21970 6096 22018 6152
rect 22074 6096 22144 6152
rect 22200 6096 22264 6152
rect 22320 6096 22370 6152
rect 21970 6050 22370 6096
rect 463 5290 863 5349
rect 463 5234 512 5290
rect 568 5234 634 5290
rect 690 5234 760 5290
rect 816 5234 863 5290
rect 463 5143 863 5234
rect 463 5087 512 5143
rect 568 5087 634 5143
rect 690 5087 760 5143
rect 816 5087 863 5143
rect 463 5006 863 5087
rect 463 4950 512 5006
rect 568 4950 634 5006
rect 690 4950 760 5006
rect 816 4950 863 5006
rect 463 4890 863 4950
rect 463 4695 865 4730
rect 463 4639 511 4695
rect 567 4639 637 4695
rect 693 4639 757 4695
rect 813 4639 865 4695
rect 463 4577 865 4639
rect 463 4521 511 4577
rect 567 4521 637 4577
rect 693 4521 757 4577
rect 813 4521 865 4577
rect 463 4475 865 4521
rect 21028 4584 21428 4619
rect 21028 4528 21076 4584
rect 21132 4528 21202 4584
rect 21258 4528 21322 4584
rect 21378 4528 21428 4584
rect 21028 4466 21428 4528
rect 21028 4410 21076 4466
rect 21132 4410 21202 4466
rect 21258 4410 21322 4466
rect 21378 4410 21428 4466
rect 21028 4364 21428 4410
rect 463 3518 863 3553
rect 463 3462 511 3518
rect 567 3462 637 3518
rect 693 3462 757 3518
rect 813 3462 863 3518
rect 463 3400 863 3462
rect 463 3344 511 3400
rect 567 3344 637 3400
rect 693 3344 757 3400
rect 813 3344 863 3400
rect 463 3298 863 3344
rect 21027 3427 21427 3462
rect 21027 3371 21076 3427
rect 21132 3371 21202 3427
rect 21258 3371 21322 3427
rect 21378 3371 21427 3427
rect 21027 3309 21427 3371
rect 21027 3253 21076 3309
rect 21132 3253 21202 3309
rect 21258 3253 21322 3309
rect 21378 3253 21427 3309
rect 21027 3207 21427 3253
rect 463 3051 863 3110
rect 463 2995 512 3051
rect 568 2995 634 3051
rect 690 2995 760 3051
rect 816 2995 863 3051
rect 463 2904 863 2995
rect 463 2848 512 2904
rect 568 2848 634 2904
rect 690 2848 760 2904
rect 816 2848 863 2904
rect 463 2767 863 2848
rect 463 2711 512 2767
rect 568 2711 634 2767
rect 690 2711 760 2767
rect 816 2711 863 2767
rect 463 2651 863 2711
rect 21970 2270 22370 2305
rect 21970 2214 22018 2270
rect 22074 2214 22144 2270
rect 22200 2214 22264 2270
rect 22320 2214 22370 2270
rect 21970 2152 22370 2214
rect 21970 2096 22018 2152
rect 22074 2096 22144 2152
rect 22200 2096 22264 2152
rect 22320 2096 22370 2152
rect 21970 2050 22370 2096
rect 463 1290 863 1349
rect 463 1234 512 1290
rect 568 1234 634 1290
rect 690 1234 760 1290
rect 816 1234 863 1290
rect 463 1143 863 1234
rect 463 1087 512 1143
rect 568 1087 634 1143
rect 690 1087 760 1143
rect 816 1087 863 1143
rect 463 1006 863 1087
rect 463 950 512 1006
rect 568 950 634 1006
rect 690 950 760 1006
rect 816 950 863 1006
rect 463 890 863 950
rect 463 695 865 730
rect 463 639 511 695
rect 567 639 637 695
rect 693 639 757 695
rect 813 639 865 695
rect 463 577 865 639
rect 463 521 511 577
rect 567 521 637 577
rect 693 521 757 577
rect 813 521 865 577
rect 463 475 865 521
rect 21028 584 21428 619
rect 21028 528 21076 584
rect 21132 528 21202 584
rect 21258 528 21322 584
rect 21378 528 21428 584
rect 21028 466 21428 528
rect 21028 410 21076 466
rect 21132 410 21202 466
rect 21258 410 21322 466
rect 21378 410 21428 466
rect 21028 364 21428 410
<< via2 >>
rect 511 75440 567 75442
rect 511 75388 513 75440
rect 513 75388 565 75440
rect 565 75388 567 75440
rect 511 75386 567 75388
rect 637 75440 693 75442
rect 637 75388 639 75440
rect 639 75388 691 75440
rect 691 75388 693 75440
rect 637 75386 693 75388
rect 757 75440 813 75442
rect 757 75388 759 75440
rect 759 75388 811 75440
rect 811 75388 813 75440
rect 757 75386 813 75388
rect 511 75322 567 75324
rect 511 75270 513 75322
rect 513 75270 565 75322
rect 565 75270 567 75322
rect 511 75268 567 75270
rect 637 75322 693 75324
rect 637 75270 639 75322
rect 639 75270 691 75322
rect 691 75270 693 75322
rect 637 75268 693 75270
rect 757 75322 813 75324
rect 757 75270 759 75322
rect 759 75270 811 75322
rect 811 75270 813 75322
rect 757 75268 813 75270
rect 21076 75480 21132 75482
rect 21076 75428 21078 75480
rect 21078 75428 21130 75480
rect 21130 75428 21132 75480
rect 21076 75426 21132 75428
rect 21202 75480 21258 75482
rect 21202 75428 21204 75480
rect 21204 75428 21256 75480
rect 21256 75428 21258 75480
rect 21202 75426 21258 75428
rect 21322 75480 21378 75482
rect 21322 75428 21324 75480
rect 21324 75428 21376 75480
rect 21376 75428 21378 75480
rect 21322 75426 21378 75428
rect 21076 75362 21132 75364
rect 21076 75310 21078 75362
rect 21078 75310 21130 75362
rect 21130 75310 21132 75362
rect 21076 75308 21132 75310
rect 21202 75362 21258 75364
rect 21202 75310 21204 75362
rect 21204 75310 21256 75362
rect 21256 75310 21258 75362
rect 21202 75308 21258 75310
rect 21322 75362 21378 75364
rect 21322 75310 21324 75362
rect 21324 75310 21376 75362
rect 21376 75310 21378 75362
rect 21322 75308 21378 75310
rect 512 75048 568 75050
rect 512 74996 514 75048
rect 514 74996 566 75048
rect 566 74996 568 75048
rect 512 74994 568 74996
rect 634 75048 690 75050
rect 634 74996 636 75048
rect 636 74996 688 75048
rect 688 74996 690 75048
rect 634 74994 690 74996
rect 760 75048 816 75050
rect 760 74996 762 75048
rect 762 74996 814 75048
rect 814 74996 816 75048
rect 760 74994 816 74996
rect 512 74901 568 74903
rect 512 74849 514 74901
rect 514 74849 566 74901
rect 566 74849 568 74901
rect 512 74847 568 74849
rect 634 74901 690 74903
rect 634 74849 636 74901
rect 636 74849 688 74901
rect 688 74849 690 74901
rect 634 74847 690 74849
rect 760 74901 816 74903
rect 760 74849 762 74901
rect 762 74849 814 74901
rect 814 74849 816 74901
rect 760 74847 816 74849
rect 512 74764 568 74766
rect 512 74712 514 74764
rect 514 74712 566 74764
rect 566 74712 568 74764
rect 512 74710 568 74712
rect 634 74764 690 74766
rect 634 74712 636 74764
rect 636 74712 688 74764
rect 688 74712 690 74764
rect 634 74710 690 74712
rect 760 74764 816 74766
rect 760 74712 762 74764
rect 762 74712 814 74764
rect 814 74712 816 74764
rect 760 74710 816 74712
rect 22018 74059 22074 74061
rect 22018 74007 22020 74059
rect 22020 74007 22072 74059
rect 22072 74007 22074 74059
rect 22018 74005 22074 74007
rect 22144 74059 22200 74061
rect 22144 74007 22146 74059
rect 22146 74007 22198 74059
rect 22198 74007 22200 74059
rect 22144 74005 22200 74007
rect 22264 74059 22320 74061
rect 22264 74007 22266 74059
rect 22266 74007 22318 74059
rect 22318 74007 22320 74059
rect 22264 74005 22320 74007
rect 22018 73941 22074 73943
rect 22018 73889 22020 73941
rect 22020 73889 22072 73941
rect 22072 73889 22074 73941
rect 22018 73887 22074 73889
rect 22144 73941 22200 73943
rect 22144 73889 22146 73941
rect 22146 73889 22198 73941
rect 22198 73889 22200 73941
rect 22144 73887 22200 73889
rect 22264 73941 22320 73943
rect 22264 73889 22266 73941
rect 22266 73889 22318 73941
rect 22318 73889 22320 73941
rect 22264 73887 22320 73889
rect 512 73288 568 73290
rect 512 73236 514 73288
rect 514 73236 566 73288
rect 566 73236 568 73288
rect 512 73234 568 73236
rect 634 73288 690 73290
rect 634 73236 636 73288
rect 636 73236 688 73288
rect 688 73236 690 73288
rect 634 73234 690 73236
rect 760 73288 816 73290
rect 760 73236 762 73288
rect 762 73236 814 73288
rect 814 73236 816 73288
rect 760 73234 816 73236
rect 512 73141 568 73143
rect 512 73089 514 73141
rect 514 73089 566 73141
rect 566 73089 568 73141
rect 512 73087 568 73089
rect 634 73141 690 73143
rect 634 73089 636 73141
rect 636 73089 688 73141
rect 688 73089 690 73141
rect 634 73087 690 73089
rect 760 73141 816 73143
rect 760 73089 762 73141
rect 762 73089 814 73141
rect 814 73089 816 73141
rect 760 73087 816 73089
rect 512 73004 568 73006
rect 512 72952 514 73004
rect 514 72952 566 73004
rect 566 72952 568 73004
rect 512 72950 568 72952
rect 634 73004 690 73006
rect 634 72952 636 73004
rect 636 72952 688 73004
rect 688 72952 690 73004
rect 634 72950 690 72952
rect 760 73004 816 73006
rect 760 72952 762 73004
rect 762 72952 814 73004
rect 814 72952 816 73004
rect 760 72950 816 72952
rect 511 72767 567 72769
rect 511 72715 513 72767
rect 513 72715 565 72767
rect 565 72715 567 72767
rect 511 72713 567 72715
rect 637 72767 693 72769
rect 637 72715 639 72767
rect 639 72715 691 72767
rect 691 72715 693 72767
rect 637 72713 693 72715
rect 757 72767 813 72769
rect 757 72715 759 72767
rect 759 72715 811 72767
rect 811 72715 813 72767
rect 757 72713 813 72715
rect 511 72649 567 72651
rect 511 72597 513 72649
rect 513 72597 565 72649
rect 565 72597 567 72649
rect 511 72595 567 72597
rect 637 72649 693 72651
rect 637 72597 639 72649
rect 639 72597 691 72649
rect 691 72597 693 72649
rect 637 72595 693 72597
rect 757 72649 813 72651
rect 757 72597 759 72649
rect 759 72597 811 72649
rect 811 72597 813 72649
rect 757 72595 813 72597
rect 21076 72683 21132 72685
rect 21076 72631 21078 72683
rect 21078 72631 21130 72683
rect 21130 72631 21132 72683
rect 21076 72629 21132 72631
rect 21202 72683 21258 72685
rect 21202 72631 21204 72683
rect 21204 72631 21256 72683
rect 21256 72631 21258 72683
rect 21202 72629 21258 72631
rect 21322 72683 21378 72685
rect 21322 72631 21324 72683
rect 21324 72631 21376 72683
rect 21376 72631 21378 72683
rect 21322 72629 21378 72631
rect 21076 72565 21132 72567
rect 21076 72513 21078 72565
rect 21078 72513 21130 72565
rect 21130 72513 21132 72565
rect 21076 72511 21132 72513
rect 21202 72565 21258 72567
rect 21202 72513 21204 72565
rect 21204 72513 21256 72565
rect 21256 72513 21258 72565
rect 21202 72511 21258 72513
rect 21322 72565 21378 72567
rect 21322 72513 21324 72565
rect 21324 72513 21376 72565
rect 21376 72513 21378 72565
rect 21322 72511 21378 72513
rect 511 71440 567 71442
rect 511 71388 513 71440
rect 513 71388 565 71440
rect 565 71388 567 71440
rect 511 71386 567 71388
rect 637 71440 693 71442
rect 637 71388 639 71440
rect 639 71388 691 71440
rect 691 71388 693 71440
rect 637 71386 693 71388
rect 757 71440 813 71442
rect 757 71388 759 71440
rect 759 71388 811 71440
rect 811 71388 813 71440
rect 757 71386 813 71388
rect 511 71322 567 71324
rect 511 71270 513 71322
rect 513 71270 565 71322
rect 565 71270 567 71322
rect 511 71268 567 71270
rect 637 71322 693 71324
rect 637 71270 639 71322
rect 639 71270 691 71322
rect 691 71270 693 71322
rect 637 71268 693 71270
rect 757 71322 813 71324
rect 757 71270 759 71322
rect 759 71270 811 71322
rect 811 71270 813 71322
rect 757 71268 813 71270
rect 21076 71480 21132 71482
rect 21076 71428 21078 71480
rect 21078 71428 21130 71480
rect 21130 71428 21132 71480
rect 21076 71426 21132 71428
rect 21202 71480 21258 71482
rect 21202 71428 21204 71480
rect 21204 71428 21256 71480
rect 21256 71428 21258 71480
rect 21202 71426 21258 71428
rect 21322 71480 21378 71482
rect 21322 71428 21324 71480
rect 21324 71428 21376 71480
rect 21376 71428 21378 71480
rect 21322 71426 21378 71428
rect 21076 71362 21132 71364
rect 21076 71310 21078 71362
rect 21078 71310 21130 71362
rect 21130 71310 21132 71362
rect 21076 71308 21132 71310
rect 21202 71362 21258 71364
rect 21202 71310 21204 71362
rect 21204 71310 21256 71362
rect 21256 71310 21258 71362
rect 21202 71308 21258 71310
rect 21322 71362 21378 71364
rect 21322 71310 21324 71362
rect 21324 71310 21376 71362
rect 21376 71310 21378 71362
rect 21322 71308 21378 71310
rect 512 71048 568 71050
rect 512 70996 514 71048
rect 514 70996 566 71048
rect 566 70996 568 71048
rect 512 70994 568 70996
rect 634 71048 690 71050
rect 634 70996 636 71048
rect 636 70996 688 71048
rect 688 70996 690 71048
rect 634 70994 690 70996
rect 760 71048 816 71050
rect 760 70996 762 71048
rect 762 70996 814 71048
rect 814 70996 816 71048
rect 760 70994 816 70996
rect 512 70901 568 70903
rect 512 70849 514 70901
rect 514 70849 566 70901
rect 566 70849 568 70901
rect 512 70847 568 70849
rect 634 70901 690 70903
rect 634 70849 636 70901
rect 636 70849 688 70901
rect 688 70849 690 70901
rect 634 70847 690 70849
rect 760 70901 816 70903
rect 760 70849 762 70901
rect 762 70849 814 70901
rect 814 70849 816 70901
rect 760 70847 816 70849
rect 512 70764 568 70766
rect 512 70712 514 70764
rect 514 70712 566 70764
rect 566 70712 568 70764
rect 512 70710 568 70712
rect 634 70764 690 70766
rect 634 70712 636 70764
rect 636 70712 688 70764
rect 688 70712 690 70764
rect 634 70710 690 70712
rect 760 70764 816 70766
rect 760 70712 762 70764
rect 762 70712 814 70764
rect 814 70712 816 70764
rect 760 70710 816 70712
rect 22018 70059 22074 70061
rect 22018 70007 22020 70059
rect 22020 70007 22072 70059
rect 22072 70007 22074 70059
rect 22018 70005 22074 70007
rect 22144 70059 22200 70061
rect 22144 70007 22146 70059
rect 22146 70007 22198 70059
rect 22198 70007 22200 70059
rect 22144 70005 22200 70007
rect 22264 70059 22320 70061
rect 22264 70007 22266 70059
rect 22266 70007 22318 70059
rect 22318 70007 22320 70059
rect 22264 70005 22320 70007
rect 22018 69941 22074 69943
rect 22018 69889 22020 69941
rect 22020 69889 22072 69941
rect 22072 69889 22074 69941
rect 22018 69887 22074 69889
rect 22144 69941 22200 69943
rect 22144 69889 22146 69941
rect 22146 69889 22198 69941
rect 22198 69889 22200 69941
rect 22144 69887 22200 69889
rect 22264 69941 22320 69943
rect 22264 69889 22266 69941
rect 22266 69889 22318 69941
rect 22318 69889 22320 69941
rect 22264 69887 22320 69889
rect 512 69288 568 69290
rect 512 69236 514 69288
rect 514 69236 566 69288
rect 566 69236 568 69288
rect 512 69234 568 69236
rect 634 69288 690 69290
rect 634 69236 636 69288
rect 636 69236 688 69288
rect 688 69236 690 69288
rect 634 69234 690 69236
rect 760 69288 816 69290
rect 760 69236 762 69288
rect 762 69236 814 69288
rect 814 69236 816 69288
rect 760 69234 816 69236
rect 512 69141 568 69143
rect 512 69089 514 69141
rect 514 69089 566 69141
rect 566 69089 568 69141
rect 512 69087 568 69089
rect 634 69141 690 69143
rect 634 69089 636 69141
rect 636 69089 688 69141
rect 688 69089 690 69141
rect 634 69087 690 69089
rect 760 69141 816 69143
rect 760 69089 762 69141
rect 762 69089 814 69141
rect 814 69089 816 69141
rect 760 69087 816 69089
rect 512 69004 568 69006
rect 512 68952 514 69004
rect 514 68952 566 69004
rect 566 68952 568 69004
rect 512 68950 568 68952
rect 634 69004 690 69006
rect 634 68952 636 69004
rect 636 68952 688 69004
rect 688 68952 690 69004
rect 634 68950 690 68952
rect 760 69004 816 69006
rect 760 68952 762 69004
rect 762 68952 814 69004
rect 814 68952 816 69004
rect 760 68950 816 68952
rect 511 68767 567 68769
rect 511 68715 513 68767
rect 513 68715 565 68767
rect 565 68715 567 68767
rect 511 68713 567 68715
rect 637 68767 693 68769
rect 637 68715 639 68767
rect 639 68715 691 68767
rect 691 68715 693 68767
rect 637 68713 693 68715
rect 757 68767 813 68769
rect 757 68715 759 68767
rect 759 68715 811 68767
rect 811 68715 813 68767
rect 757 68713 813 68715
rect 511 68649 567 68651
rect 511 68597 513 68649
rect 513 68597 565 68649
rect 565 68597 567 68649
rect 511 68595 567 68597
rect 637 68649 693 68651
rect 637 68597 639 68649
rect 639 68597 691 68649
rect 691 68597 693 68649
rect 637 68595 693 68597
rect 757 68649 813 68651
rect 757 68597 759 68649
rect 759 68597 811 68649
rect 811 68597 813 68649
rect 757 68595 813 68597
rect 21076 68683 21132 68685
rect 21076 68631 21078 68683
rect 21078 68631 21130 68683
rect 21130 68631 21132 68683
rect 21076 68629 21132 68631
rect 21202 68683 21258 68685
rect 21202 68631 21204 68683
rect 21204 68631 21256 68683
rect 21256 68631 21258 68683
rect 21202 68629 21258 68631
rect 21322 68683 21378 68685
rect 21322 68631 21324 68683
rect 21324 68631 21376 68683
rect 21376 68631 21378 68683
rect 21322 68629 21378 68631
rect 21076 68565 21132 68567
rect 21076 68513 21078 68565
rect 21078 68513 21130 68565
rect 21130 68513 21132 68565
rect 21076 68511 21132 68513
rect 21202 68565 21258 68567
rect 21202 68513 21204 68565
rect 21204 68513 21256 68565
rect 21256 68513 21258 68565
rect 21202 68511 21258 68513
rect 21322 68565 21378 68567
rect 21322 68513 21324 68565
rect 21324 68513 21376 68565
rect 21376 68513 21378 68565
rect 21322 68511 21378 68513
rect 511 67438 567 67440
rect 511 67386 513 67438
rect 513 67386 565 67438
rect 565 67386 567 67438
rect 511 67384 567 67386
rect 637 67438 693 67440
rect 637 67386 639 67438
rect 639 67386 691 67438
rect 691 67386 693 67438
rect 637 67384 693 67386
rect 757 67438 813 67440
rect 757 67386 759 67438
rect 759 67386 811 67438
rect 811 67386 813 67438
rect 757 67384 813 67386
rect 511 67320 567 67322
rect 511 67268 513 67320
rect 513 67268 565 67320
rect 565 67268 567 67320
rect 511 67266 567 67268
rect 637 67320 693 67322
rect 637 67268 639 67320
rect 639 67268 691 67320
rect 691 67268 693 67320
rect 637 67266 693 67268
rect 757 67320 813 67322
rect 757 67268 759 67320
rect 759 67268 811 67320
rect 811 67268 813 67320
rect 757 67266 813 67268
rect 21076 67480 21132 67482
rect 21076 67428 21078 67480
rect 21078 67428 21130 67480
rect 21130 67428 21132 67480
rect 21076 67426 21132 67428
rect 21202 67480 21258 67482
rect 21202 67428 21204 67480
rect 21204 67428 21256 67480
rect 21256 67428 21258 67480
rect 21202 67426 21258 67428
rect 21322 67480 21378 67482
rect 21322 67428 21324 67480
rect 21324 67428 21376 67480
rect 21376 67428 21378 67480
rect 21322 67426 21378 67428
rect 21076 67362 21132 67364
rect 21076 67310 21078 67362
rect 21078 67310 21130 67362
rect 21130 67310 21132 67362
rect 21076 67308 21132 67310
rect 21202 67362 21258 67364
rect 21202 67310 21204 67362
rect 21204 67310 21256 67362
rect 21256 67310 21258 67362
rect 21202 67308 21258 67310
rect 21322 67362 21378 67364
rect 21322 67310 21324 67362
rect 21324 67310 21376 67362
rect 21376 67310 21378 67362
rect 21322 67308 21378 67310
rect 512 67048 568 67050
rect 512 66996 514 67048
rect 514 66996 566 67048
rect 566 66996 568 67048
rect 512 66994 568 66996
rect 634 67048 690 67050
rect 634 66996 636 67048
rect 636 66996 688 67048
rect 688 66996 690 67048
rect 634 66994 690 66996
rect 760 67048 816 67050
rect 760 66996 762 67048
rect 762 66996 814 67048
rect 814 66996 816 67048
rect 760 66994 816 66996
rect 512 66901 568 66903
rect 512 66849 514 66901
rect 514 66849 566 66901
rect 566 66849 568 66901
rect 512 66847 568 66849
rect 634 66901 690 66903
rect 634 66849 636 66901
rect 636 66849 688 66901
rect 688 66849 690 66901
rect 634 66847 690 66849
rect 760 66901 816 66903
rect 760 66849 762 66901
rect 762 66849 814 66901
rect 814 66849 816 66901
rect 760 66847 816 66849
rect 512 66764 568 66766
rect 512 66712 514 66764
rect 514 66712 566 66764
rect 566 66712 568 66764
rect 512 66710 568 66712
rect 634 66764 690 66766
rect 634 66712 636 66764
rect 636 66712 688 66764
rect 688 66712 690 66764
rect 634 66710 690 66712
rect 760 66764 816 66766
rect 760 66712 762 66764
rect 762 66712 814 66764
rect 814 66712 816 66764
rect 760 66710 816 66712
rect 22018 66046 22074 66048
rect 22018 65994 22020 66046
rect 22020 65994 22072 66046
rect 22072 65994 22074 66046
rect 22018 65992 22074 65994
rect 22144 66046 22200 66048
rect 22144 65994 22146 66046
rect 22146 65994 22198 66046
rect 22198 65994 22200 66046
rect 22144 65992 22200 65994
rect 22264 66046 22320 66048
rect 22264 65994 22266 66046
rect 22266 65994 22318 66046
rect 22318 65994 22320 66046
rect 22264 65992 22320 65994
rect 22018 65928 22074 65930
rect 22018 65876 22020 65928
rect 22020 65876 22072 65928
rect 22072 65876 22074 65928
rect 22018 65874 22074 65876
rect 22144 65928 22200 65930
rect 22144 65876 22146 65928
rect 22146 65876 22198 65928
rect 22198 65876 22200 65928
rect 22144 65874 22200 65876
rect 22264 65928 22320 65930
rect 22264 65876 22266 65928
rect 22266 65876 22318 65928
rect 22318 65876 22320 65928
rect 22264 65874 22320 65876
rect 512 65289 568 65291
rect 512 65237 514 65289
rect 514 65237 566 65289
rect 566 65237 568 65289
rect 512 65235 568 65237
rect 634 65289 690 65291
rect 634 65237 636 65289
rect 636 65237 688 65289
rect 688 65237 690 65289
rect 634 65235 690 65237
rect 760 65289 816 65291
rect 760 65237 762 65289
rect 762 65237 814 65289
rect 814 65237 816 65289
rect 760 65235 816 65237
rect 512 65142 568 65144
rect 512 65090 514 65142
rect 514 65090 566 65142
rect 566 65090 568 65142
rect 512 65088 568 65090
rect 634 65142 690 65144
rect 634 65090 636 65142
rect 636 65090 688 65142
rect 688 65090 690 65142
rect 634 65088 690 65090
rect 760 65142 816 65144
rect 760 65090 762 65142
rect 762 65090 814 65142
rect 814 65090 816 65142
rect 760 65088 816 65090
rect 512 65005 568 65007
rect 512 64953 514 65005
rect 514 64953 566 65005
rect 566 64953 568 65005
rect 512 64951 568 64953
rect 634 65005 690 65007
rect 634 64953 636 65005
rect 636 64953 688 65005
rect 688 64953 690 65005
rect 634 64951 690 64953
rect 760 65005 816 65007
rect 760 64953 762 65005
rect 762 64953 814 65005
rect 814 64953 816 65005
rect 760 64951 816 64953
rect 511 64698 567 64700
rect 511 64646 513 64698
rect 513 64646 565 64698
rect 565 64646 567 64698
rect 511 64644 567 64646
rect 637 64698 693 64700
rect 637 64646 639 64698
rect 639 64646 691 64698
rect 691 64646 693 64698
rect 637 64644 693 64646
rect 757 64698 813 64700
rect 757 64646 759 64698
rect 759 64646 811 64698
rect 811 64646 813 64698
rect 757 64644 813 64646
rect 511 64580 567 64582
rect 511 64528 513 64580
rect 513 64528 565 64580
rect 565 64528 567 64580
rect 511 64526 567 64528
rect 637 64580 693 64582
rect 637 64528 639 64580
rect 639 64528 691 64580
rect 691 64528 693 64580
rect 637 64526 693 64528
rect 757 64580 813 64582
rect 757 64528 759 64580
rect 759 64528 811 64580
rect 811 64528 813 64580
rect 757 64526 813 64528
rect 21076 64683 21132 64685
rect 21076 64631 21078 64683
rect 21078 64631 21130 64683
rect 21130 64631 21132 64683
rect 21076 64629 21132 64631
rect 21202 64683 21258 64685
rect 21202 64631 21204 64683
rect 21204 64631 21256 64683
rect 21256 64631 21258 64683
rect 21202 64629 21258 64631
rect 21322 64683 21378 64685
rect 21322 64631 21324 64683
rect 21324 64631 21376 64683
rect 21376 64631 21378 64683
rect 21322 64629 21378 64631
rect 21076 64565 21132 64567
rect 21076 64513 21078 64565
rect 21078 64513 21130 64565
rect 21130 64513 21132 64565
rect 21076 64511 21132 64513
rect 21202 64565 21258 64567
rect 21202 64513 21204 64565
rect 21204 64513 21256 64565
rect 21256 64513 21258 64565
rect 21202 64511 21258 64513
rect 21322 64565 21378 64567
rect 21322 64513 21324 64565
rect 21324 64513 21376 64565
rect 21376 64513 21378 64565
rect 21322 64511 21378 64513
rect 511 63520 567 63522
rect 511 63468 513 63520
rect 513 63468 565 63520
rect 565 63468 567 63520
rect 511 63466 567 63468
rect 637 63520 693 63522
rect 637 63468 639 63520
rect 639 63468 691 63520
rect 691 63468 693 63520
rect 637 63466 693 63468
rect 757 63520 813 63522
rect 757 63468 759 63520
rect 759 63468 811 63520
rect 811 63468 813 63520
rect 757 63466 813 63468
rect 511 63402 567 63404
rect 511 63350 513 63402
rect 513 63350 565 63402
rect 565 63350 567 63402
rect 511 63348 567 63350
rect 637 63402 693 63404
rect 637 63350 639 63402
rect 639 63350 691 63402
rect 691 63350 693 63402
rect 637 63348 693 63350
rect 757 63402 813 63404
rect 757 63350 759 63402
rect 759 63350 811 63402
rect 811 63350 813 63402
rect 757 63348 813 63350
rect 21076 63480 21132 63482
rect 21076 63428 21078 63480
rect 21078 63428 21130 63480
rect 21130 63428 21132 63480
rect 21076 63426 21132 63428
rect 21202 63480 21258 63482
rect 21202 63428 21204 63480
rect 21204 63428 21256 63480
rect 21256 63428 21258 63480
rect 21202 63426 21258 63428
rect 21322 63480 21378 63482
rect 21322 63428 21324 63480
rect 21324 63428 21376 63480
rect 21376 63428 21378 63480
rect 21322 63426 21378 63428
rect 21076 63362 21132 63364
rect 21076 63310 21078 63362
rect 21078 63310 21130 63362
rect 21130 63310 21132 63362
rect 21076 63308 21132 63310
rect 21202 63362 21258 63364
rect 21202 63310 21204 63362
rect 21204 63310 21256 63362
rect 21256 63310 21258 63362
rect 21202 63308 21258 63310
rect 21322 63362 21378 63364
rect 21322 63310 21324 63362
rect 21324 63310 21376 63362
rect 21376 63310 21378 63362
rect 21322 63308 21378 63310
rect 512 63048 568 63050
rect 512 62996 514 63048
rect 514 62996 566 63048
rect 566 62996 568 63048
rect 512 62994 568 62996
rect 634 63048 690 63050
rect 634 62996 636 63048
rect 636 62996 688 63048
rect 688 62996 690 63048
rect 634 62994 690 62996
rect 760 63048 816 63050
rect 760 62996 762 63048
rect 762 62996 814 63048
rect 814 62996 816 63048
rect 760 62994 816 62996
rect 512 62901 568 62903
rect 512 62849 514 62901
rect 514 62849 566 62901
rect 566 62849 568 62901
rect 512 62847 568 62849
rect 634 62901 690 62903
rect 634 62849 636 62901
rect 636 62849 688 62901
rect 688 62849 690 62901
rect 634 62847 690 62849
rect 760 62901 816 62903
rect 760 62849 762 62901
rect 762 62849 814 62901
rect 814 62849 816 62901
rect 760 62847 816 62849
rect 512 62764 568 62766
rect 512 62712 514 62764
rect 514 62712 566 62764
rect 566 62712 568 62764
rect 512 62710 568 62712
rect 634 62764 690 62766
rect 634 62712 636 62764
rect 636 62712 688 62764
rect 688 62712 690 62764
rect 634 62710 690 62712
rect 760 62764 816 62766
rect 760 62712 762 62764
rect 762 62712 814 62764
rect 814 62712 816 62764
rect 760 62710 816 62712
rect 22018 62045 22074 62047
rect 22018 61993 22020 62045
rect 22020 61993 22072 62045
rect 22072 61993 22074 62045
rect 22018 61991 22074 61993
rect 22144 62045 22200 62047
rect 22144 61993 22146 62045
rect 22146 61993 22198 62045
rect 22198 61993 22200 62045
rect 22144 61991 22200 61993
rect 22264 62045 22320 62047
rect 22264 61993 22266 62045
rect 22266 61993 22318 62045
rect 22318 61993 22320 62045
rect 22264 61991 22320 61993
rect 22018 61927 22074 61929
rect 22018 61875 22020 61927
rect 22020 61875 22072 61927
rect 22072 61875 22074 61927
rect 22018 61873 22074 61875
rect 22144 61927 22200 61929
rect 22144 61875 22146 61927
rect 22146 61875 22198 61927
rect 22198 61875 22200 61927
rect 22144 61873 22200 61875
rect 22264 61927 22320 61929
rect 22264 61875 22266 61927
rect 22266 61875 22318 61927
rect 22318 61875 22320 61927
rect 22264 61873 22320 61875
rect 512 61289 568 61291
rect 512 61237 514 61289
rect 514 61237 566 61289
rect 566 61237 568 61289
rect 512 61235 568 61237
rect 634 61289 690 61291
rect 634 61237 636 61289
rect 636 61237 688 61289
rect 688 61237 690 61289
rect 634 61235 690 61237
rect 760 61289 816 61291
rect 760 61237 762 61289
rect 762 61237 814 61289
rect 814 61237 816 61289
rect 760 61235 816 61237
rect 512 61142 568 61144
rect 512 61090 514 61142
rect 514 61090 566 61142
rect 566 61090 568 61142
rect 512 61088 568 61090
rect 634 61142 690 61144
rect 634 61090 636 61142
rect 636 61090 688 61142
rect 688 61090 690 61142
rect 634 61088 690 61090
rect 760 61142 816 61144
rect 760 61090 762 61142
rect 762 61090 814 61142
rect 814 61090 816 61142
rect 760 61088 816 61090
rect 512 61005 568 61007
rect 512 60953 514 61005
rect 514 60953 566 61005
rect 566 60953 568 61005
rect 512 60951 568 60953
rect 634 61005 690 61007
rect 634 60953 636 61005
rect 636 60953 688 61005
rect 688 60953 690 61005
rect 634 60951 690 60953
rect 760 61005 816 61007
rect 760 60953 762 61005
rect 762 60953 814 61005
rect 814 60953 816 61005
rect 760 60951 816 60953
rect 511 60672 567 60674
rect 511 60620 513 60672
rect 513 60620 565 60672
rect 565 60620 567 60672
rect 511 60618 567 60620
rect 637 60672 693 60674
rect 637 60620 639 60672
rect 639 60620 691 60672
rect 691 60620 693 60672
rect 637 60618 693 60620
rect 757 60672 813 60674
rect 757 60620 759 60672
rect 759 60620 811 60672
rect 811 60620 813 60672
rect 757 60618 813 60620
rect 511 60554 567 60556
rect 511 60502 513 60554
rect 513 60502 565 60554
rect 565 60502 567 60554
rect 511 60500 567 60502
rect 637 60554 693 60556
rect 637 60502 639 60554
rect 639 60502 691 60554
rect 691 60502 693 60554
rect 637 60500 693 60502
rect 757 60554 813 60556
rect 757 60502 759 60554
rect 759 60502 811 60554
rect 811 60502 813 60554
rect 757 60500 813 60502
rect 21076 60683 21132 60685
rect 21076 60631 21078 60683
rect 21078 60631 21130 60683
rect 21130 60631 21132 60683
rect 21076 60629 21132 60631
rect 21202 60683 21258 60685
rect 21202 60631 21204 60683
rect 21204 60631 21256 60683
rect 21256 60631 21258 60683
rect 21202 60629 21258 60631
rect 21322 60683 21378 60685
rect 21322 60631 21324 60683
rect 21324 60631 21376 60683
rect 21376 60631 21378 60683
rect 21322 60629 21378 60631
rect 21076 60565 21132 60567
rect 21076 60513 21078 60565
rect 21078 60513 21130 60565
rect 21130 60513 21132 60565
rect 21076 60511 21132 60513
rect 21202 60565 21258 60567
rect 21202 60513 21204 60565
rect 21204 60513 21256 60565
rect 21256 60513 21258 60565
rect 21202 60511 21258 60513
rect 21322 60565 21378 60567
rect 21322 60513 21324 60565
rect 21324 60513 21376 60565
rect 21376 60513 21378 60565
rect 21322 60511 21378 60513
rect 511 59469 567 59471
rect 511 59417 513 59469
rect 513 59417 565 59469
rect 565 59417 567 59469
rect 511 59415 567 59417
rect 637 59469 693 59471
rect 637 59417 639 59469
rect 639 59417 691 59469
rect 691 59417 693 59469
rect 637 59415 693 59417
rect 757 59469 813 59471
rect 757 59417 759 59469
rect 759 59417 811 59469
rect 811 59417 813 59469
rect 757 59415 813 59417
rect 511 59351 567 59353
rect 511 59299 513 59351
rect 513 59299 565 59351
rect 565 59299 567 59351
rect 511 59297 567 59299
rect 637 59351 693 59353
rect 637 59299 639 59351
rect 639 59299 691 59351
rect 691 59299 693 59351
rect 637 59297 693 59299
rect 757 59351 813 59353
rect 757 59299 759 59351
rect 759 59299 811 59351
rect 811 59299 813 59351
rect 757 59297 813 59299
rect 21076 59534 21132 59536
rect 21076 59482 21078 59534
rect 21078 59482 21130 59534
rect 21130 59482 21132 59534
rect 21076 59480 21132 59482
rect 21202 59534 21258 59536
rect 21202 59482 21204 59534
rect 21204 59482 21256 59534
rect 21256 59482 21258 59534
rect 21202 59480 21258 59482
rect 21322 59534 21378 59536
rect 21322 59482 21324 59534
rect 21324 59482 21376 59534
rect 21376 59482 21378 59534
rect 21322 59480 21378 59482
rect 21076 59416 21132 59418
rect 21076 59364 21078 59416
rect 21078 59364 21130 59416
rect 21130 59364 21132 59416
rect 21076 59362 21132 59364
rect 21202 59416 21258 59418
rect 21202 59364 21204 59416
rect 21204 59364 21256 59416
rect 21256 59364 21258 59416
rect 21202 59362 21258 59364
rect 21322 59416 21378 59418
rect 21322 59364 21324 59416
rect 21324 59364 21376 59416
rect 21376 59364 21378 59416
rect 21322 59362 21378 59364
rect 512 59048 568 59050
rect 512 58996 514 59048
rect 514 58996 566 59048
rect 566 58996 568 59048
rect 512 58994 568 58996
rect 634 59048 690 59050
rect 634 58996 636 59048
rect 636 58996 688 59048
rect 688 58996 690 59048
rect 634 58994 690 58996
rect 760 59048 816 59050
rect 760 58996 762 59048
rect 762 58996 814 59048
rect 814 58996 816 59048
rect 760 58994 816 58996
rect 512 58901 568 58903
rect 512 58849 514 58901
rect 514 58849 566 58901
rect 566 58849 568 58901
rect 512 58847 568 58849
rect 634 58901 690 58903
rect 634 58849 636 58901
rect 636 58849 688 58901
rect 688 58849 690 58901
rect 634 58847 690 58849
rect 760 58901 816 58903
rect 760 58849 762 58901
rect 762 58849 814 58901
rect 814 58849 816 58901
rect 760 58847 816 58849
rect 512 58764 568 58766
rect 512 58712 514 58764
rect 514 58712 566 58764
rect 566 58712 568 58764
rect 512 58710 568 58712
rect 634 58764 690 58766
rect 634 58712 636 58764
rect 636 58712 688 58764
rect 688 58712 690 58764
rect 634 58710 690 58712
rect 760 58764 816 58766
rect 760 58712 762 58764
rect 762 58712 814 58764
rect 814 58712 816 58764
rect 760 58710 816 58712
rect 22018 58084 22074 58086
rect 22018 58032 22020 58084
rect 22020 58032 22072 58084
rect 22072 58032 22074 58084
rect 22018 58030 22074 58032
rect 22144 58084 22200 58086
rect 22144 58032 22146 58084
rect 22146 58032 22198 58084
rect 22198 58032 22200 58084
rect 22144 58030 22200 58032
rect 22264 58084 22320 58086
rect 22264 58032 22266 58084
rect 22266 58032 22318 58084
rect 22318 58032 22320 58084
rect 22264 58030 22320 58032
rect 22018 57966 22074 57968
rect 22018 57914 22020 57966
rect 22020 57914 22072 57966
rect 22072 57914 22074 57966
rect 22018 57912 22074 57914
rect 22144 57966 22200 57968
rect 22144 57914 22146 57966
rect 22146 57914 22198 57966
rect 22198 57914 22200 57966
rect 22144 57912 22200 57914
rect 22264 57966 22320 57968
rect 22264 57914 22266 57966
rect 22266 57914 22318 57966
rect 22318 57914 22320 57966
rect 22264 57912 22320 57914
rect 512 57287 568 57289
rect 512 57235 514 57287
rect 514 57235 566 57287
rect 566 57235 568 57287
rect 512 57233 568 57235
rect 634 57287 690 57289
rect 634 57235 636 57287
rect 636 57235 688 57287
rect 688 57235 690 57287
rect 634 57233 690 57235
rect 760 57287 816 57289
rect 760 57235 762 57287
rect 762 57235 814 57287
rect 814 57235 816 57287
rect 760 57233 816 57235
rect 512 57140 568 57142
rect 512 57088 514 57140
rect 514 57088 566 57140
rect 566 57088 568 57140
rect 512 57086 568 57088
rect 634 57140 690 57142
rect 634 57088 636 57140
rect 636 57088 688 57140
rect 688 57088 690 57140
rect 634 57086 690 57088
rect 760 57140 816 57142
rect 760 57088 762 57140
rect 762 57088 814 57140
rect 814 57088 816 57140
rect 760 57086 816 57088
rect 512 57003 568 57005
rect 512 56951 514 57003
rect 514 56951 566 57003
rect 566 56951 568 57003
rect 512 56949 568 56951
rect 634 57003 690 57005
rect 634 56951 636 57003
rect 636 56951 688 57003
rect 688 56951 690 57003
rect 634 56949 690 56951
rect 760 57003 816 57005
rect 760 56951 762 57003
rect 762 56951 814 57003
rect 814 56951 816 57003
rect 760 56949 816 56951
rect 511 56692 567 56694
rect 511 56640 513 56692
rect 513 56640 565 56692
rect 565 56640 567 56692
rect 511 56638 567 56640
rect 637 56692 693 56694
rect 637 56640 639 56692
rect 639 56640 691 56692
rect 691 56640 693 56692
rect 637 56638 693 56640
rect 757 56692 813 56694
rect 757 56640 759 56692
rect 759 56640 811 56692
rect 811 56640 813 56692
rect 757 56638 813 56640
rect 511 56574 567 56576
rect 511 56522 513 56574
rect 513 56522 565 56574
rect 565 56522 567 56574
rect 511 56520 567 56522
rect 637 56574 693 56576
rect 637 56522 639 56574
rect 639 56522 691 56574
rect 691 56522 693 56574
rect 637 56520 693 56522
rect 757 56574 813 56576
rect 757 56522 759 56574
rect 759 56522 811 56574
rect 811 56522 813 56574
rect 757 56520 813 56522
rect 21076 56618 21132 56620
rect 21076 56566 21078 56618
rect 21078 56566 21130 56618
rect 21130 56566 21132 56618
rect 21076 56564 21132 56566
rect 21202 56618 21258 56620
rect 21202 56566 21204 56618
rect 21204 56566 21256 56618
rect 21256 56566 21258 56618
rect 21202 56564 21258 56566
rect 21322 56618 21378 56620
rect 21322 56566 21324 56618
rect 21324 56566 21376 56618
rect 21376 56566 21378 56618
rect 21322 56564 21378 56566
rect 21076 56500 21132 56502
rect 21076 56448 21078 56500
rect 21078 56448 21130 56500
rect 21130 56448 21132 56500
rect 21076 56446 21132 56448
rect 21202 56500 21258 56502
rect 21202 56448 21204 56500
rect 21204 56448 21256 56500
rect 21256 56448 21258 56500
rect 21202 56446 21258 56448
rect 21322 56500 21378 56502
rect 21322 56448 21324 56500
rect 21324 56448 21376 56500
rect 21376 56448 21378 56500
rect 21322 56446 21378 56448
rect 511 55485 567 55487
rect 511 55433 513 55485
rect 513 55433 565 55485
rect 565 55433 567 55485
rect 511 55431 567 55433
rect 637 55485 693 55487
rect 637 55433 639 55485
rect 639 55433 691 55485
rect 691 55433 693 55485
rect 637 55431 693 55433
rect 757 55485 813 55487
rect 757 55433 759 55485
rect 759 55433 811 55485
rect 811 55433 813 55485
rect 757 55431 813 55433
rect 511 55367 567 55369
rect 511 55315 513 55367
rect 513 55315 565 55367
rect 565 55315 567 55367
rect 511 55313 567 55315
rect 637 55367 693 55369
rect 637 55315 639 55367
rect 639 55315 691 55367
rect 691 55315 693 55367
rect 637 55313 693 55315
rect 757 55367 813 55369
rect 757 55315 759 55367
rect 759 55315 811 55367
rect 811 55315 813 55367
rect 757 55313 813 55315
rect 21076 55435 21132 55437
rect 21076 55383 21078 55435
rect 21078 55383 21130 55435
rect 21130 55383 21132 55435
rect 21076 55381 21132 55383
rect 21202 55435 21258 55437
rect 21202 55383 21204 55435
rect 21204 55383 21256 55435
rect 21256 55383 21258 55435
rect 21202 55381 21258 55383
rect 21322 55435 21378 55437
rect 21322 55383 21324 55435
rect 21324 55383 21376 55435
rect 21376 55383 21378 55435
rect 21322 55381 21378 55383
rect 21076 55317 21132 55319
rect 21076 55265 21078 55317
rect 21078 55265 21130 55317
rect 21130 55265 21132 55317
rect 21076 55263 21132 55265
rect 21202 55317 21258 55319
rect 21202 55265 21204 55317
rect 21204 55265 21256 55317
rect 21256 55265 21258 55317
rect 21202 55263 21258 55265
rect 21322 55317 21378 55319
rect 21322 55265 21324 55317
rect 21324 55265 21376 55317
rect 21376 55265 21378 55317
rect 21322 55263 21378 55265
rect 512 55048 568 55050
rect 512 54996 514 55048
rect 514 54996 566 55048
rect 566 54996 568 55048
rect 512 54994 568 54996
rect 634 55048 690 55050
rect 634 54996 636 55048
rect 636 54996 688 55048
rect 688 54996 690 55048
rect 634 54994 690 54996
rect 760 55048 816 55050
rect 760 54996 762 55048
rect 762 54996 814 55048
rect 814 54996 816 55048
rect 760 54994 816 54996
rect 512 54901 568 54903
rect 512 54849 514 54901
rect 514 54849 566 54901
rect 566 54849 568 54901
rect 512 54847 568 54849
rect 634 54901 690 54903
rect 634 54849 636 54901
rect 636 54849 688 54901
rect 688 54849 690 54901
rect 634 54847 690 54849
rect 760 54901 816 54903
rect 760 54849 762 54901
rect 762 54849 814 54901
rect 814 54849 816 54901
rect 760 54847 816 54849
rect 512 54764 568 54766
rect 512 54712 514 54764
rect 514 54712 566 54764
rect 566 54712 568 54764
rect 512 54710 568 54712
rect 634 54764 690 54766
rect 634 54712 636 54764
rect 636 54712 688 54764
rect 688 54712 690 54764
rect 634 54710 690 54712
rect 760 54764 816 54766
rect 760 54712 762 54764
rect 762 54712 814 54764
rect 814 54712 816 54764
rect 760 54710 816 54712
rect 22018 54067 22074 54069
rect 22018 54015 22020 54067
rect 22020 54015 22072 54067
rect 22072 54015 22074 54067
rect 22018 54013 22074 54015
rect 22144 54067 22200 54069
rect 22144 54015 22146 54067
rect 22146 54015 22198 54067
rect 22198 54015 22200 54067
rect 22144 54013 22200 54015
rect 22264 54067 22320 54069
rect 22264 54015 22266 54067
rect 22266 54015 22318 54067
rect 22318 54015 22320 54067
rect 22264 54013 22320 54015
rect 22018 53949 22074 53951
rect 22018 53897 22020 53949
rect 22020 53897 22072 53949
rect 22072 53897 22074 53949
rect 22018 53895 22074 53897
rect 22144 53949 22200 53951
rect 22144 53897 22146 53949
rect 22146 53897 22198 53949
rect 22198 53897 22200 53949
rect 22144 53895 22200 53897
rect 22264 53949 22320 53951
rect 22264 53897 22266 53949
rect 22266 53897 22318 53949
rect 22318 53897 22320 53949
rect 22264 53895 22320 53897
rect 512 53289 568 53291
rect 512 53237 514 53289
rect 514 53237 566 53289
rect 566 53237 568 53289
rect 512 53235 568 53237
rect 634 53289 690 53291
rect 634 53237 636 53289
rect 636 53237 688 53289
rect 688 53237 690 53289
rect 634 53235 690 53237
rect 760 53289 816 53291
rect 760 53237 762 53289
rect 762 53237 814 53289
rect 814 53237 816 53289
rect 760 53235 816 53237
rect 512 53142 568 53144
rect 512 53090 514 53142
rect 514 53090 566 53142
rect 566 53090 568 53142
rect 512 53088 568 53090
rect 634 53142 690 53144
rect 634 53090 636 53142
rect 636 53090 688 53142
rect 688 53090 690 53142
rect 634 53088 690 53090
rect 760 53142 816 53144
rect 760 53090 762 53142
rect 762 53090 814 53142
rect 814 53090 816 53142
rect 760 53088 816 53090
rect 512 53005 568 53007
rect 512 52953 514 53005
rect 514 52953 566 53005
rect 566 52953 568 53005
rect 512 52951 568 52953
rect 634 53005 690 53007
rect 634 52953 636 53005
rect 636 52953 688 53005
rect 688 52953 690 53005
rect 634 52951 690 52953
rect 760 53005 816 53007
rect 760 52953 762 53005
rect 762 52953 814 53005
rect 814 52953 816 53005
rect 760 52951 816 52953
rect 511 52719 567 52721
rect 511 52667 513 52719
rect 513 52667 565 52719
rect 565 52667 567 52719
rect 511 52665 567 52667
rect 637 52719 693 52721
rect 637 52667 639 52719
rect 639 52667 691 52719
rect 691 52667 693 52719
rect 637 52665 693 52667
rect 757 52719 813 52721
rect 757 52667 759 52719
rect 759 52667 811 52719
rect 811 52667 813 52719
rect 757 52665 813 52667
rect 511 52601 567 52603
rect 511 52549 513 52601
rect 513 52549 565 52601
rect 565 52549 567 52601
rect 511 52547 567 52549
rect 637 52601 693 52603
rect 637 52549 639 52601
rect 639 52549 691 52601
rect 691 52549 693 52601
rect 637 52547 693 52549
rect 757 52601 813 52603
rect 757 52549 759 52601
rect 759 52549 811 52601
rect 811 52549 813 52601
rect 757 52547 813 52549
rect 21076 52563 21132 52565
rect 21076 52511 21078 52563
rect 21078 52511 21130 52563
rect 21130 52511 21132 52563
rect 21076 52509 21132 52511
rect 21202 52563 21258 52565
rect 21202 52511 21204 52563
rect 21204 52511 21256 52563
rect 21256 52511 21258 52563
rect 21202 52509 21258 52511
rect 21322 52563 21378 52565
rect 21322 52511 21324 52563
rect 21324 52511 21376 52563
rect 21376 52511 21378 52563
rect 21322 52509 21378 52511
rect 21076 52445 21132 52447
rect 21076 52393 21078 52445
rect 21078 52393 21130 52445
rect 21130 52393 21132 52445
rect 21076 52391 21132 52393
rect 21202 52445 21258 52447
rect 21202 52393 21204 52445
rect 21204 52393 21256 52445
rect 21256 52393 21258 52445
rect 21202 52391 21258 52393
rect 21322 52445 21378 52447
rect 21322 52393 21324 52445
rect 21324 52393 21376 52445
rect 21376 52393 21378 52445
rect 21322 52391 21378 52393
rect 511 51532 567 51534
rect 511 51480 513 51532
rect 513 51480 565 51532
rect 565 51480 567 51532
rect 511 51478 567 51480
rect 637 51532 693 51534
rect 637 51480 639 51532
rect 639 51480 691 51532
rect 691 51480 693 51532
rect 637 51478 693 51480
rect 757 51532 813 51534
rect 757 51480 759 51532
rect 759 51480 811 51532
rect 811 51480 813 51532
rect 757 51478 813 51480
rect 511 51414 567 51416
rect 511 51362 513 51414
rect 513 51362 565 51414
rect 565 51362 567 51414
rect 511 51360 567 51362
rect 637 51414 693 51416
rect 637 51362 639 51414
rect 639 51362 691 51414
rect 691 51362 693 51414
rect 637 51360 693 51362
rect 757 51414 813 51416
rect 757 51362 759 51414
rect 759 51362 811 51414
rect 811 51362 813 51414
rect 757 51360 813 51362
rect 21076 51428 21132 51430
rect 21076 51376 21078 51428
rect 21078 51376 21130 51428
rect 21130 51376 21132 51428
rect 21076 51374 21132 51376
rect 21202 51428 21258 51430
rect 21202 51376 21204 51428
rect 21204 51376 21256 51428
rect 21256 51376 21258 51428
rect 21202 51374 21258 51376
rect 21322 51428 21378 51430
rect 21322 51376 21324 51428
rect 21324 51376 21376 51428
rect 21376 51376 21378 51428
rect 21322 51374 21378 51376
rect 21076 51310 21132 51312
rect 21076 51258 21078 51310
rect 21078 51258 21130 51310
rect 21130 51258 21132 51310
rect 21076 51256 21132 51258
rect 21202 51310 21258 51312
rect 21202 51258 21204 51310
rect 21204 51258 21256 51310
rect 21256 51258 21258 51310
rect 21202 51256 21258 51258
rect 21322 51310 21378 51312
rect 21322 51258 21324 51310
rect 21324 51258 21376 51310
rect 21376 51258 21378 51310
rect 21322 51256 21378 51258
rect 512 51048 568 51050
rect 512 50996 514 51048
rect 514 50996 566 51048
rect 566 50996 568 51048
rect 512 50994 568 50996
rect 634 51048 690 51050
rect 634 50996 636 51048
rect 636 50996 688 51048
rect 688 50996 690 51048
rect 634 50994 690 50996
rect 760 51048 816 51050
rect 760 50996 762 51048
rect 762 50996 814 51048
rect 814 50996 816 51048
rect 760 50994 816 50996
rect 512 50901 568 50903
rect 512 50849 514 50901
rect 514 50849 566 50901
rect 566 50849 568 50901
rect 512 50847 568 50849
rect 634 50901 690 50903
rect 634 50849 636 50901
rect 636 50849 688 50901
rect 688 50849 690 50901
rect 634 50847 690 50849
rect 760 50901 816 50903
rect 760 50849 762 50901
rect 762 50849 814 50901
rect 814 50849 816 50901
rect 760 50847 816 50849
rect 512 50764 568 50766
rect 512 50712 514 50764
rect 514 50712 566 50764
rect 566 50712 568 50764
rect 512 50710 568 50712
rect 634 50764 690 50766
rect 634 50712 636 50764
rect 636 50712 688 50764
rect 688 50712 690 50764
rect 634 50710 690 50712
rect 760 50764 816 50766
rect 760 50712 762 50764
rect 762 50712 814 50764
rect 814 50712 816 50764
rect 760 50710 816 50712
rect 22018 50146 22074 50148
rect 22018 50094 22020 50146
rect 22020 50094 22072 50146
rect 22072 50094 22074 50146
rect 22018 50092 22074 50094
rect 22144 50146 22200 50148
rect 22144 50094 22146 50146
rect 22146 50094 22198 50146
rect 22198 50094 22200 50146
rect 22144 50092 22200 50094
rect 22264 50146 22320 50148
rect 22264 50094 22266 50146
rect 22266 50094 22318 50146
rect 22318 50094 22320 50146
rect 22264 50092 22320 50094
rect 22018 50028 22074 50030
rect 22018 49976 22020 50028
rect 22020 49976 22072 50028
rect 22072 49976 22074 50028
rect 22018 49974 22074 49976
rect 22144 50028 22200 50030
rect 22144 49976 22146 50028
rect 22146 49976 22198 50028
rect 22198 49976 22200 50028
rect 22144 49974 22200 49976
rect 22264 50028 22320 50030
rect 22264 49976 22266 50028
rect 22266 49976 22318 50028
rect 22318 49976 22320 50028
rect 22264 49974 22320 49976
rect 512 49289 568 49291
rect 512 49237 514 49289
rect 514 49237 566 49289
rect 566 49237 568 49289
rect 512 49235 568 49237
rect 634 49289 690 49291
rect 634 49237 636 49289
rect 636 49237 688 49289
rect 688 49237 690 49289
rect 634 49235 690 49237
rect 760 49289 816 49291
rect 760 49237 762 49289
rect 762 49237 814 49289
rect 814 49237 816 49289
rect 760 49235 816 49237
rect 512 49142 568 49144
rect 512 49090 514 49142
rect 514 49090 566 49142
rect 566 49090 568 49142
rect 512 49088 568 49090
rect 634 49142 690 49144
rect 634 49090 636 49142
rect 636 49090 688 49142
rect 688 49090 690 49142
rect 634 49088 690 49090
rect 760 49142 816 49144
rect 760 49090 762 49142
rect 762 49090 814 49142
rect 814 49090 816 49142
rect 760 49088 816 49090
rect 512 49005 568 49007
rect 512 48953 514 49005
rect 514 48953 566 49005
rect 566 48953 568 49005
rect 512 48951 568 48953
rect 634 49005 690 49007
rect 634 48953 636 49005
rect 636 48953 688 49005
rect 688 48953 690 49005
rect 634 48951 690 48953
rect 760 49005 816 49007
rect 760 48953 762 49005
rect 762 48953 814 49005
rect 814 48953 816 49005
rect 760 48951 816 48953
rect 511 48710 567 48712
rect 511 48658 513 48710
rect 513 48658 565 48710
rect 565 48658 567 48710
rect 511 48656 567 48658
rect 637 48710 693 48712
rect 637 48658 639 48710
rect 639 48658 691 48710
rect 691 48658 693 48710
rect 637 48656 693 48658
rect 757 48710 813 48712
rect 757 48658 759 48710
rect 759 48658 811 48710
rect 811 48658 813 48710
rect 757 48656 813 48658
rect 511 48592 567 48594
rect 511 48540 513 48592
rect 513 48540 565 48592
rect 565 48540 567 48592
rect 511 48538 567 48540
rect 637 48592 693 48594
rect 637 48540 639 48592
rect 639 48540 691 48592
rect 691 48540 693 48592
rect 637 48538 693 48540
rect 757 48592 813 48594
rect 757 48540 759 48592
rect 759 48540 811 48592
rect 811 48540 813 48592
rect 757 48538 813 48540
rect 21076 48669 21132 48671
rect 21076 48617 21078 48669
rect 21078 48617 21130 48669
rect 21130 48617 21132 48669
rect 21076 48615 21132 48617
rect 21202 48669 21258 48671
rect 21202 48617 21204 48669
rect 21204 48617 21256 48669
rect 21256 48617 21258 48669
rect 21202 48615 21258 48617
rect 21322 48669 21378 48671
rect 21322 48617 21324 48669
rect 21324 48617 21376 48669
rect 21376 48617 21378 48669
rect 21322 48615 21378 48617
rect 21076 48551 21132 48553
rect 21076 48499 21078 48551
rect 21078 48499 21130 48551
rect 21130 48499 21132 48551
rect 21076 48497 21132 48499
rect 21202 48551 21258 48553
rect 21202 48499 21204 48551
rect 21204 48499 21256 48551
rect 21256 48499 21258 48551
rect 21202 48497 21258 48499
rect 21322 48551 21378 48553
rect 21322 48499 21324 48551
rect 21324 48499 21376 48551
rect 21376 48499 21378 48551
rect 21322 48497 21378 48499
rect 511 47557 567 47559
rect 511 47505 513 47557
rect 513 47505 565 47557
rect 565 47505 567 47557
rect 511 47503 567 47505
rect 637 47557 693 47559
rect 637 47505 639 47557
rect 639 47505 691 47557
rect 691 47505 693 47557
rect 637 47503 693 47505
rect 757 47557 813 47559
rect 757 47505 759 47557
rect 759 47505 811 47557
rect 811 47505 813 47557
rect 757 47503 813 47505
rect 511 47439 567 47441
rect 511 47387 513 47439
rect 513 47387 565 47439
rect 565 47387 567 47439
rect 511 47385 567 47387
rect 637 47439 693 47441
rect 637 47387 639 47439
rect 639 47387 691 47439
rect 691 47387 693 47439
rect 637 47385 693 47387
rect 757 47439 813 47441
rect 757 47387 759 47439
rect 759 47387 811 47439
rect 811 47387 813 47439
rect 757 47385 813 47387
rect 21076 47516 21132 47518
rect 21076 47464 21078 47516
rect 21078 47464 21130 47516
rect 21130 47464 21132 47516
rect 21076 47462 21132 47464
rect 21202 47516 21258 47518
rect 21202 47464 21204 47516
rect 21204 47464 21256 47516
rect 21256 47464 21258 47516
rect 21202 47462 21258 47464
rect 21322 47516 21378 47518
rect 21322 47464 21324 47516
rect 21324 47464 21376 47516
rect 21376 47464 21378 47516
rect 21322 47462 21378 47464
rect 21076 47398 21132 47400
rect 21076 47346 21078 47398
rect 21078 47346 21130 47398
rect 21130 47346 21132 47398
rect 21076 47344 21132 47346
rect 21202 47398 21258 47400
rect 21202 47346 21204 47398
rect 21204 47346 21256 47398
rect 21256 47346 21258 47398
rect 21202 47344 21258 47346
rect 21322 47398 21378 47400
rect 21322 47346 21324 47398
rect 21324 47346 21376 47398
rect 21376 47346 21378 47398
rect 21322 47344 21378 47346
rect 512 47048 568 47050
rect 512 46996 514 47048
rect 514 46996 566 47048
rect 566 46996 568 47048
rect 512 46994 568 46996
rect 634 47048 690 47050
rect 634 46996 636 47048
rect 636 46996 688 47048
rect 688 46996 690 47048
rect 634 46994 690 46996
rect 760 47048 816 47050
rect 760 46996 762 47048
rect 762 46996 814 47048
rect 814 46996 816 47048
rect 760 46994 816 46996
rect 512 46901 568 46903
rect 512 46849 514 46901
rect 514 46849 566 46901
rect 566 46849 568 46901
rect 512 46847 568 46849
rect 634 46901 690 46903
rect 634 46849 636 46901
rect 636 46849 688 46901
rect 688 46849 690 46901
rect 634 46847 690 46849
rect 760 46901 816 46903
rect 760 46849 762 46901
rect 762 46849 814 46901
rect 814 46849 816 46901
rect 760 46847 816 46849
rect 512 46764 568 46766
rect 512 46712 514 46764
rect 514 46712 566 46764
rect 566 46712 568 46764
rect 512 46710 568 46712
rect 634 46764 690 46766
rect 634 46712 636 46764
rect 636 46712 688 46764
rect 688 46712 690 46764
rect 634 46710 690 46712
rect 760 46764 816 46766
rect 760 46712 762 46764
rect 762 46712 814 46764
rect 814 46712 816 46764
rect 760 46710 816 46712
rect 22018 45888 22074 45890
rect 22018 45836 22020 45888
rect 22020 45836 22072 45888
rect 22072 45836 22074 45888
rect 22018 45834 22074 45836
rect 22144 45888 22200 45890
rect 22144 45836 22146 45888
rect 22146 45836 22198 45888
rect 22198 45836 22200 45888
rect 22144 45834 22200 45836
rect 22264 45888 22320 45890
rect 22264 45836 22266 45888
rect 22266 45836 22318 45888
rect 22318 45836 22320 45888
rect 22264 45834 22320 45836
rect 22018 45770 22074 45772
rect 22018 45718 22020 45770
rect 22020 45718 22072 45770
rect 22072 45718 22074 45770
rect 22018 45716 22074 45718
rect 22144 45770 22200 45772
rect 22144 45718 22146 45770
rect 22146 45718 22198 45770
rect 22198 45718 22200 45770
rect 22144 45716 22200 45718
rect 22264 45770 22320 45772
rect 22264 45718 22266 45770
rect 22266 45718 22318 45770
rect 22318 45718 22320 45770
rect 22264 45716 22320 45718
rect 512 45288 568 45290
rect 512 45236 514 45288
rect 514 45236 566 45288
rect 566 45236 568 45288
rect 512 45234 568 45236
rect 634 45288 690 45290
rect 634 45236 636 45288
rect 636 45236 688 45288
rect 688 45236 690 45288
rect 634 45234 690 45236
rect 760 45288 816 45290
rect 760 45236 762 45288
rect 762 45236 814 45288
rect 814 45236 816 45288
rect 760 45234 816 45236
rect 512 45141 568 45143
rect 512 45089 514 45141
rect 514 45089 566 45141
rect 566 45089 568 45141
rect 512 45087 568 45089
rect 634 45141 690 45143
rect 634 45089 636 45141
rect 636 45089 688 45141
rect 688 45089 690 45141
rect 634 45087 690 45089
rect 760 45141 816 45143
rect 760 45089 762 45141
rect 762 45089 814 45141
rect 814 45089 816 45141
rect 760 45087 816 45089
rect 512 45004 568 45006
rect 512 44952 514 45004
rect 514 44952 566 45004
rect 566 44952 568 45004
rect 512 44950 568 44952
rect 634 45004 690 45006
rect 634 44952 636 45004
rect 636 44952 688 45004
rect 688 44952 690 45004
rect 634 44950 690 44952
rect 760 45004 816 45006
rect 760 44952 762 45004
rect 762 44952 814 45004
rect 814 44952 816 45004
rect 760 44950 816 44952
rect 511 44497 567 44499
rect 511 44445 513 44497
rect 513 44445 565 44497
rect 565 44445 567 44497
rect 511 44443 567 44445
rect 637 44497 693 44499
rect 637 44445 639 44497
rect 639 44445 691 44497
rect 691 44445 693 44497
rect 637 44443 693 44445
rect 757 44497 813 44499
rect 757 44445 759 44497
rect 759 44445 811 44497
rect 811 44445 813 44497
rect 757 44443 813 44445
rect 511 44379 567 44381
rect 511 44327 513 44379
rect 513 44327 565 44379
rect 565 44327 567 44379
rect 511 44325 567 44327
rect 637 44379 693 44381
rect 637 44327 639 44379
rect 639 44327 691 44379
rect 691 44327 693 44379
rect 637 44325 693 44327
rect 757 44379 813 44381
rect 757 44327 759 44379
rect 759 44327 811 44379
rect 811 44327 813 44379
rect 757 44325 813 44327
rect 21076 44400 21132 44402
rect 21076 44348 21078 44400
rect 21078 44348 21130 44400
rect 21130 44348 21132 44400
rect 21076 44346 21132 44348
rect 21202 44400 21258 44402
rect 21202 44348 21204 44400
rect 21204 44348 21256 44400
rect 21256 44348 21258 44400
rect 21202 44346 21258 44348
rect 21322 44400 21378 44402
rect 21322 44348 21324 44400
rect 21324 44348 21376 44400
rect 21376 44348 21378 44400
rect 21322 44346 21378 44348
rect 21076 44282 21132 44284
rect 21076 44230 21078 44282
rect 21078 44230 21130 44282
rect 21130 44230 21132 44282
rect 21076 44228 21132 44230
rect 21202 44282 21258 44284
rect 21202 44230 21204 44282
rect 21204 44230 21256 44282
rect 21256 44230 21258 44282
rect 21202 44228 21258 44230
rect 21322 44282 21378 44284
rect 21322 44230 21324 44282
rect 21324 44230 21376 44282
rect 21376 44230 21378 44282
rect 21322 44228 21378 44230
rect 2257 39789 2393 39925
rect 44 39727 100 39729
rect 44 39675 46 39727
rect 46 39675 98 39727
rect 98 39675 100 39727
rect 44 39673 100 39675
rect 169 39727 225 39729
rect 169 39675 171 39727
rect 171 39675 223 39727
rect 223 39675 225 39727
rect 169 39673 225 39675
rect 294 39727 350 39729
rect 294 39675 296 39727
rect 296 39675 348 39727
rect 348 39675 350 39727
rect 294 39673 350 39675
rect 44 39621 100 39623
rect 44 39569 46 39621
rect 46 39569 98 39621
rect 98 39569 100 39621
rect 44 39567 100 39569
rect 169 39621 225 39623
rect 169 39569 171 39621
rect 171 39569 223 39621
rect 223 39569 225 39621
rect 169 39567 225 39569
rect 294 39621 350 39623
rect 294 39569 296 39621
rect 296 39569 348 39621
rect 348 39569 350 39621
rect 294 39567 350 39569
rect 1416 39263 1472 39319
rect 1498 39264 1554 39320
rect 1417 39183 1473 39239
rect 1499 39184 1555 39240
rect 22044 43528 22260 43824
rect 3361 39768 3497 39904
rect 492 39117 548 39119
rect 492 39065 494 39117
rect 494 39065 546 39117
rect 546 39065 548 39117
rect 492 39063 548 39065
rect 606 39117 662 39119
rect 606 39065 608 39117
rect 608 39065 660 39117
rect 660 39065 662 39117
rect 606 39063 662 39065
rect 720 39117 776 39119
rect 720 39065 722 39117
rect 722 39065 774 39117
rect 774 39065 776 39117
rect 720 39063 776 39065
rect 29 38573 85 38575
rect 29 38521 31 38573
rect 31 38521 83 38573
rect 83 38521 85 38573
rect 29 38519 85 38521
rect 143 38573 199 38575
rect 143 38521 145 38573
rect 145 38521 197 38573
rect 197 38521 199 38573
rect 143 38519 199 38521
rect 257 38573 313 38575
rect 257 38521 259 38573
rect 259 38521 311 38573
rect 311 38521 313 38573
rect 257 38519 313 38521
rect 492 38029 548 38031
rect 492 37977 494 38029
rect 494 37977 546 38029
rect 546 37977 548 38029
rect 492 37975 548 37977
rect 606 38029 662 38031
rect 606 37977 608 38029
rect 608 37977 660 38029
rect 660 37977 662 38029
rect 606 37975 662 37977
rect 720 38029 776 38031
rect 720 37977 722 38029
rect 722 37977 774 38029
rect 774 37977 776 38029
rect 720 37975 776 37977
rect 29 37485 85 37487
rect 29 37433 31 37485
rect 31 37433 83 37485
rect 83 37433 85 37485
rect 29 37431 85 37433
rect 143 37485 199 37487
rect 143 37433 145 37485
rect 145 37433 197 37485
rect 197 37433 199 37485
rect 143 37431 199 37433
rect 257 37485 313 37487
rect 257 37433 259 37485
rect 259 37433 311 37485
rect 311 37433 313 37485
rect 257 37431 313 37433
rect 492 36941 548 36943
rect 492 36889 494 36941
rect 494 36889 546 36941
rect 546 36889 548 36941
rect 492 36887 548 36889
rect 606 36941 662 36943
rect 606 36889 608 36941
rect 608 36889 660 36941
rect 660 36889 662 36941
rect 606 36887 662 36889
rect 720 36941 776 36943
rect 720 36889 722 36941
rect 722 36889 774 36941
rect 774 36889 776 36941
rect 720 36887 776 36889
rect 2760 39262 2816 39318
rect 2840 39261 2896 39317
rect 2761 39181 2817 39237
rect 2841 39181 2897 39237
rect 21547 39712 21603 39714
rect 21547 39660 21549 39712
rect 21549 39660 21601 39712
rect 21601 39660 21603 39712
rect 21547 39658 21603 39660
rect 21672 39712 21728 39714
rect 21672 39660 21674 39712
rect 21674 39660 21726 39712
rect 21726 39660 21728 39712
rect 21672 39658 21728 39660
rect 21797 39712 21853 39714
rect 21797 39660 21799 39712
rect 21799 39660 21851 39712
rect 21851 39660 21853 39712
rect 21797 39658 21853 39660
rect 21546 39592 21602 39594
rect 21546 39540 21548 39592
rect 21548 39540 21600 39592
rect 21600 39540 21602 39592
rect 21546 39538 21602 39540
rect 21671 39592 21727 39594
rect 21671 39540 21673 39592
rect 21673 39540 21725 39592
rect 21725 39540 21727 39592
rect 21671 39538 21727 39540
rect 21796 39592 21852 39594
rect 21796 39540 21798 39592
rect 21798 39540 21850 39592
rect 21850 39540 21852 39592
rect 21796 39538 21852 39540
rect 3360 39261 3416 39317
rect 3440 39260 3496 39316
rect 3361 39180 3417 39236
rect 3441 39180 3497 39236
rect 22044 36644 22260 36940
rect 2544 36404 2600 36460
rect 2624 36404 2680 36460
rect 21073 36158 21129 36160
rect 21073 36106 21075 36158
rect 21075 36106 21127 36158
rect 21127 36106 21129 36158
rect 21073 36104 21129 36106
rect 21198 36158 21254 36160
rect 21198 36106 21200 36158
rect 21200 36106 21252 36158
rect 21252 36106 21254 36158
rect 21198 36104 21254 36106
rect 21323 36158 21379 36160
rect 21323 36106 21325 36158
rect 21325 36106 21377 36158
rect 21377 36106 21379 36158
rect 21323 36104 21379 36106
rect 21072 36038 21128 36040
rect 21072 35986 21074 36038
rect 21074 35986 21126 36038
rect 21126 35986 21128 36038
rect 21072 35984 21128 35986
rect 21197 36038 21253 36040
rect 21197 35986 21199 36038
rect 21199 35986 21251 36038
rect 21251 35986 21253 36038
rect 21197 35984 21253 35986
rect 21322 36038 21378 36040
rect 21322 35986 21324 36038
rect 21324 35986 21376 36038
rect 21376 35986 21378 36038
rect 21322 35984 21378 35986
rect 21077 35580 21133 35582
rect 21077 35528 21079 35580
rect 21079 35528 21131 35580
rect 21131 35528 21133 35580
rect 21077 35526 21133 35528
rect 21199 35580 21255 35582
rect 21199 35528 21201 35580
rect 21201 35528 21253 35580
rect 21253 35528 21255 35580
rect 21199 35526 21255 35528
rect 21325 35580 21381 35582
rect 21325 35528 21327 35580
rect 21327 35528 21379 35580
rect 21379 35528 21381 35580
rect 21325 35526 21381 35528
rect 21077 35433 21133 35435
rect 21077 35381 21079 35433
rect 21079 35381 21131 35433
rect 21131 35381 21133 35433
rect 21077 35379 21133 35381
rect 21199 35433 21255 35435
rect 21199 35381 21201 35433
rect 21201 35381 21253 35433
rect 21253 35381 21255 35433
rect 21199 35379 21255 35381
rect 21325 35433 21381 35435
rect 21325 35381 21327 35433
rect 21327 35381 21379 35433
rect 21379 35381 21381 35433
rect 21325 35379 21381 35381
rect 21077 35296 21133 35298
rect 21077 35244 21079 35296
rect 21079 35244 21131 35296
rect 21131 35244 21133 35296
rect 21077 35242 21133 35244
rect 21199 35296 21255 35298
rect 21199 35244 21201 35296
rect 21201 35244 21253 35296
rect 21253 35244 21255 35296
rect 21199 35242 21255 35244
rect 21325 35296 21381 35298
rect 21325 35244 21327 35296
rect 21327 35244 21379 35296
rect 21379 35244 21381 35296
rect 21325 35242 21381 35244
rect 20572 34662 20628 34664
rect 20572 34610 20574 34662
rect 20574 34610 20626 34662
rect 20626 34610 20628 34662
rect 20572 34608 20628 34610
rect 20697 34662 20753 34664
rect 20697 34610 20699 34662
rect 20699 34610 20751 34662
rect 20751 34610 20753 34662
rect 20697 34608 20753 34610
rect 20822 34662 20878 34664
rect 20822 34610 20824 34662
rect 20824 34610 20876 34662
rect 20876 34610 20878 34662
rect 20822 34608 20878 34610
rect 20571 34542 20627 34544
rect 20571 34490 20573 34542
rect 20573 34490 20625 34542
rect 20625 34490 20627 34542
rect 20571 34488 20627 34490
rect 20696 34542 20752 34544
rect 20696 34490 20698 34542
rect 20698 34490 20750 34542
rect 20750 34490 20752 34542
rect 20696 34488 20752 34490
rect 20821 34542 20877 34544
rect 20821 34490 20823 34542
rect 20823 34490 20875 34542
rect 20875 34490 20877 34542
rect 20821 34488 20877 34490
rect 21547 34662 21603 34664
rect 21547 34610 21549 34662
rect 21549 34610 21601 34662
rect 21601 34610 21603 34662
rect 21547 34608 21603 34610
rect 21672 34662 21728 34664
rect 21672 34610 21674 34662
rect 21674 34610 21726 34662
rect 21726 34610 21728 34662
rect 21672 34608 21728 34610
rect 21797 34662 21853 34664
rect 21797 34610 21799 34662
rect 21799 34610 21851 34662
rect 21851 34610 21853 34662
rect 21797 34608 21853 34610
rect 21546 34542 21602 34544
rect 21546 34490 21548 34542
rect 21548 34490 21600 34542
rect 21600 34490 21602 34542
rect 21546 34488 21602 34490
rect 21671 34542 21727 34544
rect 21671 34490 21673 34542
rect 21673 34490 21725 34542
rect 21725 34490 21727 34542
rect 21671 34488 21727 34490
rect 21796 34542 21852 34544
rect 21796 34490 21798 34542
rect 21798 34490 21850 34542
rect 21850 34490 21852 34542
rect 21796 34488 21852 34490
rect 21077 33820 21133 33822
rect 21077 33768 21079 33820
rect 21079 33768 21131 33820
rect 21131 33768 21133 33820
rect 21077 33766 21133 33768
rect 21199 33820 21255 33822
rect 21199 33768 21201 33820
rect 21201 33768 21253 33820
rect 21253 33768 21255 33820
rect 21199 33766 21255 33768
rect 21325 33820 21381 33822
rect 21325 33768 21327 33820
rect 21327 33768 21379 33820
rect 21379 33768 21381 33820
rect 21325 33766 21381 33768
rect 21077 33673 21133 33675
rect 21077 33621 21079 33673
rect 21079 33621 21131 33673
rect 21131 33621 21133 33673
rect 21077 33619 21133 33621
rect 21199 33673 21255 33675
rect 21199 33621 21201 33673
rect 21201 33621 21253 33673
rect 21253 33621 21255 33673
rect 21199 33619 21255 33621
rect 21325 33673 21381 33675
rect 21325 33621 21327 33673
rect 21327 33621 21379 33673
rect 21379 33621 21381 33673
rect 21325 33619 21381 33621
rect 21077 33536 21133 33538
rect 21077 33484 21079 33536
rect 21079 33484 21131 33536
rect 21131 33484 21133 33536
rect 21077 33482 21133 33484
rect 21199 33536 21255 33538
rect 21199 33484 21201 33536
rect 21201 33484 21253 33536
rect 21253 33484 21255 33536
rect 21199 33482 21255 33484
rect 21325 33536 21381 33538
rect 21325 33484 21327 33536
rect 21327 33484 21379 33536
rect 21379 33484 21381 33536
rect 21325 33482 21381 33484
rect 21072 33103 21128 33105
rect 21072 33051 21074 33103
rect 21074 33051 21126 33103
rect 21126 33051 21128 33103
rect 21072 33049 21128 33051
rect 21197 33103 21253 33105
rect 21197 33051 21199 33103
rect 21199 33051 21251 33103
rect 21251 33051 21253 33103
rect 21197 33049 21253 33051
rect 21322 33103 21378 33105
rect 21322 33051 21324 33103
rect 21324 33051 21376 33103
rect 21376 33051 21378 33103
rect 21322 33049 21378 33051
rect 21071 32983 21127 32985
rect 21071 32931 21073 32983
rect 21073 32931 21125 32983
rect 21125 32931 21127 32983
rect 21071 32929 21127 32931
rect 21196 32983 21252 32985
rect 21196 32931 21198 32983
rect 21198 32931 21250 32983
rect 21250 32931 21252 32983
rect 21196 32929 21252 32931
rect 21321 32983 21377 32985
rect 21321 32931 21323 32983
rect 21323 32931 21375 32983
rect 21375 32931 21377 32983
rect 21321 32929 21377 32931
rect 511 32290 567 32292
rect 511 32238 513 32290
rect 513 32238 565 32290
rect 565 32238 567 32290
rect 511 32236 567 32238
rect 637 32290 693 32292
rect 637 32238 639 32290
rect 639 32238 691 32290
rect 691 32238 693 32290
rect 637 32236 693 32238
rect 757 32290 813 32292
rect 757 32238 759 32290
rect 759 32238 811 32290
rect 811 32238 813 32290
rect 757 32236 813 32238
rect 511 32172 567 32174
rect 511 32120 513 32172
rect 513 32120 565 32172
rect 565 32120 567 32172
rect 511 32118 567 32120
rect 637 32172 693 32174
rect 637 32120 639 32172
rect 639 32120 691 32172
rect 691 32120 693 32172
rect 637 32118 693 32120
rect 757 32172 813 32174
rect 757 32120 759 32172
rect 759 32120 811 32172
rect 811 32120 813 32172
rect 757 32118 813 32120
rect 21076 32290 21132 32292
rect 21076 32238 21078 32290
rect 21078 32238 21130 32290
rect 21130 32238 21132 32290
rect 21076 32236 21132 32238
rect 21202 32290 21258 32292
rect 21202 32238 21204 32290
rect 21204 32238 21256 32290
rect 21256 32238 21258 32290
rect 21202 32236 21258 32238
rect 21322 32290 21378 32292
rect 21322 32238 21324 32290
rect 21324 32238 21376 32290
rect 21376 32238 21378 32290
rect 21322 32236 21378 32238
rect 21076 32172 21132 32174
rect 21076 32120 21078 32172
rect 21078 32120 21130 32172
rect 21130 32120 21132 32172
rect 21076 32118 21132 32120
rect 21202 32172 21258 32174
rect 21202 32120 21204 32172
rect 21204 32120 21256 32172
rect 21256 32120 21258 32172
rect 21202 32118 21258 32120
rect 21322 32172 21378 32174
rect 21322 32120 21324 32172
rect 21324 32120 21376 32172
rect 21376 32120 21378 32172
rect 21322 32118 21378 32120
rect 511 31508 567 31510
rect 511 31456 513 31508
rect 513 31456 565 31508
rect 565 31456 567 31508
rect 511 31454 567 31456
rect 637 31508 693 31510
rect 637 31456 639 31508
rect 639 31456 691 31508
rect 691 31456 693 31508
rect 637 31454 693 31456
rect 757 31508 813 31510
rect 757 31456 759 31508
rect 759 31456 811 31508
rect 811 31456 813 31508
rect 757 31454 813 31456
rect 511 31390 567 31392
rect 511 31338 513 31390
rect 513 31338 565 31390
rect 565 31338 567 31390
rect 511 31336 567 31338
rect 637 31390 693 31392
rect 637 31338 639 31390
rect 639 31338 691 31390
rect 691 31338 693 31390
rect 637 31336 693 31338
rect 757 31390 813 31392
rect 757 31338 759 31390
rect 759 31338 811 31390
rect 811 31338 813 31390
rect 757 31336 813 31338
rect 21076 31508 21132 31510
rect 21076 31456 21078 31508
rect 21078 31456 21130 31508
rect 21130 31456 21132 31508
rect 21076 31454 21132 31456
rect 21202 31508 21258 31510
rect 21202 31456 21204 31508
rect 21204 31456 21256 31508
rect 21256 31456 21258 31508
rect 21202 31454 21258 31456
rect 21322 31508 21378 31510
rect 21322 31456 21324 31508
rect 21324 31456 21376 31508
rect 21376 31456 21378 31508
rect 21322 31454 21378 31456
rect 21076 31390 21132 31392
rect 21076 31338 21078 31390
rect 21078 31338 21130 31390
rect 21130 31338 21132 31390
rect 21076 31336 21132 31338
rect 21202 31390 21258 31392
rect 21202 31338 21204 31390
rect 21204 31338 21256 31390
rect 21256 31338 21258 31390
rect 21202 31336 21258 31338
rect 21322 31390 21378 31392
rect 21322 31338 21324 31390
rect 21324 31338 21376 31390
rect 21376 31338 21378 31390
rect 21322 31336 21378 31338
rect 512 31049 568 31051
rect 512 30997 514 31049
rect 514 30997 566 31049
rect 566 30997 568 31049
rect 512 30995 568 30997
rect 634 31049 690 31051
rect 634 30997 636 31049
rect 636 30997 688 31049
rect 688 30997 690 31049
rect 634 30995 690 30997
rect 760 31049 816 31051
rect 760 30997 762 31049
rect 762 30997 814 31049
rect 814 30997 816 31049
rect 760 30995 816 30997
rect 512 30902 568 30904
rect 512 30850 514 30902
rect 514 30850 566 30902
rect 566 30850 568 30902
rect 512 30848 568 30850
rect 634 30902 690 30904
rect 634 30850 636 30902
rect 636 30850 688 30902
rect 688 30850 690 30902
rect 634 30848 690 30850
rect 760 30902 816 30904
rect 760 30850 762 30902
rect 762 30850 814 30902
rect 814 30850 816 30902
rect 760 30848 816 30850
rect 512 30765 568 30767
rect 512 30713 514 30765
rect 514 30713 566 30765
rect 566 30713 568 30765
rect 512 30711 568 30713
rect 634 30765 690 30767
rect 634 30713 636 30765
rect 636 30713 688 30765
rect 688 30713 690 30765
rect 634 30711 690 30713
rect 760 30765 816 30767
rect 760 30713 762 30765
rect 762 30713 814 30765
rect 814 30713 816 30765
rect 760 30711 816 30713
rect 22018 30118 22074 30120
rect 22018 30066 22020 30118
rect 22020 30066 22072 30118
rect 22072 30066 22074 30118
rect 22018 30064 22074 30066
rect 22144 30118 22200 30120
rect 22144 30066 22146 30118
rect 22146 30066 22198 30118
rect 22198 30066 22200 30118
rect 22144 30064 22200 30066
rect 22264 30118 22320 30120
rect 22264 30066 22266 30118
rect 22266 30066 22318 30118
rect 22318 30066 22320 30118
rect 22264 30064 22320 30066
rect 22018 30000 22074 30002
rect 22018 29948 22020 30000
rect 22020 29948 22072 30000
rect 22072 29948 22074 30000
rect 22018 29946 22074 29948
rect 22144 30000 22200 30002
rect 22144 29948 22146 30000
rect 22146 29948 22198 30000
rect 22198 29948 22200 30000
rect 22144 29946 22200 29948
rect 22264 30000 22320 30002
rect 22264 29948 22266 30000
rect 22266 29948 22318 30000
rect 22318 29948 22320 30000
rect 22264 29946 22320 29948
rect 512 29282 568 29284
rect 512 29230 514 29282
rect 514 29230 566 29282
rect 566 29230 568 29282
rect 512 29228 568 29230
rect 634 29282 690 29284
rect 634 29230 636 29282
rect 636 29230 688 29282
rect 688 29230 690 29282
rect 634 29228 690 29230
rect 760 29282 816 29284
rect 760 29230 762 29282
rect 762 29230 814 29282
rect 814 29230 816 29282
rect 760 29228 816 29230
rect 512 29135 568 29137
rect 512 29083 514 29135
rect 514 29083 566 29135
rect 566 29083 568 29135
rect 512 29081 568 29083
rect 634 29135 690 29137
rect 634 29083 636 29135
rect 636 29083 688 29135
rect 688 29083 690 29135
rect 634 29081 690 29083
rect 760 29135 816 29137
rect 760 29083 762 29135
rect 762 29083 814 29135
rect 814 29083 816 29135
rect 760 29081 816 29083
rect 512 28998 568 29000
rect 512 28946 514 28998
rect 514 28946 566 28998
rect 566 28946 568 28998
rect 512 28944 568 28946
rect 634 28998 690 29000
rect 634 28946 636 28998
rect 636 28946 688 28998
rect 688 28946 690 28998
rect 634 28944 690 28946
rect 760 28998 816 29000
rect 760 28946 762 28998
rect 762 28946 814 28998
rect 814 28946 816 28998
rect 760 28944 816 28946
rect 511 28596 567 28598
rect 511 28544 513 28596
rect 513 28544 565 28596
rect 565 28544 567 28596
rect 511 28542 567 28544
rect 637 28596 693 28598
rect 637 28544 639 28596
rect 639 28544 691 28596
rect 691 28544 693 28596
rect 637 28542 693 28544
rect 757 28596 813 28598
rect 757 28544 759 28596
rect 759 28544 811 28596
rect 811 28544 813 28596
rect 757 28542 813 28544
rect 511 28478 567 28480
rect 511 28426 513 28478
rect 513 28426 565 28478
rect 565 28426 567 28478
rect 511 28424 567 28426
rect 637 28478 693 28480
rect 637 28426 639 28478
rect 639 28426 691 28478
rect 691 28426 693 28478
rect 637 28424 693 28426
rect 757 28478 813 28480
rect 757 28426 759 28478
rect 759 28426 811 28478
rect 811 28426 813 28478
rect 757 28424 813 28426
rect 21076 28547 21132 28549
rect 21076 28495 21078 28547
rect 21078 28495 21130 28547
rect 21130 28495 21132 28547
rect 21076 28493 21132 28495
rect 21202 28547 21258 28549
rect 21202 28495 21204 28547
rect 21204 28495 21256 28547
rect 21256 28495 21258 28547
rect 21202 28493 21258 28495
rect 21322 28547 21378 28549
rect 21322 28495 21324 28547
rect 21324 28495 21376 28547
rect 21376 28495 21378 28547
rect 21322 28493 21378 28495
rect 21076 28429 21132 28431
rect 21076 28377 21078 28429
rect 21078 28377 21130 28429
rect 21130 28377 21132 28429
rect 21076 28375 21132 28377
rect 21202 28429 21258 28431
rect 21202 28377 21204 28429
rect 21204 28377 21256 28429
rect 21256 28377 21258 28429
rect 21202 28375 21258 28377
rect 21322 28429 21378 28431
rect 21322 28377 21324 28429
rect 21324 28377 21376 28429
rect 21376 28377 21378 28429
rect 21322 28375 21378 28377
rect 511 27592 567 27594
rect 511 27540 513 27592
rect 513 27540 565 27592
rect 565 27540 567 27592
rect 511 27538 567 27540
rect 637 27592 693 27594
rect 637 27540 639 27592
rect 639 27540 691 27592
rect 691 27540 693 27592
rect 637 27538 693 27540
rect 757 27592 813 27594
rect 757 27540 759 27592
rect 759 27540 811 27592
rect 811 27540 813 27592
rect 757 27538 813 27540
rect 511 27474 567 27476
rect 511 27422 513 27474
rect 513 27422 565 27474
rect 565 27422 567 27474
rect 511 27420 567 27422
rect 637 27474 693 27476
rect 637 27422 639 27474
rect 639 27422 691 27474
rect 691 27422 693 27474
rect 637 27420 693 27422
rect 757 27474 813 27476
rect 757 27422 759 27474
rect 759 27422 811 27474
rect 811 27422 813 27474
rect 757 27420 813 27422
rect 21076 27430 21132 27432
rect 21076 27378 21078 27430
rect 21078 27378 21130 27430
rect 21130 27378 21132 27430
rect 21076 27376 21132 27378
rect 21202 27430 21258 27432
rect 21202 27378 21204 27430
rect 21204 27378 21256 27430
rect 21256 27378 21258 27430
rect 21202 27376 21258 27378
rect 21322 27430 21378 27432
rect 21322 27378 21324 27430
rect 21324 27378 21376 27430
rect 21376 27378 21378 27430
rect 21322 27376 21378 27378
rect 21076 27312 21132 27314
rect 21076 27260 21078 27312
rect 21078 27260 21130 27312
rect 21130 27260 21132 27312
rect 21076 27258 21132 27260
rect 21202 27312 21258 27314
rect 21202 27260 21204 27312
rect 21204 27260 21256 27312
rect 21256 27260 21258 27312
rect 21202 27258 21258 27260
rect 21322 27312 21378 27314
rect 21322 27260 21324 27312
rect 21324 27260 21376 27312
rect 21376 27260 21378 27312
rect 21322 27258 21378 27260
rect 512 27048 568 27050
rect 512 26996 514 27048
rect 514 26996 566 27048
rect 566 26996 568 27048
rect 512 26994 568 26996
rect 634 27048 690 27050
rect 634 26996 636 27048
rect 636 26996 688 27048
rect 688 26996 690 27048
rect 634 26994 690 26996
rect 760 27048 816 27050
rect 760 26996 762 27048
rect 762 26996 814 27048
rect 814 26996 816 27048
rect 760 26994 816 26996
rect 512 26901 568 26903
rect 512 26849 514 26901
rect 514 26849 566 26901
rect 566 26849 568 26901
rect 512 26847 568 26849
rect 634 26901 690 26903
rect 634 26849 636 26901
rect 636 26849 688 26901
rect 688 26849 690 26901
rect 634 26847 690 26849
rect 760 26901 816 26903
rect 760 26849 762 26901
rect 762 26849 814 26901
rect 814 26849 816 26901
rect 760 26847 816 26849
rect 512 26764 568 26766
rect 512 26712 514 26764
rect 514 26712 566 26764
rect 566 26712 568 26764
rect 512 26710 568 26712
rect 634 26764 690 26766
rect 634 26712 636 26764
rect 636 26712 688 26764
rect 688 26712 690 26764
rect 634 26710 690 26712
rect 760 26764 816 26766
rect 760 26712 762 26764
rect 762 26712 814 26764
rect 814 26712 816 26764
rect 760 26710 816 26712
rect 22018 25959 22074 25961
rect 22018 25907 22020 25959
rect 22020 25907 22072 25959
rect 22072 25907 22074 25959
rect 22018 25905 22074 25907
rect 22144 25959 22200 25961
rect 22144 25907 22146 25959
rect 22146 25907 22198 25959
rect 22198 25907 22200 25959
rect 22144 25905 22200 25907
rect 22264 25959 22320 25961
rect 22264 25907 22266 25959
rect 22266 25907 22318 25959
rect 22318 25907 22320 25959
rect 22264 25905 22320 25907
rect 22018 25841 22074 25843
rect 22018 25789 22020 25841
rect 22020 25789 22072 25841
rect 22072 25789 22074 25841
rect 22018 25787 22074 25789
rect 22144 25841 22200 25843
rect 22144 25789 22146 25841
rect 22146 25789 22198 25841
rect 22198 25789 22200 25841
rect 22144 25787 22200 25789
rect 22264 25841 22320 25843
rect 22264 25789 22266 25841
rect 22266 25789 22318 25841
rect 22318 25789 22320 25841
rect 22264 25787 22320 25789
rect 512 25288 568 25290
rect 512 25236 514 25288
rect 514 25236 566 25288
rect 566 25236 568 25288
rect 512 25234 568 25236
rect 634 25288 690 25290
rect 634 25236 636 25288
rect 636 25236 688 25288
rect 688 25236 690 25288
rect 634 25234 690 25236
rect 760 25288 816 25290
rect 760 25236 762 25288
rect 762 25236 814 25288
rect 814 25236 816 25288
rect 760 25234 816 25236
rect 512 25141 568 25143
rect 512 25089 514 25141
rect 514 25089 566 25141
rect 566 25089 568 25141
rect 512 25087 568 25089
rect 634 25141 690 25143
rect 634 25089 636 25141
rect 636 25089 688 25141
rect 688 25089 690 25141
rect 634 25087 690 25089
rect 760 25141 816 25143
rect 760 25089 762 25141
rect 762 25089 814 25141
rect 814 25089 816 25141
rect 760 25087 816 25089
rect 512 25004 568 25006
rect 512 24952 514 25004
rect 514 24952 566 25004
rect 566 24952 568 25004
rect 512 24950 568 24952
rect 634 25004 690 25006
rect 634 24952 636 25004
rect 636 24952 688 25004
rect 688 24952 690 25004
rect 634 24950 690 24952
rect 760 25004 816 25006
rect 760 24952 762 25004
rect 762 24952 814 25004
rect 814 24952 816 25004
rect 760 24950 816 24952
rect 511 24614 567 24616
rect 511 24562 513 24614
rect 513 24562 565 24614
rect 565 24562 567 24614
rect 511 24560 567 24562
rect 637 24614 693 24616
rect 637 24562 639 24614
rect 639 24562 691 24614
rect 691 24562 693 24614
rect 637 24560 693 24562
rect 757 24614 813 24616
rect 757 24562 759 24614
rect 759 24562 811 24614
rect 811 24562 813 24614
rect 757 24560 813 24562
rect 511 24496 567 24498
rect 511 24444 513 24496
rect 513 24444 565 24496
rect 565 24444 567 24496
rect 511 24442 567 24444
rect 637 24496 693 24498
rect 637 24444 639 24496
rect 639 24444 691 24496
rect 691 24444 693 24496
rect 637 24442 693 24444
rect 757 24496 813 24498
rect 757 24444 759 24496
rect 759 24444 811 24496
rect 811 24444 813 24496
rect 757 24442 813 24444
rect 21076 24587 21132 24589
rect 21076 24535 21078 24587
rect 21078 24535 21130 24587
rect 21130 24535 21132 24587
rect 21076 24533 21132 24535
rect 21202 24587 21258 24589
rect 21202 24535 21204 24587
rect 21204 24535 21256 24587
rect 21256 24535 21258 24587
rect 21202 24533 21258 24535
rect 21322 24587 21378 24589
rect 21322 24535 21324 24587
rect 21324 24535 21376 24587
rect 21376 24535 21378 24587
rect 21322 24533 21378 24535
rect 21076 24469 21132 24471
rect 21076 24417 21078 24469
rect 21078 24417 21130 24469
rect 21130 24417 21132 24469
rect 21076 24415 21132 24417
rect 21202 24469 21258 24471
rect 21202 24417 21204 24469
rect 21204 24417 21256 24469
rect 21256 24417 21258 24469
rect 21202 24415 21258 24417
rect 21322 24469 21378 24471
rect 21322 24417 21324 24469
rect 21324 24417 21376 24469
rect 21376 24417 21378 24469
rect 21322 24415 21378 24417
rect 511 23532 567 23534
rect 511 23480 513 23532
rect 513 23480 565 23532
rect 565 23480 567 23532
rect 511 23478 567 23480
rect 637 23532 693 23534
rect 637 23480 639 23532
rect 639 23480 691 23532
rect 691 23480 693 23532
rect 637 23478 693 23480
rect 757 23532 813 23534
rect 757 23480 759 23532
rect 759 23480 811 23532
rect 811 23480 813 23532
rect 757 23478 813 23480
rect 511 23414 567 23416
rect 511 23362 513 23414
rect 513 23362 565 23414
rect 565 23362 567 23414
rect 511 23360 567 23362
rect 637 23414 693 23416
rect 637 23362 639 23414
rect 639 23362 691 23414
rect 691 23362 693 23414
rect 637 23360 693 23362
rect 757 23414 813 23416
rect 757 23362 759 23414
rect 759 23362 811 23414
rect 811 23362 813 23414
rect 757 23360 813 23362
rect 21076 23412 21132 23414
rect 21076 23360 21078 23412
rect 21078 23360 21130 23412
rect 21130 23360 21132 23412
rect 21076 23358 21132 23360
rect 21202 23412 21258 23414
rect 21202 23360 21204 23412
rect 21204 23360 21256 23412
rect 21256 23360 21258 23412
rect 21202 23358 21258 23360
rect 21322 23412 21378 23414
rect 21322 23360 21324 23412
rect 21324 23360 21376 23412
rect 21376 23360 21378 23412
rect 21322 23358 21378 23360
rect 21076 23294 21132 23296
rect 21076 23242 21078 23294
rect 21078 23242 21130 23294
rect 21130 23242 21132 23294
rect 21076 23240 21132 23242
rect 21202 23294 21258 23296
rect 21202 23242 21204 23294
rect 21204 23242 21256 23294
rect 21256 23242 21258 23294
rect 21202 23240 21258 23242
rect 21322 23294 21378 23296
rect 21322 23242 21324 23294
rect 21324 23242 21376 23294
rect 21376 23242 21378 23294
rect 21322 23240 21378 23242
rect 512 23048 568 23050
rect 512 22996 514 23048
rect 514 22996 566 23048
rect 566 22996 568 23048
rect 512 22994 568 22996
rect 634 23048 690 23050
rect 634 22996 636 23048
rect 636 22996 688 23048
rect 688 22996 690 23048
rect 634 22994 690 22996
rect 760 23048 816 23050
rect 760 22996 762 23048
rect 762 22996 814 23048
rect 814 22996 816 23048
rect 760 22994 816 22996
rect 512 22901 568 22903
rect 512 22849 514 22901
rect 514 22849 566 22901
rect 566 22849 568 22901
rect 512 22847 568 22849
rect 634 22901 690 22903
rect 634 22849 636 22901
rect 636 22849 688 22901
rect 688 22849 690 22901
rect 634 22847 690 22849
rect 760 22901 816 22903
rect 760 22849 762 22901
rect 762 22849 814 22901
rect 814 22849 816 22901
rect 760 22847 816 22849
rect 512 22764 568 22766
rect 512 22712 514 22764
rect 514 22712 566 22764
rect 566 22712 568 22764
rect 512 22710 568 22712
rect 634 22764 690 22766
rect 634 22712 636 22764
rect 636 22712 688 22764
rect 688 22712 690 22764
rect 634 22710 690 22712
rect 760 22764 816 22766
rect 760 22712 762 22764
rect 762 22712 814 22764
rect 814 22712 816 22764
rect 760 22710 816 22712
rect 22018 22169 22074 22171
rect 22018 22117 22020 22169
rect 22020 22117 22072 22169
rect 22072 22117 22074 22169
rect 22018 22115 22074 22117
rect 22144 22169 22200 22171
rect 22144 22117 22146 22169
rect 22146 22117 22198 22169
rect 22198 22117 22200 22169
rect 22144 22115 22200 22117
rect 22264 22169 22320 22171
rect 22264 22117 22266 22169
rect 22266 22117 22318 22169
rect 22318 22117 22320 22169
rect 22264 22115 22320 22117
rect 22018 22051 22074 22053
rect 22018 21999 22020 22051
rect 22020 21999 22072 22051
rect 22072 21999 22074 22051
rect 22018 21997 22074 21999
rect 22144 22051 22200 22053
rect 22144 21999 22146 22051
rect 22146 21999 22198 22051
rect 22198 21999 22200 22051
rect 22144 21997 22200 21999
rect 22264 22051 22320 22053
rect 22264 21999 22266 22051
rect 22266 21999 22318 22051
rect 22318 21999 22320 22051
rect 22264 21997 22320 21999
rect 512 21289 568 21291
rect 512 21237 514 21289
rect 514 21237 566 21289
rect 566 21237 568 21289
rect 512 21235 568 21237
rect 634 21289 690 21291
rect 634 21237 636 21289
rect 636 21237 688 21289
rect 688 21237 690 21289
rect 634 21235 690 21237
rect 760 21289 816 21291
rect 760 21237 762 21289
rect 762 21237 814 21289
rect 814 21237 816 21289
rect 760 21235 816 21237
rect 512 21142 568 21144
rect 512 21090 514 21142
rect 514 21090 566 21142
rect 566 21090 568 21142
rect 512 21088 568 21090
rect 634 21142 690 21144
rect 634 21090 636 21142
rect 636 21090 688 21142
rect 688 21090 690 21142
rect 634 21088 690 21090
rect 760 21142 816 21144
rect 760 21090 762 21142
rect 762 21090 814 21142
rect 814 21090 816 21142
rect 760 21088 816 21090
rect 512 21005 568 21007
rect 512 20953 514 21005
rect 514 20953 566 21005
rect 566 20953 568 21005
rect 512 20951 568 20953
rect 634 21005 690 21007
rect 634 20953 636 21005
rect 636 20953 688 21005
rect 688 20953 690 21005
rect 634 20951 690 20953
rect 760 21005 816 21007
rect 760 20953 762 21005
rect 762 20953 814 21005
rect 814 20953 816 21005
rect 760 20951 816 20953
rect 511 20657 567 20659
rect 511 20605 513 20657
rect 513 20605 565 20657
rect 565 20605 567 20657
rect 511 20603 567 20605
rect 637 20657 693 20659
rect 637 20605 639 20657
rect 639 20605 691 20657
rect 691 20605 693 20657
rect 637 20603 693 20605
rect 757 20657 813 20659
rect 757 20605 759 20657
rect 759 20605 811 20657
rect 811 20605 813 20657
rect 757 20603 813 20605
rect 511 20539 567 20541
rect 511 20487 513 20539
rect 513 20487 565 20539
rect 565 20487 567 20539
rect 511 20485 567 20487
rect 637 20539 693 20541
rect 637 20487 639 20539
rect 639 20487 691 20539
rect 691 20487 693 20539
rect 637 20485 693 20487
rect 757 20539 813 20541
rect 757 20487 759 20539
rect 759 20487 811 20539
rect 811 20487 813 20539
rect 757 20485 813 20487
rect 21076 20571 21132 20573
rect 21076 20519 21078 20571
rect 21078 20519 21130 20571
rect 21130 20519 21132 20571
rect 21076 20517 21132 20519
rect 21202 20571 21258 20573
rect 21202 20519 21204 20571
rect 21204 20519 21256 20571
rect 21256 20519 21258 20571
rect 21202 20517 21258 20519
rect 21322 20571 21378 20573
rect 21322 20519 21324 20571
rect 21324 20519 21376 20571
rect 21376 20519 21378 20571
rect 21322 20517 21378 20519
rect 21076 20453 21132 20455
rect 21076 20401 21078 20453
rect 21078 20401 21130 20453
rect 21130 20401 21132 20453
rect 21076 20399 21132 20401
rect 21202 20453 21258 20455
rect 21202 20401 21204 20453
rect 21204 20401 21256 20453
rect 21256 20401 21258 20453
rect 21202 20399 21258 20401
rect 21322 20453 21378 20455
rect 21322 20401 21324 20453
rect 21324 20401 21376 20453
rect 21376 20401 21378 20453
rect 21322 20399 21378 20401
rect 511 19556 567 19558
rect 511 19504 513 19556
rect 513 19504 565 19556
rect 565 19504 567 19556
rect 511 19502 567 19504
rect 637 19556 693 19558
rect 637 19504 639 19556
rect 639 19504 691 19556
rect 691 19504 693 19556
rect 637 19502 693 19504
rect 757 19556 813 19558
rect 757 19504 759 19556
rect 759 19504 811 19556
rect 811 19504 813 19556
rect 757 19502 813 19504
rect 511 19438 567 19440
rect 511 19386 513 19438
rect 513 19386 565 19438
rect 565 19386 567 19438
rect 511 19384 567 19386
rect 637 19438 693 19440
rect 637 19386 639 19438
rect 639 19386 691 19438
rect 691 19386 693 19438
rect 637 19384 693 19386
rect 757 19438 813 19440
rect 757 19386 759 19438
rect 759 19386 811 19438
rect 811 19386 813 19438
rect 757 19384 813 19386
rect 21076 19400 21132 19402
rect 21076 19348 21078 19400
rect 21078 19348 21130 19400
rect 21130 19348 21132 19400
rect 21076 19346 21132 19348
rect 21202 19400 21258 19402
rect 21202 19348 21204 19400
rect 21204 19348 21256 19400
rect 21256 19348 21258 19400
rect 21202 19346 21258 19348
rect 21322 19400 21378 19402
rect 21322 19348 21324 19400
rect 21324 19348 21376 19400
rect 21376 19348 21378 19400
rect 21322 19346 21378 19348
rect 21076 19282 21132 19284
rect 21076 19230 21078 19282
rect 21078 19230 21130 19282
rect 21130 19230 21132 19282
rect 21076 19228 21132 19230
rect 21202 19282 21258 19284
rect 21202 19230 21204 19282
rect 21204 19230 21256 19282
rect 21256 19230 21258 19282
rect 21202 19228 21258 19230
rect 21322 19282 21378 19284
rect 21322 19230 21324 19282
rect 21324 19230 21376 19282
rect 21376 19230 21378 19282
rect 21322 19228 21378 19230
rect 512 19048 568 19050
rect 512 18996 514 19048
rect 514 18996 566 19048
rect 566 18996 568 19048
rect 512 18994 568 18996
rect 634 19048 690 19050
rect 634 18996 636 19048
rect 636 18996 688 19048
rect 688 18996 690 19048
rect 634 18994 690 18996
rect 760 19048 816 19050
rect 760 18996 762 19048
rect 762 18996 814 19048
rect 814 18996 816 19048
rect 760 18994 816 18996
rect 512 18901 568 18903
rect 512 18849 514 18901
rect 514 18849 566 18901
rect 566 18849 568 18901
rect 512 18847 568 18849
rect 634 18901 690 18903
rect 634 18849 636 18901
rect 636 18849 688 18901
rect 688 18849 690 18901
rect 634 18847 690 18849
rect 760 18901 816 18903
rect 760 18849 762 18901
rect 762 18849 814 18901
rect 814 18849 816 18901
rect 760 18847 816 18849
rect 512 18764 568 18766
rect 512 18712 514 18764
rect 514 18712 566 18764
rect 566 18712 568 18764
rect 512 18710 568 18712
rect 634 18764 690 18766
rect 634 18712 636 18764
rect 636 18712 688 18764
rect 688 18712 690 18764
rect 634 18710 690 18712
rect 760 18764 816 18766
rect 760 18712 762 18764
rect 762 18712 814 18764
rect 814 18712 816 18764
rect 760 18710 816 18712
rect 22018 18062 22074 18064
rect 22018 18010 22020 18062
rect 22020 18010 22072 18062
rect 22072 18010 22074 18062
rect 22018 18008 22074 18010
rect 22144 18062 22200 18064
rect 22144 18010 22146 18062
rect 22146 18010 22198 18062
rect 22198 18010 22200 18062
rect 22144 18008 22200 18010
rect 22264 18062 22320 18064
rect 22264 18010 22266 18062
rect 22266 18010 22318 18062
rect 22318 18010 22320 18062
rect 22264 18008 22320 18010
rect 22018 17944 22074 17946
rect 22018 17892 22020 17944
rect 22020 17892 22072 17944
rect 22072 17892 22074 17944
rect 22018 17890 22074 17892
rect 22144 17944 22200 17946
rect 22144 17892 22146 17944
rect 22146 17892 22198 17944
rect 22198 17892 22200 17944
rect 22144 17890 22200 17892
rect 22264 17944 22320 17946
rect 22264 17892 22266 17944
rect 22266 17892 22318 17944
rect 22318 17892 22320 17944
rect 22264 17890 22320 17892
rect 512 17288 568 17290
rect 512 17236 514 17288
rect 514 17236 566 17288
rect 566 17236 568 17288
rect 512 17234 568 17236
rect 634 17288 690 17290
rect 634 17236 636 17288
rect 636 17236 688 17288
rect 688 17236 690 17288
rect 634 17234 690 17236
rect 760 17288 816 17290
rect 760 17236 762 17288
rect 762 17236 814 17288
rect 814 17236 816 17288
rect 760 17234 816 17236
rect 512 17141 568 17143
rect 512 17089 514 17141
rect 514 17089 566 17141
rect 566 17089 568 17141
rect 512 17087 568 17089
rect 634 17141 690 17143
rect 634 17089 636 17141
rect 636 17089 688 17141
rect 688 17089 690 17141
rect 634 17087 690 17089
rect 760 17141 816 17143
rect 760 17089 762 17141
rect 762 17089 814 17141
rect 814 17089 816 17141
rect 760 17087 816 17089
rect 512 17004 568 17006
rect 512 16952 514 17004
rect 514 16952 566 17004
rect 566 16952 568 17004
rect 512 16950 568 16952
rect 634 17004 690 17006
rect 634 16952 636 17004
rect 636 16952 688 17004
rect 688 16952 690 17004
rect 634 16950 690 16952
rect 760 17004 816 17006
rect 760 16952 762 17004
rect 762 16952 814 17004
rect 814 16952 816 17004
rect 760 16950 816 16952
rect 511 16690 567 16692
rect 511 16638 513 16690
rect 513 16638 565 16690
rect 565 16638 567 16690
rect 511 16636 567 16638
rect 637 16690 693 16692
rect 637 16638 639 16690
rect 639 16638 691 16690
rect 691 16638 693 16690
rect 637 16636 693 16638
rect 757 16690 813 16692
rect 757 16638 759 16690
rect 759 16638 811 16690
rect 811 16638 813 16690
rect 757 16636 813 16638
rect 511 16572 567 16574
rect 511 16520 513 16572
rect 513 16520 565 16572
rect 565 16520 567 16572
rect 511 16518 567 16520
rect 637 16572 693 16574
rect 637 16520 639 16572
rect 639 16520 691 16572
rect 691 16520 693 16572
rect 637 16518 693 16520
rect 757 16572 813 16574
rect 757 16520 759 16572
rect 759 16520 811 16572
rect 811 16520 813 16572
rect 757 16518 813 16520
rect 21076 16639 21132 16641
rect 21076 16587 21078 16639
rect 21078 16587 21130 16639
rect 21130 16587 21132 16639
rect 21076 16585 21132 16587
rect 21202 16639 21258 16641
rect 21202 16587 21204 16639
rect 21204 16587 21256 16639
rect 21256 16587 21258 16639
rect 21202 16585 21258 16587
rect 21322 16639 21378 16641
rect 21322 16587 21324 16639
rect 21324 16587 21376 16639
rect 21376 16587 21378 16639
rect 21322 16585 21378 16587
rect 21076 16521 21132 16523
rect 21076 16469 21078 16521
rect 21078 16469 21130 16521
rect 21130 16469 21132 16521
rect 21076 16467 21132 16469
rect 21202 16521 21258 16523
rect 21202 16469 21204 16521
rect 21204 16469 21256 16521
rect 21256 16469 21258 16521
rect 21202 16467 21258 16469
rect 21322 16521 21378 16523
rect 21322 16469 21324 16521
rect 21324 16469 21376 16521
rect 21376 16469 21378 16521
rect 21322 16467 21378 16469
rect 511 15474 567 15476
rect 511 15422 513 15474
rect 513 15422 565 15474
rect 565 15422 567 15474
rect 511 15420 567 15422
rect 637 15474 693 15476
rect 637 15422 639 15474
rect 639 15422 691 15474
rect 691 15422 693 15474
rect 637 15420 693 15422
rect 757 15474 813 15476
rect 757 15422 759 15474
rect 759 15422 811 15474
rect 811 15422 813 15474
rect 757 15420 813 15422
rect 511 15356 567 15358
rect 511 15304 513 15356
rect 513 15304 565 15356
rect 565 15304 567 15356
rect 511 15302 567 15304
rect 637 15356 693 15358
rect 637 15304 639 15356
rect 639 15304 691 15356
rect 691 15304 693 15356
rect 637 15302 693 15304
rect 757 15356 813 15358
rect 757 15304 759 15356
rect 759 15304 811 15356
rect 811 15304 813 15356
rect 757 15302 813 15304
rect 21076 15425 21132 15427
rect 21076 15373 21078 15425
rect 21078 15373 21130 15425
rect 21130 15373 21132 15425
rect 21076 15371 21132 15373
rect 21202 15425 21258 15427
rect 21202 15373 21204 15425
rect 21204 15373 21256 15425
rect 21256 15373 21258 15425
rect 21202 15371 21258 15373
rect 21322 15425 21378 15427
rect 21322 15373 21324 15425
rect 21324 15373 21376 15425
rect 21376 15373 21378 15425
rect 21322 15371 21378 15373
rect 21076 15307 21132 15309
rect 21076 15255 21078 15307
rect 21078 15255 21130 15307
rect 21130 15255 21132 15307
rect 21076 15253 21132 15255
rect 21202 15307 21258 15309
rect 21202 15255 21204 15307
rect 21204 15255 21256 15307
rect 21256 15255 21258 15307
rect 21202 15253 21258 15255
rect 21322 15307 21378 15309
rect 21322 15255 21324 15307
rect 21324 15255 21376 15307
rect 21376 15255 21378 15307
rect 21322 15253 21378 15255
rect 512 15048 568 15050
rect 512 14996 514 15048
rect 514 14996 566 15048
rect 566 14996 568 15048
rect 512 14994 568 14996
rect 634 15048 690 15050
rect 634 14996 636 15048
rect 636 14996 688 15048
rect 688 14996 690 15048
rect 634 14994 690 14996
rect 760 15048 816 15050
rect 760 14996 762 15048
rect 762 14996 814 15048
rect 814 14996 816 15048
rect 760 14994 816 14996
rect 512 14901 568 14903
rect 512 14849 514 14901
rect 514 14849 566 14901
rect 566 14849 568 14901
rect 512 14847 568 14849
rect 634 14901 690 14903
rect 634 14849 636 14901
rect 636 14849 688 14901
rect 688 14849 690 14901
rect 634 14847 690 14849
rect 760 14901 816 14903
rect 760 14849 762 14901
rect 762 14849 814 14901
rect 814 14849 816 14901
rect 760 14847 816 14849
rect 512 14764 568 14766
rect 512 14712 514 14764
rect 514 14712 566 14764
rect 566 14712 568 14764
rect 512 14710 568 14712
rect 634 14764 690 14766
rect 634 14712 636 14764
rect 636 14712 688 14764
rect 688 14712 690 14764
rect 634 14710 690 14712
rect 760 14764 816 14766
rect 760 14712 762 14764
rect 762 14712 814 14764
rect 814 14712 816 14764
rect 760 14710 816 14712
rect 22018 14244 22074 14246
rect 22018 14192 22020 14244
rect 22020 14192 22072 14244
rect 22072 14192 22074 14244
rect 22018 14190 22074 14192
rect 22144 14244 22200 14246
rect 22144 14192 22146 14244
rect 22146 14192 22198 14244
rect 22198 14192 22200 14244
rect 22144 14190 22200 14192
rect 22264 14244 22320 14246
rect 22264 14192 22266 14244
rect 22266 14192 22318 14244
rect 22318 14192 22320 14244
rect 22264 14190 22320 14192
rect 22018 14126 22074 14128
rect 22018 14074 22020 14126
rect 22020 14074 22072 14126
rect 22072 14074 22074 14126
rect 22018 14072 22074 14074
rect 22144 14126 22200 14128
rect 22144 14074 22146 14126
rect 22146 14074 22198 14126
rect 22198 14074 22200 14126
rect 22144 14072 22200 14074
rect 22264 14126 22320 14128
rect 22264 14074 22266 14126
rect 22266 14074 22318 14126
rect 22318 14074 22320 14126
rect 22264 14072 22320 14074
rect 512 13288 568 13290
rect 512 13236 514 13288
rect 514 13236 566 13288
rect 566 13236 568 13288
rect 512 13234 568 13236
rect 634 13288 690 13290
rect 634 13236 636 13288
rect 636 13236 688 13288
rect 688 13236 690 13288
rect 634 13234 690 13236
rect 760 13288 816 13290
rect 760 13236 762 13288
rect 762 13236 814 13288
rect 814 13236 816 13288
rect 760 13234 816 13236
rect 512 13141 568 13143
rect 512 13089 514 13141
rect 514 13089 566 13141
rect 566 13089 568 13141
rect 512 13087 568 13089
rect 634 13141 690 13143
rect 634 13089 636 13141
rect 636 13089 688 13141
rect 688 13089 690 13141
rect 634 13087 690 13089
rect 760 13141 816 13143
rect 760 13089 762 13141
rect 762 13089 814 13141
rect 814 13089 816 13141
rect 760 13087 816 13089
rect 512 13004 568 13006
rect 512 12952 514 13004
rect 514 12952 566 13004
rect 566 12952 568 13004
rect 512 12950 568 12952
rect 634 13004 690 13006
rect 634 12952 636 13004
rect 636 12952 688 13004
rect 688 12952 690 13004
rect 634 12950 690 12952
rect 760 13004 816 13006
rect 760 12952 762 13004
rect 762 12952 814 13004
rect 814 12952 816 13004
rect 760 12950 816 12952
rect 511 12609 567 12611
rect 511 12557 513 12609
rect 513 12557 565 12609
rect 565 12557 567 12609
rect 511 12555 567 12557
rect 637 12609 693 12611
rect 637 12557 639 12609
rect 639 12557 691 12609
rect 691 12557 693 12609
rect 637 12555 693 12557
rect 757 12609 813 12611
rect 757 12557 759 12609
rect 759 12557 811 12609
rect 811 12557 813 12609
rect 757 12555 813 12557
rect 511 12491 567 12493
rect 511 12439 513 12491
rect 513 12439 565 12491
rect 565 12439 567 12491
rect 511 12437 567 12439
rect 637 12491 693 12493
rect 637 12439 639 12491
rect 639 12439 691 12491
rect 691 12439 693 12491
rect 637 12437 693 12439
rect 757 12491 813 12493
rect 757 12439 759 12491
rect 759 12439 811 12491
rect 811 12439 813 12491
rect 757 12437 813 12439
rect 21076 12582 21132 12584
rect 21076 12530 21078 12582
rect 21078 12530 21130 12582
rect 21130 12530 21132 12582
rect 21076 12528 21132 12530
rect 21202 12582 21258 12584
rect 21202 12530 21204 12582
rect 21204 12530 21256 12582
rect 21256 12530 21258 12582
rect 21202 12528 21258 12530
rect 21322 12582 21378 12584
rect 21322 12530 21324 12582
rect 21324 12530 21376 12582
rect 21376 12530 21378 12582
rect 21322 12528 21378 12530
rect 21076 12464 21132 12466
rect 21076 12412 21078 12464
rect 21078 12412 21130 12464
rect 21130 12412 21132 12464
rect 21076 12410 21132 12412
rect 21202 12464 21258 12466
rect 21202 12412 21204 12464
rect 21204 12412 21256 12464
rect 21256 12412 21258 12464
rect 21202 12410 21258 12412
rect 21322 12464 21378 12466
rect 21322 12412 21324 12464
rect 21324 12412 21376 12464
rect 21376 12412 21378 12464
rect 21322 12410 21378 12412
rect 511 11487 567 11489
rect 511 11435 513 11487
rect 513 11435 565 11487
rect 565 11435 567 11487
rect 511 11433 567 11435
rect 637 11487 693 11489
rect 637 11435 639 11487
rect 639 11435 691 11487
rect 691 11435 693 11487
rect 637 11433 693 11435
rect 757 11487 813 11489
rect 757 11435 759 11487
rect 759 11435 811 11487
rect 811 11435 813 11487
rect 757 11433 813 11435
rect 511 11369 567 11371
rect 511 11317 513 11369
rect 513 11317 565 11369
rect 565 11317 567 11369
rect 511 11315 567 11317
rect 637 11369 693 11371
rect 637 11317 639 11369
rect 639 11317 691 11369
rect 691 11317 693 11369
rect 637 11315 693 11317
rect 757 11369 813 11371
rect 757 11317 759 11369
rect 759 11317 811 11369
rect 811 11317 813 11369
rect 757 11315 813 11317
rect 21076 11425 21132 11427
rect 21076 11373 21078 11425
rect 21078 11373 21130 11425
rect 21130 11373 21132 11425
rect 21076 11371 21132 11373
rect 21202 11425 21258 11427
rect 21202 11373 21204 11425
rect 21204 11373 21256 11425
rect 21256 11373 21258 11425
rect 21202 11371 21258 11373
rect 21322 11425 21378 11427
rect 21322 11373 21324 11425
rect 21324 11373 21376 11425
rect 21376 11373 21378 11425
rect 21322 11371 21378 11373
rect 21076 11307 21132 11309
rect 21076 11255 21078 11307
rect 21078 11255 21130 11307
rect 21130 11255 21132 11307
rect 21076 11253 21132 11255
rect 21202 11307 21258 11309
rect 21202 11255 21204 11307
rect 21204 11255 21256 11307
rect 21256 11255 21258 11307
rect 21202 11253 21258 11255
rect 21322 11307 21378 11309
rect 21322 11255 21324 11307
rect 21324 11255 21376 11307
rect 21376 11255 21378 11307
rect 21322 11253 21378 11255
rect 512 11049 568 11051
rect 512 10997 514 11049
rect 514 10997 566 11049
rect 566 10997 568 11049
rect 512 10995 568 10997
rect 634 11049 690 11051
rect 634 10997 636 11049
rect 636 10997 688 11049
rect 688 10997 690 11049
rect 634 10995 690 10997
rect 760 11049 816 11051
rect 760 10997 762 11049
rect 762 10997 814 11049
rect 814 10997 816 11049
rect 760 10995 816 10997
rect 512 10902 568 10904
rect 512 10850 514 10902
rect 514 10850 566 10902
rect 566 10850 568 10902
rect 512 10848 568 10850
rect 634 10902 690 10904
rect 634 10850 636 10902
rect 636 10850 688 10902
rect 688 10850 690 10902
rect 634 10848 690 10850
rect 760 10902 816 10904
rect 760 10850 762 10902
rect 762 10850 814 10902
rect 814 10850 816 10902
rect 760 10848 816 10850
rect 512 10765 568 10767
rect 512 10713 514 10765
rect 514 10713 566 10765
rect 566 10713 568 10765
rect 512 10711 568 10713
rect 634 10765 690 10767
rect 634 10713 636 10765
rect 636 10713 688 10765
rect 688 10713 690 10765
rect 634 10711 690 10713
rect 760 10765 816 10767
rect 760 10713 762 10765
rect 762 10713 814 10765
rect 814 10713 816 10765
rect 760 10711 816 10713
rect 22018 10280 22074 10282
rect 22018 10228 22020 10280
rect 22020 10228 22072 10280
rect 22072 10228 22074 10280
rect 22018 10226 22074 10228
rect 22144 10280 22200 10282
rect 22144 10228 22146 10280
rect 22146 10228 22198 10280
rect 22198 10228 22200 10280
rect 22144 10226 22200 10228
rect 22264 10280 22320 10282
rect 22264 10228 22266 10280
rect 22266 10228 22318 10280
rect 22318 10228 22320 10280
rect 22264 10226 22320 10228
rect 22018 10162 22074 10164
rect 22018 10110 22020 10162
rect 22020 10110 22072 10162
rect 22072 10110 22074 10162
rect 22018 10108 22074 10110
rect 22144 10162 22200 10164
rect 22144 10110 22146 10162
rect 22146 10110 22198 10162
rect 22198 10110 22200 10162
rect 22144 10108 22200 10110
rect 22264 10162 22320 10164
rect 22264 10110 22266 10162
rect 22266 10110 22318 10162
rect 22318 10110 22320 10162
rect 22264 10108 22320 10110
rect 512 9287 568 9289
rect 512 9235 514 9287
rect 514 9235 566 9287
rect 566 9235 568 9287
rect 512 9233 568 9235
rect 634 9287 690 9289
rect 634 9235 636 9287
rect 636 9235 688 9287
rect 688 9235 690 9287
rect 634 9233 690 9235
rect 760 9287 816 9289
rect 760 9235 762 9287
rect 762 9235 814 9287
rect 814 9235 816 9287
rect 760 9233 816 9235
rect 512 9140 568 9142
rect 512 9088 514 9140
rect 514 9088 566 9140
rect 566 9088 568 9140
rect 512 9086 568 9088
rect 634 9140 690 9142
rect 634 9088 636 9140
rect 636 9088 688 9140
rect 688 9088 690 9140
rect 634 9086 690 9088
rect 760 9140 816 9142
rect 760 9088 762 9140
rect 762 9088 814 9140
rect 814 9088 816 9140
rect 760 9086 816 9088
rect 512 9003 568 9005
rect 512 8951 514 9003
rect 514 8951 566 9003
rect 566 8951 568 9003
rect 512 8949 568 8951
rect 634 9003 690 9005
rect 634 8951 636 9003
rect 636 8951 688 9003
rect 688 8951 690 9003
rect 634 8949 690 8951
rect 760 9003 816 9005
rect 760 8951 762 9003
rect 762 8951 814 9003
rect 814 8951 816 9003
rect 760 8949 816 8951
rect 511 8627 567 8629
rect 511 8575 513 8627
rect 513 8575 565 8627
rect 565 8575 567 8627
rect 511 8573 567 8575
rect 637 8627 693 8629
rect 637 8575 639 8627
rect 639 8575 691 8627
rect 691 8575 693 8627
rect 637 8573 693 8575
rect 757 8627 813 8629
rect 757 8575 759 8627
rect 759 8575 811 8627
rect 811 8575 813 8627
rect 757 8573 813 8575
rect 511 8509 567 8511
rect 511 8457 513 8509
rect 513 8457 565 8509
rect 565 8457 567 8509
rect 511 8455 567 8457
rect 637 8509 693 8511
rect 637 8457 639 8509
rect 639 8457 691 8509
rect 691 8457 693 8509
rect 637 8455 693 8457
rect 757 8509 813 8511
rect 757 8457 759 8509
rect 759 8457 811 8509
rect 811 8457 813 8509
rect 757 8455 813 8457
rect 21076 8582 21132 8584
rect 21076 8530 21078 8582
rect 21078 8530 21130 8582
rect 21130 8530 21132 8582
rect 21076 8528 21132 8530
rect 21202 8582 21258 8584
rect 21202 8530 21204 8582
rect 21204 8530 21256 8582
rect 21256 8530 21258 8582
rect 21202 8528 21258 8530
rect 21322 8582 21378 8584
rect 21322 8530 21324 8582
rect 21324 8530 21376 8582
rect 21376 8530 21378 8582
rect 21322 8528 21378 8530
rect 21076 8464 21132 8466
rect 21076 8412 21078 8464
rect 21078 8412 21130 8464
rect 21130 8412 21132 8464
rect 21076 8410 21132 8412
rect 21202 8464 21258 8466
rect 21202 8412 21204 8464
rect 21204 8412 21256 8464
rect 21256 8412 21258 8464
rect 21202 8410 21258 8412
rect 21322 8464 21378 8466
rect 21322 8412 21324 8464
rect 21324 8412 21376 8464
rect 21376 8412 21378 8464
rect 21322 8410 21378 8412
rect 511 7516 567 7518
rect 511 7464 513 7516
rect 513 7464 565 7516
rect 565 7464 567 7516
rect 511 7462 567 7464
rect 637 7516 693 7518
rect 637 7464 639 7516
rect 639 7464 691 7516
rect 691 7464 693 7516
rect 637 7462 693 7464
rect 757 7516 813 7518
rect 757 7464 759 7516
rect 759 7464 811 7516
rect 811 7464 813 7516
rect 757 7462 813 7464
rect 511 7398 567 7400
rect 511 7346 513 7398
rect 513 7346 565 7398
rect 565 7346 567 7398
rect 511 7344 567 7346
rect 637 7398 693 7400
rect 637 7346 639 7398
rect 639 7346 691 7398
rect 691 7346 693 7398
rect 637 7344 693 7346
rect 757 7398 813 7400
rect 757 7346 759 7398
rect 759 7346 811 7398
rect 811 7346 813 7398
rect 757 7344 813 7346
rect 21076 7425 21132 7427
rect 21076 7373 21078 7425
rect 21078 7373 21130 7425
rect 21130 7373 21132 7425
rect 21076 7371 21132 7373
rect 21202 7425 21258 7427
rect 21202 7373 21204 7425
rect 21204 7373 21256 7425
rect 21256 7373 21258 7425
rect 21202 7371 21258 7373
rect 21322 7425 21378 7427
rect 21322 7373 21324 7425
rect 21324 7373 21376 7425
rect 21376 7373 21378 7425
rect 21322 7371 21378 7373
rect 21076 7307 21132 7309
rect 21076 7255 21078 7307
rect 21078 7255 21130 7307
rect 21130 7255 21132 7307
rect 21076 7253 21132 7255
rect 21202 7307 21258 7309
rect 21202 7255 21204 7307
rect 21204 7255 21256 7307
rect 21256 7255 21258 7307
rect 21202 7253 21258 7255
rect 21322 7307 21378 7309
rect 21322 7255 21324 7307
rect 21324 7255 21376 7307
rect 21376 7255 21378 7307
rect 21322 7253 21378 7255
rect 512 7049 568 7051
rect 512 6997 514 7049
rect 514 6997 566 7049
rect 566 6997 568 7049
rect 512 6995 568 6997
rect 634 7049 690 7051
rect 634 6997 636 7049
rect 636 6997 688 7049
rect 688 6997 690 7049
rect 634 6995 690 6997
rect 760 7049 816 7051
rect 760 6997 762 7049
rect 762 6997 814 7049
rect 814 6997 816 7049
rect 760 6995 816 6997
rect 512 6902 568 6904
rect 512 6850 514 6902
rect 514 6850 566 6902
rect 566 6850 568 6902
rect 512 6848 568 6850
rect 634 6902 690 6904
rect 634 6850 636 6902
rect 636 6850 688 6902
rect 688 6850 690 6902
rect 634 6848 690 6850
rect 760 6902 816 6904
rect 760 6850 762 6902
rect 762 6850 814 6902
rect 814 6850 816 6902
rect 760 6848 816 6850
rect 512 6765 568 6767
rect 512 6713 514 6765
rect 514 6713 566 6765
rect 566 6713 568 6765
rect 512 6711 568 6713
rect 634 6765 690 6767
rect 634 6713 636 6765
rect 636 6713 688 6765
rect 688 6713 690 6765
rect 634 6711 690 6713
rect 760 6765 816 6767
rect 760 6713 762 6765
rect 762 6713 814 6765
rect 814 6713 816 6765
rect 760 6711 816 6713
rect 22018 6268 22074 6270
rect 22018 6216 22020 6268
rect 22020 6216 22072 6268
rect 22072 6216 22074 6268
rect 22018 6214 22074 6216
rect 22144 6268 22200 6270
rect 22144 6216 22146 6268
rect 22146 6216 22198 6268
rect 22198 6216 22200 6268
rect 22144 6214 22200 6216
rect 22264 6268 22320 6270
rect 22264 6216 22266 6268
rect 22266 6216 22318 6268
rect 22318 6216 22320 6268
rect 22264 6214 22320 6216
rect 22018 6150 22074 6152
rect 22018 6098 22020 6150
rect 22020 6098 22072 6150
rect 22072 6098 22074 6150
rect 22018 6096 22074 6098
rect 22144 6150 22200 6152
rect 22144 6098 22146 6150
rect 22146 6098 22198 6150
rect 22198 6098 22200 6150
rect 22144 6096 22200 6098
rect 22264 6150 22320 6152
rect 22264 6098 22266 6150
rect 22266 6098 22318 6150
rect 22318 6098 22320 6150
rect 22264 6096 22320 6098
rect 512 5288 568 5290
rect 512 5236 514 5288
rect 514 5236 566 5288
rect 566 5236 568 5288
rect 512 5234 568 5236
rect 634 5288 690 5290
rect 634 5236 636 5288
rect 636 5236 688 5288
rect 688 5236 690 5288
rect 634 5234 690 5236
rect 760 5288 816 5290
rect 760 5236 762 5288
rect 762 5236 814 5288
rect 814 5236 816 5288
rect 760 5234 816 5236
rect 512 5141 568 5143
rect 512 5089 514 5141
rect 514 5089 566 5141
rect 566 5089 568 5141
rect 512 5087 568 5089
rect 634 5141 690 5143
rect 634 5089 636 5141
rect 636 5089 688 5141
rect 688 5089 690 5141
rect 634 5087 690 5089
rect 760 5141 816 5143
rect 760 5089 762 5141
rect 762 5089 814 5141
rect 814 5089 816 5141
rect 760 5087 816 5089
rect 512 5004 568 5006
rect 512 4952 514 5004
rect 514 4952 566 5004
rect 566 4952 568 5004
rect 512 4950 568 4952
rect 634 5004 690 5006
rect 634 4952 636 5004
rect 636 4952 688 5004
rect 688 4952 690 5004
rect 634 4950 690 4952
rect 760 5004 816 5006
rect 760 4952 762 5004
rect 762 4952 814 5004
rect 814 4952 816 5004
rect 760 4950 816 4952
rect 511 4693 567 4695
rect 511 4641 513 4693
rect 513 4641 565 4693
rect 565 4641 567 4693
rect 511 4639 567 4641
rect 637 4693 693 4695
rect 637 4641 639 4693
rect 639 4641 691 4693
rect 691 4641 693 4693
rect 637 4639 693 4641
rect 757 4693 813 4695
rect 757 4641 759 4693
rect 759 4641 811 4693
rect 811 4641 813 4693
rect 757 4639 813 4641
rect 511 4575 567 4577
rect 511 4523 513 4575
rect 513 4523 565 4575
rect 565 4523 567 4575
rect 511 4521 567 4523
rect 637 4575 693 4577
rect 637 4523 639 4575
rect 639 4523 691 4575
rect 691 4523 693 4575
rect 637 4521 693 4523
rect 757 4575 813 4577
rect 757 4523 759 4575
rect 759 4523 811 4575
rect 811 4523 813 4575
rect 757 4521 813 4523
rect 21076 4582 21132 4584
rect 21076 4530 21078 4582
rect 21078 4530 21130 4582
rect 21130 4530 21132 4582
rect 21076 4528 21132 4530
rect 21202 4582 21258 4584
rect 21202 4530 21204 4582
rect 21204 4530 21256 4582
rect 21256 4530 21258 4582
rect 21202 4528 21258 4530
rect 21322 4582 21378 4584
rect 21322 4530 21324 4582
rect 21324 4530 21376 4582
rect 21376 4530 21378 4582
rect 21322 4528 21378 4530
rect 21076 4464 21132 4466
rect 21076 4412 21078 4464
rect 21078 4412 21130 4464
rect 21130 4412 21132 4464
rect 21076 4410 21132 4412
rect 21202 4464 21258 4466
rect 21202 4412 21204 4464
rect 21204 4412 21256 4464
rect 21256 4412 21258 4464
rect 21202 4410 21258 4412
rect 21322 4464 21378 4466
rect 21322 4412 21324 4464
rect 21324 4412 21376 4464
rect 21376 4412 21378 4464
rect 21322 4410 21378 4412
rect 511 3516 567 3518
rect 511 3464 513 3516
rect 513 3464 565 3516
rect 565 3464 567 3516
rect 511 3462 567 3464
rect 637 3516 693 3518
rect 637 3464 639 3516
rect 639 3464 691 3516
rect 691 3464 693 3516
rect 637 3462 693 3464
rect 757 3516 813 3518
rect 757 3464 759 3516
rect 759 3464 811 3516
rect 811 3464 813 3516
rect 757 3462 813 3464
rect 511 3398 567 3400
rect 511 3346 513 3398
rect 513 3346 565 3398
rect 565 3346 567 3398
rect 511 3344 567 3346
rect 637 3398 693 3400
rect 637 3346 639 3398
rect 639 3346 691 3398
rect 691 3346 693 3398
rect 637 3344 693 3346
rect 757 3398 813 3400
rect 757 3346 759 3398
rect 759 3346 811 3398
rect 811 3346 813 3398
rect 757 3344 813 3346
rect 21076 3425 21132 3427
rect 21076 3373 21078 3425
rect 21078 3373 21130 3425
rect 21130 3373 21132 3425
rect 21076 3371 21132 3373
rect 21202 3425 21258 3427
rect 21202 3373 21204 3425
rect 21204 3373 21256 3425
rect 21256 3373 21258 3425
rect 21202 3371 21258 3373
rect 21322 3425 21378 3427
rect 21322 3373 21324 3425
rect 21324 3373 21376 3425
rect 21376 3373 21378 3425
rect 21322 3371 21378 3373
rect 21076 3307 21132 3309
rect 21076 3255 21078 3307
rect 21078 3255 21130 3307
rect 21130 3255 21132 3307
rect 21076 3253 21132 3255
rect 21202 3307 21258 3309
rect 21202 3255 21204 3307
rect 21204 3255 21256 3307
rect 21256 3255 21258 3307
rect 21202 3253 21258 3255
rect 21322 3307 21378 3309
rect 21322 3255 21324 3307
rect 21324 3255 21376 3307
rect 21376 3255 21378 3307
rect 21322 3253 21378 3255
rect 512 3049 568 3051
rect 512 2997 514 3049
rect 514 2997 566 3049
rect 566 2997 568 3049
rect 512 2995 568 2997
rect 634 3049 690 3051
rect 634 2997 636 3049
rect 636 2997 688 3049
rect 688 2997 690 3049
rect 634 2995 690 2997
rect 760 3049 816 3051
rect 760 2997 762 3049
rect 762 2997 814 3049
rect 814 2997 816 3049
rect 760 2995 816 2997
rect 512 2902 568 2904
rect 512 2850 514 2902
rect 514 2850 566 2902
rect 566 2850 568 2902
rect 512 2848 568 2850
rect 634 2902 690 2904
rect 634 2850 636 2902
rect 636 2850 688 2902
rect 688 2850 690 2902
rect 634 2848 690 2850
rect 760 2902 816 2904
rect 760 2850 762 2902
rect 762 2850 814 2902
rect 814 2850 816 2902
rect 760 2848 816 2850
rect 512 2765 568 2767
rect 512 2713 514 2765
rect 514 2713 566 2765
rect 566 2713 568 2765
rect 512 2711 568 2713
rect 634 2765 690 2767
rect 634 2713 636 2765
rect 636 2713 688 2765
rect 688 2713 690 2765
rect 634 2711 690 2713
rect 760 2765 816 2767
rect 760 2713 762 2765
rect 762 2713 814 2765
rect 814 2713 816 2765
rect 760 2711 816 2713
rect 22018 2268 22074 2270
rect 22018 2216 22020 2268
rect 22020 2216 22072 2268
rect 22072 2216 22074 2268
rect 22018 2214 22074 2216
rect 22144 2268 22200 2270
rect 22144 2216 22146 2268
rect 22146 2216 22198 2268
rect 22198 2216 22200 2268
rect 22144 2214 22200 2216
rect 22264 2268 22320 2270
rect 22264 2216 22266 2268
rect 22266 2216 22318 2268
rect 22318 2216 22320 2268
rect 22264 2214 22320 2216
rect 22018 2150 22074 2152
rect 22018 2098 22020 2150
rect 22020 2098 22072 2150
rect 22072 2098 22074 2150
rect 22018 2096 22074 2098
rect 22144 2150 22200 2152
rect 22144 2098 22146 2150
rect 22146 2098 22198 2150
rect 22198 2098 22200 2150
rect 22144 2096 22200 2098
rect 22264 2150 22320 2152
rect 22264 2098 22266 2150
rect 22266 2098 22318 2150
rect 22318 2098 22320 2150
rect 22264 2096 22320 2098
rect 512 1288 568 1290
rect 512 1236 514 1288
rect 514 1236 566 1288
rect 566 1236 568 1288
rect 512 1234 568 1236
rect 634 1288 690 1290
rect 634 1236 636 1288
rect 636 1236 688 1288
rect 688 1236 690 1288
rect 634 1234 690 1236
rect 760 1288 816 1290
rect 760 1236 762 1288
rect 762 1236 814 1288
rect 814 1236 816 1288
rect 760 1234 816 1236
rect 512 1141 568 1143
rect 512 1089 514 1141
rect 514 1089 566 1141
rect 566 1089 568 1141
rect 512 1087 568 1089
rect 634 1141 690 1143
rect 634 1089 636 1141
rect 636 1089 688 1141
rect 688 1089 690 1141
rect 634 1087 690 1089
rect 760 1141 816 1143
rect 760 1089 762 1141
rect 762 1089 814 1141
rect 814 1089 816 1141
rect 760 1087 816 1089
rect 512 1004 568 1006
rect 512 952 514 1004
rect 514 952 566 1004
rect 566 952 568 1004
rect 512 950 568 952
rect 634 1004 690 1006
rect 634 952 636 1004
rect 636 952 688 1004
rect 688 952 690 1004
rect 634 950 690 952
rect 760 1004 816 1006
rect 760 952 762 1004
rect 762 952 814 1004
rect 814 952 816 1004
rect 760 950 816 952
rect 511 693 567 695
rect 511 641 513 693
rect 513 641 565 693
rect 565 641 567 693
rect 511 639 567 641
rect 637 693 693 695
rect 637 641 639 693
rect 639 641 691 693
rect 691 641 693 693
rect 637 639 693 641
rect 757 693 813 695
rect 757 641 759 693
rect 759 641 811 693
rect 811 641 813 693
rect 757 639 813 641
rect 511 575 567 577
rect 511 523 513 575
rect 513 523 565 575
rect 565 523 567 575
rect 511 521 567 523
rect 637 575 693 577
rect 637 523 639 575
rect 639 523 691 575
rect 691 523 693 575
rect 637 521 693 523
rect 757 575 813 577
rect 757 523 759 575
rect 759 523 811 575
rect 811 523 813 575
rect 757 521 813 523
rect 21076 582 21132 584
rect 21076 530 21078 582
rect 21078 530 21130 582
rect 21130 530 21132 582
rect 21076 528 21132 530
rect 21202 582 21258 584
rect 21202 530 21204 582
rect 21204 530 21256 582
rect 21256 530 21258 582
rect 21202 528 21258 530
rect 21322 582 21378 584
rect 21322 530 21324 582
rect 21324 530 21376 582
rect 21376 530 21378 582
rect 21322 528 21378 530
rect 21076 464 21132 466
rect 21076 412 21078 464
rect 21078 412 21130 464
rect 21130 412 21132 464
rect 21076 410 21132 412
rect 21202 464 21258 466
rect 21202 412 21204 464
rect 21204 412 21256 464
rect 21256 412 21258 464
rect 21202 410 21258 412
rect 21322 464 21378 466
rect 21322 412 21324 464
rect 21324 412 21376 464
rect 21376 412 21378 464
rect 21322 410 21378 412
<< metal3 >>
rect 21026 75486 21426 75517
rect 463 75446 864 75477
rect 463 75382 507 75446
rect 571 75382 633 75446
rect 697 75382 753 75446
rect 817 75382 864 75446
rect 463 75328 864 75382
rect 463 75264 507 75328
rect 571 75264 633 75328
rect 697 75264 753 75328
rect 817 75264 864 75328
rect 463 75222 864 75264
rect 21026 75422 21072 75486
rect 21136 75422 21198 75486
rect 21262 75422 21318 75486
rect 21382 75422 21426 75486
rect 21026 75368 21426 75422
rect 21026 75304 21072 75368
rect 21136 75304 21198 75368
rect 21262 75304 21318 75368
rect 21382 75304 21426 75368
rect 21026 75262 21426 75304
rect 463 75054 863 75109
rect 463 74990 508 75054
rect 572 74990 630 75054
rect 694 74990 756 75054
rect 820 74990 863 75054
rect 463 74907 863 74990
rect 463 74843 508 74907
rect 572 74843 630 74907
rect 694 74843 756 74907
rect 820 74843 863 74907
rect 463 74770 863 74843
rect 463 74706 508 74770
rect 572 74706 630 74770
rect 694 74706 756 74770
rect 820 74706 863 74770
rect 463 74650 863 74706
rect 21970 74065 22370 74096
rect 21970 74001 22014 74065
rect 22078 74001 22140 74065
rect 22204 74001 22260 74065
rect 22324 74001 22370 74065
rect 21970 73947 22370 74001
rect 21970 73883 22014 73947
rect 22078 73883 22140 73947
rect 22204 73883 22260 73947
rect 22324 73883 22370 73947
rect 21970 73841 22370 73883
rect 463 73294 863 73349
rect 463 73230 508 73294
rect 572 73230 630 73294
rect 694 73230 756 73294
rect 820 73230 863 73294
rect 463 73147 863 73230
rect 463 73083 508 73147
rect 572 73083 630 73147
rect 694 73083 756 73147
rect 820 73083 863 73147
rect 463 73010 863 73083
rect 463 72946 508 73010
rect 572 72946 630 73010
rect 694 72946 756 73010
rect 820 72946 863 73010
rect 463 72890 863 72946
rect 463 72773 864 72804
rect 463 72709 507 72773
rect 571 72709 633 72773
rect 697 72709 753 72773
rect 817 72709 864 72773
rect 463 72655 864 72709
rect 463 72591 507 72655
rect 571 72591 633 72655
rect 697 72591 753 72655
rect 817 72591 864 72655
rect 463 72549 864 72591
rect 21028 72689 21428 72720
rect 21028 72625 21072 72689
rect 21136 72625 21198 72689
rect 21262 72625 21318 72689
rect 21382 72625 21428 72689
rect 21028 72571 21428 72625
rect 21028 72507 21072 72571
rect 21136 72507 21198 72571
rect 21262 72507 21318 72571
rect 21382 72507 21428 72571
rect 21028 72465 21428 72507
rect 21026 71486 21426 71517
rect 463 71446 864 71477
rect 463 71382 507 71446
rect 571 71382 633 71446
rect 697 71382 753 71446
rect 817 71382 864 71446
rect 463 71328 864 71382
rect 463 71264 507 71328
rect 571 71264 633 71328
rect 697 71264 753 71328
rect 817 71264 864 71328
rect 463 71222 864 71264
rect 21026 71422 21072 71486
rect 21136 71422 21198 71486
rect 21262 71422 21318 71486
rect 21382 71422 21426 71486
rect 21026 71368 21426 71422
rect 21026 71304 21072 71368
rect 21136 71304 21198 71368
rect 21262 71304 21318 71368
rect 21382 71304 21426 71368
rect 21026 71262 21426 71304
rect 463 71054 863 71109
rect 463 70990 508 71054
rect 572 70990 630 71054
rect 694 70990 756 71054
rect 820 70990 863 71054
rect 463 70907 863 70990
rect 463 70843 508 70907
rect 572 70843 630 70907
rect 694 70843 756 70907
rect 820 70843 863 70907
rect 463 70770 863 70843
rect 463 70706 508 70770
rect 572 70706 630 70770
rect 694 70706 756 70770
rect 820 70706 863 70770
rect 463 70650 863 70706
rect 21970 70065 22370 70096
rect 21970 70001 22014 70065
rect 22078 70001 22140 70065
rect 22204 70001 22260 70065
rect 22324 70001 22370 70065
rect 21970 69947 22370 70001
rect 21970 69883 22014 69947
rect 22078 69883 22140 69947
rect 22204 69883 22260 69947
rect 22324 69883 22370 69947
rect 21970 69841 22370 69883
rect 463 69294 863 69349
rect 463 69230 508 69294
rect 572 69230 630 69294
rect 694 69230 756 69294
rect 820 69230 863 69294
rect 463 69147 863 69230
rect 463 69083 508 69147
rect 572 69083 630 69147
rect 694 69083 756 69147
rect 820 69083 863 69147
rect 463 69010 863 69083
rect 463 68946 508 69010
rect 572 68946 630 69010
rect 694 68946 756 69010
rect 820 68946 863 69010
rect 463 68890 863 68946
rect 463 68773 864 68804
rect 463 68709 507 68773
rect 571 68709 633 68773
rect 697 68709 753 68773
rect 817 68709 864 68773
rect 463 68655 864 68709
rect 463 68591 507 68655
rect 571 68591 633 68655
rect 697 68591 753 68655
rect 817 68591 864 68655
rect 463 68549 864 68591
rect 21028 68689 21428 68720
rect 21028 68625 21072 68689
rect 21136 68625 21198 68689
rect 21262 68625 21318 68689
rect 21382 68625 21428 68689
rect 21028 68571 21428 68625
rect 21028 68507 21072 68571
rect 21136 68507 21198 68571
rect 21262 68507 21318 68571
rect 21382 68507 21428 68571
rect 21028 68465 21428 68507
rect 21026 67486 21426 67517
rect 463 67444 864 67475
rect 463 67380 507 67444
rect 571 67380 633 67444
rect 697 67380 753 67444
rect 817 67380 864 67444
rect 463 67326 864 67380
rect 463 67262 507 67326
rect 571 67262 633 67326
rect 697 67262 753 67326
rect 817 67262 864 67326
rect 21026 67422 21072 67486
rect 21136 67422 21198 67486
rect 21262 67422 21318 67486
rect 21382 67422 21426 67486
rect 21026 67368 21426 67422
rect 21026 67304 21072 67368
rect 21136 67304 21198 67368
rect 21262 67304 21318 67368
rect 21382 67304 21426 67368
rect 21026 67262 21426 67304
rect 463 67220 864 67262
rect 463 67054 863 67109
rect 463 66990 508 67054
rect 572 66990 630 67054
rect 694 66990 756 67054
rect 820 66990 863 67054
rect 463 66907 863 66990
rect 463 66843 508 66907
rect 572 66843 630 66907
rect 694 66843 756 66907
rect 820 66843 863 66907
rect 463 66770 863 66843
rect 463 66706 508 66770
rect 572 66706 630 66770
rect 694 66706 756 66770
rect 820 66706 863 66770
rect 463 66650 863 66706
rect 21970 66052 22370 66083
rect 21970 65988 22014 66052
rect 22078 65988 22140 66052
rect 22204 65988 22260 66052
rect 22324 65988 22370 66052
rect 21970 65934 22370 65988
rect 21970 65870 22014 65934
rect 22078 65870 22140 65934
rect 22204 65870 22260 65934
rect 22324 65870 22370 65934
rect 21970 65828 22370 65870
rect 463 65295 863 65350
rect 463 65231 508 65295
rect 572 65231 630 65295
rect 694 65231 756 65295
rect 820 65231 863 65295
rect 463 65148 863 65231
rect 463 65084 508 65148
rect 572 65084 630 65148
rect 694 65084 756 65148
rect 820 65084 863 65148
rect 463 65011 863 65084
rect 463 64947 508 65011
rect 572 64947 630 65011
rect 694 64947 756 65011
rect 820 64947 863 65011
rect 463 64891 863 64947
rect 463 64704 864 64735
rect 463 64640 507 64704
rect 571 64640 633 64704
rect 697 64640 753 64704
rect 817 64640 864 64704
rect 463 64586 864 64640
rect 463 64522 507 64586
rect 571 64522 633 64586
rect 697 64522 753 64586
rect 817 64522 864 64586
rect 463 64480 864 64522
rect 21028 64689 21428 64720
rect 21028 64625 21072 64689
rect 21136 64625 21198 64689
rect 21262 64625 21318 64689
rect 21382 64625 21428 64689
rect 21028 64571 21428 64625
rect 21028 64507 21072 64571
rect 21136 64507 21198 64571
rect 21262 64507 21318 64571
rect 21382 64507 21428 64571
rect 21028 64465 21428 64507
rect 463 63526 864 63557
rect 463 63462 507 63526
rect 571 63462 633 63526
rect 697 63462 753 63526
rect 817 63462 864 63526
rect 463 63408 864 63462
rect 463 63344 507 63408
rect 571 63344 633 63408
rect 697 63344 753 63408
rect 817 63344 864 63408
rect 463 63302 864 63344
rect 21026 63486 21426 63517
rect 21026 63422 21072 63486
rect 21136 63422 21198 63486
rect 21262 63422 21318 63486
rect 21382 63422 21426 63486
rect 21026 63368 21426 63422
rect 21026 63304 21072 63368
rect 21136 63304 21198 63368
rect 21262 63304 21318 63368
rect 21382 63304 21426 63368
rect 21026 63262 21426 63304
rect 464 63068 864 63109
rect 463 63054 864 63068
rect 463 62990 508 63054
rect 572 62990 630 63054
rect 694 62990 756 63054
rect 820 62990 864 63054
rect 463 62907 864 62990
rect 463 62843 508 62907
rect 572 62843 630 62907
rect 694 62843 756 62907
rect 820 62843 864 62907
rect 463 62770 864 62843
rect 463 62706 508 62770
rect 572 62706 630 62770
rect 694 62706 756 62770
rect 820 62706 864 62770
rect 463 62650 864 62706
rect 21970 62051 22370 62082
rect 21970 61987 22014 62051
rect 22078 61987 22140 62051
rect 22204 61987 22260 62051
rect 22324 61987 22370 62051
rect 21970 61933 22370 61987
rect 21970 61869 22014 61933
rect 22078 61869 22140 61933
rect 22204 61869 22260 61933
rect 22324 61869 22370 61933
rect 21970 61827 22370 61869
rect 463 61295 863 61350
rect 463 61231 508 61295
rect 572 61231 630 61295
rect 694 61231 756 61295
rect 820 61231 863 61295
rect 463 61148 863 61231
rect 463 61084 508 61148
rect 572 61084 630 61148
rect 694 61084 756 61148
rect 820 61084 863 61148
rect 463 61011 863 61084
rect 463 60947 508 61011
rect 572 60947 630 61011
rect 694 60947 756 61011
rect 820 60947 863 61011
rect 463 60891 863 60947
rect 463 60678 866 60709
rect 463 60614 507 60678
rect 571 60614 633 60678
rect 697 60614 753 60678
rect 817 60614 866 60678
rect 463 60560 866 60614
rect 463 60496 507 60560
rect 571 60496 633 60560
rect 697 60496 753 60560
rect 817 60496 866 60560
rect 463 60454 866 60496
rect 21028 60689 21428 60720
rect 21028 60625 21072 60689
rect 21136 60625 21198 60689
rect 21262 60625 21318 60689
rect 21382 60625 21428 60689
rect 21028 60571 21428 60625
rect 21028 60507 21072 60571
rect 21136 60507 21198 60571
rect 21262 60507 21318 60571
rect 21382 60507 21428 60571
rect 21028 60465 21428 60507
rect 21027 59540 21427 59571
rect 463 59475 864 59506
rect 463 59411 507 59475
rect 571 59411 633 59475
rect 697 59411 753 59475
rect 817 59411 864 59475
rect 463 59357 864 59411
rect 463 59293 507 59357
rect 571 59293 633 59357
rect 697 59293 753 59357
rect 817 59293 864 59357
rect 21027 59476 21072 59540
rect 21136 59476 21198 59540
rect 21262 59476 21318 59540
rect 21382 59476 21427 59540
rect 21027 59422 21427 59476
rect 21027 59358 21072 59422
rect 21136 59358 21198 59422
rect 21262 59358 21318 59422
rect 21382 59358 21427 59422
rect 21027 59316 21427 59358
rect 463 59251 864 59293
rect 464 59068 864 59109
rect 463 59054 864 59068
rect 463 58990 508 59054
rect 572 58990 630 59054
rect 694 58990 756 59054
rect 820 58990 864 59054
rect 463 58907 864 58990
rect 463 58843 508 58907
rect 572 58843 630 58907
rect 694 58843 756 58907
rect 820 58843 864 58907
rect 463 58770 864 58843
rect 463 58706 508 58770
rect 572 58706 630 58770
rect 694 58706 756 58770
rect 820 58706 864 58770
rect 463 58650 864 58706
rect 21970 58090 22370 58121
rect 21970 58026 22014 58090
rect 22078 58026 22140 58090
rect 22204 58026 22260 58090
rect 22324 58026 22370 58090
rect 21970 57972 22370 58026
rect 21970 57908 22014 57972
rect 22078 57908 22140 57972
rect 22204 57908 22260 57972
rect 22324 57908 22370 57972
rect 21970 57866 22370 57908
rect 463 57293 863 57348
rect 463 57229 508 57293
rect 572 57229 630 57293
rect 694 57229 756 57293
rect 820 57229 863 57293
rect 463 57146 863 57229
rect 463 57082 508 57146
rect 572 57082 630 57146
rect 694 57082 756 57146
rect 820 57082 863 57146
rect 463 57009 863 57082
rect 463 56945 508 57009
rect 572 56945 630 57009
rect 694 56945 756 57009
rect 820 56945 863 57009
rect 463 56889 863 56945
rect 463 56698 864 56729
rect 463 56634 507 56698
rect 571 56634 633 56698
rect 697 56634 753 56698
rect 817 56634 864 56698
rect 463 56580 864 56634
rect 463 56516 507 56580
rect 571 56516 633 56580
rect 697 56516 753 56580
rect 817 56516 864 56580
rect 463 56474 864 56516
rect 21028 56624 21428 56655
rect 21028 56560 21072 56624
rect 21136 56560 21198 56624
rect 21262 56560 21318 56624
rect 21382 56560 21428 56624
rect 21028 56506 21428 56560
rect 21028 56442 21072 56506
rect 21136 56442 21198 56506
rect 21262 56442 21318 56506
rect 21382 56442 21428 56506
rect 21028 56400 21428 56442
rect 463 55491 866 55522
rect 463 55427 507 55491
rect 571 55427 633 55491
rect 697 55427 753 55491
rect 817 55427 866 55491
rect 463 55373 866 55427
rect 463 55309 507 55373
rect 571 55309 633 55373
rect 697 55309 753 55373
rect 817 55309 866 55373
rect 463 55267 866 55309
rect 21027 55441 21427 55472
rect 21027 55377 21072 55441
rect 21136 55377 21198 55441
rect 21262 55377 21318 55441
rect 21382 55377 21427 55441
rect 21027 55323 21427 55377
rect 21027 55259 21072 55323
rect 21136 55259 21198 55323
rect 21262 55259 21318 55323
rect 21382 55259 21427 55323
rect 21027 55217 21427 55259
rect 463 55054 863 55109
rect 463 54990 508 55054
rect 572 54990 630 55054
rect 694 54990 756 55054
rect 820 54990 863 55054
rect 463 54907 863 54990
rect 463 54843 508 54907
rect 572 54843 630 54907
rect 694 54843 756 54907
rect 820 54843 863 54907
rect 463 54770 863 54843
rect 463 54706 508 54770
rect 572 54706 630 54770
rect 694 54706 756 54770
rect 820 54706 863 54770
rect 463 54650 863 54706
rect 21970 54073 22370 54104
rect 21970 54009 22014 54073
rect 22078 54009 22140 54073
rect 22204 54009 22260 54073
rect 22324 54009 22370 54073
rect 21970 53955 22370 54009
rect 21970 53891 22014 53955
rect 22078 53891 22140 53955
rect 22204 53891 22260 53955
rect 22324 53891 22370 53955
rect 21970 53849 22370 53891
rect 463 53295 863 53350
rect 463 53231 508 53295
rect 572 53231 630 53295
rect 694 53231 756 53295
rect 820 53231 863 53295
rect 463 53148 863 53231
rect 463 53084 508 53148
rect 572 53084 630 53148
rect 694 53084 756 53148
rect 820 53084 863 53148
rect 463 53011 863 53084
rect 463 52947 508 53011
rect 572 52947 630 53011
rect 694 52947 756 53011
rect 820 52947 863 53011
rect 463 52891 863 52947
rect 463 52725 864 52756
rect 463 52661 507 52725
rect 571 52661 633 52725
rect 697 52661 753 52725
rect 817 52661 864 52725
rect 463 52607 864 52661
rect 463 52543 507 52607
rect 571 52543 633 52607
rect 697 52543 753 52607
rect 817 52543 864 52607
rect 463 52501 864 52543
rect 21028 52569 21428 52600
rect 21028 52505 21072 52569
rect 21136 52505 21198 52569
rect 21262 52505 21318 52569
rect 21382 52505 21428 52569
rect 21028 52451 21428 52505
rect 21028 52387 21072 52451
rect 21136 52387 21198 52451
rect 21262 52387 21318 52451
rect 21382 52387 21428 52451
rect 21028 52345 21428 52387
rect 463 51538 864 51569
rect 463 51474 507 51538
rect 571 51474 633 51538
rect 697 51474 753 51538
rect 817 51474 864 51538
rect 463 51420 864 51474
rect 463 51356 507 51420
rect 571 51356 633 51420
rect 697 51356 753 51420
rect 817 51356 864 51420
rect 463 51314 864 51356
rect 21028 51434 21428 51465
rect 21028 51370 21072 51434
rect 21136 51370 21198 51434
rect 21262 51370 21318 51434
rect 21382 51370 21428 51434
rect 21028 51316 21428 51370
rect 21028 51252 21072 51316
rect 21136 51252 21198 51316
rect 21262 51252 21318 51316
rect 21382 51252 21428 51316
rect 21028 51210 21428 51252
rect 463 51054 863 51109
rect 463 50990 508 51054
rect 572 50990 630 51054
rect 694 50990 756 51054
rect 820 50990 863 51054
rect 463 50907 863 50990
rect 463 50843 508 50907
rect 572 50843 630 50907
rect 694 50843 756 50907
rect 820 50843 863 50907
rect 463 50770 863 50843
rect 463 50706 508 50770
rect 572 50706 630 50770
rect 694 50706 756 50770
rect 820 50706 863 50770
rect 463 50650 863 50706
rect 21970 50152 22370 50183
rect 21970 50088 22014 50152
rect 22078 50088 22140 50152
rect 22204 50088 22260 50152
rect 22324 50088 22370 50152
rect 21970 50034 22370 50088
rect 21970 49970 22014 50034
rect 22078 49970 22140 50034
rect 22204 49970 22260 50034
rect 22324 49970 22370 50034
rect 21970 49928 22370 49970
rect 463 49295 863 49350
rect 463 49231 508 49295
rect 572 49231 630 49295
rect 694 49231 756 49295
rect 820 49231 863 49295
rect 463 49148 863 49231
rect 463 49084 508 49148
rect 572 49084 630 49148
rect 694 49084 756 49148
rect 820 49084 863 49148
rect 463 49011 863 49084
rect 463 48947 508 49011
rect 572 48947 630 49011
rect 694 48947 756 49011
rect 820 48947 863 49011
rect 463 48891 863 48947
rect 463 48716 864 48747
rect 463 48652 507 48716
rect 571 48652 633 48716
rect 697 48652 753 48716
rect 817 48652 864 48716
rect 463 48598 864 48652
rect 463 48534 507 48598
rect 571 48534 633 48598
rect 697 48534 753 48598
rect 817 48534 864 48598
rect 463 48492 864 48534
rect 21028 48675 21428 48706
rect 21028 48611 21072 48675
rect 21136 48611 21198 48675
rect 21262 48611 21318 48675
rect 21382 48611 21428 48675
rect 21028 48557 21428 48611
rect 21028 48493 21072 48557
rect 21136 48493 21198 48557
rect 21262 48493 21318 48557
rect 21382 48493 21428 48557
rect 21028 48451 21428 48493
rect 463 47563 864 47594
rect 463 47499 507 47563
rect 571 47499 633 47563
rect 697 47499 753 47563
rect 817 47499 864 47563
rect 463 47445 864 47499
rect 463 47381 507 47445
rect 571 47381 633 47445
rect 697 47381 753 47445
rect 817 47381 864 47445
rect 463 47339 864 47381
rect 21028 47522 21428 47553
rect 21028 47458 21072 47522
rect 21136 47458 21198 47522
rect 21262 47458 21318 47522
rect 21382 47458 21428 47522
rect 21028 47404 21428 47458
rect 21028 47340 21072 47404
rect 21136 47340 21198 47404
rect 21262 47340 21318 47404
rect 21382 47340 21428 47404
rect 21028 47298 21428 47340
rect 463 47054 863 47109
rect 463 46990 508 47054
rect 572 46990 630 47054
rect 694 46990 756 47054
rect 820 46990 863 47054
rect 463 46907 863 46990
rect 463 46843 508 46907
rect 572 46843 630 46907
rect 694 46843 756 46907
rect 820 46843 863 46907
rect 463 46770 863 46843
rect 463 46706 508 46770
rect 572 46706 630 46770
rect 694 46706 756 46770
rect 820 46706 863 46770
rect 463 46650 863 46706
rect 21970 45894 22370 45925
rect 21970 45830 22014 45894
rect 22078 45830 22140 45894
rect 22204 45830 22260 45894
rect 22324 45830 22370 45894
rect 21970 45776 22370 45830
rect 21970 45712 22014 45776
rect 22078 45712 22140 45776
rect 22204 45712 22260 45776
rect 22324 45712 22370 45776
rect 21970 45670 22370 45712
rect 463 45294 863 45350
rect 463 45230 508 45294
rect 572 45230 630 45294
rect 694 45230 756 45294
rect 820 45230 863 45294
rect 463 45147 863 45230
rect 463 45083 508 45147
rect 572 45083 630 45147
rect 694 45083 756 45147
rect 820 45083 863 45147
rect 463 45010 863 45083
rect 463 44946 508 45010
rect 572 44946 630 45010
rect 694 44946 756 45010
rect 820 44946 863 45010
rect 463 44891 863 44946
rect 463 44890 836 44891
rect 463 44503 863 44534
rect 463 44439 507 44503
rect 571 44439 633 44503
rect 697 44439 753 44503
rect 817 44439 863 44503
rect 463 44385 863 44439
rect 463 44321 507 44385
rect 571 44321 633 44385
rect 697 44321 753 44385
rect 817 44321 863 44385
rect 463 44279 863 44321
rect 21028 44406 21428 44437
rect 21028 44342 21072 44406
rect 21136 44342 21198 44406
rect 21262 44342 21318 44406
rect 21382 44342 21428 44406
rect 21028 44288 21428 44342
rect 21028 44224 21072 44288
rect 21136 44224 21198 44288
rect 21262 44224 21318 44288
rect 21382 44224 21428 44288
rect 21028 44182 21428 44224
rect 21970 43828 22370 43870
rect 21970 43524 22040 43828
rect 22264 43524 22370 43828
rect 21970 43480 22370 43524
rect 2248 39925 2401 39940
rect 2248 39861 2249 39925
rect 2248 39845 2257 39861
rect 2393 39845 2401 39861
rect 2248 39781 2249 39845
rect 2313 39781 2337 39789
rect 2248 39775 2401 39781
rect 3352 39905 4345 39920
rect 3352 39904 4192 39905
rect 3352 39768 3361 39904
rect 3497 39841 4192 39904
rect 4256 39841 4280 39905
rect 4344 39841 4345 39905
rect 3497 39825 4345 39841
rect 3497 39768 4192 39825
rect 3352 39761 4192 39768
rect 4256 39761 4280 39825
rect 4344 39761 4345 39825
rect 3352 39754 4345 39761
rect 0 39733 400 39752
rect 0 39669 39 39733
rect 103 39669 164 39733
rect 228 39669 290 39733
rect 354 39669 400 39733
rect 0 39627 400 39669
rect 0 39563 39 39627
rect 103 39563 164 39627
rect 228 39563 290 39627
rect 354 39563 400 39627
rect 0 39528 400 39563
rect 21502 39718 21902 39752
rect 21502 39654 21543 39718
rect 21607 39654 21668 39718
rect 21732 39654 21793 39718
rect 21857 39654 21902 39718
rect 21502 39598 21902 39654
rect 21502 39534 21542 39598
rect 21606 39534 21667 39598
rect 21731 39534 21792 39598
rect 21856 39534 21902 39598
rect 21502 39497 21902 39534
rect 2689 39333 3502 39334
rect 1411 39320 3502 39333
rect 1411 39319 1498 39320
rect 1411 39263 1416 39319
rect 1472 39264 1498 39319
rect 1554 39318 3502 39320
rect 1554 39264 2760 39318
rect 1472 39263 2760 39264
rect 1411 39262 2760 39263
rect 2816 39317 3502 39318
rect 2816 39262 2840 39317
rect 1411 39261 2840 39262
rect 2896 39261 3360 39317
rect 3416 39316 3502 39317
rect 3416 39261 3440 39316
rect 1411 39260 3440 39261
rect 3496 39260 3502 39316
rect 1411 39240 3502 39260
rect 1411 39239 1499 39240
rect 1411 39183 1417 39239
rect 1473 39184 1499 39239
rect 1555 39237 3502 39240
rect 1555 39184 2761 39237
rect 1473 39183 2761 39184
rect 1411 39181 2761 39183
rect 2817 39181 2841 39237
rect 2897 39236 3502 39237
rect 2897 39181 3361 39236
rect 1411 39180 3361 39181
rect 3417 39180 3441 39236
rect 3497 39180 3502 39236
rect 1411 39169 3502 39180
rect 463 39123 805 39139
rect 463 39059 488 39123
rect 552 39059 602 39123
rect 666 39059 716 39123
rect 780 39059 805 39123
rect 463 39043 805 39059
rect 0 38579 342 38595
rect 0 38515 25 38579
rect 89 38515 139 38579
rect 203 38515 253 38579
rect 317 38515 342 38579
rect 0 38499 342 38515
rect 463 38035 805 38051
rect 463 37971 488 38035
rect 552 37971 602 38035
rect 666 37971 716 38035
rect 780 37971 805 38035
rect 463 37955 805 37971
rect 0 37491 342 37507
rect 0 37427 25 37491
rect 89 37427 139 37491
rect 203 37427 253 37491
rect 317 37427 342 37491
rect 0 37411 342 37427
rect 463 36947 805 36963
rect 463 36883 488 36947
rect 552 36883 602 36947
rect 666 36883 716 36947
rect 780 36883 805 36947
rect 463 36867 805 36883
rect 21970 36944 22370 36986
rect 21970 36640 22040 36944
rect 22264 36640 22370 36944
rect 21970 36596 22370 36640
rect 2535 36475 2688 36476
rect 2535 36463 2689 36475
rect 2535 36399 2536 36463
rect 2600 36399 2624 36463
rect 2688 36399 2689 36463
rect 2535 36391 2689 36399
rect 21028 36164 21428 36198
rect 21028 36100 21069 36164
rect 21133 36100 21194 36164
rect 21258 36100 21319 36164
rect 21383 36100 21428 36164
rect 21028 36044 21428 36100
rect 21028 35980 21068 36044
rect 21132 35980 21193 36044
rect 21257 35980 21318 36044
rect 21382 35980 21428 36044
rect 21028 35943 21428 35980
rect 21028 35586 21428 35642
rect 21028 35522 21073 35586
rect 21137 35522 21195 35586
rect 21259 35522 21321 35586
rect 21385 35522 21428 35586
rect 21028 35439 21428 35522
rect 21028 35375 21073 35439
rect 21137 35375 21195 35439
rect 21259 35375 21321 35439
rect 21385 35375 21428 35439
rect 21028 35302 21428 35375
rect 21028 35238 21073 35302
rect 21137 35238 21195 35302
rect 21259 35238 21321 35302
rect 21385 35238 21428 35302
rect 21028 35183 21428 35238
rect 21028 35182 21401 35183
rect 20527 34668 20927 34702
rect 20527 34604 20568 34668
rect 20632 34604 20693 34668
rect 20757 34604 20818 34668
rect 20882 34604 20927 34668
rect 20527 34548 20927 34604
rect 20527 34484 20567 34548
rect 20631 34484 20692 34548
rect 20756 34484 20817 34548
rect 20881 34484 20927 34548
rect 20527 34447 20927 34484
rect 21502 34668 21902 34702
rect 21502 34604 21543 34668
rect 21607 34604 21668 34668
rect 21732 34604 21793 34668
rect 21857 34604 21902 34668
rect 21502 34548 21902 34604
rect 21502 34484 21542 34548
rect 21606 34484 21667 34548
rect 21731 34484 21792 34548
rect 21856 34484 21902 34548
rect 21502 34447 21902 34484
rect 21028 33826 21428 33882
rect 21028 33762 21073 33826
rect 21137 33762 21195 33826
rect 21259 33762 21321 33826
rect 21385 33762 21428 33826
rect 21028 33679 21428 33762
rect 21028 33615 21073 33679
rect 21137 33615 21195 33679
rect 21259 33615 21321 33679
rect 21385 33615 21428 33679
rect 21028 33542 21428 33615
rect 21028 33478 21073 33542
rect 21137 33478 21195 33542
rect 21259 33478 21321 33542
rect 21385 33478 21428 33542
rect 21028 33423 21428 33478
rect 21028 33422 21401 33423
rect 21027 33109 21427 33143
rect 21027 33045 21068 33109
rect 21132 33045 21193 33109
rect 21257 33045 21318 33109
rect 21382 33045 21427 33109
rect 21027 32989 21427 33045
rect 21027 32925 21067 32989
rect 21131 32925 21192 32989
rect 21256 32925 21317 32989
rect 21381 32925 21427 32989
rect 21027 32888 21427 32925
rect 463 32296 866 32360
rect 463 32232 507 32296
rect 571 32232 633 32296
rect 697 32232 753 32296
rect 817 32232 866 32296
rect 463 32178 866 32232
rect 463 32114 507 32178
rect 571 32114 633 32178
rect 697 32114 753 32178
rect 817 32114 866 32178
rect 463 32072 866 32114
rect 21025 32296 21428 32360
rect 21025 32232 21072 32296
rect 21136 32232 21198 32296
rect 21262 32232 21318 32296
rect 21382 32232 21428 32296
rect 21025 32178 21428 32232
rect 21025 32114 21072 32178
rect 21136 32114 21198 32178
rect 21262 32114 21318 32178
rect 21382 32114 21428 32178
rect 21025 32072 21428 32114
rect 463 31514 863 31545
rect 463 31450 507 31514
rect 571 31450 633 31514
rect 697 31450 753 31514
rect 817 31450 863 31514
rect 463 31396 863 31450
rect 463 31332 507 31396
rect 571 31332 633 31396
rect 697 31332 753 31396
rect 817 31332 863 31396
rect 463 31290 863 31332
rect 21028 31514 21428 31545
rect 21028 31450 21072 31514
rect 21136 31450 21198 31514
rect 21262 31450 21318 31514
rect 21382 31450 21428 31514
rect 21028 31396 21428 31450
rect 21028 31332 21072 31396
rect 21136 31332 21198 31396
rect 21262 31332 21318 31396
rect 21382 31332 21428 31396
rect 21028 31290 21428 31332
rect 463 31055 863 31111
rect 463 30991 508 31055
rect 572 30991 630 31055
rect 694 30991 756 31055
rect 820 30991 863 31055
rect 463 30908 863 30991
rect 463 30844 508 30908
rect 572 30844 630 30908
rect 694 30844 756 30908
rect 820 30844 863 30908
rect 463 30771 863 30844
rect 463 30707 508 30771
rect 572 30707 630 30771
rect 694 30707 756 30771
rect 820 30707 863 30771
rect 463 30651 863 30707
rect 21970 30124 22370 30155
rect 21970 30060 22014 30124
rect 22078 30060 22140 30124
rect 22204 30060 22260 30124
rect 22324 30060 22370 30124
rect 21970 30006 22370 30060
rect 21970 29942 22014 30006
rect 22078 29942 22140 30006
rect 22204 29942 22260 30006
rect 22324 29942 22370 30006
rect 21970 29900 22370 29942
rect 463 29288 863 29349
rect 463 29224 508 29288
rect 572 29224 630 29288
rect 694 29224 756 29288
rect 820 29224 863 29288
rect 463 29141 863 29224
rect 463 29077 508 29141
rect 572 29077 630 29141
rect 694 29077 756 29141
rect 820 29077 863 29141
rect 463 29004 863 29077
rect 463 28940 508 29004
rect 572 28940 630 29004
rect 694 28940 756 29004
rect 820 28940 863 29004
rect 463 28890 863 28940
rect 463 28602 863 28633
rect 463 28538 507 28602
rect 571 28538 633 28602
rect 697 28538 753 28602
rect 817 28538 863 28602
rect 463 28484 863 28538
rect 463 28420 507 28484
rect 571 28420 633 28484
rect 697 28420 753 28484
rect 817 28420 863 28484
rect 463 28378 863 28420
rect 21028 28553 21428 28584
rect 21028 28489 21072 28553
rect 21136 28489 21198 28553
rect 21262 28489 21318 28553
rect 21382 28489 21428 28553
rect 21028 28435 21428 28489
rect 21028 28371 21072 28435
rect 21136 28371 21198 28435
rect 21262 28371 21318 28435
rect 21382 28371 21428 28435
rect 21028 28329 21428 28371
rect 463 27598 863 27629
rect 463 27534 507 27598
rect 571 27534 633 27598
rect 697 27534 753 27598
rect 817 27534 863 27598
rect 463 27480 863 27534
rect 463 27416 507 27480
rect 571 27416 633 27480
rect 697 27416 753 27480
rect 817 27416 863 27480
rect 463 27374 863 27416
rect 21027 27436 21427 27467
rect 21027 27372 21072 27436
rect 21136 27372 21198 27436
rect 21262 27372 21318 27436
rect 21382 27372 21427 27436
rect 21027 27318 21427 27372
rect 21027 27254 21072 27318
rect 21136 27254 21198 27318
rect 21262 27254 21318 27318
rect 21382 27254 21427 27318
rect 21027 27212 21427 27254
rect 463 27054 863 27109
rect 463 26990 508 27054
rect 572 26990 630 27054
rect 694 26990 756 27054
rect 820 26990 863 27054
rect 463 26907 863 26990
rect 463 26843 508 26907
rect 572 26843 630 26907
rect 694 26843 756 26907
rect 820 26843 863 26907
rect 463 26770 863 26843
rect 463 26706 508 26770
rect 572 26706 630 26770
rect 694 26706 756 26770
rect 820 26706 863 26770
rect 463 26650 863 26706
rect 21970 25965 22370 25996
rect 21970 25901 22014 25965
rect 22078 25901 22140 25965
rect 22204 25901 22260 25965
rect 22324 25901 22370 25965
rect 21970 25847 22370 25901
rect 21970 25783 22014 25847
rect 22078 25783 22140 25847
rect 22204 25783 22260 25847
rect 22324 25783 22370 25847
rect 21970 25741 22370 25783
rect 463 25294 863 25349
rect 463 25230 508 25294
rect 572 25230 630 25294
rect 694 25230 756 25294
rect 820 25230 863 25294
rect 463 25147 863 25230
rect 463 25083 508 25147
rect 572 25083 630 25147
rect 694 25083 756 25147
rect 820 25083 863 25147
rect 463 25010 863 25083
rect 463 24946 508 25010
rect 572 24946 630 25010
rect 694 24946 756 25010
rect 820 24946 863 25010
rect 463 24890 863 24946
rect 463 24620 864 24651
rect 463 24556 507 24620
rect 571 24556 633 24620
rect 697 24556 753 24620
rect 817 24556 864 24620
rect 463 24502 864 24556
rect 463 24438 507 24502
rect 571 24438 633 24502
rect 697 24438 753 24502
rect 817 24438 864 24502
rect 463 24396 864 24438
rect 21028 24593 21428 24624
rect 21028 24529 21072 24593
rect 21136 24529 21198 24593
rect 21262 24529 21318 24593
rect 21382 24529 21428 24593
rect 21028 24475 21428 24529
rect 21028 24411 21072 24475
rect 21136 24411 21198 24475
rect 21262 24411 21318 24475
rect 21382 24411 21428 24475
rect 21028 24369 21428 24411
rect 463 23538 864 23569
rect 463 23474 507 23538
rect 571 23474 633 23538
rect 697 23474 753 23538
rect 817 23474 864 23538
rect 463 23420 864 23474
rect 463 23356 507 23420
rect 571 23356 633 23420
rect 697 23356 753 23420
rect 817 23356 864 23420
rect 463 23314 864 23356
rect 21028 23418 21428 23449
rect 21028 23354 21072 23418
rect 21136 23354 21198 23418
rect 21262 23354 21318 23418
rect 21382 23354 21428 23418
rect 21028 23300 21428 23354
rect 21028 23236 21072 23300
rect 21136 23236 21198 23300
rect 21262 23236 21318 23300
rect 21382 23236 21428 23300
rect 21028 23194 21428 23236
rect 463 23054 863 23109
rect 463 22990 508 23054
rect 572 22990 630 23054
rect 694 22990 756 23054
rect 820 22990 863 23054
rect 463 22907 863 22990
rect 463 22843 508 22907
rect 572 22843 630 22907
rect 694 22843 756 22907
rect 820 22843 863 22907
rect 463 22770 863 22843
rect 463 22706 508 22770
rect 572 22706 630 22770
rect 694 22706 756 22770
rect 820 22706 863 22770
rect 463 22650 863 22706
rect 21970 22175 22370 22206
rect 21970 22111 22014 22175
rect 22078 22111 22140 22175
rect 22204 22111 22260 22175
rect 22324 22111 22370 22175
rect 21970 22057 22370 22111
rect 21970 21993 22014 22057
rect 22078 21993 22140 22057
rect 22204 21993 22260 22057
rect 22324 21993 22370 22057
rect 21970 21951 22370 21993
rect 463 21295 863 21350
rect 463 21231 508 21295
rect 572 21231 630 21295
rect 694 21231 756 21295
rect 820 21231 863 21295
rect 463 21148 863 21231
rect 463 21084 508 21148
rect 572 21084 630 21148
rect 694 21084 756 21148
rect 820 21084 863 21148
rect 463 21011 863 21084
rect 463 20947 508 21011
rect 572 20947 630 21011
rect 694 20947 756 21011
rect 820 20947 863 21011
rect 463 20891 863 20947
rect 463 20663 864 20694
rect 463 20599 507 20663
rect 571 20599 633 20663
rect 697 20599 753 20663
rect 817 20599 864 20663
rect 463 20545 864 20599
rect 463 20481 507 20545
rect 571 20481 633 20545
rect 697 20481 753 20545
rect 817 20481 864 20545
rect 463 20439 864 20481
rect 21027 20577 21427 20608
rect 21027 20513 21072 20577
rect 21136 20513 21198 20577
rect 21262 20513 21318 20577
rect 21382 20513 21427 20577
rect 21027 20459 21427 20513
rect 21027 20395 21072 20459
rect 21136 20395 21198 20459
rect 21262 20395 21318 20459
rect 21382 20395 21427 20459
rect 21027 20353 21427 20395
rect 463 19562 864 19593
rect 463 19498 507 19562
rect 571 19498 633 19562
rect 697 19498 753 19562
rect 817 19498 864 19562
rect 463 19444 864 19498
rect 463 19380 507 19444
rect 571 19380 633 19444
rect 697 19380 753 19444
rect 817 19380 864 19444
rect 463 19338 864 19380
rect 21027 19406 21427 19437
rect 21027 19342 21072 19406
rect 21136 19342 21198 19406
rect 21262 19342 21318 19406
rect 21382 19342 21427 19406
rect 21027 19288 21427 19342
rect 21027 19224 21072 19288
rect 21136 19224 21198 19288
rect 21262 19224 21318 19288
rect 21382 19224 21427 19288
rect 21027 19182 21427 19224
rect 463 19054 863 19109
rect 463 18990 508 19054
rect 572 18990 630 19054
rect 694 18990 756 19054
rect 820 18990 863 19054
rect 463 18907 863 18990
rect 463 18843 508 18907
rect 572 18843 630 18907
rect 694 18843 756 18907
rect 820 18843 863 18907
rect 463 18770 863 18843
rect 463 18706 508 18770
rect 572 18706 630 18770
rect 694 18706 756 18770
rect 820 18706 863 18770
rect 463 18650 863 18706
rect 21970 18068 22370 18099
rect 21970 18004 22014 18068
rect 22078 18004 22140 18068
rect 22204 18004 22260 18068
rect 22324 18004 22370 18068
rect 21970 17950 22370 18004
rect 21970 17886 22014 17950
rect 22078 17886 22140 17950
rect 22204 17886 22260 17950
rect 22324 17886 22370 17950
rect 21970 17844 22370 17886
rect 463 17294 863 17349
rect 463 17230 508 17294
rect 572 17230 630 17294
rect 694 17230 756 17294
rect 820 17230 863 17294
rect 463 17147 863 17230
rect 463 17083 508 17147
rect 572 17083 630 17147
rect 694 17083 756 17147
rect 820 17083 863 17147
rect 463 17010 863 17083
rect 463 16946 508 17010
rect 572 16946 630 17010
rect 694 16946 756 17010
rect 820 16946 863 17010
rect 463 16890 863 16946
rect 463 16696 865 16727
rect 463 16632 507 16696
rect 571 16632 633 16696
rect 697 16632 753 16696
rect 817 16632 865 16696
rect 463 16578 865 16632
rect 463 16514 507 16578
rect 571 16514 633 16578
rect 697 16514 753 16578
rect 817 16514 865 16578
rect 463 16472 865 16514
rect 21027 16645 21427 16676
rect 21027 16581 21072 16645
rect 21136 16581 21198 16645
rect 21262 16581 21318 16645
rect 21382 16581 21427 16645
rect 21027 16527 21427 16581
rect 21027 16463 21072 16527
rect 21136 16463 21198 16527
rect 21262 16463 21318 16527
rect 21382 16463 21427 16527
rect 21027 16421 21427 16463
rect 463 15480 866 15511
rect 463 15416 507 15480
rect 571 15416 633 15480
rect 697 15416 753 15480
rect 817 15416 866 15480
rect 463 15362 866 15416
rect 463 15298 507 15362
rect 571 15298 633 15362
rect 697 15298 753 15362
rect 817 15298 866 15362
rect 463 15256 866 15298
rect 21027 15431 21427 15462
rect 21027 15367 21072 15431
rect 21136 15367 21198 15431
rect 21262 15367 21318 15431
rect 21382 15367 21427 15431
rect 21027 15313 21427 15367
rect 21027 15249 21072 15313
rect 21136 15249 21198 15313
rect 21262 15249 21318 15313
rect 21382 15249 21427 15313
rect 21027 15207 21427 15249
rect 463 15054 863 15109
rect 463 14990 508 15054
rect 572 14990 630 15054
rect 694 14990 756 15054
rect 820 14990 863 15054
rect 463 14907 863 14990
rect 463 14843 508 14907
rect 572 14843 630 14907
rect 694 14843 756 14907
rect 820 14843 863 14907
rect 463 14770 863 14843
rect 463 14706 508 14770
rect 572 14706 630 14770
rect 694 14706 756 14770
rect 820 14706 863 14770
rect 463 14650 863 14706
rect 21970 14250 22370 14281
rect 21970 14186 22014 14250
rect 22078 14186 22140 14250
rect 22204 14186 22260 14250
rect 22324 14186 22370 14250
rect 21970 14132 22370 14186
rect 21970 14068 22014 14132
rect 22078 14068 22140 14132
rect 22204 14068 22260 14132
rect 22324 14068 22370 14132
rect 21970 14026 22370 14068
rect 463 13294 863 13349
rect 463 13230 508 13294
rect 572 13230 630 13294
rect 694 13230 756 13294
rect 820 13230 863 13294
rect 463 13147 863 13230
rect 463 13083 508 13147
rect 572 13083 630 13147
rect 694 13083 756 13147
rect 820 13083 863 13147
rect 463 13010 863 13083
rect 463 12946 508 13010
rect 572 12946 630 13010
rect 694 12946 756 13010
rect 820 12946 863 13010
rect 463 12890 863 12946
rect 463 12615 864 12646
rect 463 12551 507 12615
rect 571 12551 633 12615
rect 697 12551 753 12615
rect 817 12551 864 12615
rect 463 12497 864 12551
rect 463 12433 507 12497
rect 571 12433 633 12497
rect 697 12433 753 12497
rect 817 12433 864 12497
rect 463 12391 864 12433
rect 21028 12588 21428 12619
rect 21028 12524 21072 12588
rect 21136 12524 21198 12588
rect 21262 12524 21318 12588
rect 21382 12524 21428 12588
rect 21028 12470 21428 12524
rect 21028 12406 21072 12470
rect 21136 12406 21198 12470
rect 21262 12406 21318 12470
rect 21382 12406 21428 12470
rect 21028 12364 21428 12406
rect 463 11493 864 11524
rect 463 11429 507 11493
rect 571 11429 633 11493
rect 697 11429 753 11493
rect 817 11429 864 11493
rect 463 11375 864 11429
rect 463 11311 507 11375
rect 571 11311 633 11375
rect 697 11311 753 11375
rect 817 11311 864 11375
rect 463 11269 864 11311
rect 21027 11431 21427 11462
rect 21027 11367 21072 11431
rect 21136 11367 21198 11431
rect 21262 11367 21318 11431
rect 21382 11367 21427 11431
rect 21027 11313 21427 11367
rect 21027 11249 21072 11313
rect 21136 11249 21198 11313
rect 21262 11249 21318 11313
rect 21382 11249 21427 11313
rect 21027 11207 21427 11249
rect 463 11055 863 11110
rect 463 10991 508 11055
rect 572 10991 630 11055
rect 694 10991 756 11055
rect 820 10991 863 11055
rect 463 10908 863 10991
rect 463 10844 508 10908
rect 572 10844 630 10908
rect 694 10844 756 10908
rect 820 10844 863 10908
rect 463 10771 863 10844
rect 463 10707 508 10771
rect 572 10707 630 10771
rect 694 10707 756 10771
rect 820 10707 863 10771
rect 463 10651 863 10707
rect 21970 10286 22370 10317
rect 21970 10222 22014 10286
rect 22078 10222 22140 10286
rect 22204 10222 22260 10286
rect 22324 10222 22370 10286
rect 21970 10168 22370 10222
rect 21970 10104 22014 10168
rect 22078 10104 22140 10168
rect 22204 10104 22260 10168
rect 22324 10104 22370 10168
rect 21970 10062 22370 10104
rect 463 9293 863 9348
rect 463 9229 508 9293
rect 572 9229 630 9293
rect 694 9229 756 9293
rect 820 9229 863 9293
rect 463 9146 863 9229
rect 463 9082 508 9146
rect 572 9082 630 9146
rect 694 9082 756 9146
rect 820 9082 863 9146
rect 463 9009 863 9082
rect 463 8945 508 9009
rect 572 8945 630 9009
rect 694 8945 756 9009
rect 820 8945 863 9009
rect 463 8889 863 8945
rect 463 8633 863 8664
rect 463 8569 507 8633
rect 571 8569 633 8633
rect 697 8569 753 8633
rect 817 8569 863 8633
rect 463 8515 863 8569
rect 463 8451 507 8515
rect 571 8451 633 8515
rect 697 8451 753 8515
rect 817 8451 863 8515
rect 463 8409 863 8451
rect 21028 8588 21428 8619
rect 21028 8524 21072 8588
rect 21136 8524 21198 8588
rect 21262 8524 21318 8588
rect 21382 8524 21428 8588
rect 21028 8470 21428 8524
rect 21028 8406 21072 8470
rect 21136 8406 21198 8470
rect 21262 8406 21318 8470
rect 21382 8406 21428 8470
rect 21028 8364 21428 8406
rect 463 7522 863 7553
rect 463 7458 507 7522
rect 571 7458 633 7522
rect 697 7458 753 7522
rect 817 7458 863 7522
rect 463 7404 863 7458
rect 463 7340 507 7404
rect 571 7340 633 7404
rect 697 7340 753 7404
rect 817 7340 863 7404
rect 463 7298 863 7340
rect 21027 7431 21427 7462
rect 21027 7367 21072 7431
rect 21136 7367 21198 7431
rect 21262 7367 21318 7431
rect 21382 7367 21427 7431
rect 21027 7313 21427 7367
rect 21027 7249 21072 7313
rect 21136 7249 21198 7313
rect 21262 7249 21318 7313
rect 21382 7249 21427 7313
rect 21027 7207 21427 7249
rect 463 7055 863 7110
rect 463 6991 508 7055
rect 572 6991 630 7055
rect 694 6991 756 7055
rect 820 6991 863 7055
rect 463 6908 863 6991
rect 463 6844 508 6908
rect 572 6844 630 6908
rect 694 6844 756 6908
rect 820 6844 863 6908
rect 463 6771 863 6844
rect 463 6707 508 6771
rect 572 6707 630 6771
rect 694 6707 756 6771
rect 820 6707 863 6771
rect 463 6651 863 6707
rect 21970 6274 22370 6305
rect 21970 6210 22014 6274
rect 22078 6210 22140 6274
rect 22204 6210 22260 6274
rect 22324 6210 22370 6274
rect 21970 6156 22370 6210
rect 21970 6092 22014 6156
rect 22078 6092 22140 6156
rect 22204 6092 22260 6156
rect 22324 6092 22370 6156
rect 21970 6050 22370 6092
rect 463 5294 863 5349
rect 463 5230 508 5294
rect 572 5230 630 5294
rect 694 5230 756 5294
rect 820 5230 863 5294
rect 463 5147 863 5230
rect 463 5083 508 5147
rect 572 5083 630 5147
rect 694 5083 756 5147
rect 820 5083 863 5147
rect 463 5010 863 5083
rect 463 4946 508 5010
rect 572 4946 630 5010
rect 694 4946 756 5010
rect 820 4946 863 5010
rect 463 4890 863 4946
rect 463 4699 865 4730
rect 463 4635 507 4699
rect 571 4635 633 4699
rect 697 4635 753 4699
rect 817 4635 865 4699
rect 463 4581 865 4635
rect 463 4517 507 4581
rect 571 4517 633 4581
rect 697 4517 753 4581
rect 817 4517 865 4581
rect 463 4475 865 4517
rect 21028 4588 21428 4619
rect 21028 4524 21072 4588
rect 21136 4524 21198 4588
rect 21262 4524 21318 4588
rect 21382 4524 21428 4588
rect 21028 4470 21428 4524
rect 21028 4406 21072 4470
rect 21136 4406 21198 4470
rect 21262 4406 21318 4470
rect 21382 4406 21428 4470
rect 21028 4364 21428 4406
rect 463 3522 863 3553
rect 463 3458 507 3522
rect 571 3458 633 3522
rect 697 3458 753 3522
rect 817 3458 863 3522
rect 463 3404 863 3458
rect 463 3340 507 3404
rect 571 3340 633 3404
rect 697 3340 753 3404
rect 817 3340 863 3404
rect 463 3298 863 3340
rect 21027 3431 21427 3462
rect 21027 3367 21072 3431
rect 21136 3367 21198 3431
rect 21262 3367 21318 3431
rect 21382 3367 21427 3431
rect 21027 3313 21427 3367
rect 21027 3249 21072 3313
rect 21136 3249 21198 3313
rect 21262 3249 21318 3313
rect 21382 3249 21427 3313
rect 21027 3207 21427 3249
rect 463 3055 863 3110
rect 463 2991 508 3055
rect 572 2991 630 3055
rect 694 2991 756 3055
rect 820 2991 863 3055
rect 463 2908 863 2991
rect 463 2844 508 2908
rect 572 2844 630 2908
rect 694 2844 756 2908
rect 820 2844 863 2908
rect 463 2771 863 2844
rect 463 2707 508 2771
rect 572 2707 630 2771
rect 694 2707 756 2771
rect 820 2707 863 2771
rect 463 2651 863 2707
rect 21970 2274 22370 2305
rect 21970 2210 22014 2274
rect 22078 2210 22140 2274
rect 22204 2210 22260 2274
rect 22324 2210 22370 2274
rect 21970 2156 22370 2210
rect 21970 2092 22014 2156
rect 22078 2092 22140 2156
rect 22204 2092 22260 2156
rect 22324 2092 22370 2156
rect 21970 2050 22370 2092
rect 463 1294 863 1349
rect 463 1230 508 1294
rect 572 1230 630 1294
rect 694 1230 756 1294
rect 820 1230 863 1294
rect 463 1147 863 1230
rect 463 1083 508 1147
rect 572 1083 630 1147
rect 694 1083 756 1147
rect 820 1083 863 1147
rect 463 1010 863 1083
rect 463 946 508 1010
rect 572 946 630 1010
rect 694 946 756 1010
rect 820 946 863 1010
rect 463 890 863 946
rect 463 699 865 730
rect 463 635 507 699
rect 571 635 633 699
rect 697 635 753 699
rect 817 635 865 699
rect 463 581 865 635
rect 463 517 507 581
rect 571 517 633 581
rect 697 517 753 581
rect 817 517 865 581
rect 463 475 865 517
rect 21028 588 21428 619
rect 21028 524 21072 588
rect 21136 524 21198 588
rect 21262 524 21318 588
rect 21382 524 21428 588
rect 21028 470 21428 524
rect 21028 406 21072 470
rect 21136 406 21198 470
rect 21262 406 21318 470
rect 21382 406 21428 470
rect 21028 364 21428 406
<< via3 >>
rect 507 75442 571 75446
rect 507 75386 511 75442
rect 511 75386 567 75442
rect 567 75386 571 75442
rect 507 75382 571 75386
rect 633 75442 697 75446
rect 633 75386 637 75442
rect 637 75386 693 75442
rect 693 75386 697 75442
rect 633 75382 697 75386
rect 753 75442 817 75446
rect 753 75386 757 75442
rect 757 75386 813 75442
rect 813 75386 817 75442
rect 753 75382 817 75386
rect 507 75324 571 75328
rect 507 75268 511 75324
rect 511 75268 567 75324
rect 567 75268 571 75324
rect 507 75264 571 75268
rect 633 75324 697 75328
rect 633 75268 637 75324
rect 637 75268 693 75324
rect 693 75268 697 75324
rect 633 75264 697 75268
rect 753 75324 817 75328
rect 753 75268 757 75324
rect 757 75268 813 75324
rect 813 75268 817 75324
rect 753 75264 817 75268
rect 21072 75482 21136 75486
rect 21072 75426 21076 75482
rect 21076 75426 21132 75482
rect 21132 75426 21136 75482
rect 21072 75422 21136 75426
rect 21198 75482 21262 75486
rect 21198 75426 21202 75482
rect 21202 75426 21258 75482
rect 21258 75426 21262 75482
rect 21198 75422 21262 75426
rect 21318 75482 21382 75486
rect 21318 75426 21322 75482
rect 21322 75426 21378 75482
rect 21378 75426 21382 75482
rect 21318 75422 21382 75426
rect 21072 75364 21136 75368
rect 21072 75308 21076 75364
rect 21076 75308 21132 75364
rect 21132 75308 21136 75364
rect 21072 75304 21136 75308
rect 21198 75364 21262 75368
rect 21198 75308 21202 75364
rect 21202 75308 21258 75364
rect 21258 75308 21262 75364
rect 21198 75304 21262 75308
rect 21318 75364 21382 75368
rect 21318 75308 21322 75364
rect 21322 75308 21378 75364
rect 21378 75308 21382 75364
rect 21318 75304 21382 75308
rect 508 75050 572 75054
rect 508 74994 512 75050
rect 512 74994 568 75050
rect 568 74994 572 75050
rect 508 74990 572 74994
rect 630 75050 694 75054
rect 630 74994 634 75050
rect 634 74994 690 75050
rect 690 74994 694 75050
rect 630 74990 694 74994
rect 756 75050 820 75054
rect 756 74994 760 75050
rect 760 74994 816 75050
rect 816 74994 820 75050
rect 756 74990 820 74994
rect 508 74903 572 74907
rect 508 74847 512 74903
rect 512 74847 568 74903
rect 568 74847 572 74903
rect 508 74843 572 74847
rect 630 74903 694 74907
rect 630 74847 634 74903
rect 634 74847 690 74903
rect 690 74847 694 74903
rect 630 74843 694 74847
rect 756 74903 820 74907
rect 756 74847 760 74903
rect 760 74847 816 74903
rect 816 74847 820 74903
rect 756 74843 820 74847
rect 508 74766 572 74770
rect 508 74710 512 74766
rect 512 74710 568 74766
rect 568 74710 572 74766
rect 508 74706 572 74710
rect 630 74766 694 74770
rect 630 74710 634 74766
rect 634 74710 690 74766
rect 690 74710 694 74766
rect 630 74706 694 74710
rect 756 74766 820 74770
rect 756 74710 760 74766
rect 760 74710 816 74766
rect 816 74710 820 74766
rect 756 74706 820 74710
rect 22014 74061 22078 74065
rect 22014 74005 22018 74061
rect 22018 74005 22074 74061
rect 22074 74005 22078 74061
rect 22014 74001 22078 74005
rect 22140 74061 22204 74065
rect 22140 74005 22144 74061
rect 22144 74005 22200 74061
rect 22200 74005 22204 74061
rect 22140 74001 22204 74005
rect 22260 74061 22324 74065
rect 22260 74005 22264 74061
rect 22264 74005 22320 74061
rect 22320 74005 22324 74061
rect 22260 74001 22324 74005
rect 22014 73943 22078 73947
rect 22014 73887 22018 73943
rect 22018 73887 22074 73943
rect 22074 73887 22078 73943
rect 22014 73883 22078 73887
rect 22140 73943 22204 73947
rect 22140 73887 22144 73943
rect 22144 73887 22200 73943
rect 22200 73887 22204 73943
rect 22140 73883 22204 73887
rect 22260 73943 22324 73947
rect 22260 73887 22264 73943
rect 22264 73887 22320 73943
rect 22320 73887 22324 73943
rect 22260 73883 22324 73887
rect 508 73290 572 73294
rect 508 73234 512 73290
rect 512 73234 568 73290
rect 568 73234 572 73290
rect 508 73230 572 73234
rect 630 73290 694 73294
rect 630 73234 634 73290
rect 634 73234 690 73290
rect 690 73234 694 73290
rect 630 73230 694 73234
rect 756 73290 820 73294
rect 756 73234 760 73290
rect 760 73234 816 73290
rect 816 73234 820 73290
rect 756 73230 820 73234
rect 508 73143 572 73147
rect 508 73087 512 73143
rect 512 73087 568 73143
rect 568 73087 572 73143
rect 508 73083 572 73087
rect 630 73143 694 73147
rect 630 73087 634 73143
rect 634 73087 690 73143
rect 690 73087 694 73143
rect 630 73083 694 73087
rect 756 73143 820 73147
rect 756 73087 760 73143
rect 760 73087 816 73143
rect 816 73087 820 73143
rect 756 73083 820 73087
rect 508 73006 572 73010
rect 508 72950 512 73006
rect 512 72950 568 73006
rect 568 72950 572 73006
rect 508 72946 572 72950
rect 630 73006 694 73010
rect 630 72950 634 73006
rect 634 72950 690 73006
rect 690 72950 694 73006
rect 630 72946 694 72950
rect 756 73006 820 73010
rect 756 72950 760 73006
rect 760 72950 816 73006
rect 816 72950 820 73006
rect 756 72946 820 72950
rect 507 72769 571 72773
rect 507 72713 511 72769
rect 511 72713 567 72769
rect 567 72713 571 72769
rect 507 72709 571 72713
rect 633 72769 697 72773
rect 633 72713 637 72769
rect 637 72713 693 72769
rect 693 72713 697 72769
rect 633 72709 697 72713
rect 753 72769 817 72773
rect 753 72713 757 72769
rect 757 72713 813 72769
rect 813 72713 817 72769
rect 753 72709 817 72713
rect 507 72651 571 72655
rect 507 72595 511 72651
rect 511 72595 567 72651
rect 567 72595 571 72651
rect 507 72591 571 72595
rect 633 72651 697 72655
rect 633 72595 637 72651
rect 637 72595 693 72651
rect 693 72595 697 72651
rect 633 72591 697 72595
rect 753 72651 817 72655
rect 753 72595 757 72651
rect 757 72595 813 72651
rect 813 72595 817 72651
rect 753 72591 817 72595
rect 21072 72685 21136 72689
rect 21072 72629 21076 72685
rect 21076 72629 21132 72685
rect 21132 72629 21136 72685
rect 21072 72625 21136 72629
rect 21198 72685 21262 72689
rect 21198 72629 21202 72685
rect 21202 72629 21258 72685
rect 21258 72629 21262 72685
rect 21198 72625 21262 72629
rect 21318 72685 21382 72689
rect 21318 72629 21322 72685
rect 21322 72629 21378 72685
rect 21378 72629 21382 72685
rect 21318 72625 21382 72629
rect 21072 72567 21136 72571
rect 21072 72511 21076 72567
rect 21076 72511 21132 72567
rect 21132 72511 21136 72567
rect 21072 72507 21136 72511
rect 21198 72567 21262 72571
rect 21198 72511 21202 72567
rect 21202 72511 21258 72567
rect 21258 72511 21262 72567
rect 21198 72507 21262 72511
rect 21318 72567 21382 72571
rect 21318 72511 21322 72567
rect 21322 72511 21378 72567
rect 21378 72511 21382 72567
rect 21318 72507 21382 72511
rect 507 71442 571 71446
rect 507 71386 511 71442
rect 511 71386 567 71442
rect 567 71386 571 71442
rect 507 71382 571 71386
rect 633 71442 697 71446
rect 633 71386 637 71442
rect 637 71386 693 71442
rect 693 71386 697 71442
rect 633 71382 697 71386
rect 753 71442 817 71446
rect 753 71386 757 71442
rect 757 71386 813 71442
rect 813 71386 817 71442
rect 753 71382 817 71386
rect 507 71324 571 71328
rect 507 71268 511 71324
rect 511 71268 567 71324
rect 567 71268 571 71324
rect 507 71264 571 71268
rect 633 71324 697 71328
rect 633 71268 637 71324
rect 637 71268 693 71324
rect 693 71268 697 71324
rect 633 71264 697 71268
rect 753 71324 817 71328
rect 753 71268 757 71324
rect 757 71268 813 71324
rect 813 71268 817 71324
rect 753 71264 817 71268
rect 21072 71482 21136 71486
rect 21072 71426 21076 71482
rect 21076 71426 21132 71482
rect 21132 71426 21136 71482
rect 21072 71422 21136 71426
rect 21198 71482 21262 71486
rect 21198 71426 21202 71482
rect 21202 71426 21258 71482
rect 21258 71426 21262 71482
rect 21198 71422 21262 71426
rect 21318 71482 21382 71486
rect 21318 71426 21322 71482
rect 21322 71426 21378 71482
rect 21378 71426 21382 71482
rect 21318 71422 21382 71426
rect 21072 71364 21136 71368
rect 21072 71308 21076 71364
rect 21076 71308 21132 71364
rect 21132 71308 21136 71364
rect 21072 71304 21136 71308
rect 21198 71364 21262 71368
rect 21198 71308 21202 71364
rect 21202 71308 21258 71364
rect 21258 71308 21262 71364
rect 21198 71304 21262 71308
rect 21318 71364 21382 71368
rect 21318 71308 21322 71364
rect 21322 71308 21378 71364
rect 21378 71308 21382 71364
rect 21318 71304 21382 71308
rect 508 71050 572 71054
rect 508 70994 512 71050
rect 512 70994 568 71050
rect 568 70994 572 71050
rect 508 70990 572 70994
rect 630 71050 694 71054
rect 630 70994 634 71050
rect 634 70994 690 71050
rect 690 70994 694 71050
rect 630 70990 694 70994
rect 756 71050 820 71054
rect 756 70994 760 71050
rect 760 70994 816 71050
rect 816 70994 820 71050
rect 756 70990 820 70994
rect 508 70903 572 70907
rect 508 70847 512 70903
rect 512 70847 568 70903
rect 568 70847 572 70903
rect 508 70843 572 70847
rect 630 70903 694 70907
rect 630 70847 634 70903
rect 634 70847 690 70903
rect 690 70847 694 70903
rect 630 70843 694 70847
rect 756 70903 820 70907
rect 756 70847 760 70903
rect 760 70847 816 70903
rect 816 70847 820 70903
rect 756 70843 820 70847
rect 508 70766 572 70770
rect 508 70710 512 70766
rect 512 70710 568 70766
rect 568 70710 572 70766
rect 508 70706 572 70710
rect 630 70766 694 70770
rect 630 70710 634 70766
rect 634 70710 690 70766
rect 690 70710 694 70766
rect 630 70706 694 70710
rect 756 70766 820 70770
rect 756 70710 760 70766
rect 760 70710 816 70766
rect 816 70710 820 70766
rect 756 70706 820 70710
rect 22014 70061 22078 70065
rect 22014 70005 22018 70061
rect 22018 70005 22074 70061
rect 22074 70005 22078 70061
rect 22014 70001 22078 70005
rect 22140 70061 22204 70065
rect 22140 70005 22144 70061
rect 22144 70005 22200 70061
rect 22200 70005 22204 70061
rect 22140 70001 22204 70005
rect 22260 70061 22324 70065
rect 22260 70005 22264 70061
rect 22264 70005 22320 70061
rect 22320 70005 22324 70061
rect 22260 70001 22324 70005
rect 22014 69943 22078 69947
rect 22014 69887 22018 69943
rect 22018 69887 22074 69943
rect 22074 69887 22078 69943
rect 22014 69883 22078 69887
rect 22140 69943 22204 69947
rect 22140 69887 22144 69943
rect 22144 69887 22200 69943
rect 22200 69887 22204 69943
rect 22140 69883 22204 69887
rect 22260 69943 22324 69947
rect 22260 69887 22264 69943
rect 22264 69887 22320 69943
rect 22320 69887 22324 69943
rect 22260 69883 22324 69887
rect 508 69290 572 69294
rect 508 69234 512 69290
rect 512 69234 568 69290
rect 568 69234 572 69290
rect 508 69230 572 69234
rect 630 69290 694 69294
rect 630 69234 634 69290
rect 634 69234 690 69290
rect 690 69234 694 69290
rect 630 69230 694 69234
rect 756 69290 820 69294
rect 756 69234 760 69290
rect 760 69234 816 69290
rect 816 69234 820 69290
rect 756 69230 820 69234
rect 508 69143 572 69147
rect 508 69087 512 69143
rect 512 69087 568 69143
rect 568 69087 572 69143
rect 508 69083 572 69087
rect 630 69143 694 69147
rect 630 69087 634 69143
rect 634 69087 690 69143
rect 690 69087 694 69143
rect 630 69083 694 69087
rect 756 69143 820 69147
rect 756 69087 760 69143
rect 760 69087 816 69143
rect 816 69087 820 69143
rect 756 69083 820 69087
rect 508 69006 572 69010
rect 508 68950 512 69006
rect 512 68950 568 69006
rect 568 68950 572 69006
rect 508 68946 572 68950
rect 630 69006 694 69010
rect 630 68950 634 69006
rect 634 68950 690 69006
rect 690 68950 694 69006
rect 630 68946 694 68950
rect 756 69006 820 69010
rect 756 68950 760 69006
rect 760 68950 816 69006
rect 816 68950 820 69006
rect 756 68946 820 68950
rect 507 68769 571 68773
rect 507 68713 511 68769
rect 511 68713 567 68769
rect 567 68713 571 68769
rect 507 68709 571 68713
rect 633 68769 697 68773
rect 633 68713 637 68769
rect 637 68713 693 68769
rect 693 68713 697 68769
rect 633 68709 697 68713
rect 753 68769 817 68773
rect 753 68713 757 68769
rect 757 68713 813 68769
rect 813 68713 817 68769
rect 753 68709 817 68713
rect 507 68651 571 68655
rect 507 68595 511 68651
rect 511 68595 567 68651
rect 567 68595 571 68651
rect 507 68591 571 68595
rect 633 68651 697 68655
rect 633 68595 637 68651
rect 637 68595 693 68651
rect 693 68595 697 68651
rect 633 68591 697 68595
rect 753 68651 817 68655
rect 753 68595 757 68651
rect 757 68595 813 68651
rect 813 68595 817 68651
rect 753 68591 817 68595
rect 21072 68685 21136 68689
rect 21072 68629 21076 68685
rect 21076 68629 21132 68685
rect 21132 68629 21136 68685
rect 21072 68625 21136 68629
rect 21198 68685 21262 68689
rect 21198 68629 21202 68685
rect 21202 68629 21258 68685
rect 21258 68629 21262 68685
rect 21198 68625 21262 68629
rect 21318 68685 21382 68689
rect 21318 68629 21322 68685
rect 21322 68629 21378 68685
rect 21378 68629 21382 68685
rect 21318 68625 21382 68629
rect 21072 68567 21136 68571
rect 21072 68511 21076 68567
rect 21076 68511 21132 68567
rect 21132 68511 21136 68567
rect 21072 68507 21136 68511
rect 21198 68567 21262 68571
rect 21198 68511 21202 68567
rect 21202 68511 21258 68567
rect 21258 68511 21262 68567
rect 21198 68507 21262 68511
rect 21318 68567 21382 68571
rect 21318 68511 21322 68567
rect 21322 68511 21378 68567
rect 21378 68511 21382 68567
rect 21318 68507 21382 68511
rect 507 67440 571 67444
rect 507 67384 511 67440
rect 511 67384 567 67440
rect 567 67384 571 67440
rect 507 67380 571 67384
rect 633 67440 697 67444
rect 633 67384 637 67440
rect 637 67384 693 67440
rect 693 67384 697 67440
rect 633 67380 697 67384
rect 753 67440 817 67444
rect 753 67384 757 67440
rect 757 67384 813 67440
rect 813 67384 817 67440
rect 753 67380 817 67384
rect 507 67322 571 67326
rect 507 67266 511 67322
rect 511 67266 567 67322
rect 567 67266 571 67322
rect 507 67262 571 67266
rect 633 67322 697 67326
rect 633 67266 637 67322
rect 637 67266 693 67322
rect 693 67266 697 67322
rect 633 67262 697 67266
rect 753 67322 817 67326
rect 753 67266 757 67322
rect 757 67266 813 67322
rect 813 67266 817 67322
rect 753 67262 817 67266
rect 21072 67482 21136 67486
rect 21072 67426 21076 67482
rect 21076 67426 21132 67482
rect 21132 67426 21136 67482
rect 21072 67422 21136 67426
rect 21198 67482 21262 67486
rect 21198 67426 21202 67482
rect 21202 67426 21258 67482
rect 21258 67426 21262 67482
rect 21198 67422 21262 67426
rect 21318 67482 21382 67486
rect 21318 67426 21322 67482
rect 21322 67426 21378 67482
rect 21378 67426 21382 67482
rect 21318 67422 21382 67426
rect 21072 67364 21136 67368
rect 21072 67308 21076 67364
rect 21076 67308 21132 67364
rect 21132 67308 21136 67364
rect 21072 67304 21136 67308
rect 21198 67364 21262 67368
rect 21198 67308 21202 67364
rect 21202 67308 21258 67364
rect 21258 67308 21262 67364
rect 21198 67304 21262 67308
rect 21318 67364 21382 67368
rect 21318 67308 21322 67364
rect 21322 67308 21378 67364
rect 21378 67308 21382 67364
rect 21318 67304 21382 67308
rect 508 67050 572 67054
rect 508 66994 512 67050
rect 512 66994 568 67050
rect 568 66994 572 67050
rect 508 66990 572 66994
rect 630 67050 694 67054
rect 630 66994 634 67050
rect 634 66994 690 67050
rect 690 66994 694 67050
rect 630 66990 694 66994
rect 756 67050 820 67054
rect 756 66994 760 67050
rect 760 66994 816 67050
rect 816 66994 820 67050
rect 756 66990 820 66994
rect 508 66903 572 66907
rect 508 66847 512 66903
rect 512 66847 568 66903
rect 568 66847 572 66903
rect 508 66843 572 66847
rect 630 66903 694 66907
rect 630 66847 634 66903
rect 634 66847 690 66903
rect 690 66847 694 66903
rect 630 66843 694 66847
rect 756 66903 820 66907
rect 756 66847 760 66903
rect 760 66847 816 66903
rect 816 66847 820 66903
rect 756 66843 820 66847
rect 508 66766 572 66770
rect 508 66710 512 66766
rect 512 66710 568 66766
rect 568 66710 572 66766
rect 508 66706 572 66710
rect 630 66766 694 66770
rect 630 66710 634 66766
rect 634 66710 690 66766
rect 690 66710 694 66766
rect 630 66706 694 66710
rect 756 66766 820 66770
rect 756 66710 760 66766
rect 760 66710 816 66766
rect 816 66710 820 66766
rect 756 66706 820 66710
rect 22014 66048 22078 66052
rect 22014 65992 22018 66048
rect 22018 65992 22074 66048
rect 22074 65992 22078 66048
rect 22014 65988 22078 65992
rect 22140 66048 22204 66052
rect 22140 65992 22144 66048
rect 22144 65992 22200 66048
rect 22200 65992 22204 66048
rect 22140 65988 22204 65992
rect 22260 66048 22324 66052
rect 22260 65992 22264 66048
rect 22264 65992 22320 66048
rect 22320 65992 22324 66048
rect 22260 65988 22324 65992
rect 22014 65930 22078 65934
rect 22014 65874 22018 65930
rect 22018 65874 22074 65930
rect 22074 65874 22078 65930
rect 22014 65870 22078 65874
rect 22140 65930 22204 65934
rect 22140 65874 22144 65930
rect 22144 65874 22200 65930
rect 22200 65874 22204 65930
rect 22140 65870 22204 65874
rect 22260 65930 22324 65934
rect 22260 65874 22264 65930
rect 22264 65874 22320 65930
rect 22320 65874 22324 65930
rect 22260 65870 22324 65874
rect 508 65291 572 65295
rect 508 65235 512 65291
rect 512 65235 568 65291
rect 568 65235 572 65291
rect 508 65231 572 65235
rect 630 65291 694 65295
rect 630 65235 634 65291
rect 634 65235 690 65291
rect 690 65235 694 65291
rect 630 65231 694 65235
rect 756 65291 820 65295
rect 756 65235 760 65291
rect 760 65235 816 65291
rect 816 65235 820 65291
rect 756 65231 820 65235
rect 508 65144 572 65148
rect 508 65088 512 65144
rect 512 65088 568 65144
rect 568 65088 572 65144
rect 508 65084 572 65088
rect 630 65144 694 65148
rect 630 65088 634 65144
rect 634 65088 690 65144
rect 690 65088 694 65144
rect 630 65084 694 65088
rect 756 65144 820 65148
rect 756 65088 760 65144
rect 760 65088 816 65144
rect 816 65088 820 65144
rect 756 65084 820 65088
rect 508 65007 572 65011
rect 508 64951 512 65007
rect 512 64951 568 65007
rect 568 64951 572 65007
rect 508 64947 572 64951
rect 630 65007 694 65011
rect 630 64951 634 65007
rect 634 64951 690 65007
rect 690 64951 694 65007
rect 630 64947 694 64951
rect 756 65007 820 65011
rect 756 64951 760 65007
rect 760 64951 816 65007
rect 816 64951 820 65007
rect 756 64947 820 64951
rect 507 64700 571 64704
rect 507 64644 511 64700
rect 511 64644 567 64700
rect 567 64644 571 64700
rect 507 64640 571 64644
rect 633 64700 697 64704
rect 633 64644 637 64700
rect 637 64644 693 64700
rect 693 64644 697 64700
rect 633 64640 697 64644
rect 753 64700 817 64704
rect 753 64644 757 64700
rect 757 64644 813 64700
rect 813 64644 817 64700
rect 753 64640 817 64644
rect 507 64582 571 64586
rect 507 64526 511 64582
rect 511 64526 567 64582
rect 567 64526 571 64582
rect 507 64522 571 64526
rect 633 64582 697 64586
rect 633 64526 637 64582
rect 637 64526 693 64582
rect 693 64526 697 64582
rect 633 64522 697 64526
rect 753 64582 817 64586
rect 753 64526 757 64582
rect 757 64526 813 64582
rect 813 64526 817 64582
rect 753 64522 817 64526
rect 21072 64685 21136 64689
rect 21072 64629 21076 64685
rect 21076 64629 21132 64685
rect 21132 64629 21136 64685
rect 21072 64625 21136 64629
rect 21198 64685 21262 64689
rect 21198 64629 21202 64685
rect 21202 64629 21258 64685
rect 21258 64629 21262 64685
rect 21198 64625 21262 64629
rect 21318 64685 21382 64689
rect 21318 64629 21322 64685
rect 21322 64629 21378 64685
rect 21378 64629 21382 64685
rect 21318 64625 21382 64629
rect 21072 64567 21136 64571
rect 21072 64511 21076 64567
rect 21076 64511 21132 64567
rect 21132 64511 21136 64567
rect 21072 64507 21136 64511
rect 21198 64567 21262 64571
rect 21198 64511 21202 64567
rect 21202 64511 21258 64567
rect 21258 64511 21262 64567
rect 21198 64507 21262 64511
rect 21318 64567 21382 64571
rect 21318 64511 21322 64567
rect 21322 64511 21378 64567
rect 21378 64511 21382 64567
rect 21318 64507 21382 64511
rect 507 63522 571 63526
rect 507 63466 511 63522
rect 511 63466 567 63522
rect 567 63466 571 63522
rect 507 63462 571 63466
rect 633 63522 697 63526
rect 633 63466 637 63522
rect 637 63466 693 63522
rect 693 63466 697 63522
rect 633 63462 697 63466
rect 753 63522 817 63526
rect 753 63466 757 63522
rect 757 63466 813 63522
rect 813 63466 817 63522
rect 753 63462 817 63466
rect 507 63404 571 63408
rect 507 63348 511 63404
rect 511 63348 567 63404
rect 567 63348 571 63404
rect 507 63344 571 63348
rect 633 63404 697 63408
rect 633 63348 637 63404
rect 637 63348 693 63404
rect 693 63348 697 63404
rect 633 63344 697 63348
rect 753 63404 817 63408
rect 753 63348 757 63404
rect 757 63348 813 63404
rect 813 63348 817 63404
rect 753 63344 817 63348
rect 21072 63482 21136 63486
rect 21072 63426 21076 63482
rect 21076 63426 21132 63482
rect 21132 63426 21136 63482
rect 21072 63422 21136 63426
rect 21198 63482 21262 63486
rect 21198 63426 21202 63482
rect 21202 63426 21258 63482
rect 21258 63426 21262 63482
rect 21198 63422 21262 63426
rect 21318 63482 21382 63486
rect 21318 63426 21322 63482
rect 21322 63426 21378 63482
rect 21378 63426 21382 63482
rect 21318 63422 21382 63426
rect 21072 63364 21136 63368
rect 21072 63308 21076 63364
rect 21076 63308 21132 63364
rect 21132 63308 21136 63364
rect 21072 63304 21136 63308
rect 21198 63364 21262 63368
rect 21198 63308 21202 63364
rect 21202 63308 21258 63364
rect 21258 63308 21262 63364
rect 21198 63304 21262 63308
rect 21318 63364 21382 63368
rect 21318 63308 21322 63364
rect 21322 63308 21378 63364
rect 21378 63308 21382 63364
rect 21318 63304 21382 63308
rect 508 63050 572 63054
rect 508 62994 512 63050
rect 512 62994 568 63050
rect 568 62994 572 63050
rect 508 62990 572 62994
rect 630 63050 694 63054
rect 630 62994 634 63050
rect 634 62994 690 63050
rect 690 62994 694 63050
rect 630 62990 694 62994
rect 756 63050 820 63054
rect 756 62994 760 63050
rect 760 62994 816 63050
rect 816 62994 820 63050
rect 756 62990 820 62994
rect 508 62903 572 62907
rect 508 62847 512 62903
rect 512 62847 568 62903
rect 568 62847 572 62903
rect 508 62843 572 62847
rect 630 62903 694 62907
rect 630 62847 634 62903
rect 634 62847 690 62903
rect 690 62847 694 62903
rect 630 62843 694 62847
rect 756 62903 820 62907
rect 756 62847 760 62903
rect 760 62847 816 62903
rect 816 62847 820 62903
rect 756 62843 820 62847
rect 508 62766 572 62770
rect 508 62710 512 62766
rect 512 62710 568 62766
rect 568 62710 572 62766
rect 508 62706 572 62710
rect 630 62766 694 62770
rect 630 62710 634 62766
rect 634 62710 690 62766
rect 690 62710 694 62766
rect 630 62706 694 62710
rect 756 62766 820 62770
rect 756 62710 760 62766
rect 760 62710 816 62766
rect 816 62710 820 62766
rect 756 62706 820 62710
rect 22014 62047 22078 62051
rect 22014 61991 22018 62047
rect 22018 61991 22074 62047
rect 22074 61991 22078 62047
rect 22014 61987 22078 61991
rect 22140 62047 22204 62051
rect 22140 61991 22144 62047
rect 22144 61991 22200 62047
rect 22200 61991 22204 62047
rect 22140 61987 22204 61991
rect 22260 62047 22324 62051
rect 22260 61991 22264 62047
rect 22264 61991 22320 62047
rect 22320 61991 22324 62047
rect 22260 61987 22324 61991
rect 22014 61929 22078 61933
rect 22014 61873 22018 61929
rect 22018 61873 22074 61929
rect 22074 61873 22078 61929
rect 22014 61869 22078 61873
rect 22140 61929 22204 61933
rect 22140 61873 22144 61929
rect 22144 61873 22200 61929
rect 22200 61873 22204 61929
rect 22140 61869 22204 61873
rect 22260 61929 22324 61933
rect 22260 61873 22264 61929
rect 22264 61873 22320 61929
rect 22320 61873 22324 61929
rect 22260 61869 22324 61873
rect 508 61291 572 61295
rect 508 61235 512 61291
rect 512 61235 568 61291
rect 568 61235 572 61291
rect 508 61231 572 61235
rect 630 61291 694 61295
rect 630 61235 634 61291
rect 634 61235 690 61291
rect 690 61235 694 61291
rect 630 61231 694 61235
rect 756 61291 820 61295
rect 756 61235 760 61291
rect 760 61235 816 61291
rect 816 61235 820 61291
rect 756 61231 820 61235
rect 508 61144 572 61148
rect 508 61088 512 61144
rect 512 61088 568 61144
rect 568 61088 572 61144
rect 508 61084 572 61088
rect 630 61144 694 61148
rect 630 61088 634 61144
rect 634 61088 690 61144
rect 690 61088 694 61144
rect 630 61084 694 61088
rect 756 61144 820 61148
rect 756 61088 760 61144
rect 760 61088 816 61144
rect 816 61088 820 61144
rect 756 61084 820 61088
rect 508 61007 572 61011
rect 508 60951 512 61007
rect 512 60951 568 61007
rect 568 60951 572 61007
rect 508 60947 572 60951
rect 630 61007 694 61011
rect 630 60951 634 61007
rect 634 60951 690 61007
rect 690 60951 694 61007
rect 630 60947 694 60951
rect 756 61007 820 61011
rect 756 60951 760 61007
rect 760 60951 816 61007
rect 816 60951 820 61007
rect 756 60947 820 60951
rect 507 60674 571 60678
rect 507 60618 511 60674
rect 511 60618 567 60674
rect 567 60618 571 60674
rect 507 60614 571 60618
rect 633 60674 697 60678
rect 633 60618 637 60674
rect 637 60618 693 60674
rect 693 60618 697 60674
rect 633 60614 697 60618
rect 753 60674 817 60678
rect 753 60618 757 60674
rect 757 60618 813 60674
rect 813 60618 817 60674
rect 753 60614 817 60618
rect 507 60556 571 60560
rect 507 60500 511 60556
rect 511 60500 567 60556
rect 567 60500 571 60556
rect 507 60496 571 60500
rect 633 60556 697 60560
rect 633 60500 637 60556
rect 637 60500 693 60556
rect 693 60500 697 60556
rect 633 60496 697 60500
rect 753 60556 817 60560
rect 753 60500 757 60556
rect 757 60500 813 60556
rect 813 60500 817 60556
rect 753 60496 817 60500
rect 21072 60685 21136 60689
rect 21072 60629 21076 60685
rect 21076 60629 21132 60685
rect 21132 60629 21136 60685
rect 21072 60625 21136 60629
rect 21198 60685 21262 60689
rect 21198 60629 21202 60685
rect 21202 60629 21258 60685
rect 21258 60629 21262 60685
rect 21198 60625 21262 60629
rect 21318 60685 21382 60689
rect 21318 60629 21322 60685
rect 21322 60629 21378 60685
rect 21378 60629 21382 60685
rect 21318 60625 21382 60629
rect 21072 60567 21136 60571
rect 21072 60511 21076 60567
rect 21076 60511 21132 60567
rect 21132 60511 21136 60567
rect 21072 60507 21136 60511
rect 21198 60567 21262 60571
rect 21198 60511 21202 60567
rect 21202 60511 21258 60567
rect 21258 60511 21262 60567
rect 21198 60507 21262 60511
rect 21318 60567 21382 60571
rect 21318 60511 21322 60567
rect 21322 60511 21378 60567
rect 21378 60511 21382 60567
rect 21318 60507 21382 60511
rect 507 59471 571 59475
rect 507 59415 511 59471
rect 511 59415 567 59471
rect 567 59415 571 59471
rect 507 59411 571 59415
rect 633 59471 697 59475
rect 633 59415 637 59471
rect 637 59415 693 59471
rect 693 59415 697 59471
rect 633 59411 697 59415
rect 753 59471 817 59475
rect 753 59415 757 59471
rect 757 59415 813 59471
rect 813 59415 817 59471
rect 753 59411 817 59415
rect 507 59353 571 59357
rect 507 59297 511 59353
rect 511 59297 567 59353
rect 567 59297 571 59353
rect 507 59293 571 59297
rect 633 59353 697 59357
rect 633 59297 637 59353
rect 637 59297 693 59353
rect 693 59297 697 59353
rect 633 59293 697 59297
rect 753 59353 817 59357
rect 753 59297 757 59353
rect 757 59297 813 59353
rect 813 59297 817 59353
rect 753 59293 817 59297
rect 21072 59536 21136 59540
rect 21072 59480 21076 59536
rect 21076 59480 21132 59536
rect 21132 59480 21136 59536
rect 21072 59476 21136 59480
rect 21198 59536 21262 59540
rect 21198 59480 21202 59536
rect 21202 59480 21258 59536
rect 21258 59480 21262 59536
rect 21198 59476 21262 59480
rect 21318 59536 21382 59540
rect 21318 59480 21322 59536
rect 21322 59480 21378 59536
rect 21378 59480 21382 59536
rect 21318 59476 21382 59480
rect 21072 59418 21136 59422
rect 21072 59362 21076 59418
rect 21076 59362 21132 59418
rect 21132 59362 21136 59418
rect 21072 59358 21136 59362
rect 21198 59418 21262 59422
rect 21198 59362 21202 59418
rect 21202 59362 21258 59418
rect 21258 59362 21262 59418
rect 21198 59358 21262 59362
rect 21318 59418 21382 59422
rect 21318 59362 21322 59418
rect 21322 59362 21378 59418
rect 21378 59362 21382 59418
rect 21318 59358 21382 59362
rect 508 59050 572 59054
rect 508 58994 512 59050
rect 512 58994 568 59050
rect 568 58994 572 59050
rect 508 58990 572 58994
rect 630 59050 694 59054
rect 630 58994 634 59050
rect 634 58994 690 59050
rect 690 58994 694 59050
rect 630 58990 694 58994
rect 756 59050 820 59054
rect 756 58994 760 59050
rect 760 58994 816 59050
rect 816 58994 820 59050
rect 756 58990 820 58994
rect 508 58903 572 58907
rect 508 58847 512 58903
rect 512 58847 568 58903
rect 568 58847 572 58903
rect 508 58843 572 58847
rect 630 58903 694 58907
rect 630 58847 634 58903
rect 634 58847 690 58903
rect 690 58847 694 58903
rect 630 58843 694 58847
rect 756 58903 820 58907
rect 756 58847 760 58903
rect 760 58847 816 58903
rect 816 58847 820 58903
rect 756 58843 820 58847
rect 508 58766 572 58770
rect 508 58710 512 58766
rect 512 58710 568 58766
rect 568 58710 572 58766
rect 508 58706 572 58710
rect 630 58766 694 58770
rect 630 58710 634 58766
rect 634 58710 690 58766
rect 690 58710 694 58766
rect 630 58706 694 58710
rect 756 58766 820 58770
rect 756 58710 760 58766
rect 760 58710 816 58766
rect 816 58710 820 58766
rect 756 58706 820 58710
rect 22014 58086 22078 58090
rect 22014 58030 22018 58086
rect 22018 58030 22074 58086
rect 22074 58030 22078 58086
rect 22014 58026 22078 58030
rect 22140 58086 22204 58090
rect 22140 58030 22144 58086
rect 22144 58030 22200 58086
rect 22200 58030 22204 58086
rect 22140 58026 22204 58030
rect 22260 58086 22324 58090
rect 22260 58030 22264 58086
rect 22264 58030 22320 58086
rect 22320 58030 22324 58086
rect 22260 58026 22324 58030
rect 22014 57968 22078 57972
rect 22014 57912 22018 57968
rect 22018 57912 22074 57968
rect 22074 57912 22078 57968
rect 22014 57908 22078 57912
rect 22140 57968 22204 57972
rect 22140 57912 22144 57968
rect 22144 57912 22200 57968
rect 22200 57912 22204 57968
rect 22140 57908 22204 57912
rect 22260 57968 22324 57972
rect 22260 57912 22264 57968
rect 22264 57912 22320 57968
rect 22320 57912 22324 57968
rect 22260 57908 22324 57912
rect 508 57289 572 57293
rect 508 57233 512 57289
rect 512 57233 568 57289
rect 568 57233 572 57289
rect 508 57229 572 57233
rect 630 57289 694 57293
rect 630 57233 634 57289
rect 634 57233 690 57289
rect 690 57233 694 57289
rect 630 57229 694 57233
rect 756 57289 820 57293
rect 756 57233 760 57289
rect 760 57233 816 57289
rect 816 57233 820 57289
rect 756 57229 820 57233
rect 508 57142 572 57146
rect 508 57086 512 57142
rect 512 57086 568 57142
rect 568 57086 572 57142
rect 508 57082 572 57086
rect 630 57142 694 57146
rect 630 57086 634 57142
rect 634 57086 690 57142
rect 690 57086 694 57142
rect 630 57082 694 57086
rect 756 57142 820 57146
rect 756 57086 760 57142
rect 760 57086 816 57142
rect 816 57086 820 57142
rect 756 57082 820 57086
rect 508 57005 572 57009
rect 508 56949 512 57005
rect 512 56949 568 57005
rect 568 56949 572 57005
rect 508 56945 572 56949
rect 630 57005 694 57009
rect 630 56949 634 57005
rect 634 56949 690 57005
rect 690 56949 694 57005
rect 630 56945 694 56949
rect 756 57005 820 57009
rect 756 56949 760 57005
rect 760 56949 816 57005
rect 816 56949 820 57005
rect 756 56945 820 56949
rect 507 56694 571 56698
rect 507 56638 511 56694
rect 511 56638 567 56694
rect 567 56638 571 56694
rect 507 56634 571 56638
rect 633 56694 697 56698
rect 633 56638 637 56694
rect 637 56638 693 56694
rect 693 56638 697 56694
rect 633 56634 697 56638
rect 753 56694 817 56698
rect 753 56638 757 56694
rect 757 56638 813 56694
rect 813 56638 817 56694
rect 753 56634 817 56638
rect 507 56576 571 56580
rect 507 56520 511 56576
rect 511 56520 567 56576
rect 567 56520 571 56576
rect 507 56516 571 56520
rect 633 56576 697 56580
rect 633 56520 637 56576
rect 637 56520 693 56576
rect 693 56520 697 56576
rect 633 56516 697 56520
rect 753 56576 817 56580
rect 753 56520 757 56576
rect 757 56520 813 56576
rect 813 56520 817 56576
rect 753 56516 817 56520
rect 21072 56620 21136 56624
rect 21072 56564 21076 56620
rect 21076 56564 21132 56620
rect 21132 56564 21136 56620
rect 21072 56560 21136 56564
rect 21198 56620 21262 56624
rect 21198 56564 21202 56620
rect 21202 56564 21258 56620
rect 21258 56564 21262 56620
rect 21198 56560 21262 56564
rect 21318 56620 21382 56624
rect 21318 56564 21322 56620
rect 21322 56564 21378 56620
rect 21378 56564 21382 56620
rect 21318 56560 21382 56564
rect 21072 56502 21136 56506
rect 21072 56446 21076 56502
rect 21076 56446 21132 56502
rect 21132 56446 21136 56502
rect 21072 56442 21136 56446
rect 21198 56502 21262 56506
rect 21198 56446 21202 56502
rect 21202 56446 21258 56502
rect 21258 56446 21262 56502
rect 21198 56442 21262 56446
rect 21318 56502 21382 56506
rect 21318 56446 21322 56502
rect 21322 56446 21378 56502
rect 21378 56446 21382 56502
rect 21318 56442 21382 56446
rect 507 55487 571 55491
rect 507 55431 511 55487
rect 511 55431 567 55487
rect 567 55431 571 55487
rect 507 55427 571 55431
rect 633 55487 697 55491
rect 633 55431 637 55487
rect 637 55431 693 55487
rect 693 55431 697 55487
rect 633 55427 697 55431
rect 753 55487 817 55491
rect 753 55431 757 55487
rect 757 55431 813 55487
rect 813 55431 817 55487
rect 753 55427 817 55431
rect 507 55369 571 55373
rect 507 55313 511 55369
rect 511 55313 567 55369
rect 567 55313 571 55369
rect 507 55309 571 55313
rect 633 55369 697 55373
rect 633 55313 637 55369
rect 637 55313 693 55369
rect 693 55313 697 55369
rect 633 55309 697 55313
rect 753 55369 817 55373
rect 753 55313 757 55369
rect 757 55313 813 55369
rect 813 55313 817 55369
rect 753 55309 817 55313
rect 21072 55437 21136 55441
rect 21072 55381 21076 55437
rect 21076 55381 21132 55437
rect 21132 55381 21136 55437
rect 21072 55377 21136 55381
rect 21198 55437 21262 55441
rect 21198 55381 21202 55437
rect 21202 55381 21258 55437
rect 21258 55381 21262 55437
rect 21198 55377 21262 55381
rect 21318 55437 21382 55441
rect 21318 55381 21322 55437
rect 21322 55381 21378 55437
rect 21378 55381 21382 55437
rect 21318 55377 21382 55381
rect 21072 55319 21136 55323
rect 21072 55263 21076 55319
rect 21076 55263 21132 55319
rect 21132 55263 21136 55319
rect 21072 55259 21136 55263
rect 21198 55319 21262 55323
rect 21198 55263 21202 55319
rect 21202 55263 21258 55319
rect 21258 55263 21262 55319
rect 21198 55259 21262 55263
rect 21318 55319 21382 55323
rect 21318 55263 21322 55319
rect 21322 55263 21378 55319
rect 21378 55263 21382 55319
rect 21318 55259 21382 55263
rect 508 55050 572 55054
rect 508 54994 512 55050
rect 512 54994 568 55050
rect 568 54994 572 55050
rect 508 54990 572 54994
rect 630 55050 694 55054
rect 630 54994 634 55050
rect 634 54994 690 55050
rect 690 54994 694 55050
rect 630 54990 694 54994
rect 756 55050 820 55054
rect 756 54994 760 55050
rect 760 54994 816 55050
rect 816 54994 820 55050
rect 756 54990 820 54994
rect 508 54903 572 54907
rect 508 54847 512 54903
rect 512 54847 568 54903
rect 568 54847 572 54903
rect 508 54843 572 54847
rect 630 54903 694 54907
rect 630 54847 634 54903
rect 634 54847 690 54903
rect 690 54847 694 54903
rect 630 54843 694 54847
rect 756 54903 820 54907
rect 756 54847 760 54903
rect 760 54847 816 54903
rect 816 54847 820 54903
rect 756 54843 820 54847
rect 508 54766 572 54770
rect 508 54710 512 54766
rect 512 54710 568 54766
rect 568 54710 572 54766
rect 508 54706 572 54710
rect 630 54766 694 54770
rect 630 54710 634 54766
rect 634 54710 690 54766
rect 690 54710 694 54766
rect 630 54706 694 54710
rect 756 54766 820 54770
rect 756 54710 760 54766
rect 760 54710 816 54766
rect 816 54710 820 54766
rect 756 54706 820 54710
rect 22014 54069 22078 54073
rect 22014 54013 22018 54069
rect 22018 54013 22074 54069
rect 22074 54013 22078 54069
rect 22014 54009 22078 54013
rect 22140 54069 22204 54073
rect 22140 54013 22144 54069
rect 22144 54013 22200 54069
rect 22200 54013 22204 54069
rect 22140 54009 22204 54013
rect 22260 54069 22324 54073
rect 22260 54013 22264 54069
rect 22264 54013 22320 54069
rect 22320 54013 22324 54069
rect 22260 54009 22324 54013
rect 22014 53951 22078 53955
rect 22014 53895 22018 53951
rect 22018 53895 22074 53951
rect 22074 53895 22078 53951
rect 22014 53891 22078 53895
rect 22140 53951 22204 53955
rect 22140 53895 22144 53951
rect 22144 53895 22200 53951
rect 22200 53895 22204 53951
rect 22140 53891 22204 53895
rect 22260 53951 22324 53955
rect 22260 53895 22264 53951
rect 22264 53895 22320 53951
rect 22320 53895 22324 53951
rect 22260 53891 22324 53895
rect 508 53291 572 53295
rect 508 53235 512 53291
rect 512 53235 568 53291
rect 568 53235 572 53291
rect 508 53231 572 53235
rect 630 53291 694 53295
rect 630 53235 634 53291
rect 634 53235 690 53291
rect 690 53235 694 53291
rect 630 53231 694 53235
rect 756 53291 820 53295
rect 756 53235 760 53291
rect 760 53235 816 53291
rect 816 53235 820 53291
rect 756 53231 820 53235
rect 508 53144 572 53148
rect 508 53088 512 53144
rect 512 53088 568 53144
rect 568 53088 572 53144
rect 508 53084 572 53088
rect 630 53144 694 53148
rect 630 53088 634 53144
rect 634 53088 690 53144
rect 690 53088 694 53144
rect 630 53084 694 53088
rect 756 53144 820 53148
rect 756 53088 760 53144
rect 760 53088 816 53144
rect 816 53088 820 53144
rect 756 53084 820 53088
rect 508 53007 572 53011
rect 508 52951 512 53007
rect 512 52951 568 53007
rect 568 52951 572 53007
rect 508 52947 572 52951
rect 630 53007 694 53011
rect 630 52951 634 53007
rect 634 52951 690 53007
rect 690 52951 694 53007
rect 630 52947 694 52951
rect 756 53007 820 53011
rect 756 52951 760 53007
rect 760 52951 816 53007
rect 816 52951 820 53007
rect 756 52947 820 52951
rect 507 52721 571 52725
rect 507 52665 511 52721
rect 511 52665 567 52721
rect 567 52665 571 52721
rect 507 52661 571 52665
rect 633 52721 697 52725
rect 633 52665 637 52721
rect 637 52665 693 52721
rect 693 52665 697 52721
rect 633 52661 697 52665
rect 753 52721 817 52725
rect 753 52665 757 52721
rect 757 52665 813 52721
rect 813 52665 817 52721
rect 753 52661 817 52665
rect 507 52603 571 52607
rect 507 52547 511 52603
rect 511 52547 567 52603
rect 567 52547 571 52603
rect 507 52543 571 52547
rect 633 52603 697 52607
rect 633 52547 637 52603
rect 637 52547 693 52603
rect 693 52547 697 52603
rect 633 52543 697 52547
rect 753 52603 817 52607
rect 753 52547 757 52603
rect 757 52547 813 52603
rect 813 52547 817 52603
rect 753 52543 817 52547
rect 21072 52565 21136 52569
rect 21072 52509 21076 52565
rect 21076 52509 21132 52565
rect 21132 52509 21136 52565
rect 21072 52505 21136 52509
rect 21198 52565 21262 52569
rect 21198 52509 21202 52565
rect 21202 52509 21258 52565
rect 21258 52509 21262 52565
rect 21198 52505 21262 52509
rect 21318 52565 21382 52569
rect 21318 52509 21322 52565
rect 21322 52509 21378 52565
rect 21378 52509 21382 52565
rect 21318 52505 21382 52509
rect 21072 52447 21136 52451
rect 21072 52391 21076 52447
rect 21076 52391 21132 52447
rect 21132 52391 21136 52447
rect 21072 52387 21136 52391
rect 21198 52447 21262 52451
rect 21198 52391 21202 52447
rect 21202 52391 21258 52447
rect 21258 52391 21262 52447
rect 21198 52387 21262 52391
rect 21318 52447 21382 52451
rect 21318 52391 21322 52447
rect 21322 52391 21378 52447
rect 21378 52391 21382 52447
rect 21318 52387 21382 52391
rect 507 51534 571 51538
rect 507 51478 511 51534
rect 511 51478 567 51534
rect 567 51478 571 51534
rect 507 51474 571 51478
rect 633 51534 697 51538
rect 633 51478 637 51534
rect 637 51478 693 51534
rect 693 51478 697 51534
rect 633 51474 697 51478
rect 753 51534 817 51538
rect 753 51478 757 51534
rect 757 51478 813 51534
rect 813 51478 817 51534
rect 753 51474 817 51478
rect 507 51416 571 51420
rect 507 51360 511 51416
rect 511 51360 567 51416
rect 567 51360 571 51416
rect 507 51356 571 51360
rect 633 51416 697 51420
rect 633 51360 637 51416
rect 637 51360 693 51416
rect 693 51360 697 51416
rect 633 51356 697 51360
rect 753 51416 817 51420
rect 753 51360 757 51416
rect 757 51360 813 51416
rect 813 51360 817 51416
rect 753 51356 817 51360
rect 21072 51430 21136 51434
rect 21072 51374 21076 51430
rect 21076 51374 21132 51430
rect 21132 51374 21136 51430
rect 21072 51370 21136 51374
rect 21198 51430 21262 51434
rect 21198 51374 21202 51430
rect 21202 51374 21258 51430
rect 21258 51374 21262 51430
rect 21198 51370 21262 51374
rect 21318 51430 21382 51434
rect 21318 51374 21322 51430
rect 21322 51374 21378 51430
rect 21378 51374 21382 51430
rect 21318 51370 21382 51374
rect 21072 51312 21136 51316
rect 21072 51256 21076 51312
rect 21076 51256 21132 51312
rect 21132 51256 21136 51312
rect 21072 51252 21136 51256
rect 21198 51312 21262 51316
rect 21198 51256 21202 51312
rect 21202 51256 21258 51312
rect 21258 51256 21262 51312
rect 21198 51252 21262 51256
rect 21318 51312 21382 51316
rect 21318 51256 21322 51312
rect 21322 51256 21378 51312
rect 21378 51256 21382 51312
rect 21318 51252 21382 51256
rect 508 51050 572 51054
rect 508 50994 512 51050
rect 512 50994 568 51050
rect 568 50994 572 51050
rect 508 50990 572 50994
rect 630 51050 694 51054
rect 630 50994 634 51050
rect 634 50994 690 51050
rect 690 50994 694 51050
rect 630 50990 694 50994
rect 756 51050 820 51054
rect 756 50994 760 51050
rect 760 50994 816 51050
rect 816 50994 820 51050
rect 756 50990 820 50994
rect 508 50903 572 50907
rect 508 50847 512 50903
rect 512 50847 568 50903
rect 568 50847 572 50903
rect 508 50843 572 50847
rect 630 50903 694 50907
rect 630 50847 634 50903
rect 634 50847 690 50903
rect 690 50847 694 50903
rect 630 50843 694 50847
rect 756 50903 820 50907
rect 756 50847 760 50903
rect 760 50847 816 50903
rect 816 50847 820 50903
rect 756 50843 820 50847
rect 508 50766 572 50770
rect 508 50710 512 50766
rect 512 50710 568 50766
rect 568 50710 572 50766
rect 508 50706 572 50710
rect 630 50766 694 50770
rect 630 50710 634 50766
rect 634 50710 690 50766
rect 690 50710 694 50766
rect 630 50706 694 50710
rect 756 50766 820 50770
rect 756 50710 760 50766
rect 760 50710 816 50766
rect 816 50710 820 50766
rect 756 50706 820 50710
rect 22014 50148 22078 50152
rect 22014 50092 22018 50148
rect 22018 50092 22074 50148
rect 22074 50092 22078 50148
rect 22014 50088 22078 50092
rect 22140 50148 22204 50152
rect 22140 50092 22144 50148
rect 22144 50092 22200 50148
rect 22200 50092 22204 50148
rect 22140 50088 22204 50092
rect 22260 50148 22324 50152
rect 22260 50092 22264 50148
rect 22264 50092 22320 50148
rect 22320 50092 22324 50148
rect 22260 50088 22324 50092
rect 22014 50030 22078 50034
rect 22014 49974 22018 50030
rect 22018 49974 22074 50030
rect 22074 49974 22078 50030
rect 22014 49970 22078 49974
rect 22140 50030 22204 50034
rect 22140 49974 22144 50030
rect 22144 49974 22200 50030
rect 22200 49974 22204 50030
rect 22140 49970 22204 49974
rect 22260 50030 22324 50034
rect 22260 49974 22264 50030
rect 22264 49974 22320 50030
rect 22320 49974 22324 50030
rect 22260 49970 22324 49974
rect 508 49291 572 49295
rect 508 49235 512 49291
rect 512 49235 568 49291
rect 568 49235 572 49291
rect 508 49231 572 49235
rect 630 49291 694 49295
rect 630 49235 634 49291
rect 634 49235 690 49291
rect 690 49235 694 49291
rect 630 49231 694 49235
rect 756 49291 820 49295
rect 756 49235 760 49291
rect 760 49235 816 49291
rect 816 49235 820 49291
rect 756 49231 820 49235
rect 508 49144 572 49148
rect 508 49088 512 49144
rect 512 49088 568 49144
rect 568 49088 572 49144
rect 508 49084 572 49088
rect 630 49144 694 49148
rect 630 49088 634 49144
rect 634 49088 690 49144
rect 690 49088 694 49144
rect 630 49084 694 49088
rect 756 49144 820 49148
rect 756 49088 760 49144
rect 760 49088 816 49144
rect 816 49088 820 49144
rect 756 49084 820 49088
rect 508 49007 572 49011
rect 508 48951 512 49007
rect 512 48951 568 49007
rect 568 48951 572 49007
rect 508 48947 572 48951
rect 630 49007 694 49011
rect 630 48951 634 49007
rect 634 48951 690 49007
rect 690 48951 694 49007
rect 630 48947 694 48951
rect 756 49007 820 49011
rect 756 48951 760 49007
rect 760 48951 816 49007
rect 816 48951 820 49007
rect 756 48947 820 48951
rect 507 48712 571 48716
rect 507 48656 511 48712
rect 511 48656 567 48712
rect 567 48656 571 48712
rect 507 48652 571 48656
rect 633 48712 697 48716
rect 633 48656 637 48712
rect 637 48656 693 48712
rect 693 48656 697 48712
rect 633 48652 697 48656
rect 753 48712 817 48716
rect 753 48656 757 48712
rect 757 48656 813 48712
rect 813 48656 817 48712
rect 753 48652 817 48656
rect 507 48594 571 48598
rect 507 48538 511 48594
rect 511 48538 567 48594
rect 567 48538 571 48594
rect 507 48534 571 48538
rect 633 48594 697 48598
rect 633 48538 637 48594
rect 637 48538 693 48594
rect 693 48538 697 48594
rect 633 48534 697 48538
rect 753 48594 817 48598
rect 753 48538 757 48594
rect 757 48538 813 48594
rect 813 48538 817 48594
rect 753 48534 817 48538
rect 21072 48671 21136 48675
rect 21072 48615 21076 48671
rect 21076 48615 21132 48671
rect 21132 48615 21136 48671
rect 21072 48611 21136 48615
rect 21198 48671 21262 48675
rect 21198 48615 21202 48671
rect 21202 48615 21258 48671
rect 21258 48615 21262 48671
rect 21198 48611 21262 48615
rect 21318 48671 21382 48675
rect 21318 48615 21322 48671
rect 21322 48615 21378 48671
rect 21378 48615 21382 48671
rect 21318 48611 21382 48615
rect 21072 48553 21136 48557
rect 21072 48497 21076 48553
rect 21076 48497 21132 48553
rect 21132 48497 21136 48553
rect 21072 48493 21136 48497
rect 21198 48553 21262 48557
rect 21198 48497 21202 48553
rect 21202 48497 21258 48553
rect 21258 48497 21262 48553
rect 21198 48493 21262 48497
rect 21318 48553 21382 48557
rect 21318 48497 21322 48553
rect 21322 48497 21378 48553
rect 21378 48497 21382 48553
rect 21318 48493 21382 48497
rect 507 47559 571 47563
rect 507 47503 511 47559
rect 511 47503 567 47559
rect 567 47503 571 47559
rect 507 47499 571 47503
rect 633 47559 697 47563
rect 633 47503 637 47559
rect 637 47503 693 47559
rect 693 47503 697 47559
rect 633 47499 697 47503
rect 753 47559 817 47563
rect 753 47503 757 47559
rect 757 47503 813 47559
rect 813 47503 817 47559
rect 753 47499 817 47503
rect 507 47441 571 47445
rect 507 47385 511 47441
rect 511 47385 567 47441
rect 567 47385 571 47441
rect 507 47381 571 47385
rect 633 47441 697 47445
rect 633 47385 637 47441
rect 637 47385 693 47441
rect 693 47385 697 47441
rect 633 47381 697 47385
rect 753 47441 817 47445
rect 753 47385 757 47441
rect 757 47385 813 47441
rect 813 47385 817 47441
rect 753 47381 817 47385
rect 21072 47518 21136 47522
rect 21072 47462 21076 47518
rect 21076 47462 21132 47518
rect 21132 47462 21136 47518
rect 21072 47458 21136 47462
rect 21198 47518 21262 47522
rect 21198 47462 21202 47518
rect 21202 47462 21258 47518
rect 21258 47462 21262 47518
rect 21198 47458 21262 47462
rect 21318 47518 21382 47522
rect 21318 47462 21322 47518
rect 21322 47462 21378 47518
rect 21378 47462 21382 47518
rect 21318 47458 21382 47462
rect 21072 47400 21136 47404
rect 21072 47344 21076 47400
rect 21076 47344 21132 47400
rect 21132 47344 21136 47400
rect 21072 47340 21136 47344
rect 21198 47400 21262 47404
rect 21198 47344 21202 47400
rect 21202 47344 21258 47400
rect 21258 47344 21262 47400
rect 21198 47340 21262 47344
rect 21318 47400 21382 47404
rect 21318 47344 21322 47400
rect 21322 47344 21378 47400
rect 21378 47344 21382 47400
rect 21318 47340 21382 47344
rect 508 47050 572 47054
rect 508 46994 512 47050
rect 512 46994 568 47050
rect 568 46994 572 47050
rect 508 46990 572 46994
rect 630 47050 694 47054
rect 630 46994 634 47050
rect 634 46994 690 47050
rect 690 46994 694 47050
rect 630 46990 694 46994
rect 756 47050 820 47054
rect 756 46994 760 47050
rect 760 46994 816 47050
rect 816 46994 820 47050
rect 756 46990 820 46994
rect 508 46903 572 46907
rect 508 46847 512 46903
rect 512 46847 568 46903
rect 568 46847 572 46903
rect 508 46843 572 46847
rect 630 46903 694 46907
rect 630 46847 634 46903
rect 634 46847 690 46903
rect 690 46847 694 46903
rect 630 46843 694 46847
rect 756 46903 820 46907
rect 756 46847 760 46903
rect 760 46847 816 46903
rect 816 46847 820 46903
rect 756 46843 820 46847
rect 508 46766 572 46770
rect 508 46710 512 46766
rect 512 46710 568 46766
rect 568 46710 572 46766
rect 508 46706 572 46710
rect 630 46766 694 46770
rect 630 46710 634 46766
rect 634 46710 690 46766
rect 690 46710 694 46766
rect 630 46706 694 46710
rect 756 46766 820 46770
rect 756 46710 760 46766
rect 760 46710 816 46766
rect 816 46710 820 46766
rect 756 46706 820 46710
rect 22014 45890 22078 45894
rect 22014 45834 22018 45890
rect 22018 45834 22074 45890
rect 22074 45834 22078 45890
rect 22014 45830 22078 45834
rect 22140 45890 22204 45894
rect 22140 45834 22144 45890
rect 22144 45834 22200 45890
rect 22200 45834 22204 45890
rect 22140 45830 22204 45834
rect 22260 45890 22324 45894
rect 22260 45834 22264 45890
rect 22264 45834 22320 45890
rect 22320 45834 22324 45890
rect 22260 45830 22324 45834
rect 22014 45772 22078 45776
rect 22014 45716 22018 45772
rect 22018 45716 22074 45772
rect 22074 45716 22078 45772
rect 22014 45712 22078 45716
rect 22140 45772 22204 45776
rect 22140 45716 22144 45772
rect 22144 45716 22200 45772
rect 22200 45716 22204 45772
rect 22140 45712 22204 45716
rect 22260 45772 22324 45776
rect 22260 45716 22264 45772
rect 22264 45716 22320 45772
rect 22320 45716 22324 45772
rect 22260 45712 22324 45716
rect 508 45290 572 45294
rect 508 45234 512 45290
rect 512 45234 568 45290
rect 568 45234 572 45290
rect 508 45230 572 45234
rect 630 45290 694 45294
rect 630 45234 634 45290
rect 634 45234 690 45290
rect 690 45234 694 45290
rect 630 45230 694 45234
rect 756 45290 820 45294
rect 756 45234 760 45290
rect 760 45234 816 45290
rect 816 45234 820 45290
rect 756 45230 820 45234
rect 508 45143 572 45147
rect 508 45087 512 45143
rect 512 45087 568 45143
rect 568 45087 572 45143
rect 508 45083 572 45087
rect 630 45143 694 45147
rect 630 45087 634 45143
rect 634 45087 690 45143
rect 690 45087 694 45143
rect 630 45083 694 45087
rect 756 45143 820 45147
rect 756 45087 760 45143
rect 760 45087 816 45143
rect 816 45087 820 45143
rect 756 45083 820 45087
rect 508 45006 572 45010
rect 508 44950 512 45006
rect 512 44950 568 45006
rect 568 44950 572 45006
rect 508 44946 572 44950
rect 630 45006 694 45010
rect 630 44950 634 45006
rect 634 44950 690 45006
rect 690 44950 694 45006
rect 630 44946 694 44950
rect 756 45006 820 45010
rect 756 44950 760 45006
rect 760 44950 816 45006
rect 816 44950 820 45006
rect 756 44946 820 44950
rect 507 44499 571 44503
rect 507 44443 511 44499
rect 511 44443 567 44499
rect 567 44443 571 44499
rect 507 44439 571 44443
rect 633 44499 697 44503
rect 633 44443 637 44499
rect 637 44443 693 44499
rect 693 44443 697 44499
rect 633 44439 697 44443
rect 753 44499 817 44503
rect 753 44443 757 44499
rect 757 44443 813 44499
rect 813 44443 817 44499
rect 753 44439 817 44443
rect 507 44381 571 44385
rect 507 44325 511 44381
rect 511 44325 567 44381
rect 567 44325 571 44381
rect 507 44321 571 44325
rect 633 44381 697 44385
rect 633 44325 637 44381
rect 637 44325 693 44381
rect 693 44325 697 44381
rect 633 44321 697 44325
rect 753 44381 817 44385
rect 753 44325 757 44381
rect 757 44325 813 44381
rect 813 44325 817 44381
rect 753 44321 817 44325
rect 21072 44402 21136 44406
rect 21072 44346 21076 44402
rect 21076 44346 21132 44402
rect 21132 44346 21136 44402
rect 21072 44342 21136 44346
rect 21198 44402 21262 44406
rect 21198 44346 21202 44402
rect 21202 44346 21258 44402
rect 21258 44346 21262 44402
rect 21198 44342 21262 44346
rect 21318 44402 21382 44406
rect 21318 44346 21322 44402
rect 21322 44346 21378 44402
rect 21378 44346 21382 44402
rect 21318 44342 21382 44346
rect 21072 44284 21136 44288
rect 21072 44228 21076 44284
rect 21076 44228 21132 44284
rect 21132 44228 21136 44284
rect 21072 44224 21136 44228
rect 21198 44284 21262 44288
rect 21198 44228 21202 44284
rect 21202 44228 21258 44284
rect 21258 44228 21262 44284
rect 21198 44224 21262 44228
rect 21318 44284 21382 44288
rect 21318 44228 21322 44284
rect 21322 44228 21378 44284
rect 21378 44228 21382 44284
rect 21318 44224 21382 44228
rect 22040 43824 22264 43828
rect 22040 43528 22044 43824
rect 22044 43528 22260 43824
rect 22260 43528 22264 43824
rect 22040 43524 22264 43528
rect 2249 39861 2257 39925
rect 2257 39861 2313 39925
rect 2337 39861 2393 39925
rect 2393 39861 2401 39925
rect 2249 39789 2257 39845
rect 2257 39789 2313 39845
rect 2337 39789 2393 39845
rect 2393 39789 2401 39845
rect 2249 39781 2313 39789
rect 2337 39781 2401 39789
rect 4192 39841 4256 39905
rect 4280 39841 4344 39905
rect 4192 39761 4256 39825
rect 4280 39761 4344 39825
rect 39 39729 103 39733
rect 39 39673 44 39729
rect 44 39673 100 39729
rect 100 39673 103 39729
rect 39 39669 103 39673
rect 164 39729 228 39733
rect 164 39673 169 39729
rect 169 39673 225 39729
rect 225 39673 228 39729
rect 164 39669 228 39673
rect 290 39729 354 39733
rect 290 39673 294 39729
rect 294 39673 350 39729
rect 350 39673 354 39729
rect 290 39669 354 39673
rect 39 39623 103 39627
rect 39 39567 44 39623
rect 44 39567 100 39623
rect 100 39567 103 39623
rect 39 39563 103 39567
rect 164 39623 228 39627
rect 164 39567 169 39623
rect 169 39567 225 39623
rect 225 39567 228 39623
rect 164 39563 228 39567
rect 290 39623 354 39627
rect 290 39567 294 39623
rect 294 39567 350 39623
rect 350 39567 354 39623
rect 290 39563 354 39567
rect 21543 39714 21607 39718
rect 21543 39658 21547 39714
rect 21547 39658 21603 39714
rect 21603 39658 21607 39714
rect 21543 39654 21607 39658
rect 21668 39714 21732 39718
rect 21668 39658 21672 39714
rect 21672 39658 21728 39714
rect 21728 39658 21732 39714
rect 21668 39654 21732 39658
rect 21793 39714 21857 39718
rect 21793 39658 21797 39714
rect 21797 39658 21853 39714
rect 21853 39658 21857 39714
rect 21793 39654 21857 39658
rect 21542 39594 21606 39598
rect 21542 39538 21546 39594
rect 21546 39538 21602 39594
rect 21602 39538 21606 39594
rect 21542 39534 21606 39538
rect 21667 39594 21731 39598
rect 21667 39538 21671 39594
rect 21671 39538 21727 39594
rect 21727 39538 21731 39594
rect 21667 39534 21731 39538
rect 21792 39594 21856 39598
rect 21792 39538 21796 39594
rect 21796 39538 21852 39594
rect 21852 39538 21856 39594
rect 21792 39534 21856 39538
rect 488 39119 552 39123
rect 488 39063 492 39119
rect 492 39063 548 39119
rect 548 39063 552 39119
rect 488 39059 552 39063
rect 602 39119 666 39123
rect 602 39063 606 39119
rect 606 39063 662 39119
rect 662 39063 666 39119
rect 602 39059 666 39063
rect 716 39119 780 39123
rect 716 39063 720 39119
rect 720 39063 776 39119
rect 776 39063 780 39119
rect 716 39059 780 39063
rect 25 38575 89 38579
rect 25 38519 29 38575
rect 29 38519 85 38575
rect 85 38519 89 38575
rect 25 38515 89 38519
rect 139 38575 203 38579
rect 139 38519 143 38575
rect 143 38519 199 38575
rect 199 38519 203 38575
rect 139 38515 203 38519
rect 253 38575 317 38579
rect 253 38519 257 38575
rect 257 38519 313 38575
rect 313 38519 317 38575
rect 253 38515 317 38519
rect 488 38031 552 38035
rect 488 37975 492 38031
rect 492 37975 548 38031
rect 548 37975 552 38031
rect 488 37971 552 37975
rect 602 38031 666 38035
rect 602 37975 606 38031
rect 606 37975 662 38031
rect 662 37975 666 38031
rect 602 37971 666 37975
rect 716 38031 780 38035
rect 716 37975 720 38031
rect 720 37975 776 38031
rect 776 37975 780 38031
rect 716 37971 780 37975
rect 25 37487 89 37491
rect 25 37431 29 37487
rect 29 37431 85 37487
rect 85 37431 89 37487
rect 25 37427 89 37431
rect 139 37487 203 37491
rect 139 37431 143 37487
rect 143 37431 199 37487
rect 199 37431 203 37487
rect 139 37427 203 37431
rect 253 37487 317 37491
rect 253 37431 257 37487
rect 257 37431 313 37487
rect 313 37431 317 37487
rect 253 37427 317 37431
rect 488 36943 552 36947
rect 488 36887 492 36943
rect 492 36887 548 36943
rect 548 36887 552 36943
rect 488 36883 552 36887
rect 602 36943 666 36947
rect 602 36887 606 36943
rect 606 36887 662 36943
rect 662 36887 666 36943
rect 602 36883 666 36887
rect 716 36943 780 36947
rect 716 36887 720 36943
rect 720 36887 776 36943
rect 776 36887 780 36943
rect 716 36883 780 36887
rect 22040 36940 22264 36944
rect 22040 36644 22044 36940
rect 22044 36644 22260 36940
rect 22260 36644 22264 36940
rect 22040 36640 22264 36644
rect 2536 36460 2600 36463
rect 2536 36404 2544 36460
rect 2544 36404 2600 36460
rect 2536 36399 2600 36404
rect 2624 36460 2688 36463
rect 2624 36404 2680 36460
rect 2680 36404 2688 36460
rect 2624 36399 2688 36404
rect 21069 36160 21133 36164
rect 21069 36104 21073 36160
rect 21073 36104 21129 36160
rect 21129 36104 21133 36160
rect 21069 36100 21133 36104
rect 21194 36160 21258 36164
rect 21194 36104 21198 36160
rect 21198 36104 21254 36160
rect 21254 36104 21258 36160
rect 21194 36100 21258 36104
rect 21319 36160 21383 36164
rect 21319 36104 21323 36160
rect 21323 36104 21379 36160
rect 21379 36104 21383 36160
rect 21319 36100 21383 36104
rect 21068 36040 21132 36044
rect 21068 35984 21072 36040
rect 21072 35984 21128 36040
rect 21128 35984 21132 36040
rect 21068 35980 21132 35984
rect 21193 36040 21257 36044
rect 21193 35984 21197 36040
rect 21197 35984 21253 36040
rect 21253 35984 21257 36040
rect 21193 35980 21257 35984
rect 21318 36040 21382 36044
rect 21318 35984 21322 36040
rect 21322 35984 21378 36040
rect 21378 35984 21382 36040
rect 21318 35980 21382 35984
rect 21073 35582 21137 35586
rect 21073 35526 21077 35582
rect 21077 35526 21133 35582
rect 21133 35526 21137 35582
rect 21073 35522 21137 35526
rect 21195 35582 21259 35586
rect 21195 35526 21199 35582
rect 21199 35526 21255 35582
rect 21255 35526 21259 35582
rect 21195 35522 21259 35526
rect 21321 35582 21385 35586
rect 21321 35526 21325 35582
rect 21325 35526 21381 35582
rect 21381 35526 21385 35582
rect 21321 35522 21385 35526
rect 21073 35435 21137 35439
rect 21073 35379 21077 35435
rect 21077 35379 21133 35435
rect 21133 35379 21137 35435
rect 21073 35375 21137 35379
rect 21195 35435 21259 35439
rect 21195 35379 21199 35435
rect 21199 35379 21255 35435
rect 21255 35379 21259 35435
rect 21195 35375 21259 35379
rect 21321 35435 21385 35439
rect 21321 35379 21325 35435
rect 21325 35379 21381 35435
rect 21381 35379 21385 35435
rect 21321 35375 21385 35379
rect 21073 35298 21137 35302
rect 21073 35242 21077 35298
rect 21077 35242 21133 35298
rect 21133 35242 21137 35298
rect 21073 35238 21137 35242
rect 21195 35298 21259 35302
rect 21195 35242 21199 35298
rect 21199 35242 21255 35298
rect 21255 35242 21259 35298
rect 21195 35238 21259 35242
rect 21321 35298 21385 35302
rect 21321 35242 21325 35298
rect 21325 35242 21381 35298
rect 21381 35242 21385 35298
rect 21321 35238 21385 35242
rect 20568 34664 20632 34668
rect 20568 34608 20572 34664
rect 20572 34608 20628 34664
rect 20628 34608 20632 34664
rect 20568 34604 20632 34608
rect 20693 34664 20757 34668
rect 20693 34608 20697 34664
rect 20697 34608 20753 34664
rect 20753 34608 20757 34664
rect 20693 34604 20757 34608
rect 20818 34664 20882 34668
rect 20818 34608 20822 34664
rect 20822 34608 20878 34664
rect 20878 34608 20882 34664
rect 20818 34604 20882 34608
rect 20567 34544 20631 34548
rect 20567 34488 20571 34544
rect 20571 34488 20627 34544
rect 20627 34488 20631 34544
rect 20567 34484 20631 34488
rect 20692 34544 20756 34548
rect 20692 34488 20696 34544
rect 20696 34488 20752 34544
rect 20752 34488 20756 34544
rect 20692 34484 20756 34488
rect 20817 34544 20881 34548
rect 20817 34488 20821 34544
rect 20821 34488 20877 34544
rect 20877 34488 20881 34544
rect 20817 34484 20881 34488
rect 21543 34664 21607 34668
rect 21543 34608 21547 34664
rect 21547 34608 21603 34664
rect 21603 34608 21607 34664
rect 21543 34604 21607 34608
rect 21668 34664 21732 34668
rect 21668 34608 21672 34664
rect 21672 34608 21728 34664
rect 21728 34608 21732 34664
rect 21668 34604 21732 34608
rect 21793 34664 21857 34668
rect 21793 34608 21797 34664
rect 21797 34608 21853 34664
rect 21853 34608 21857 34664
rect 21793 34604 21857 34608
rect 21542 34544 21606 34548
rect 21542 34488 21546 34544
rect 21546 34488 21602 34544
rect 21602 34488 21606 34544
rect 21542 34484 21606 34488
rect 21667 34544 21731 34548
rect 21667 34488 21671 34544
rect 21671 34488 21727 34544
rect 21727 34488 21731 34544
rect 21667 34484 21731 34488
rect 21792 34544 21856 34548
rect 21792 34488 21796 34544
rect 21796 34488 21852 34544
rect 21852 34488 21856 34544
rect 21792 34484 21856 34488
rect 21073 33822 21137 33826
rect 21073 33766 21077 33822
rect 21077 33766 21133 33822
rect 21133 33766 21137 33822
rect 21073 33762 21137 33766
rect 21195 33822 21259 33826
rect 21195 33766 21199 33822
rect 21199 33766 21255 33822
rect 21255 33766 21259 33822
rect 21195 33762 21259 33766
rect 21321 33822 21385 33826
rect 21321 33766 21325 33822
rect 21325 33766 21381 33822
rect 21381 33766 21385 33822
rect 21321 33762 21385 33766
rect 21073 33675 21137 33679
rect 21073 33619 21077 33675
rect 21077 33619 21133 33675
rect 21133 33619 21137 33675
rect 21073 33615 21137 33619
rect 21195 33675 21259 33679
rect 21195 33619 21199 33675
rect 21199 33619 21255 33675
rect 21255 33619 21259 33675
rect 21195 33615 21259 33619
rect 21321 33675 21385 33679
rect 21321 33619 21325 33675
rect 21325 33619 21381 33675
rect 21381 33619 21385 33675
rect 21321 33615 21385 33619
rect 21073 33538 21137 33542
rect 21073 33482 21077 33538
rect 21077 33482 21133 33538
rect 21133 33482 21137 33538
rect 21073 33478 21137 33482
rect 21195 33538 21259 33542
rect 21195 33482 21199 33538
rect 21199 33482 21255 33538
rect 21255 33482 21259 33538
rect 21195 33478 21259 33482
rect 21321 33538 21385 33542
rect 21321 33482 21325 33538
rect 21325 33482 21381 33538
rect 21381 33482 21385 33538
rect 21321 33478 21385 33482
rect 21068 33105 21132 33109
rect 21068 33049 21072 33105
rect 21072 33049 21128 33105
rect 21128 33049 21132 33105
rect 21068 33045 21132 33049
rect 21193 33105 21257 33109
rect 21193 33049 21197 33105
rect 21197 33049 21253 33105
rect 21253 33049 21257 33105
rect 21193 33045 21257 33049
rect 21318 33105 21382 33109
rect 21318 33049 21322 33105
rect 21322 33049 21378 33105
rect 21378 33049 21382 33105
rect 21318 33045 21382 33049
rect 21067 32985 21131 32989
rect 21067 32929 21071 32985
rect 21071 32929 21127 32985
rect 21127 32929 21131 32985
rect 21067 32925 21131 32929
rect 21192 32985 21256 32989
rect 21192 32929 21196 32985
rect 21196 32929 21252 32985
rect 21252 32929 21256 32985
rect 21192 32925 21256 32929
rect 21317 32985 21381 32989
rect 21317 32929 21321 32985
rect 21321 32929 21377 32985
rect 21377 32929 21381 32985
rect 21317 32925 21381 32929
rect 507 32292 571 32296
rect 507 32236 511 32292
rect 511 32236 567 32292
rect 567 32236 571 32292
rect 507 32232 571 32236
rect 633 32292 697 32296
rect 633 32236 637 32292
rect 637 32236 693 32292
rect 693 32236 697 32292
rect 633 32232 697 32236
rect 753 32292 817 32296
rect 753 32236 757 32292
rect 757 32236 813 32292
rect 813 32236 817 32292
rect 753 32232 817 32236
rect 507 32174 571 32178
rect 507 32118 511 32174
rect 511 32118 567 32174
rect 567 32118 571 32174
rect 507 32114 571 32118
rect 633 32174 697 32178
rect 633 32118 637 32174
rect 637 32118 693 32174
rect 693 32118 697 32174
rect 633 32114 697 32118
rect 753 32174 817 32178
rect 753 32118 757 32174
rect 757 32118 813 32174
rect 813 32118 817 32174
rect 753 32114 817 32118
rect 21072 32292 21136 32296
rect 21072 32236 21076 32292
rect 21076 32236 21132 32292
rect 21132 32236 21136 32292
rect 21072 32232 21136 32236
rect 21198 32292 21262 32296
rect 21198 32236 21202 32292
rect 21202 32236 21258 32292
rect 21258 32236 21262 32292
rect 21198 32232 21262 32236
rect 21318 32292 21382 32296
rect 21318 32236 21322 32292
rect 21322 32236 21378 32292
rect 21378 32236 21382 32292
rect 21318 32232 21382 32236
rect 21072 32174 21136 32178
rect 21072 32118 21076 32174
rect 21076 32118 21132 32174
rect 21132 32118 21136 32174
rect 21072 32114 21136 32118
rect 21198 32174 21262 32178
rect 21198 32118 21202 32174
rect 21202 32118 21258 32174
rect 21258 32118 21262 32174
rect 21198 32114 21262 32118
rect 21318 32174 21382 32178
rect 21318 32118 21322 32174
rect 21322 32118 21378 32174
rect 21378 32118 21382 32174
rect 21318 32114 21382 32118
rect 507 31510 571 31514
rect 507 31454 511 31510
rect 511 31454 567 31510
rect 567 31454 571 31510
rect 507 31450 571 31454
rect 633 31510 697 31514
rect 633 31454 637 31510
rect 637 31454 693 31510
rect 693 31454 697 31510
rect 633 31450 697 31454
rect 753 31510 817 31514
rect 753 31454 757 31510
rect 757 31454 813 31510
rect 813 31454 817 31510
rect 753 31450 817 31454
rect 507 31392 571 31396
rect 507 31336 511 31392
rect 511 31336 567 31392
rect 567 31336 571 31392
rect 507 31332 571 31336
rect 633 31392 697 31396
rect 633 31336 637 31392
rect 637 31336 693 31392
rect 693 31336 697 31392
rect 633 31332 697 31336
rect 753 31392 817 31396
rect 753 31336 757 31392
rect 757 31336 813 31392
rect 813 31336 817 31392
rect 753 31332 817 31336
rect 21072 31510 21136 31514
rect 21072 31454 21076 31510
rect 21076 31454 21132 31510
rect 21132 31454 21136 31510
rect 21072 31450 21136 31454
rect 21198 31510 21262 31514
rect 21198 31454 21202 31510
rect 21202 31454 21258 31510
rect 21258 31454 21262 31510
rect 21198 31450 21262 31454
rect 21318 31510 21382 31514
rect 21318 31454 21322 31510
rect 21322 31454 21378 31510
rect 21378 31454 21382 31510
rect 21318 31450 21382 31454
rect 21072 31392 21136 31396
rect 21072 31336 21076 31392
rect 21076 31336 21132 31392
rect 21132 31336 21136 31392
rect 21072 31332 21136 31336
rect 21198 31392 21262 31396
rect 21198 31336 21202 31392
rect 21202 31336 21258 31392
rect 21258 31336 21262 31392
rect 21198 31332 21262 31336
rect 21318 31392 21382 31396
rect 21318 31336 21322 31392
rect 21322 31336 21378 31392
rect 21378 31336 21382 31392
rect 21318 31332 21382 31336
rect 508 31051 572 31055
rect 508 30995 512 31051
rect 512 30995 568 31051
rect 568 30995 572 31051
rect 508 30991 572 30995
rect 630 31051 694 31055
rect 630 30995 634 31051
rect 634 30995 690 31051
rect 690 30995 694 31051
rect 630 30991 694 30995
rect 756 31051 820 31055
rect 756 30995 760 31051
rect 760 30995 816 31051
rect 816 30995 820 31051
rect 756 30991 820 30995
rect 508 30904 572 30908
rect 508 30848 512 30904
rect 512 30848 568 30904
rect 568 30848 572 30904
rect 508 30844 572 30848
rect 630 30904 694 30908
rect 630 30848 634 30904
rect 634 30848 690 30904
rect 690 30848 694 30904
rect 630 30844 694 30848
rect 756 30904 820 30908
rect 756 30848 760 30904
rect 760 30848 816 30904
rect 816 30848 820 30904
rect 756 30844 820 30848
rect 508 30767 572 30771
rect 508 30711 512 30767
rect 512 30711 568 30767
rect 568 30711 572 30767
rect 508 30707 572 30711
rect 630 30767 694 30771
rect 630 30711 634 30767
rect 634 30711 690 30767
rect 690 30711 694 30767
rect 630 30707 694 30711
rect 756 30767 820 30771
rect 756 30711 760 30767
rect 760 30711 816 30767
rect 816 30711 820 30767
rect 756 30707 820 30711
rect 22014 30120 22078 30124
rect 22014 30064 22018 30120
rect 22018 30064 22074 30120
rect 22074 30064 22078 30120
rect 22014 30060 22078 30064
rect 22140 30120 22204 30124
rect 22140 30064 22144 30120
rect 22144 30064 22200 30120
rect 22200 30064 22204 30120
rect 22140 30060 22204 30064
rect 22260 30120 22324 30124
rect 22260 30064 22264 30120
rect 22264 30064 22320 30120
rect 22320 30064 22324 30120
rect 22260 30060 22324 30064
rect 22014 30002 22078 30006
rect 22014 29946 22018 30002
rect 22018 29946 22074 30002
rect 22074 29946 22078 30002
rect 22014 29942 22078 29946
rect 22140 30002 22204 30006
rect 22140 29946 22144 30002
rect 22144 29946 22200 30002
rect 22200 29946 22204 30002
rect 22140 29942 22204 29946
rect 22260 30002 22324 30006
rect 22260 29946 22264 30002
rect 22264 29946 22320 30002
rect 22320 29946 22324 30002
rect 22260 29942 22324 29946
rect 508 29284 572 29288
rect 508 29228 512 29284
rect 512 29228 568 29284
rect 568 29228 572 29284
rect 508 29224 572 29228
rect 630 29284 694 29288
rect 630 29228 634 29284
rect 634 29228 690 29284
rect 690 29228 694 29284
rect 630 29224 694 29228
rect 756 29284 820 29288
rect 756 29228 760 29284
rect 760 29228 816 29284
rect 816 29228 820 29284
rect 756 29224 820 29228
rect 508 29137 572 29141
rect 508 29081 512 29137
rect 512 29081 568 29137
rect 568 29081 572 29137
rect 508 29077 572 29081
rect 630 29137 694 29141
rect 630 29081 634 29137
rect 634 29081 690 29137
rect 690 29081 694 29137
rect 630 29077 694 29081
rect 756 29137 820 29141
rect 756 29081 760 29137
rect 760 29081 816 29137
rect 816 29081 820 29137
rect 756 29077 820 29081
rect 508 29000 572 29004
rect 508 28944 512 29000
rect 512 28944 568 29000
rect 568 28944 572 29000
rect 508 28940 572 28944
rect 630 29000 694 29004
rect 630 28944 634 29000
rect 634 28944 690 29000
rect 690 28944 694 29000
rect 630 28940 694 28944
rect 756 29000 820 29004
rect 756 28944 760 29000
rect 760 28944 816 29000
rect 816 28944 820 29000
rect 756 28940 820 28944
rect 507 28598 571 28602
rect 507 28542 511 28598
rect 511 28542 567 28598
rect 567 28542 571 28598
rect 507 28538 571 28542
rect 633 28598 697 28602
rect 633 28542 637 28598
rect 637 28542 693 28598
rect 693 28542 697 28598
rect 633 28538 697 28542
rect 753 28598 817 28602
rect 753 28542 757 28598
rect 757 28542 813 28598
rect 813 28542 817 28598
rect 753 28538 817 28542
rect 507 28480 571 28484
rect 507 28424 511 28480
rect 511 28424 567 28480
rect 567 28424 571 28480
rect 507 28420 571 28424
rect 633 28480 697 28484
rect 633 28424 637 28480
rect 637 28424 693 28480
rect 693 28424 697 28480
rect 633 28420 697 28424
rect 753 28480 817 28484
rect 753 28424 757 28480
rect 757 28424 813 28480
rect 813 28424 817 28480
rect 753 28420 817 28424
rect 21072 28549 21136 28553
rect 21072 28493 21076 28549
rect 21076 28493 21132 28549
rect 21132 28493 21136 28549
rect 21072 28489 21136 28493
rect 21198 28549 21262 28553
rect 21198 28493 21202 28549
rect 21202 28493 21258 28549
rect 21258 28493 21262 28549
rect 21198 28489 21262 28493
rect 21318 28549 21382 28553
rect 21318 28493 21322 28549
rect 21322 28493 21378 28549
rect 21378 28493 21382 28549
rect 21318 28489 21382 28493
rect 21072 28431 21136 28435
rect 21072 28375 21076 28431
rect 21076 28375 21132 28431
rect 21132 28375 21136 28431
rect 21072 28371 21136 28375
rect 21198 28431 21262 28435
rect 21198 28375 21202 28431
rect 21202 28375 21258 28431
rect 21258 28375 21262 28431
rect 21198 28371 21262 28375
rect 21318 28431 21382 28435
rect 21318 28375 21322 28431
rect 21322 28375 21378 28431
rect 21378 28375 21382 28431
rect 21318 28371 21382 28375
rect 507 27594 571 27598
rect 507 27538 511 27594
rect 511 27538 567 27594
rect 567 27538 571 27594
rect 507 27534 571 27538
rect 633 27594 697 27598
rect 633 27538 637 27594
rect 637 27538 693 27594
rect 693 27538 697 27594
rect 633 27534 697 27538
rect 753 27594 817 27598
rect 753 27538 757 27594
rect 757 27538 813 27594
rect 813 27538 817 27594
rect 753 27534 817 27538
rect 507 27476 571 27480
rect 507 27420 511 27476
rect 511 27420 567 27476
rect 567 27420 571 27476
rect 507 27416 571 27420
rect 633 27476 697 27480
rect 633 27420 637 27476
rect 637 27420 693 27476
rect 693 27420 697 27476
rect 633 27416 697 27420
rect 753 27476 817 27480
rect 753 27420 757 27476
rect 757 27420 813 27476
rect 813 27420 817 27476
rect 753 27416 817 27420
rect 21072 27432 21136 27436
rect 21072 27376 21076 27432
rect 21076 27376 21132 27432
rect 21132 27376 21136 27432
rect 21072 27372 21136 27376
rect 21198 27432 21262 27436
rect 21198 27376 21202 27432
rect 21202 27376 21258 27432
rect 21258 27376 21262 27432
rect 21198 27372 21262 27376
rect 21318 27432 21382 27436
rect 21318 27376 21322 27432
rect 21322 27376 21378 27432
rect 21378 27376 21382 27432
rect 21318 27372 21382 27376
rect 21072 27314 21136 27318
rect 21072 27258 21076 27314
rect 21076 27258 21132 27314
rect 21132 27258 21136 27314
rect 21072 27254 21136 27258
rect 21198 27314 21262 27318
rect 21198 27258 21202 27314
rect 21202 27258 21258 27314
rect 21258 27258 21262 27314
rect 21198 27254 21262 27258
rect 21318 27314 21382 27318
rect 21318 27258 21322 27314
rect 21322 27258 21378 27314
rect 21378 27258 21382 27314
rect 21318 27254 21382 27258
rect 508 27050 572 27054
rect 508 26994 512 27050
rect 512 26994 568 27050
rect 568 26994 572 27050
rect 508 26990 572 26994
rect 630 27050 694 27054
rect 630 26994 634 27050
rect 634 26994 690 27050
rect 690 26994 694 27050
rect 630 26990 694 26994
rect 756 27050 820 27054
rect 756 26994 760 27050
rect 760 26994 816 27050
rect 816 26994 820 27050
rect 756 26990 820 26994
rect 508 26903 572 26907
rect 508 26847 512 26903
rect 512 26847 568 26903
rect 568 26847 572 26903
rect 508 26843 572 26847
rect 630 26903 694 26907
rect 630 26847 634 26903
rect 634 26847 690 26903
rect 690 26847 694 26903
rect 630 26843 694 26847
rect 756 26903 820 26907
rect 756 26847 760 26903
rect 760 26847 816 26903
rect 816 26847 820 26903
rect 756 26843 820 26847
rect 508 26766 572 26770
rect 508 26710 512 26766
rect 512 26710 568 26766
rect 568 26710 572 26766
rect 508 26706 572 26710
rect 630 26766 694 26770
rect 630 26710 634 26766
rect 634 26710 690 26766
rect 690 26710 694 26766
rect 630 26706 694 26710
rect 756 26766 820 26770
rect 756 26710 760 26766
rect 760 26710 816 26766
rect 816 26710 820 26766
rect 756 26706 820 26710
rect 22014 25961 22078 25965
rect 22014 25905 22018 25961
rect 22018 25905 22074 25961
rect 22074 25905 22078 25961
rect 22014 25901 22078 25905
rect 22140 25961 22204 25965
rect 22140 25905 22144 25961
rect 22144 25905 22200 25961
rect 22200 25905 22204 25961
rect 22140 25901 22204 25905
rect 22260 25961 22324 25965
rect 22260 25905 22264 25961
rect 22264 25905 22320 25961
rect 22320 25905 22324 25961
rect 22260 25901 22324 25905
rect 22014 25843 22078 25847
rect 22014 25787 22018 25843
rect 22018 25787 22074 25843
rect 22074 25787 22078 25843
rect 22014 25783 22078 25787
rect 22140 25843 22204 25847
rect 22140 25787 22144 25843
rect 22144 25787 22200 25843
rect 22200 25787 22204 25843
rect 22140 25783 22204 25787
rect 22260 25843 22324 25847
rect 22260 25787 22264 25843
rect 22264 25787 22320 25843
rect 22320 25787 22324 25843
rect 22260 25783 22324 25787
rect 508 25290 572 25294
rect 508 25234 512 25290
rect 512 25234 568 25290
rect 568 25234 572 25290
rect 508 25230 572 25234
rect 630 25290 694 25294
rect 630 25234 634 25290
rect 634 25234 690 25290
rect 690 25234 694 25290
rect 630 25230 694 25234
rect 756 25290 820 25294
rect 756 25234 760 25290
rect 760 25234 816 25290
rect 816 25234 820 25290
rect 756 25230 820 25234
rect 508 25143 572 25147
rect 508 25087 512 25143
rect 512 25087 568 25143
rect 568 25087 572 25143
rect 508 25083 572 25087
rect 630 25143 694 25147
rect 630 25087 634 25143
rect 634 25087 690 25143
rect 690 25087 694 25143
rect 630 25083 694 25087
rect 756 25143 820 25147
rect 756 25087 760 25143
rect 760 25087 816 25143
rect 816 25087 820 25143
rect 756 25083 820 25087
rect 508 25006 572 25010
rect 508 24950 512 25006
rect 512 24950 568 25006
rect 568 24950 572 25006
rect 508 24946 572 24950
rect 630 25006 694 25010
rect 630 24950 634 25006
rect 634 24950 690 25006
rect 690 24950 694 25006
rect 630 24946 694 24950
rect 756 25006 820 25010
rect 756 24950 760 25006
rect 760 24950 816 25006
rect 816 24950 820 25006
rect 756 24946 820 24950
rect 507 24616 571 24620
rect 507 24560 511 24616
rect 511 24560 567 24616
rect 567 24560 571 24616
rect 507 24556 571 24560
rect 633 24616 697 24620
rect 633 24560 637 24616
rect 637 24560 693 24616
rect 693 24560 697 24616
rect 633 24556 697 24560
rect 753 24616 817 24620
rect 753 24560 757 24616
rect 757 24560 813 24616
rect 813 24560 817 24616
rect 753 24556 817 24560
rect 507 24498 571 24502
rect 507 24442 511 24498
rect 511 24442 567 24498
rect 567 24442 571 24498
rect 507 24438 571 24442
rect 633 24498 697 24502
rect 633 24442 637 24498
rect 637 24442 693 24498
rect 693 24442 697 24498
rect 633 24438 697 24442
rect 753 24498 817 24502
rect 753 24442 757 24498
rect 757 24442 813 24498
rect 813 24442 817 24498
rect 753 24438 817 24442
rect 21072 24589 21136 24593
rect 21072 24533 21076 24589
rect 21076 24533 21132 24589
rect 21132 24533 21136 24589
rect 21072 24529 21136 24533
rect 21198 24589 21262 24593
rect 21198 24533 21202 24589
rect 21202 24533 21258 24589
rect 21258 24533 21262 24589
rect 21198 24529 21262 24533
rect 21318 24589 21382 24593
rect 21318 24533 21322 24589
rect 21322 24533 21378 24589
rect 21378 24533 21382 24589
rect 21318 24529 21382 24533
rect 21072 24471 21136 24475
rect 21072 24415 21076 24471
rect 21076 24415 21132 24471
rect 21132 24415 21136 24471
rect 21072 24411 21136 24415
rect 21198 24471 21262 24475
rect 21198 24415 21202 24471
rect 21202 24415 21258 24471
rect 21258 24415 21262 24471
rect 21198 24411 21262 24415
rect 21318 24471 21382 24475
rect 21318 24415 21322 24471
rect 21322 24415 21378 24471
rect 21378 24415 21382 24471
rect 21318 24411 21382 24415
rect 507 23534 571 23538
rect 507 23478 511 23534
rect 511 23478 567 23534
rect 567 23478 571 23534
rect 507 23474 571 23478
rect 633 23534 697 23538
rect 633 23478 637 23534
rect 637 23478 693 23534
rect 693 23478 697 23534
rect 633 23474 697 23478
rect 753 23534 817 23538
rect 753 23478 757 23534
rect 757 23478 813 23534
rect 813 23478 817 23534
rect 753 23474 817 23478
rect 507 23416 571 23420
rect 507 23360 511 23416
rect 511 23360 567 23416
rect 567 23360 571 23416
rect 507 23356 571 23360
rect 633 23416 697 23420
rect 633 23360 637 23416
rect 637 23360 693 23416
rect 693 23360 697 23416
rect 633 23356 697 23360
rect 753 23416 817 23420
rect 753 23360 757 23416
rect 757 23360 813 23416
rect 813 23360 817 23416
rect 753 23356 817 23360
rect 21072 23414 21136 23418
rect 21072 23358 21076 23414
rect 21076 23358 21132 23414
rect 21132 23358 21136 23414
rect 21072 23354 21136 23358
rect 21198 23414 21262 23418
rect 21198 23358 21202 23414
rect 21202 23358 21258 23414
rect 21258 23358 21262 23414
rect 21198 23354 21262 23358
rect 21318 23414 21382 23418
rect 21318 23358 21322 23414
rect 21322 23358 21378 23414
rect 21378 23358 21382 23414
rect 21318 23354 21382 23358
rect 21072 23296 21136 23300
rect 21072 23240 21076 23296
rect 21076 23240 21132 23296
rect 21132 23240 21136 23296
rect 21072 23236 21136 23240
rect 21198 23296 21262 23300
rect 21198 23240 21202 23296
rect 21202 23240 21258 23296
rect 21258 23240 21262 23296
rect 21198 23236 21262 23240
rect 21318 23296 21382 23300
rect 21318 23240 21322 23296
rect 21322 23240 21378 23296
rect 21378 23240 21382 23296
rect 21318 23236 21382 23240
rect 508 23050 572 23054
rect 508 22994 512 23050
rect 512 22994 568 23050
rect 568 22994 572 23050
rect 508 22990 572 22994
rect 630 23050 694 23054
rect 630 22994 634 23050
rect 634 22994 690 23050
rect 690 22994 694 23050
rect 630 22990 694 22994
rect 756 23050 820 23054
rect 756 22994 760 23050
rect 760 22994 816 23050
rect 816 22994 820 23050
rect 756 22990 820 22994
rect 508 22903 572 22907
rect 508 22847 512 22903
rect 512 22847 568 22903
rect 568 22847 572 22903
rect 508 22843 572 22847
rect 630 22903 694 22907
rect 630 22847 634 22903
rect 634 22847 690 22903
rect 690 22847 694 22903
rect 630 22843 694 22847
rect 756 22903 820 22907
rect 756 22847 760 22903
rect 760 22847 816 22903
rect 816 22847 820 22903
rect 756 22843 820 22847
rect 508 22766 572 22770
rect 508 22710 512 22766
rect 512 22710 568 22766
rect 568 22710 572 22766
rect 508 22706 572 22710
rect 630 22766 694 22770
rect 630 22710 634 22766
rect 634 22710 690 22766
rect 690 22710 694 22766
rect 630 22706 694 22710
rect 756 22766 820 22770
rect 756 22710 760 22766
rect 760 22710 816 22766
rect 816 22710 820 22766
rect 756 22706 820 22710
rect 22014 22171 22078 22175
rect 22014 22115 22018 22171
rect 22018 22115 22074 22171
rect 22074 22115 22078 22171
rect 22014 22111 22078 22115
rect 22140 22171 22204 22175
rect 22140 22115 22144 22171
rect 22144 22115 22200 22171
rect 22200 22115 22204 22171
rect 22140 22111 22204 22115
rect 22260 22171 22324 22175
rect 22260 22115 22264 22171
rect 22264 22115 22320 22171
rect 22320 22115 22324 22171
rect 22260 22111 22324 22115
rect 22014 22053 22078 22057
rect 22014 21997 22018 22053
rect 22018 21997 22074 22053
rect 22074 21997 22078 22053
rect 22014 21993 22078 21997
rect 22140 22053 22204 22057
rect 22140 21997 22144 22053
rect 22144 21997 22200 22053
rect 22200 21997 22204 22053
rect 22140 21993 22204 21997
rect 22260 22053 22324 22057
rect 22260 21997 22264 22053
rect 22264 21997 22320 22053
rect 22320 21997 22324 22053
rect 22260 21993 22324 21997
rect 508 21291 572 21295
rect 508 21235 512 21291
rect 512 21235 568 21291
rect 568 21235 572 21291
rect 508 21231 572 21235
rect 630 21291 694 21295
rect 630 21235 634 21291
rect 634 21235 690 21291
rect 690 21235 694 21291
rect 630 21231 694 21235
rect 756 21291 820 21295
rect 756 21235 760 21291
rect 760 21235 816 21291
rect 816 21235 820 21291
rect 756 21231 820 21235
rect 508 21144 572 21148
rect 508 21088 512 21144
rect 512 21088 568 21144
rect 568 21088 572 21144
rect 508 21084 572 21088
rect 630 21144 694 21148
rect 630 21088 634 21144
rect 634 21088 690 21144
rect 690 21088 694 21144
rect 630 21084 694 21088
rect 756 21144 820 21148
rect 756 21088 760 21144
rect 760 21088 816 21144
rect 816 21088 820 21144
rect 756 21084 820 21088
rect 508 21007 572 21011
rect 508 20951 512 21007
rect 512 20951 568 21007
rect 568 20951 572 21007
rect 508 20947 572 20951
rect 630 21007 694 21011
rect 630 20951 634 21007
rect 634 20951 690 21007
rect 690 20951 694 21007
rect 630 20947 694 20951
rect 756 21007 820 21011
rect 756 20951 760 21007
rect 760 20951 816 21007
rect 816 20951 820 21007
rect 756 20947 820 20951
rect 507 20659 571 20663
rect 507 20603 511 20659
rect 511 20603 567 20659
rect 567 20603 571 20659
rect 507 20599 571 20603
rect 633 20659 697 20663
rect 633 20603 637 20659
rect 637 20603 693 20659
rect 693 20603 697 20659
rect 633 20599 697 20603
rect 753 20659 817 20663
rect 753 20603 757 20659
rect 757 20603 813 20659
rect 813 20603 817 20659
rect 753 20599 817 20603
rect 507 20541 571 20545
rect 507 20485 511 20541
rect 511 20485 567 20541
rect 567 20485 571 20541
rect 507 20481 571 20485
rect 633 20541 697 20545
rect 633 20485 637 20541
rect 637 20485 693 20541
rect 693 20485 697 20541
rect 633 20481 697 20485
rect 753 20541 817 20545
rect 753 20485 757 20541
rect 757 20485 813 20541
rect 813 20485 817 20541
rect 753 20481 817 20485
rect 21072 20573 21136 20577
rect 21072 20517 21076 20573
rect 21076 20517 21132 20573
rect 21132 20517 21136 20573
rect 21072 20513 21136 20517
rect 21198 20573 21262 20577
rect 21198 20517 21202 20573
rect 21202 20517 21258 20573
rect 21258 20517 21262 20573
rect 21198 20513 21262 20517
rect 21318 20573 21382 20577
rect 21318 20517 21322 20573
rect 21322 20517 21378 20573
rect 21378 20517 21382 20573
rect 21318 20513 21382 20517
rect 21072 20455 21136 20459
rect 21072 20399 21076 20455
rect 21076 20399 21132 20455
rect 21132 20399 21136 20455
rect 21072 20395 21136 20399
rect 21198 20455 21262 20459
rect 21198 20399 21202 20455
rect 21202 20399 21258 20455
rect 21258 20399 21262 20455
rect 21198 20395 21262 20399
rect 21318 20455 21382 20459
rect 21318 20399 21322 20455
rect 21322 20399 21378 20455
rect 21378 20399 21382 20455
rect 21318 20395 21382 20399
rect 507 19558 571 19562
rect 507 19502 511 19558
rect 511 19502 567 19558
rect 567 19502 571 19558
rect 507 19498 571 19502
rect 633 19558 697 19562
rect 633 19502 637 19558
rect 637 19502 693 19558
rect 693 19502 697 19558
rect 633 19498 697 19502
rect 753 19558 817 19562
rect 753 19502 757 19558
rect 757 19502 813 19558
rect 813 19502 817 19558
rect 753 19498 817 19502
rect 507 19440 571 19444
rect 507 19384 511 19440
rect 511 19384 567 19440
rect 567 19384 571 19440
rect 507 19380 571 19384
rect 633 19440 697 19444
rect 633 19384 637 19440
rect 637 19384 693 19440
rect 693 19384 697 19440
rect 633 19380 697 19384
rect 753 19440 817 19444
rect 753 19384 757 19440
rect 757 19384 813 19440
rect 813 19384 817 19440
rect 753 19380 817 19384
rect 21072 19402 21136 19406
rect 21072 19346 21076 19402
rect 21076 19346 21132 19402
rect 21132 19346 21136 19402
rect 21072 19342 21136 19346
rect 21198 19402 21262 19406
rect 21198 19346 21202 19402
rect 21202 19346 21258 19402
rect 21258 19346 21262 19402
rect 21198 19342 21262 19346
rect 21318 19402 21382 19406
rect 21318 19346 21322 19402
rect 21322 19346 21378 19402
rect 21378 19346 21382 19402
rect 21318 19342 21382 19346
rect 21072 19284 21136 19288
rect 21072 19228 21076 19284
rect 21076 19228 21132 19284
rect 21132 19228 21136 19284
rect 21072 19224 21136 19228
rect 21198 19284 21262 19288
rect 21198 19228 21202 19284
rect 21202 19228 21258 19284
rect 21258 19228 21262 19284
rect 21198 19224 21262 19228
rect 21318 19284 21382 19288
rect 21318 19228 21322 19284
rect 21322 19228 21378 19284
rect 21378 19228 21382 19284
rect 21318 19224 21382 19228
rect 508 19050 572 19054
rect 508 18994 512 19050
rect 512 18994 568 19050
rect 568 18994 572 19050
rect 508 18990 572 18994
rect 630 19050 694 19054
rect 630 18994 634 19050
rect 634 18994 690 19050
rect 690 18994 694 19050
rect 630 18990 694 18994
rect 756 19050 820 19054
rect 756 18994 760 19050
rect 760 18994 816 19050
rect 816 18994 820 19050
rect 756 18990 820 18994
rect 508 18903 572 18907
rect 508 18847 512 18903
rect 512 18847 568 18903
rect 568 18847 572 18903
rect 508 18843 572 18847
rect 630 18903 694 18907
rect 630 18847 634 18903
rect 634 18847 690 18903
rect 690 18847 694 18903
rect 630 18843 694 18847
rect 756 18903 820 18907
rect 756 18847 760 18903
rect 760 18847 816 18903
rect 816 18847 820 18903
rect 756 18843 820 18847
rect 508 18766 572 18770
rect 508 18710 512 18766
rect 512 18710 568 18766
rect 568 18710 572 18766
rect 508 18706 572 18710
rect 630 18766 694 18770
rect 630 18710 634 18766
rect 634 18710 690 18766
rect 690 18710 694 18766
rect 630 18706 694 18710
rect 756 18766 820 18770
rect 756 18710 760 18766
rect 760 18710 816 18766
rect 816 18710 820 18766
rect 756 18706 820 18710
rect 22014 18064 22078 18068
rect 22014 18008 22018 18064
rect 22018 18008 22074 18064
rect 22074 18008 22078 18064
rect 22014 18004 22078 18008
rect 22140 18064 22204 18068
rect 22140 18008 22144 18064
rect 22144 18008 22200 18064
rect 22200 18008 22204 18064
rect 22140 18004 22204 18008
rect 22260 18064 22324 18068
rect 22260 18008 22264 18064
rect 22264 18008 22320 18064
rect 22320 18008 22324 18064
rect 22260 18004 22324 18008
rect 22014 17946 22078 17950
rect 22014 17890 22018 17946
rect 22018 17890 22074 17946
rect 22074 17890 22078 17946
rect 22014 17886 22078 17890
rect 22140 17946 22204 17950
rect 22140 17890 22144 17946
rect 22144 17890 22200 17946
rect 22200 17890 22204 17946
rect 22140 17886 22204 17890
rect 22260 17946 22324 17950
rect 22260 17890 22264 17946
rect 22264 17890 22320 17946
rect 22320 17890 22324 17946
rect 22260 17886 22324 17890
rect 508 17290 572 17294
rect 508 17234 512 17290
rect 512 17234 568 17290
rect 568 17234 572 17290
rect 508 17230 572 17234
rect 630 17290 694 17294
rect 630 17234 634 17290
rect 634 17234 690 17290
rect 690 17234 694 17290
rect 630 17230 694 17234
rect 756 17290 820 17294
rect 756 17234 760 17290
rect 760 17234 816 17290
rect 816 17234 820 17290
rect 756 17230 820 17234
rect 508 17143 572 17147
rect 508 17087 512 17143
rect 512 17087 568 17143
rect 568 17087 572 17143
rect 508 17083 572 17087
rect 630 17143 694 17147
rect 630 17087 634 17143
rect 634 17087 690 17143
rect 690 17087 694 17143
rect 630 17083 694 17087
rect 756 17143 820 17147
rect 756 17087 760 17143
rect 760 17087 816 17143
rect 816 17087 820 17143
rect 756 17083 820 17087
rect 508 17006 572 17010
rect 508 16950 512 17006
rect 512 16950 568 17006
rect 568 16950 572 17006
rect 508 16946 572 16950
rect 630 17006 694 17010
rect 630 16950 634 17006
rect 634 16950 690 17006
rect 690 16950 694 17006
rect 630 16946 694 16950
rect 756 17006 820 17010
rect 756 16950 760 17006
rect 760 16950 816 17006
rect 816 16950 820 17006
rect 756 16946 820 16950
rect 507 16692 571 16696
rect 507 16636 511 16692
rect 511 16636 567 16692
rect 567 16636 571 16692
rect 507 16632 571 16636
rect 633 16692 697 16696
rect 633 16636 637 16692
rect 637 16636 693 16692
rect 693 16636 697 16692
rect 633 16632 697 16636
rect 753 16692 817 16696
rect 753 16636 757 16692
rect 757 16636 813 16692
rect 813 16636 817 16692
rect 753 16632 817 16636
rect 507 16574 571 16578
rect 507 16518 511 16574
rect 511 16518 567 16574
rect 567 16518 571 16574
rect 507 16514 571 16518
rect 633 16574 697 16578
rect 633 16518 637 16574
rect 637 16518 693 16574
rect 693 16518 697 16574
rect 633 16514 697 16518
rect 753 16574 817 16578
rect 753 16518 757 16574
rect 757 16518 813 16574
rect 813 16518 817 16574
rect 753 16514 817 16518
rect 21072 16641 21136 16645
rect 21072 16585 21076 16641
rect 21076 16585 21132 16641
rect 21132 16585 21136 16641
rect 21072 16581 21136 16585
rect 21198 16641 21262 16645
rect 21198 16585 21202 16641
rect 21202 16585 21258 16641
rect 21258 16585 21262 16641
rect 21198 16581 21262 16585
rect 21318 16641 21382 16645
rect 21318 16585 21322 16641
rect 21322 16585 21378 16641
rect 21378 16585 21382 16641
rect 21318 16581 21382 16585
rect 21072 16523 21136 16527
rect 21072 16467 21076 16523
rect 21076 16467 21132 16523
rect 21132 16467 21136 16523
rect 21072 16463 21136 16467
rect 21198 16523 21262 16527
rect 21198 16467 21202 16523
rect 21202 16467 21258 16523
rect 21258 16467 21262 16523
rect 21198 16463 21262 16467
rect 21318 16523 21382 16527
rect 21318 16467 21322 16523
rect 21322 16467 21378 16523
rect 21378 16467 21382 16523
rect 21318 16463 21382 16467
rect 507 15476 571 15480
rect 507 15420 511 15476
rect 511 15420 567 15476
rect 567 15420 571 15476
rect 507 15416 571 15420
rect 633 15476 697 15480
rect 633 15420 637 15476
rect 637 15420 693 15476
rect 693 15420 697 15476
rect 633 15416 697 15420
rect 753 15476 817 15480
rect 753 15420 757 15476
rect 757 15420 813 15476
rect 813 15420 817 15476
rect 753 15416 817 15420
rect 507 15358 571 15362
rect 507 15302 511 15358
rect 511 15302 567 15358
rect 567 15302 571 15358
rect 507 15298 571 15302
rect 633 15358 697 15362
rect 633 15302 637 15358
rect 637 15302 693 15358
rect 693 15302 697 15358
rect 633 15298 697 15302
rect 753 15358 817 15362
rect 753 15302 757 15358
rect 757 15302 813 15358
rect 813 15302 817 15358
rect 753 15298 817 15302
rect 21072 15427 21136 15431
rect 21072 15371 21076 15427
rect 21076 15371 21132 15427
rect 21132 15371 21136 15427
rect 21072 15367 21136 15371
rect 21198 15427 21262 15431
rect 21198 15371 21202 15427
rect 21202 15371 21258 15427
rect 21258 15371 21262 15427
rect 21198 15367 21262 15371
rect 21318 15427 21382 15431
rect 21318 15371 21322 15427
rect 21322 15371 21378 15427
rect 21378 15371 21382 15427
rect 21318 15367 21382 15371
rect 21072 15309 21136 15313
rect 21072 15253 21076 15309
rect 21076 15253 21132 15309
rect 21132 15253 21136 15309
rect 21072 15249 21136 15253
rect 21198 15309 21262 15313
rect 21198 15253 21202 15309
rect 21202 15253 21258 15309
rect 21258 15253 21262 15309
rect 21198 15249 21262 15253
rect 21318 15309 21382 15313
rect 21318 15253 21322 15309
rect 21322 15253 21378 15309
rect 21378 15253 21382 15309
rect 21318 15249 21382 15253
rect 508 15050 572 15054
rect 508 14994 512 15050
rect 512 14994 568 15050
rect 568 14994 572 15050
rect 508 14990 572 14994
rect 630 15050 694 15054
rect 630 14994 634 15050
rect 634 14994 690 15050
rect 690 14994 694 15050
rect 630 14990 694 14994
rect 756 15050 820 15054
rect 756 14994 760 15050
rect 760 14994 816 15050
rect 816 14994 820 15050
rect 756 14990 820 14994
rect 508 14903 572 14907
rect 508 14847 512 14903
rect 512 14847 568 14903
rect 568 14847 572 14903
rect 508 14843 572 14847
rect 630 14903 694 14907
rect 630 14847 634 14903
rect 634 14847 690 14903
rect 690 14847 694 14903
rect 630 14843 694 14847
rect 756 14903 820 14907
rect 756 14847 760 14903
rect 760 14847 816 14903
rect 816 14847 820 14903
rect 756 14843 820 14847
rect 508 14766 572 14770
rect 508 14710 512 14766
rect 512 14710 568 14766
rect 568 14710 572 14766
rect 508 14706 572 14710
rect 630 14766 694 14770
rect 630 14710 634 14766
rect 634 14710 690 14766
rect 690 14710 694 14766
rect 630 14706 694 14710
rect 756 14766 820 14770
rect 756 14710 760 14766
rect 760 14710 816 14766
rect 816 14710 820 14766
rect 756 14706 820 14710
rect 22014 14246 22078 14250
rect 22014 14190 22018 14246
rect 22018 14190 22074 14246
rect 22074 14190 22078 14246
rect 22014 14186 22078 14190
rect 22140 14246 22204 14250
rect 22140 14190 22144 14246
rect 22144 14190 22200 14246
rect 22200 14190 22204 14246
rect 22140 14186 22204 14190
rect 22260 14246 22324 14250
rect 22260 14190 22264 14246
rect 22264 14190 22320 14246
rect 22320 14190 22324 14246
rect 22260 14186 22324 14190
rect 22014 14128 22078 14132
rect 22014 14072 22018 14128
rect 22018 14072 22074 14128
rect 22074 14072 22078 14128
rect 22014 14068 22078 14072
rect 22140 14128 22204 14132
rect 22140 14072 22144 14128
rect 22144 14072 22200 14128
rect 22200 14072 22204 14128
rect 22140 14068 22204 14072
rect 22260 14128 22324 14132
rect 22260 14072 22264 14128
rect 22264 14072 22320 14128
rect 22320 14072 22324 14128
rect 22260 14068 22324 14072
rect 508 13290 572 13294
rect 508 13234 512 13290
rect 512 13234 568 13290
rect 568 13234 572 13290
rect 508 13230 572 13234
rect 630 13290 694 13294
rect 630 13234 634 13290
rect 634 13234 690 13290
rect 690 13234 694 13290
rect 630 13230 694 13234
rect 756 13290 820 13294
rect 756 13234 760 13290
rect 760 13234 816 13290
rect 816 13234 820 13290
rect 756 13230 820 13234
rect 508 13143 572 13147
rect 508 13087 512 13143
rect 512 13087 568 13143
rect 568 13087 572 13143
rect 508 13083 572 13087
rect 630 13143 694 13147
rect 630 13087 634 13143
rect 634 13087 690 13143
rect 690 13087 694 13143
rect 630 13083 694 13087
rect 756 13143 820 13147
rect 756 13087 760 13143
rect 760 13087 816 13143
rect 816 13087 820 13143
rect 756 13083 820 13087
rect 508 13006 572 13010
rect 508 12950 512 13006
rect 512 12950 568 13006
rect 568 12950 572 13006
rect 508 12946 572 12950
rect 630 13006 694 13010
rect 630 12950 634 13006
rect 634 12950 690 13006
rect 690 12950 694 13006
rect 630 12946 694 12950
rect 756 13006 820 13010
rect 756 12950 760 13006
rect 760 12950 816 13006
rect 816 12950 820 13006
rect 756 12946 820 12950
rect 507 12611 571 12615
rect 507 12555 511 12611
rect 511 12555 567 12611
rect 567 12555 571 12611
rect 507 12551 571 12555
rect 633 12611 697 12615
rect 633 12555 637 12611
rect 637 12555 693 12611
rect 693 12555 697 12611
rect 633 12551 697 12555
rect 753 12611 817 12615
rect 753 12555 757 12611
rect 757 12555 813 12611
rect 813 12555 817 12611
rect 753 12551 817 12555
rect 507 12493 571 12497
rect 507 12437 511 12493
rect 511 12437 567 12493
rect 567 12437 571 12493
rect 507 12433 571 12437
rect 633 12493 697 12497
rect 633 12437 637 12493
rect 637 12437 693 12493
rect 693 12437 697 12493
rect 633 12433 697 12437
rect 753 12493 817 12497
rect 753 12437 757 12493
rect 757 12437 813 12493
rect 813 12437 817 12493
rect 753 12433 817 12437
rect 21072 12584 21136 12588
rect 21072 12528 21076 12584
rect 21076 12528 21132 12584
rect 21132 12528 21136 12584
rect 21072 12524 21136 12528
rect 21198 12584 21262 12588
rect 21198 12528 21202 12584
rect 21202 12528 21258 12584
rect 21258 12528 21262 12584
rect 21198 12524 21262 12528
rect 21318 12584 21382 12588
rect 21318 12528 21322 12584
rect 21322 12528 21378 12584
rect 21378 12528 21382 12584
rect 21318 12524 21382 12528
rect 21072 12466 21136 12470
rect 21072 12410 21076 12466
rect 21076 12410 21132 12466
rect 21132 12410 21136 12466
rect 21072 12406 21136 12410
rect 21198 12466 21262 12470
rect 21198 12410 21202 12466
rect 21202 12410 21258 12466
rect 21258 12410 21262 12466
rect 21198 12406 21262 12410
rect 21318 12466 21382 12470
rect 21318 12410 21322 12466
rect 21322 12410 21378 12466
rect 21378 12410 21382 12466
rect 21318 12406 21382 12410
rect 507 11489 571 11493
rect 507 11433 511 11489
rect 511 11433 567 11489
rect 567 11433 571 11489
rect 507 11429 571 11433
rect 633 11489 697 11493
rect 633 11433 637 11489
rect 637 11433 693 11489
rect 693 11433 697 11489
rect 633 11429 697 11433
rect 753 11489 817 11493
rect 753 11433 757 11489
rect 757 11433 813 11489
rect 813 11433 817 11489
rect 753 11429 817 11433
rect 507 11371 571 11375
rect 507 11315 511 11371
rect 511 11315 567 11371
rect 567 11315 571 11371
rect 507 11311 571 11315
rect 633 11371 697 11375
rect 633 11315 637 11371
rect 637 11315 693 11371
rect 693 11315 697 11371
rect 633 11311 697 11315
rect 753 11371 817 11375
rect 753 11315 757 11371
rect 757 11315 813 11371
rect 813 11315 817 11371
rect 753 11311 817 11315
rect 21072 11427 21136 11431
rect 21072 11371 21076 11427
rect 21076 11371 21132 11427
rect 21132 11371 21136 11427
rect 21072 11367 21136 11371
rect 21198 11427 21262 11431
rect 21198 11371 21202 11427
rect 21202 11371 21258 11427
rect 21258 11371 21262 11427
rect 21198 11367 21262 11371
rect 21318 11427 21382 11431
rect 21318 11371 21322 11427
rect 21322 11371 21378 11427
rect 21378 11371 21382 11427
rect 21318 11367 21382 11371
rect 21072 11309 21136 11313
rect 21072 11253 21076 11309
rect 21076 11253 21132 11309
rect 21132 11253 21136 11309
rect 21072 11249 21136 11253
rect 21198 11309 21262 11313
rect 21198 11253 21202 11309
rect 21202 11253 21258 11309
rect 21258 11253 21262 11309
rect 21198 11249 21262 11253
rect 21318 11309 21382 11313
rect 21318 11253 21322 11309
rect 21322 11253 21378 11309
rect 21378 11253 21382 11309
rect 21318 11249 21382 11253
rect 508 11051 572 11055
rect 508 10995 512 11051
rect 512 10995 568 11051
rect 568 10995 572 11051
rect 508 10991 572 10995
rect 630 11051 694 11055
rect 630 10995 634 11051
rect 634 10995 690 11051
rect 690 10995 694 11051
rect 630 10991 694 10995
rect 756 11051 820 11055
rect 756 10995 760 11051
rect 760 10995 816 11051
rect 816 10995 820 11051
rect 756 10991 820 10995
rect 508 10904 572 10908
rect 508 10848 512 10904
rect 512 10848 568 10904
rect 568 10848 572 10904
rect 508 10844 572 10848
rect 630 10904 694 10908
rect 630 10848 634 10904
rect 634 10848 690 10904
rect 690 10848 694 10904
rect 630 10844 694 10848
rect 756 10904 820 10908
rect 756 10848 760 10904
rect 760 10848 816 10904
rect 816 10848 820 10904
rect 756 10844 820 10848
rect 508 10767 572 10771
rect 508 10711 512 10767
rect 512 10711 568 10767
rect 568 10711 572 10767
rect 508 10707 572 10711
rect 630 10767 694 10771
rect 630 10711 634 10767
rect 634 10711 690 10767
rect 690 10711 694 10767
rect 630 10707 694 10711
rect 756 10767 820 10771
rect 756 10711 760 10767
rect 760 10711 816 10767
rect 816 10711 820 10767
rect 756 10707 820 10711
rect 22014 10282 22078 10286
rect 22014 10226 22018 10282
rect 22018 10226 22074 10282
rect 22074 10226 22078 10282
rect 22014 10222 22078 10226
rect 22140 10282 22204 10286
rect 22140 10226 22144 10282
rect 22144 10226 22200 10282
rect 22200 10226 22204 10282
rect 22140 10222 22204 10226
rect 22260 10282 22324 10286
rect 22260 10226 22264 10282
rect 22264 10226 22320 10282
rect 22320 10226 22324 10282
rect 22260 10222 22324 10226
rect 22014 10164 22078 10168
rect 22014 10108 22018 10164
rect 22018 10108 22074 10164
rect 22074 10108 22078 10164
rect 22014 10104 22078 10108
rect 22140 10164 22204 10168
rect 22140 10108 22144 10164
rect 22144 10108 22200 10164
rect 22200 10108 22204 10164
rect 22140 10104 22204 10108
rect 22260 10164 22324 10168
rect 22260 10108 22264 10164
rect 22264 10108 22320 10164
rect 22320 10108 22324 10164
rect 22260 10104 22324 10108
rect 508 9289 572 9293
rect 508 9233 512 9289
rect 512 9233 568 9289
rect 568 9233 572 9289
rect 508 9229 572 9233
rect 630 9289 694 9293
rect 630 9233 634 9289
rect 634 9233 690 9289
rect 690 9233 694 9289
rect 630 9229 694 9233
rect 756 9289 820 9293
rect 756 9233 760 9289
rect 760 9233 816 9289
rect 816 9233 820 9289
rect 756 9229 820 9233
rect 508 9142 572 9146
rect 508 9086 512 9142
rect 512 9086 568 9142
rect 568 9086 572 9142
rect 508 9082 572 9086
rect 630 9142 694 9146
rect 630 9086 634 9142
rect 634 9086 690 9142
rect 690 9086 694 9142
rect 630 9082 694 9086
rect 756 9142 820 9146
rect 756 9086 760 9142
rect 760 9086 816 9142
rect 816 9086 820 9142
rect 756 9082 820 9086
rect 508 9005 572 9009
rect 508 8949 512 9005
rect 512 8949 568 9005
rect 568 8949 572 9005
rect 508 8945 572 8949
rect 630 9005 694 9009
rect 630 8949 634 9005
rect 634 8949 690 9005
rect 690 8949 694 9005
rect 630 8945 694 8949
rect 756 9005 820 9009
rect 756 8949 760 9005
rect 760 8949 816 9005
rect 816 8949 820 9005
rect 756 8945 820 8949
rect 507 8629 571 8633
rect 507 8573 511 8629
rect 511 8573 567 8629
rect 567 8573 571 8629
rect 507 8569 571 8573
rect 633 8629 697 8633
rect 633 8573 637 8629
rect 637 8573 693 8629
rect 693 8573 697 8629
rect 633 8569 697 8573
rect 753 8629 817 8633
rect 753 8573 757 8629
rect 757 8573 813 8629
rect 813 8573 817 8629
rect 753 8569 817 8573
rect 507 8511 571 8515
rect 507 8455 511 8511
rect 511 8455 567 8511
rect 567 8455 571 8511
rect 507 8451 571 8455
rect 633 8511 697 8515
rect 633 8455 637 8511
rect 637 8455 693 8511
rect 693 8455 697 8511
rect 633 8451 697 8455
rect 753 8511 817 8515
rect 753 8455 757 8511
rect 757 8455 813 8511
rect 813 8455 817 8511
rect 753 8451 817 8455
rect 21072 8584 21136 8588
rect 21072 8528 21076 8584
rect 21076 8528 21132 8584
rect 21132 8528 21136 8584
rect 21072 8524 21136 8528
rect 21198 8584 21262 8588
rect 21198 8528 21202 8584
rect 21202 8528 21258 8584
rect 21258 8528 21262 8584
rect 21198 8524 21262 8528
rect 21318 8584 21382 8588
rect 21318 8528 21322 8584
rect 21322 8528 21378 8584
rect 21378 8528 21382 8584
rect 21318 8524 21382 8528
rect 21072 8466 21136 8470
rect 21072 8410 21076 8466
rect 21076 8410 21132 8466
rect 21132 8410 21136 8466
rect 21072 8406 21136 8410
rect 21198 8466 21262 8470
rect 21198 8410 21202 8466
rect 21202 8410 21258 8466
rect 21258 8410 21262 8466
rect 21198 8406 21262 8410
rect 21318 8466 21382 8470
rect 21318 8410 21322 8466
rect 21322 8410 21378 8466
rect 21378 8410 21382 8466
rect 21318 8406 21382 8410
rect 507 7518 571 7522
rect 507 7462 511 7518
rect 511 7462 567 7518
rect 567 7462 571 7518
rect 507 7458 571 7462
rect 633 7518 697 7522
rect 633 7462 637 7518
rect 637 7462 693 7518
rect 693 7462 697 7518
rect 633 7458 697 7462
rect 753 7518 817 7522
rect 753 7462 757 7518
rect 757 7462 813 7518
rect 813 7462 817 7518
rect 753 7458 817 7462
rect 507 7400 571 7404
rect 507 7344 511 7400
rect 511 7344 567 7400
rect 567 7344 571 7400
rect 507 7340 571 7344
rect 633 7400 697 7404
rect 633 7344 637 7400
rect 637 7344 693 7400
rect 693 7344 697 7400
rect 633 7340 697 7344
rect 753 7400 817 7404
rect 753 7344 757 7400
rect 757 7344 813 7400
rect 813 7344 817 7400
rect 753 7340 817 7344
rect 21072 7427 21136 7431
rect 21072 7371 21076 7427
rect 21076 7371 21132 7427
rect 21132 7371 21136 7427
rect 21072 7367 21136 7371
rect 21198 7427 21262 7431
rect 21198 7371 21202 7427
rect 21202 7371 21258 7427
rect 21258 7371 21262 7427
rect 21198 7367 21262 7371
rect 21318 7427 21382 7431
rect 21318 7371 21322 7427
rect 21322 7371 21378 7427
rect 21378 7371 21382 7427
rect 21318 7367 21382 7371
rect 21072 7309 21136 7313
rect 21072 7253 21076 7309
rect 21076 7253 21132 7309
rect 21132 7253 21136 7309
rect 21072 7249 21136 7253
rect 21198 7309 21262 7313
rect 21198 7253 21202 7309
rect 21202 7253 21258 7309
rect 21258 7253 21262 7309
rect 21198 7249 21262 7253
rect 21318 7309 21382 7313
rect 21318 7253 21322 7309
rect 21322 7253 21378 7309
rect 21378 7253 21382 7309
rect 21318 7249 21382 7253
rect 508 7051 572 7055
rect 508 6995 512 7051
rect 512 6995 568 7051
rect 568 6995 572 7051
rect 508 6991 572 6995
rect 630 7051 694 7055
rect 630 6995 634 7051
rect 634 6995 690 7051
rect 690 6995 694 7051
rect 630 6991 694 6995
rect 756 7051 820 7055
rect 756 6995 760 7051
rect 760 6995 816 7051
rect 816 6995 820 7051
rect 756 6991 820 6995
rect 508 6904 572 6908
rect 508 6848 512 6904
rect 512 6848 568 6904
rect 568 6848 572 6904
rect 508 6844 572 6848
rect 630 6904 694 6908
rect 630 6848 634 6904
rect 634 6848 690 6904
rect 690 6848 694 6904
rect 630 6844 694 6848
rect 756 6904 820 6908
rect 756 6848 760 6904
rect 760 6848 816 6904
rect 816 6848 820 6904
rect 756 6844 820 6848
rect 508 6767 572 6771
rect 508 6711 512 6767
rect 512 6711 568 6767
rect 568 6711 572 6767
rect 508 6707 572 6711
rect 630 6767 694 6771
rect 630 6711 634 6767
rect 634 6711 690 6767
rect 690 6711 694 6767
rect 630 6707 694 6711
rect 756 6767 820 6771
rect 756 6711 760 6767
rect 760 6711 816 6767
rect 816 6711 820 6767
rect 756 6707 820 6711
rect 22014 6270 22078 6274
rect 22014 6214 22018 6270
rect 22018 6214 22074 6270
rect 22074 6214 22078 6270
rect 22014 6210 22078 6214
rect 22140 6270 22204 6274
rect 22140 6214 22144 6270
rect 22144 6214 22200 6270
rect 22200 6214 22204 6270
rect 22140 6210 22204 6214
rect 22260 6270 22324 6274
rect 22260 6214 22264 6270
rect 22264 6214 22320 6270
rect 22320 6214 22324 6270
rect 22260 6210 22324 6214
rect 22014 6152 22078 6156
rect 22014 6096 22018 6152
rect 22018 6096 22074 6152
rect 22074 6096 22078 6152
rect 22014 6092 22078 6096
rect 22140 6152 22204 6156
rect 22140 6096 22144 6152
rect 22144 6096 22200 6152
rect 22200 6096 22204 6152
rect 22140 6092 22204 6096
rect 22260 6152 22324 6156
rect 22260 6096 22264 6152
rect 22264 6096 22320 6152
rect 22320 6096 22324 6152
rect 22260 6092 22324 6096
rect 508 5290 572 5294
rect 508 5234 512 5290
rect 512 5234 568 5290
rect 568 5234 572 5290
rect 508 5230 572 5234
rect 630 5290 694 5294
rect 630 5234 634 5290
rect 634 5234 690 5290
rect 690 5234 694 5290
rect 630 5230 694 5234
rect 756 5290 820 5294
rect 756 5234 760 5290
rect 760 5234 816 5290
rect 816 5234 820 5290
rect 756 5230 820 5234
rect 508 5143 572 5147
rect 508 5087 512 5143
rect 512 5087 568 5143
rect 568 5087 572 5143
rect 508 5083 572 5087
rect 630 5143 694 5147
rect 630 5087 634 5143
rect 634 5087 690 5143
rect 690 5087 694 5143
rect 630 5083 694 5087
rect 756 5143 820 5147
rect 756 5087 760 5143
rect 760 5087 816 5143
rect 816 5087 820 5143
rect 756 5083 820 5087
rect 508 5006 572 5010
rect 508 4950 512 5006
rect 512 4950 568 5006
rect 568 4950 572 5006
rect 508 4946 572 4950
rect 630 5006 694 5010
rect 630 4950 634 5006
rect 634 4950 690 5006
rect 690 4950 694 5006
rect 630 4946 694 4950
rect 756 5006 820 5010
rect 756 4950 760 5006
rect 760 4950 816 5006
rect 816 4950 820 5006
rect 756 4946 820 4950
rect 507 4695 571 4699
rect 507 4639 511 4695
rect 511 4639 567 4695
rect 567 4639 571 4695
rect 507 4635 571 4639
rect 633 4695 697 4699
rect 633 4639 637 4695
rect 637 4639 693 4695
rect 693 4639 697 4695
rect 633 4635 697 4639
rect 753 4695 817 4699
rect 753 4639 757 4695
rect 757 4639 813 4695
rect 813 4639 817 4695
rect 753 4635 817 4639
rect 507 4577 571 4581
rect 507 4521 511 4577
rect 511 4521 567 4577
rect 567 4521 571 4577
rect 507 4517 571 4521
rect 633 4577 697 4581
rect 633 4521 637 4577
rect 637 4521 693 4577
rect 693 4521 697 4577
rect 633 4517 697 4521
rect 753 4577 817 4581
rect 753 4521 757 4577
rect 757 4521 813 4577
rect 813 4521 817 4577
rect 753 4517 817 4521
rect 21072 4584 21136 4588
rect 21072 4528 21076 4584
rect 21076 4528 21132 4584
rect 21132 4528 21136 4584
rect 21072 4524 21136 4528
rect 21198 4584 21262 4588
rect 21198 4528 21202 4584
rect 21202 4528 21258 4584
rect 21258 4528 21262 4584
rect 21198 4524 21262 4528
rect 21318 4584 21382 4588
rect 21318 4528 21322 4584
rect 21322 4528 21378 4584
rect 21378 4528 21382 4584
rect 21318 4524 21382 4528
rect 21072 4466 21136 4470
rect 21072 4410 21076 4466
rect 21076 4410 21132 4466
rect 21132 4410 21136 4466
rect 21072 4406 21136 4410
rect 21198 4466 21262 4470
rect 21198 4410 21202 4466
rect 21202 4410 21258 4466
rect 21258 4410 21262 4466
rect 21198 4406 21262 4410
rect 21318 4466 21382 4470
rect 21318 4410 21322 4466
rect 21322 4410 21378 4466
rect 21378 4410 21382 4466
rect 21318 4406 21382 4410
rect 507 3518 571 3522
rect 507 3462 511 3518
rect 511 3462 567 3518
rect 567 3462 571 3518
rect 507 3458 571 3462
rect 633 3518 697 3522
rect 633 3462 637 3518
rect 637 3462 693 3518
rect 693 3462 697 3518
rect 633 3458 697 3462
rect 753 3518 817 3522
rect 753 3462 757 3518
rect 757 3462 813 3518
rect 813 3462 817 3518
rect 753 3458 817 3462
rect 507 3400 571 3404
rect 507 3344 511 3400
rect 511 3344 567 3400
rect 567 3344 571 3400
rect 507 3340 571 3344
rect 633 3400 697 3404
rect 633 3344 637 3400
rect 637 3344 693 3400
rect 693 3344 697 3400
rect 633 3340 697 3344
rect 753 3400 817 3404
rect 753 3344 757 3400
rect 757 3344 813 3400
rect 813 3344 817 3400
rect 753 3340 817 3344
rect 21072 3427 21136 3431
rect 21072 3371 21076 3427
rect 21076 3371 21132 3427
rect 21132 3371 21136 3427
rect 21072 3367 21136 3371
rect 21198 3427 21262 3431
rect 21198 3371 21202 3427
rect 21202 3371 21258 3427
rect 21258 3371 21262 3427
rect 21198 3367 21262 3371
rect 21318 3427 21382 3431
rect 21318 3371 21322 3427
rect 21322 3371 21378 3427
rect 21378 3371 21382 3427
rect 21318 3367 21382 3371
rect 21072 3309 21136 3313
rect 21072 3253 21076 3309
rect 21076 3253 21132 3309
rect 21132 3253 21136 3309
rect 21072 3249 21136 3253
rect 21198 3309 21262 3313
rect 21198 3253 21202 3309
rect 21202 3253 21258 3309
rect 21258 3253 21262 3309
rect 21198 3249 21262 3253
rect 21318 3309 21382 3313
rect 21318 3253 21322 3309
rect 21322 3253 21378 3309
rect 21378 3253 21382 3309
rect 21318 3249 21382 3253
rect 508 3051 572 3055
rect 508 2995 512 3051
rect 512 2995 568 3051
rect 568 2995 572 3051
rect 508 2991 572 2995
rect 630 3051 694 3055
rect 630 2995 634 3051
rect 634 2995 690 3051
rect 690 2995 694 3051
rect 630 2991 694 2995
rect 756 3051 820 3055
rect 756 2995 760 3051
rect 760 2995 816 3051
rect 816 2995 820 3051
rect 756 2991 820 2995
rect 508 2904 572 2908
rect 508 2848 512 2904
rect 512 2848 568 2904
rect 568 2848 572 2904
rect 508 2844 572 2848
rect 630 2904 694 2908
rect 630 2848 634 2904
rect 634 2848 690 2904
rect 690 2848 694 2904
rect 630 2844 694 2848
rect 756 2904 820 2908
rect 756 2848 760 2904
rect 760 2848 816 2904
rect 816 2848 820 2904
rect 756 2844 820 2848
rect 508 2767 572 2771
rect 508 2711 512 2767
rect 512 2711 568 2767
rect 568 2711 572 2767
rect 508 2707 572 2711
rect 630 2767 694 2771
rect 630 2711 634 2767
rect 634 2711 690 2767
rect 690 2711 694 2767
rect 630 2707 694 2711
rect 756 2767 820 2771
rect 756 2711 760 2767
rect 760 2711 816 2767
rect 816 2711 820 2767
rect 756 2707 820 2711
rect 22014 2270 22078 2274
rect 22014 2214 22018 2270
rect 22018 2214 22074 2270
rect 22074 2214 22078 2270
rect 22014 2210 22078 2214
rect 22140 2270 22204 2274
rect 22140 2214 22144 2270
rect 22144 2214 22200 2270
rect 22200 2214 22204 2270
rect 22140 2210 22204 2214
rect 22260 2270 22324 2274
rect 22260 2214 22264 2270
rect 22264 2214 22320 2270
rect 22320 2214 22324 2270
rect 22260 2210 22324 2214
rect 22014 2152 22078 2156
rect 22014 2096 22018 2152
rect 22018 2096 22074 2152
rect 22074 2096 22078 2152
rect 22014 2092 22078 2096
rect 22140 2152 22204 2156
rect 22140 2096 22144 2152
rect 22144 2096 22200 2152
rect 22200 2096 22204 2152
rect 22140 2092 22204 2096
rect 22260 2152 22324 2156
rect 22260 2096 22264 2152
rect 22264 2096 22320 2152
rect 22320 2096 22324 2152
rect 22260 2092 22324 2096
rect 508 1290 572 1294
rect 508 1234 512 1290
rect 512 1234 568 1290
rect 568 1234 572 1290
rect 508 1230 572 1234
rect 630 1290 694 1294
rect 630 1234 634 1290
rect 634 1234 690 1290
rect 690 1234 694 1290
rect 630 1230 694 1234
rect 756 1290 820 1294
rect 756 1234 760 1290
rect 760 1234 816 1290
rect 816 1234 820 1290
rect 756 1230 820 1234
rect 508 1143 572 1147
rect 508 1087 512 1143
rect 512 1087 568 1143
rect 568 1087 572 1143
rect 508 1083 572 1087
rect 630 1143 694 1147
rect 630 1087 634 1143
rect 634 1087 690 1143
rect 690 1087 694 1143
rect 630 1083 694 1087
rect 756 1143 820 1147
rect 756 1087 760 1143
rect 760 1087 816 1143
rect 816 1087 820 1143
rect 756 1083 820 1087
rect 508 1006 572 1010
rect 508 950 512 1006
rect 512 950 568 1006
rect 568 950 572 1006
rect 508 946 572 950
rect 630 1006 694 1010
rect 630 950 634 1006
rect 634 950 690 1006
rect 690 950 694 1006
rect 630 946 694 950
rect 756 1006 820 1010
rect 756 950 760 1006
rect 760 950 816 1006
rect 816 950 820 1006
rect 756 946 820 950
rect 507 695 571 699
rect 507 639 511 695
rect 511 639 567 695
rect 567 639 571 695
rect 507 635 571 639
rect 633 695 697 699
rect 633 639 637 695
rect 637 639 693 695
rect 693 639 697 695
rect 633 635 697 639
rect 753 695 817 699
rect 753 639 757 695
rect 757 639 813 695
rect 813 639 817 695
rect 753 635 817 639
rect 507 577 571 581
rect 507 521 511 577
rect 511 521 567 577
rect 567 521 571 577
rect 507 517 571 521
rect 633 577 697 581
rect 633 521 637 577
rect 637 521 693 577
rect 693 521 697 577
rect 633 517 697 521
rect 753 577 817 581
rect 753 521 757 577
rect 757 521 813 577
rect 813 521 817 577
rect 753 517 817 521
rect 21072 584 21136 588
rect 21072 528 21076 584
rect 21076 528 21132 584
rect 21132 528 21136 584
rect 21072 524 21136 528
rect 21198 584 21262 588
rect 21198 528 21202 584
rect 21202 528 21258 584
rect 21258 528 21262 584
rect 21198 524 21262 528
rect 21318 584 21382 588
rect 21318 528 21322 584
rect 21322 528 21378 584
rect 21378 528 21382 584
rect 21318 524 21382 528
rect 21072 466 21136 470
rect 21072 410 21076 466
rect 21076 410 21132 466
rect 21132 410 21136 466
rect 21072 406 21136 410
rect 21198 466 21262 470
rect 21198 410 21202 466
rect 21202 410 21258 466
rect 21258 410 21262 466
rect 21198 406 21262 410
rect 21318 466 21382 470
rect 21318 410 21322 466
rect 21322 410 21378 466
rect 21378 410 21382 466
rect 21318 406 21382 410
<< metal4 >>
rect 0 39733 400 76000
rect 0 39669 39 39733
rect 103 39669 164 39733
rect 228 39669 290 39733
rect 354 39669 400 39733
rect 0 39627 400 39669
rect 0 39563 39 39627
rect 103 39563 164 39627
rect 228 39563 290 39627
rect 354 39563 400 39627
rect 0 38579 400 39563
rect 0 38515 25 38579
rect 89 38515 139 38579
rect 203 38515 253 38579
rect 317 38515 400 38579
rect 0 37491 400 38515
rect 0 37427 25 37491
rect 89 37427 139 37491
rect 203 37427 253 37491
rect 317 37427 400 37491
rect 0 0 400 37427
rect 463 75477 863 76000
rect 21028 75517 21428 76000
rect 21026 75486 21428 75517
rect 463 75446 864 75477
rect 463 75382 507 75446
rect 571 75382 633 75446
rect 697 75382 753 75446
rect 817 75382 864 75446
rect 463 75328 864 75382
rect 463 75264 507 75328
rect 571 75264 633 75328
rect 697 75264 753 75328
rect 817 75264 864 75328
rect 463 75222 864 75264
rect 21026 75422 21072 75486
rect 21136 75422 21198 75486
rect 21262 75422 21318 75486
rect 21382 75422 21428 75486
rect 21026 75368 21428 75422
rect 21026 75304 21072 75368
rect 21136 75304 21198 75368
rect 21262 75304 21318 75368
rect 21382 75304 21428 75368
rect 21026 75262 21428 75304
rect 463 75054 863 75222
rect 463 74990 508 75054
rect 572 74990 630 75054
rect 694 74990 756 75054
rect 820 74990 863 75054
rect 463 74907 863 74990
rect 463 74843 508 74907
rect 572 74843 630 74907
rect 694 74843 756 74907
rect 820 74843 863 74907
rect 463 74770 863 74843
rect 463 74706 508 74770
rect 572 74706 630 74770
rect 694 74706 756 74770
rect 820 74706 863 74770
rect 463 73294 863 74706
rect 463 73230 508 73294
rect 572 73230 630 73294
rect 694 73230 756 73294
rect 820 73230 863 73294
rect 463 73147 863 73230
rect 463 73083 508 73147
rect 572 73083 630 73147
rect 694 73083 756 73147
rect 820 73083 863 73147
rect 463 73010 863 73083
rect 463 72946 508 73010
rect 572 72946 630 73010
rect 694 72946 756 73010
rect 820 72946 863 73010
rect 463 72804 863 72946
rect 463 72773 864 72804
rect 463 72709 507 72773
rect 571 72709 633 72773
rect 697 72709 753 72773
rect 817 72709 864 72773
rect 463 72655 864 72709
rect 463 72591 507 72655
rect 571 72591 633 72655
rect 697 72591 753 72655
rect 817 72591 864 72655
rect 463 72549 864 72591
rect 21028 72689 21428 75262
rect 21028 72625 21072 72689
rect 21136 72625 21198 72689
rect 21262 72625 21318 72689
rect 21382 72625 21428 72689
rect 21028 72571 21428 72625
rect 463 71477 863 72549
rect 21028 72507 21072 72571
rect 21136 72507 21198 72571
rect 21262 72507 21318 72571
rect 21382 72507 21428 72571
rect 21028 71517 21428 72507
rect 21026 71486 21428 71517
rect 463 71446 864 71477
rect 463 71382 507 71446
rect 571 71382 633 71446
rect 697 71382 753 71446
rect 817 71382 864 71446
rect 463 71328 864 71382
rect 463 71264 507 71328
rect 571 71264 633 71328
rect 697 71264 753 71328
rect 817 71264 864 71328
rect 463 71222 864 71264
rect 21026 71422 21072 71486
rect 21136 71422 21198 71486
rect 21262 71422 21318 71486
rect 21382 71422 21428 71486
rect 21026 71368 21428 71422
rect 21026 71304 21072 71368
rect 21136 71304 21198 71368
rect 21262 71304 21318 71368
rect 21382 71304 21428 71368
rect 21026 71262 21428 71304
rect 463 71054 863 71222
rect 463 70990 508 71054
rect 572 70990 630 71054
rect 694 70990 756 71054
rect 820 70990 863 71054
rect 463 70907 863 70990
rect 463 70843 508 70907
rect 572 70843 630 70907
rect 694 70843 756 70907
rect 820 70843 863 70907
rect 463 70770 863 70843
rect 463 70706 508 70770
rect 572 70706 630 70770
rect 694 70706 756 70770
rect 820 70706 863 70770
rect 463 69294 863 70706
rect 463 69230 508 69294
rect 572 69230 630 69294
rect 694 69230 756 69294
rect 820 69230 863 69294
rect 463 69147 863 69230
rect 463 69083 508 69147
rect 572 69083 630 69147
rect 694 69083 756 69147
rect 820 69083 863 69147
rect 463 69010 863 69083
rect 463 68946 508 69010
rect 572 68946 630 69010
rect 694 68946 756 69010
rect 820 68946 863 69010
rect 463 68804 863 68946
rect 463 68773 864 68804
rect 463 68709 507 68773
rect 571 68709 633 68773
rect 697 68709 753 68773
rect 817 68709 864 68773
rect 463 68655 864 68709
rect 463 68591 507 68655
rect 571 68591 633 68655
rect 697 68591 753 68655
rect 817 68591 864 68655
rect 463 68549 864 68591
rect 21028 68689 21428 71262
rect 21028 68625 21072 68689
rect 21136 68625 21198 68689
rect 21262 68625 21318 68689
rect 21382 68625 21428 68689
rect 21028 68571 21428 68625
rect 463 67475 863 68549
rect 21028 68507 21072 68571
rect 21136 68507 21198 68571
rect 21262 68507 21318 68571
rect 21382 68507 21428 68571
rect 21028 67517 21428 68507
rect 21026 67486 21428 67517
rect 463 67444 864 67475
rect 463 67380 507 67444
rect 571 67380 633 67444
rect 697 67380 753 67444
rect 817 67380 864 67444
rect 463 67326 864 67380
rect 463 67262 507 67326
rect 571 67262 633 67326
rect 697 67262 753 67326
rect 817 67262 864 67326
rect 21026 67422 21072 67486
rect 21136 67422 21198 67486
rect 21262 67422 21318 67486
rect 21382 67422 21428 67486
rect 21026 67368 21428 67422
rect 21026 67304 21072 67368
rect 21136 67304 21198 67368
rect 21262 67304 21318 67368
rect 21382 67304 21428 67368
rect 21026 67262 21428 67304
rect 463 67220 864 67262
rect 463 67054 863 67220
rect 463 66990 508 67054
rect 572 66990 630 67054
rect 694 66990 756 67054
rect 820 66990 863 67054
rect 463 66907 863 66990
rect 463 66843 508 66907
rect 572 66843 630 66907
rect 694 66843 756 66907
rect 820 66843 863 66907
rect 463 66770 863 66843
rect 463 66706 508 66770
rect 572 66706 630 66770
rect 694 66706 756 66770
rect 820 66706 863 66770
rect 463 65295 863 66706
rect 463 65231 508 65295
rect 572 65231 630 65295
rect 694 65231 756 65295
rect 820 65231 863 65295
rect 463 65148 863 65231
rect 463 65084 508 65148
rect 572 65084 630 65148
rect 694 65084 756 65148
rect 820 65084 863 65148
rect 463 65011 863 65084
rect 463 64947 508 65011
rect 572 64947 630 65011
rect 694 64947 756 65011
rect 820 64947 863 65011
rect 463 64735 863 64947
rect 463 64704 864 64735
rect 463 64640 507 64704
rect 571 64640 633 64704
rect 697 64640 753 64704
rect 817 64640 864 64704
rect 463 64586 864 64640
rect 463 64522 507 64586
rect 571 64522 633 64586
rect 697 64522 753 64586
rect 817 64522 864 64586
rect 463 64480 864 64522
rect 21028 64689 21428 67262
rect 21028 64625 21072 64689
rect 21136 64625 21198 64689
rect 21262 64625 21318 64689
rect 21382 64625 21428 64689
rect 21028 64571 21428 64625
rect 21028 64507 21072 64571
rect 21136 64507 21198 64571
rect 21262 64507 21318 64571
rect 21382 64507 21428 64571
rect 463 63557 863 64480
rect 463 63526 864 63557
rect 463 63462 507 63526
rect 571 63462 633 63526
rect 697 63462 753 63526
rect 817 63462 864 63526
rect 21028 63517 21428 64507
rect 463 63408 864 63462
rect 463 63344 507 63408
rect 571 63344 633 63408
rect 697 63344 753 63408
rect 817 63344 864 63408
rect 463 63302 864 63344
rect 21026 63486 21428 63517
rect 21026 63422 21072 63486
rect 21136 63422 21198 63486
rect 21262 63422 21318 63486
rect 21382 63422 21428 63486
rect 21026 63368 21428 63422
rect 21026 63304 21072 63368
rect 21136 63304 21198 63368
rect 21262 63304 21318 63368
rect 21382 63304 21428 63368
rect 463 63109 863 63302
rect 21026 63262 21428 63304
rect 463 63054 864 63109
rect 463 62990 508 63054
rect 572 62990 630 63054
rect 694 62990 756 63054
rect 820 62990 864 63054
rect 463 62907 864 62990
rect 463 62843 508 62907
rect 572 62843 630 62907
rect 694 62843 756 62907
rect 820 62843 864 62907
rect 463 62770 864 62843
rect 463 62706 508 62770
rect 572 62706 630 62770
rect 694 62706 756 62770
rect 820 62706 864 62770
rect 463 62650 864 62706
rect 463 61295 863 62650
rect 463 61231 508 61295
rect 572 61231 630 61295
rect 694 61231 756 61295
rect 820 61231 863 61295
rect 463 61148 863 61231
rect 463 61084 508 61148
rect 572 61084 630 61148
rect 694 61084 756 61148
rect 820 61084 863 61148
rect 463 61011 863 61084
rect 463 60947 508 61011
rect 572 60947 630 61011
rect 694 60947 756 61011
rect 820 60947 863 61011
rect 463 60709 863 60947
rect 463 60678 866 60709
rect 463 60614 507 60678
rect 571 60614 633 60678
rect 697 60614 753 60678
rect 817 60614 866 60678
rect 463 60560 866 60614
rect 463 60496 507 60560
rect 571 60496 633 60560
rect 697 60496 753 60560
rect 817 60496 866 60560
rect 463 60454 866 60496
rect 21028 60689 21428 63262
rect 21028 60625 21072 60689
rect 21136 60625 21198 60689
rect 21262 60625 21318 60689
rect 21382 60625 21428 60689
rect 21028 60571 21428 60625
rect 21028 60507 21072 60571
rect 21136 60507 21198 60571
rect 21262 60507 21318 60571
rect 21382 60507 21428 60571
rect 463 59506 863 60454
rect 21028 59571 21428 60507
rect 21027 59540 21428 59571
rect 463 59475 864 59506
rect 463 59411 507 59475
rect 571 59411 633 59475
rect 697 59411 753 59475
rect 817 59411 864 59475
rect 463 59357 864 59411
rect 463 59293 507 59357
rect 571 59293 633 59357
rect 697 59293 753 59357
rect 817 59293 864 59357
rect 21027 59476 21072 59540
rect 21136 59476 21198 59540
rect 21262 59476 21318 59540
rect 21382 59476 21428 59540
rect 21027 59422 21428 59476
rect 21027 59358 21072 59422
rect 21136 59358 21198 59422
rect 21262 59358 21318 59422
rect 21382 59358 21428 59422
rect 21027 59316 21428 59358
rect 463 59251 864 59293
rect 463 59109 863 59251
rect 463 59054 864 59109
rect 463 58990 508 59054
rect 572 58990 630 59054
rect 694 58990 756 59054
rect 820 58990 864 59054
rect 463 58907 864 58990
rect 463 58843 508 58907
rect 572 58843 630 58907
rect 694 58843 756 58907
rect 820 58843 864 58907
rect 463 58770 864 58843
rect 463 58706 508 58770
rect 572 58706 630 58770
rect 694 58706 756 58770
rect 820 58706 864 58770
rect 463 58650 864 58706
rect 463 57293 863 58650
rect 463 57229 508 57293
rect 572 57229 630 57293
rect 694 57229 756 57293
rect 820 57229 863 57293
rect 463 57146 863 57229
rect 463 57082 508 57146
rect 572 57082 630 57146
rect 694 57082 756 57146
rect 820 57082 863 57146
rect 463 57009 863 57082
rect 463 56945 508 57009
rect 572 56945 630 57009
rect 694 56945 756 57009
rect 820 56945 863 57009
rect 463 56729 863 56945
rect 463 56698 864 56729
rect 463 56634 507 56698
rect 571 56634 633 56698
rect 697 56634 753 56698
rect 817 56634 864 56698
rect 463 56580 864 56634
rect 463 56516 507 56580
rect 571 56516 633 56580
rect 697 56516 753 56580
rect 817 56516 864 56580
rect 463 56474 864 56516
rect 21028 56624 21428 59316
rect 21028 56560 21072 56624
rect 21136 56560 21198 56624
rect 21262 56560 21318 56624
rect 21382 56560 21428 56624
rect 21028 56506 21428 56560
rect 463 55522 863 56474
rect 21028 56442 21072 56506
rect 21136 56442 21198 56506
rect 21262 56442 21318 56506
rect 21382 56442 21428 56506
rect 463 55491 866 55522
rect 463 55427 507 55491
rect 571 55427 633 55491
rect 697 55427 753 55491
rect 817 55427 866 55491
rect 21028 55472 21428 56442
rect 463 55373 866 55427
rect 463 55309 507 55373
rect 571 55309 633 55373
rect 697 55309 753 55373
rect 817 55309 866 55373
rect 463 55267 866 55309
rect 21027 55441 21428 55472
rect 21027 55377 21072 55441
rect 21136 55377 21198 55441
rect 21262 55377 21318 55441
rect 21382 55377 21428 55441
rect 21027 55323 21428 55377
rect 463 55054 863 55267
rect 21027 55259 21072 55323
rect 21136 55259 21198 55323
rect 21262 55259 21318 55323
rect 21382 55259 21428 55323
rect 21027 55217 21428 55259
rect 463 54990 508 55054
rect 572 54990 630 55054
rect 694 54990 756 55054
rect 820 54990 863 55054
rect 463 54907 863 54990
rect 463 54843 508 54907
rect 572 54843 630 54907
rect 694 54843 756 54907
rect 820 54843 863 54907
rect 463 54770 863 54843
rect 463 54706 508 54770
rect 572 54706 630 54770
rect 694 54706 756 54770
rect 820 54706 863 54770
rect 463 53295 863 54706
rect 463 53231 508 53295
rect 572 53231 630 53295
rect 694 53231 756 53295
rect 820 53231 863 53295
rect 463 53148 863 53231
rect 463 53084 508 53148
rect 572 53084 630 53148
rect 694 53084 756 53148
rect 820 53084 863 53148
rect 463 53011 863 53084
rect 463 52947 508 53011
rect 572 52947 630 53011
rect 694 52947 756 53011
rect 820 52947 863 53011
rect 463 52756 863 52947
rect 463 52725 864 52756
rect 463 52661 507 52725
rect 571 52661 633 52725
rect 697 52661 753 52725
rect 817 52661 864 52725
rect 463 52607 864 52661
rect 463 52543 507 52607
rect 571 52543 633 52607
rect 697 52543 753 52607
rect 817 52543 864 52607
rect 463 52501 864 52543
rect 21028 52569 21428 55217
rect 21028 52505 21072 52569
rect 21136 52505 21198 52569
rect 21262 52505 21318 52569
rect 21382 52505 21428 52569
rect 463 51569 863 52501
rect 21028 52451 21428 52505
rect 21028 52387 21072 52451
rect 21136 52387 21198 52451
rect 21262 52387 21318 52451
rect 21382 52387 21428 52451
rect 463 51538 864 51569
rect 463 51474 507 51538
rect 571 51474 633 51538
rect 697 51474 753 51538
rect 817 51474 864 51538
rect 463 51420 864 51474
rect 463 51356 507 51420
rect 571 51356 633 51420
rect 697 51356 753 51420
rect 817 51356 864 51420
rect 463 51314 864 51356
rect 21028 51434 21428 52387
rect 21028 51370 21072 51434
rect 21136 51370 21198 51434
rect 21262 51370 21318 51434
rect 21382 51370 21428 51434
rect 21028 51316 21428 51370
rect 463 51054 863 51314
rect 463 50990 508 51054
rect 572 50990 630 51054
rect 694 50990 756 51054
rect 820 50990 863 51054
rect 463 50907 863 50990
rect 463 50843 508 50907
rect 572 50843 630 50907
rect 694 50843 756 50907
rect 820 50843 863 50907
rect 463 50770 863 50843
rect 463 50706 508 50770
rect 572 50706 630 50770
rect 694 50706 756 50770
rect 820 50706 863 50770
rect 463 49295 863 50706
rect 463 49231 508 49295
rect 572 49231 630 49295
rect 694 49231 756 49295
rect 820 49231 863 49295
rect 463 49148 863 49231
rect 463 49084 508 49148
rect 572 49084 630 49148
rect 694 49084 756 49148
rect 820 49084 863 49148
rect 463 49011 863 49084
rect 463 48947 508 49011
rect 572 48947 630 49011
rect 694 48947 756 49011
rect 820 48947 863 49011
rect 463 48747 863 48947
rect 21028 51252 21072 51316
rect 21136 51252 21198 51316
rect 21262 51252 21318 51316
rect 21382 51252 21428 51316
rect 463 48716 864 48747
rect 463 48652 507 48716
rect 571 48652 633 48716
rect 697 48652 753 48716
rect 817 48652 864 48716
rect 463 48598 864 48652
rect 463 48534 507 48598
rect 571 48534 633 48598
rect 697 48534 753 48598
rect 817 48534 864 48598
rect 463 48492 864 48534
rect 21028 48675 21428 51252
rect 21028 48611 21072 48675
rect 21136 48611 21198 48675
rect 21262 48611 21318 48675
rect 21382 48611 21428 48675
rect 21028 48557 21428 48611
rect 21028 48493 21072 48557
rect 21136 48493 21198 48557
rect 21262 48493 21318 48557
rect 21382 48493 21428 48557
rect 463 47594 863 48492
rect 463 47563 864 47594
rect 463 47499 507 47563
rect 571 47499 633 47563
rect 697 47499 753 47563
rect 817 47499 864 47563
rect 463 47445 864 47499
rect 463 47381 507 47445
rect 571 47381 633 47445
rect 697 47381 753 47445
rect 817 47381 864 47445
rect 463 47339 864 47381
rect 21028 47522 21428 48493
rect 21028 47458 21072 47522
rect 21136 47458 21198 47522
rect 21262 47458 21318 47522
rect 21382 47458 21428 47522
rect 21028 47404 21428 47458
rect 21028 47340 21072 47404
rect 21136 47340 21198 47404
rect 21262 47340 21318 47404
rect 21382 47340 21428 47404
rect 463 47054 863 47339
rect 463 46990 508 47054
rect 572 46990 630 47054
rect 694 46990 756 47054
rect 820 46990 863 47054
rect 463 46907 863 46990
rect 463 46843 508 46907
rect 572 46843 630 46907
rect 694 46843 756 46907
rect 820 46843 863 46907
rect 463 46770 863 46843
rect 463 46706 508 46770
rect 572 46706 630 46770
rect 694 46706 756 46770
rect 820 46706 863 46770
rect 463 45294 863 46706
rect 463 45230 508 45294
rect 572 45230 630 45294
rect 694 45230 756 45294
rect 820 45230 863 45294
rect 463 45147 863 45230
rect 463 45083 508 45147
rect 572 45083 630 45147
rect 694 45083 756 45147
rect 820 45083 863 45147
rect 463 45010 863 45083
rect 463 44946 508 45010
rect 572 44946 630 45010
rect 694 44946 756 45010
rect 820 44946 863 45010
rect 463 44503 863 44946
rect 463 44439 507 44503
rect 571 44439 633 44503
rect 697 44439 753 44503
rect 817 44439 863 44503
rect 463 44385 863 44439
rect 463 44321 507 44385
rect 571 44321 633 44385
rect 697 44321 753 44385
rect 817 44321 863 44385
rect 463 39123 863 44321
rect 21028 44406 21428 47340
rect 21028 44342 21072 44406
rect 21136 44342 21198 44406
rect 21262 44342 21318 44406
rect 21382 44342 21428 44406
rect 21028 44288 21428 44342
rect 21028 44224 21072 44288
rect 21136 44224 21198 44288
rect 21262 44224 21318 44288
rect 21382 44224 21428 44288
rect 2306 39942 2868 44002
rect 2246 39925 2868 39942
rect 2246 39861 2249 39925
rect 2313 39861 2337 39925
rect 2401 39861 2868 39925
rect 2246 39845 2868 39861
rect 2246 39781 2249 39845
rect 2313 39781 2337 39845
rect 2401 39781 2868 39845
rect 2246 39775 2868 39781
rect 2306 39774 2868 39775
rect 4119 39905 4490 44000
rect 4119 39841 4192 39905
rect 4256 39841 4280 39905
rect 4344 39841 4490 39905
rect 4119 39825 4490 39841
rect 4119 39761 4192 39825
rect 4256 39761 4280 39825
rect 4344 39761 4490 39825
rect 4119 39754 4490 39761
rect 463 39059 488 39123
rect 552 39059 602 39123
rect 666 39059 716 39123
rect 780 39059 863 39123
rect 463 38035 863 39059
rect 463 37971 488 38035
rect 552 37971 602 38035
rect 666 37971 716 38035
rect 780 37971 863 38035
rect 463 36947 863 37971
rect 463 36883 488 36947
rect 552 36883 602 36947
rect 666 36883 716 36947
rect 780 36883 863 36947
rect 463 32360 863 36883
rect 2306 36463 2738 36476
rect 2306 36399 2536 36463
rect 2600 36399 2624 36463
rect 2688 36399 2738 36463
rect 463 32296 866 32360
rect 463 32232 507 32296
rect 571 32232 633 32296
rect 697 32232 753 32296
rect 817 32232 866 32296
rect 463 32178 866 32232
rect 463 32114 507 32178
rect 571 32114 633 32178
rect 697 32114 753 32178
rect 817 32114 866 32178
rect 463 32072 866 32114
rect 463 32000 863 32072
rect 2306 32000 2738 36399
rect 21028 36198 21428 44224
rect 20527 36164 21428 36198
rect 20527 36100 21069 36164
rect 21133 36100 21194 36164
rect 21258 36100 21319 36164
rect 21383 36100 21428 36164
rect 20527 36044 21428 36100
rect 20527 35980 21068 36044
rect 21132 35980 21193 36044
rect 21257 35980 21318 36044
rect 21382 35980 21428 36044
rect 20527 35943 21428 35980
rect 21028 35586 21428 35943
rect 21028 35522 21073 35586
rect 21137 35522 21195 35586
rect 21259 35522 21321 35586
rect 21385 35522 21428 35586
rect 21028 35439 21428 35522
rect 21028 35375 21073 35439
rect 21137 35375 21195 35439
rect 21259 35375 21321 35439
rect 21385 35375 21428 35439
rect 21028 35302 21428 35375
rect 21028 35238 21073 35302
rect 21137 35238 21195 35302
rect 21259 35238 21321 35302
rect 21385 35238 21428 35302
rect 20527 34668 20927 34702
rect 20527 34604 20568 34668
rect 20632 34604 20693 34668
rect 20757 34604 20818 34668
rect 20882 34604 20927 34668
rect 20527 34548 20927 34604
rect 20527 34484 20567 34548
rect 20631 34484 20692 34548
rect 20756 34484 20817 34548
rect 20881 34484 20927 34548
rect 20527 34447 20927 34484
rect 21028 33826 21428 35238
rect 21028 33762 21073 33826
rect 21137 33762 21195 33826
rect 21259 33762 21321 33826
rect 21385 33762 21428 33826
rect 21028 33679 21428 33762
rect 21028 33615 21073 33679
rect 21137 33615 21195 33679
rect 21259 33615 21321 33679
rect 21385 33615 21428 33679
rect 21028 33542 21428 33615
rect 21028 33478 21073 33542
rect 21137 33478 21195 33542
rect 21259 33478 21321 33542
rect 21385 33478 21428 33542
rect 21028 33143 21428 33478
rect 20514 33109 21428 33143
rect 20514 33045 21068 33109
rect 21132 33045 21193 33109
rect 21257 33045 21318 33109
rect 21382 33045 21428 33109
rect 20514 32989 21428 33045
rect 20514 32925 21067 32989
rect 21131 32925 21192 32989
rect 21256 32925 21317 32989
rect 21381 32925 21428 32989
rect 20514 32888 21428 32925
rect 21028 32360 21428 32888
rect 21025 32296 21428 32360
rect 21025 32232 21072 32296
rect 21136 32232 21198 32296
rect 21262 32232 21318 32296
rect 21382 32232 21428 32296
rect 21025 32178 21428 32232
rect 21025 32114 21072 32178
rect 21136 32114 21198 32178
rect 21262 32114 21318 32178
rect 21382 32114 21428 32178
rect 21025 32072 21428 32114
rect 463 31760 946 32000
rect 463 31514 863 31760
rect 463 31450 507 31514
rect 571 31450 633 31514
rect 697 31450 753 31514
rect 817 31450 863 31514
rect 463 31396 863 31450
rect 463 31332 507 31396
rect 571 31332 633 31396
rect 697 31332 753 31396
rect 817 31332 863 31396
rect 463 31055 863 31332
rect 21028 31514 21428 32072
rect 21028 31450 21072 31514
rect 21136 31450 21198 31514
rect 21262 31450 21318 31514
rect 21382 31450 21428 31514
rect 21028 31396 21428 31450
rect 21028 31332 21072 31396
rect 21136 31332 21198 31396
rect 21262 31332 21318 31396
rect 21382 31332 21428 31396
rect 953 31120 1155 31121
rect 463 30991 508 31055
rect 572 30991 630 31055
rect 694 30991 756 31055
rect 820 30991 863 31055
rect 463 30908 863 30991
rect 463 30844 508 30908
rect 572 30844 630 30908
rect 694 30844 756 30908
rect 820 30844 863 30908
rect 463 30771 863 30844
rect 463 30707 508 30771
rect 572 30707 630 30771
rect 694 30707 756 30771
rect 820 30707 863 30771
rect 463 29288 863 30707
rect 463 29224 508 29288
rect 572 29224 630 29288
rect 694 29224 756 29288
rect 820 29224 863 29288
rect 463 29141 863 29224
rect 463 29077 508 29141
rect 572 29077 630 29141
rect 694 29077 756 29141
rect 820 29077 863 29141
rect 463 29004 863 29077
rect 463 28940 508 29004
rect 572 28940 630 29004
rect 694 28940 756 29004
rect 820 28940 863 29004
rect 463 28602 863 28940
rect 463 28538 507 28602
rect 571 28538 633 28602
rect 697 28538 753 28602
rect 817 28538 863 28602
rect 463 28484 863 28538
rect 463 28420 507 28484
rect 571 28420 633 28484
rect 697 28420 753 28484
rect 817 28420 863 28484
rect 463 28238 863 28420
rect 21028 28553 21428 31332
rect 21028 28489 21072 28553
rect 21136 28489 21198 28553
rect 21262 28489 21318 28553
rect 21382 28489 21428 28553
rect 21028 28435 21428 28489
rect 21028 28371 21072 28435
rect 21136 28371 21198 28435
rect 21262 28371 21318 28435
rect 21382 28371 21428 28435
rect 463 28209 946 28238
rect 21028 28232 21428 28371
rect 462 27979 946 28209
rect 463 27760 946 27979
rect 20946 27766 21428 28232
rect 463 27598 863 27760
rect 463 27534 507 27598
rect 571 27534 633 27598
rect 697 27534 753 27598
rect 817 27534 863 27598
rect 463 27480 863 27534
rect 463 27416 507 27480
rect 571 27416 633 27480
rect 697 27416 753 27480
rect 817 27416 863 27480
rect 21028 27467 21428 27766
rect 463 27054 863 27416
rect 21027 27436 21428 27467
rect 21027 27372 21072 27436
rect 21136 27372 21198 27436
rect 21262 27372 21318 27436
rect 21382 27372 21428 27436
rect 21027 27318 21428 27372
rect 21027 27254 21072 27318
rect 21136 27254 21198 27318
rect 21262 27254 21318 27318
rect 21382 27254 21428 27318
rect 21027 27212 21428 27254
rect 463 26990 508 27054
rect 572 26990 630 27054
rect 694 26990 756 27054
rect 820 26990 863 27054
rect 463 26907 863 26990
rect 463 26843 508 26907
rect 572 26843 630 26907
rect 694 26843 756 26907
rect 820 26843 863 26907
rect 463 26770 863 26843
rect 463 26706 508 26770
rect 572 26706 630 26770
rect 694 26706 756 26770
rect 820 26706 863 26770
rect 463 25294 863 26706
rect 463 25230 508 25294
rect 572 25230 630 25294
rect 694 25230 756 25294
rect 820 25230 863 25294
rect 463 25147 863 25230
rect 463 25083 508 25147
rect 572 25083 630 25147
rect 694 25083 756 25147
rect 820 25083 863 25147
rect 463 25010 863 25083
rect 463 24946 508 25010
rect 572 24946 630 25010
rect 694 24946 756 25010
rect 820 24946 863 25010
rect 463 24651 863 24946
rect 463 24620 864 24651
rect 463 24556 507 24620
rect 571 24556 633 24620
rect 697 24556 753 24620
rect 817 24556 864 24620
rect 463 24502 864 24556
rect 463 24438 507 24502
rect 571 24438 633 24502
rect 697 24438 753 24502
rect 817 24438 864 24502
rect 463 24396 864 24438
rect 21028 24593 21428 27212
rect 21028 24529 21072 24593
rect 21136 24529 21198 24593
rect 21262 24529 21318 24593
rect 21382 24529 21428 24593
rect 21028 24475 21428 24529
rect 21028 24411 21072 24475
rect 21136 24411 21198 24475
rect 21262 24411 21318 24475
rect 21382 24411 21428 24475
rect 463 24239 863 24396
rect 463 23759 947 24239
rect 21028 24232 21428 24411
rect 20946 23767 21428 24232
rect 463 23569 863 23759
rect 463 23538 864 23569
rect 463 23474 507 23538
rect 571 23474 633 23538
rect 697 23474 753 23538
rect 817 23474 864 23538
rect 463 23420 864 23474
rect 463 23356 507 23420
rect 571 23356 633 23420
rect 697 23356 753 23420
rect 817 23356 864 23420
rect 463 23314 864 23356
rect 21028 23418 21428 23767
rect 21028 23354 21072 23418
rect 21136 23354 21198 23418
rect 21262 23354 21318 23418
rect 21382 23354 21428 23418
rect 463 23054 863 23314
rect 463 22990 508 23054
rect 572 22990 630 23054
rect 694 22990 756 23054
rect 820 22990 863 23054
rect 463 22907 863 22990
rect 463 22843 508 22907
rect 572 22843 630 22907
rect 694 22843 756 22907
rect 820 22843 863 22907
rect 463 22770 863 22843
rect 463 22706 508 22770
rect 572 22706 630 22770
rect 694 22706 756 22770
rect 820 22706 863 22770
rect 463 21295 863 22706
rect 463 21231 508 21295
rect 572 21231 630 21295
rect 694 21231 756 21295
rect 820 21231 863 21295
rect 463 21148 863 21231
rect 463 21084 508 21148
rect 572 21084 630 21148
rect 694 21084 756 21148
rect 820 21084 863 21148
rect 463 21011 863 21084
rect 463 20947 508 21011
rect 572 20947 630 21011
rect 694 20947 756 21011
rect 820 20947 863 21011
rect 463 20694 863 20947
rect 21028 23300 21428 23354
rect 21028 23236 21072 23300
rect 21136 23236 21198 23300
rect 21262 23236 21318 23300
rect 21382 23236 21428 23300
rect 463 20663 864 20694
rect 463 20599 507 20663
rect 571 20599 633 20663
rect 697 20599 753 20663
rect 817 20599 864 20663
rect 21028 20608 21428 23236
rect 463 20545 864 20599
rect 463 20481 507 20545
rect 571 20481 633 20545
rect 697 20481 753 20545
rect 817 20481 864 20545
rect 463 20439 864 20481
rect 21027 20577 21428 20608
rect 21027 20513 21072 20577
rect 21136 20513 21198 20577
rect 21262 20513 21318 20577
rect 21382 20513 21428 20577
rect 21027 20459 21428 20513
rect 463 20240 863 20439
rect 21027 20395 21072 20459
rect 21136 20395 21198 20459
rect 21262 20395 21318 20459
rect 21382 20395 21428 20459
rect 21027 20353 21428 20395
rect 463 19760 946 20240
rect 21028 20233 21428 20353
rect 20946 19768 21428 20233
rect 463 19593 863 19760
rect 463 19562 864 19593
rect 463 19498 507 19562
rect 571 19498 633 19562
rect 697 19498 753 19562
rect 817 19498 864 19562
rect 463 19444 864 19498
rect 463 19380 507 19444
rect 571 19380 633 19444
rect 697 19380 753 19444
rect 817 19380 864 19444
rect 21028 19437 21428 19768
rect 463 19338 864 19380
rect 21027 19406 21428 19437
rect 21027 19342 21072 19406
rect 21136 19342 21198 19406
rect 21262 19342 21318 19406
rect 21382 19342 21428 19406
rect 463 19054 863 19338
rect 21027 19288 21428 19342
rect 21027 19224 21072 19288
rect 21136 19224 21198 19288
rect 21262 19224 21318 19288
rect 21382 19224 21428 19288
rect 21027 19182 21428 19224
rect 463 18990 508 19054
rect 572 18990 630 19054
rect 694 18990 756 19054
rect 820 18990 863 19054
rect 463 18907 863 18990
rect 463 18843 508 18907
rect 572 18843 630 18907
rect 694 18843 756 18907
rect 820 18843 863 18907
rect 463 18770 863 18843
rect 463 18706 508 18770
rect 572 18706 630 18770
rect 694 18706 756 18770
rect 820 18706 863 18770
rect 463 17294 863 18706
rect 463 17230 508 17294
rect 572 17230 630 17294
rect 694 17230 756 17294
rect 820 17230 863 17294
rect 463 17147 863 17230
rect 463 17083 508 17147
rect 572 17083 630 17147
rect 694 17083 756 17147
rect 820 17083 863 17147
rect 463 17010 863 17083
rect 463 16946 508 17010
rect 572 16946 630 17010
rect 694 16946 756 17010
rect 820 16946 863 17010
rect 463 16727 863 16946
rect 463 16696 865 16727
rect 463 16632 507 16696
rect 571 16632 633 16696
rect 697 16632 753 16696
rect 817 16632 865 16696
rect 21028 16676 21428 19182
rect 463 16578 865 16632
rect 463 16514 507 16578
rect 571 16514 633 16578
rect 697 16514 753 16578
rect 817 16514 865 16578
rect 463 16472 865 16514
rect 21027 16645 21428 16676
rect 21027 16581 21072 16645
rect 21136 16581 21198 16645
rect 21262 16581 21318 16645
rect 21382 16581 21428 16645
rect 21027 16527 21428 16581
rect 463 16239 863 16472
rect 21027 16463 21072 16527
rect 21136 16463 21198 16527
rect 21262 16463 21318 16527
rect 21382 16463 21428 16527
rect 21027 16421 21428 16463
rect 463 15759 946 16239
rect 21028 16232 21428 16421
rect 20946 15766 21428 16232
rect 463 15511 863 15759
rect 463 15480 866 15511
rect 463 15416 507 15480
rect 571 15416 633 15480
rect 697 15416 753 15480
rect 817 15416 866 15480
rect 21028 15462 21428 15766
rect 463 15362 866 15416
rect 463 15298 507 15362
rect 571 15298 633 15362
rect 697 15298 753 15362
rect 817 15298 866 15362
rect 463 15256 866 15298
rect 21027 15431 21428 15462
rect 21027 15367 21072 15431
rect 21136 15367 21198 15431
rect 21262 15367 21318 15431
rect 21382 15367 21428 15431
rect 21027 15313 21428 15367
rect 463 15054 863 15256
rect 21027 15249 21072 15313
rect 21136 15249 21198 15313
rect 21262 15249 21318 15313
rect 21382 15249 21428 15313
rect 21027 15207 21428 15249
rect 463 14990 508 15054
rect 572 14990 630 15054
rect 694 14990 756 15054
rect 820 14990 863 15054
rect 463 14907 863 14990
rect 463 14843 508 14907
rect 572 14843 630 14907
rect 694 14843 756 14907
rect 820 14843 863 14907
rect 463 14770 863 14843
rect 463 14706 508 14770
rect 572 14706 630 14770
rect 694 14706 756 14770
rect 820 14706 863 14770
rect 463 13294 863 14706
rect 463 13230 508 13294
rect 572 13230 630 13294
rect 694 13230 756 13294
rect 820 13230 863 13294
rect 463 13147 863 13230
rect 463 13083 508 13147
rect 572 13083 630 13147
rect 694 13083 756 13147
rect 820 13083 863 13147
rect 463 13010 863 13083
rect 463 12946 508 13010
rect 572 12946 630 13010
rect 694 12946 756 13010
rect 820 12946 863 13010
rect 463 12646 863 12946
rect 463 12615 864 12646
rect 463 12551 507 12615
rect 571 12551 633 12615
rect 697 12551 753 12615
rect 817 12551 864 12615
rect 463 12497 864 12551
rect 463 12433 507 12497
rect 571 12433 633 12497
rect 697 12433 753 12497
rect 817 12433 864 12497
rect 463 12391 864 12433
rect 21028 12588 21428 15207
rect 21028 12524 21072 12588
rect 21136 12524 21198 12588
rect 21262 12524 21318 12588
rect 21382 12524 21428 12588
rect 21028 12470 21428 12524
rect 21028 12406 21072 12470
rect 21136 12406 21198 12470
rect 21262 12406 21318 12470
rect 21382 12406 21428 12470
rect 463 12238 863 12391
rect 463 11998 947 12238
rect 21028 12233 21428 12406
rect 463 11758 946 11998
rect 20946 11766 21428 12233
rect 463 11524 863 11758
rect 463 11493 864 11524
rect 463 11429 507 11493
rect 571 11429 633 11493
rect 697 11429 753 11493
rect 817 11429 864 11493
rect 21028 11462 21428 11766
rect 463 11375 864 11429
rect 463 11311 507 11375
rect 571 11311 633 11375
rect 697 11311 753 11375
rect 817 11311 864 11375
rect 463 11269 864 11311
rect 21027 11431 21428 11462
rect 21027 11367 21072 11431
rect 21136 11367 21198 11431
rect 21262 11367 21318 11431
rect 21382 11367 21428 11431
rect 21027 11313 21428 11367
rect 463 11055 863 11269
rect 21027 11249 21072 11313
rect 21136 11249 21198 11313
rect 21262 11249 21318 11313
rect 21382 11249 21428 11313
rect 21027 11207 21428 11249
rect 463 10991 508 11055
rect 572 10991 630 11055
rect 694 10991 756 11055
rect 820 10991 863 11055
rect 463 10908 863 10991
rect 463 10844 508 10908
rect 572 10844 630 10908
rect 694 10844 756 10908
rect 820 10844 863 10908
rect 463 10771 863 10844
rect 463 10707 508 10771
rect 572 10707 630 10771
rect 694 10707 756 10771
rect 820 10707 863 10771
rect 463 9293 863 10707
rect 463 9229 508 9293
rect 572 9229 630 9293
rect 694 9229 756 9293
rect 820 9229 863 9293
rect 463 9146 863 9229
rect 463 9082 508 9146
rect 572 9082 630 9146
rect 694 9082 756 9146
rect 820 9082 863 9146
rect 463 9009 863 9082
rect 463 8945 508 9009
rect 572 8945 630 9009
rect 694 8945 756 9009
rect 820 8945 863 9009
rect 463 8633 863 8945
rect 463 8569 507 8633
rect 571 8569 633 8633
rect 697 8569 753 8633
rect 817 8569 863 8633
rect 463 8515 863 8569
rect 463 8451 507 8515
rect 571 8451 633 8515
rect 697 8451 753 8515
rect 817 8451 863 8515
rect 463 8238 863 8451
rect 21028 8588 21428 11207
rect 21028 8524 21072 8588
rect 21136 8524 21198 8588
rect 21262 8524 21318 8588
rect 21382 8524 21428 8588
rect 21028 8470 21428 8524
rect 21028 8406 21072 8470
rect 21136 8406 21198 8470
rect 21262 8406 21318 8470
rect 21382 8406 21428 8470
rect 463 8000 946 8238
rect 21028 8233 21428 8406
rect 463 7760 947 8000
rect 20946 7766 21428 8233
rect 463 7522 863 7760
rect 463 7458 507 7522
rect 571 7458 633 7522
rect 697 7458 753 7522
rect 817 7458 863 7522
rect 21028 7462 21428 7766
rect 463 7404 863 7458
rect 463 7340 507 7404
rect 571 7340 633 7404
rect 697 7340 753 7404
rect 817 7340 863 7404
rect 463 7055 863 7340
rect 21027 7431 21428 7462
rect 21027 7367 21072 7431
rect 21136 7367 21198 7431
rect 21262 7367 21318 7431
rect 21382 7367 21428 7431
rect 21027 7313 21428 7367
rect 21027 7249 21072 7313
rect 21136 7249 21198 7313
rect 21262 7249 21318 7313
rect 21382 7249 21428 7313
rect 21027 7207 21428 7249
rect 463 6991 508 7055
rect 572 6991 630 7055
rect 694 6991 756 7055
rect 820 6991 863 7055
rect 463 6908 863 6991
rect 463 6844 508 6908
rect 572 6844 630 6908
rect 694 6844 756 6908
rect 820 6844 863 6908
rect 463 6771 863 6844
rect 463 6707 508 6771
rect 572 6707 630 6771
rect 694 6707 756 6771
rect 820 6707 863 6771
rect 463 5294 863 6707
rect 463 5230 508 5294
rect 572 5230 630 5294
rect 694 5230 756 5294
rect 820 5230 863 5294
rect 463 5147 863 5230
rect 463 5083 508 5147
rect 572 5083 630 5147
rect 694 5083 756 5147
rect 820 5083 863 5147
rect 463 5010 863 5083
rect 463 4946 508 5010
rect 572 4946 630 5010
rect 694 4946 756 5010
rect 820 4946 863 5010
rect 463 4730 863 4946
rect 463 4699 865 4730
rect 463 4635 507 4699
rect 571 4635 633 4699
rect 697 4635 753 4699
rect 817 4635 865 4699
rect 463 4581 865 4635
rect 463 4517 507 4581
rect 571 4517 633 4581
rect 697 4517 753 4581
rect 817 4517 865 4581
rect 463 4475 865 4517
rect 21028 4588 21428 7207
rect 21028 4524 21072 4588
rect 21136 4524 21198 4588
rect 21262 4524 21318 4588
rect 21382 4524 21428 4588
rect 463 4239 863 4475
rect 21028 4470 21428 4524
rect 21028 4406 21072 4470
rect 21136 4406 21198 4470
rect 21262 4406 21318 4470
rect 21382 4406 21428 4470
rect 463 4000 947 4239
rect 21028 4233 21428 4406
rect 463 3760 946 4000
rect 20946 3766 21428 4233
rect 463 3522 863 3760
rect 463 3458 507 3522
rect 571 3458 633 3522
rect 697 3458 753 3522
rect 817 3458 863 3522
rect 21028 3462 21428 3766
rect 463 3404 863 3458
rect 463 3340 507 3404
rect 571 3340 633 3404
rect 697 3340 753 3404
rect 817 3340 863 3404
rect 463 3055 863 3340
rect 21027 3431 21428 3462
rect 21027 3367 21072 3431
rect 21136 3367 21198 3431
rect 21262 3367 21318 3431
rect 21382 3367 21428 3431
rect 21027 3313 21428 3367
rect 21027 3249 21072 3313
rect 21136 3249 21198 3313
rect 21262 3249 21318 3313
rect 21382 3249 21428 3313
rect 21027 3207 21428 3249
rect 463 2991 508 3055
rect 572 2991 630 3055
rect 694 2991 756 3055
rect 820 2991 863 3055
rect 463 2908 863 2991
rect 463 2844 508 2908
rect 572 2844 630 2908
rect 694 2844 756 2908
rect 820 2844 863 2908
rect 463 2771 863 2844
rect 463 2707 508 2771
rect 572 2707 630 2771
rect 694 2707 756 2771
rect 820 2707 863 2771
rect 463 1294 863 2707
rect 463 1230 508 1294
rect 572 1230 630 1294
rect 694 1230 756 1294
rect 820 1230 863 1294
rect 463 1147 863 1230
rect 463 1083 508 1147
rect 572 1083 630 1147
rect 694 1083 756 1147
rect 820 1083 863 1147
rect 463 1010 863 1083
rect 463 946 508 1010
rect 572 946 630 1010
rect 694 946 756 1010
rect 820 946 863 1010
rect 463 730 863 946
rect 463 699 865 730
rect 463 635 507 699
rect 571 635 633 699
rect 697 635 753 699
rect 817 635 865 699
rect 463 581 865 635
rect 463 517 507 581
rect 571 517 633 581
rect 697 517 753 581
rect 817 517 865 581
rect 463 475 865 517
rect 21028 588 21428 3207
rect 21028 524 21072 588
rect 21136 524 21198 588
rect 21262 524 21318 588
rect 21382 524 21428 588
rect 463 239 863 475
rect 21028 470 21428 524
rect 21028 406 21072 470
rect 21136 406 21198 470
rect 21262 406 21318 470
rect 21382 406 21428 470
rect 463 0 946 239
rect 21028 233 21428 406
rect 20946 0 21428 233
rect 21502 39718 21902 76000
rect 21502 39654 21543 39718
rect 21607 39654 21668 39718
rect 21732 39654 21793 39718
rect 21857 39654 21902 39718
rect 21502 39598 21902 39654
rect 21502 39534 21542 39598
rect 21606 39534 21667 39598
rect 21731 39534 21792 39598
rect 21856 39534 21902 39598
rect 21502 34668 21902 39534
rect 21502 34604 21543 34668
rect 21607 34604 21668 34668
rect 21732 34604 21793 34668
rect 21857 34604 21902 34668
rect 21502 34548 21902 34604
rect 21502 34484 21542 34548
rect 21606 34484 21667 34548
rect 21731 34484 21792 34548
rect 21856 34484 21902 34548
rect 21502 0 21902 34484
rect 21970 74065 22370 76000
rect 21970 74001 22014 74065
rect 22078 74001 22140 74065
rect 22204 74001 22260 74065
rect 22324 74001 22370 74065
rect 21970 73947 22370 74001
rect 21970 73883 22014 73947
rect 22078 73883 22140 73947
rect 22204 73883 22260 73947
rect 22324 73883 22370 73947
rect 21970 70065 22370 73883
rect 21970 70001 22014 70065
rect 22078 70001 22140 70065
rect 22204 70001 22260 70065
rect 22324 70001 22370 70065
rect 21970 69947 22370 70001
rect 21970 69883 22014 69947
rect 22078 69883 22140 69947
rect 22204 69883 22260 69947
rect 22324 69883 22370 69947
rect 21970 66052 22370 69883
rect 21970 65988 22014 66052
rect 22078 65988 22140 66052
rect 22204 65988 22260 66052
rect 22324 65988 22370 66052
rect 21970 65934 22370 65988
rect 21970 65870 22014 65934
rect 22078 65870 22140 65934
rect 22204 65870 22260 65934
rect 22324 65870 22370 65934
rect 21970 62051 22370 65870
rect 21970 61987 22014 62051
rect 22078 61987 22140 62051
rect 22204 61987 22260 62051
rect 22324 61987 22370 62051
rect 21970 61933 22370 61987
rect 21970 61869 22014 61933
rect 22078 61869 22140 61933
rect 22204 61869 22260 61933
rect 22324 61869 22370 61933
rect 21970 58090 22370 61869
rect 21970 58026 22014 58090
rect 22078 58026 22140 58090
rect 22204 58026 22260 58090
rect 22324 58026 22370 58090
rect 21970 57972 22370 58026
rect 21970 57908 22014 57972
rect 22078 57908 22140 57972
rect 22204 57908 22260 57972
rect 22324 57908 22370 57972
rect 21970 54073 22370 57908
rect 21970 54009 22014 54073
rect 22078 54009 22140 54073
rect 22204 54009 22260 54073
rect 22324 54009 22370 54073
rect 21970 53955 22370 54009
rect 21970 53891 22014 53955
rect 22078 53891 22140 53955
rect 22204 53891 22260 53955
rect 22324 53891 22370 53955
rect 21970 50152 22370 53891
rect 21970 50088 22014 50152
rect 22078 50088 22140 50152
rect 22204 50088 22260 50152
rect 22324 50088 22370 50152
rect 21970 50034 22370 50088
rect 21970 49970 22014 50034
rect 22078 49970 22140 50034
rect 22204 49970 22260 50034
rect 22324 49970 22370 50034
rect 21970 45894 22370 49970
rect 21970 45830 22014 45894
rect 22078 45830 22140 45894
rect 22204 45830 22260 45894
rect 22324 45830 22370 45894
rect 21970 45776 22370 45830
rect 21970 45712 22014 45776
rect 22078 45712 22140 45776
rect 22204 45712 22260 45776
rect 22324 45712 22370 45776
rect 21970 43828 22370 45712
rect 21970 43524 22040 43828
rect 22264 43524 22370 43828
rect 21970 36944 22370 43524
rect 21970 36640 22040 36944
rect 22264 36640 22370 36944
rect 21970 30124 22370 36640
rect 21970 30060 22014 30124
rect 22078 30060 22140 30124
rect 22204 30060 22260 30124
rect 22324 30060 22370 30124
rect 21970 30006 22370 30060
rect 21970 29942 22014 30006
rect 22078 29942 22140 30006
rect 22204 29942 22260 30006
rect 22324 29942 22370 30006
rect 21970 25965 22370 29942
rect 21970 25901 22014 25965
rect 22078 25901 22140 25965
rect 22204 25901 22260 25965
rect 22324 25901 22370 25965
rect 21970 25847 22370 25901
rect 21970 25783 22014 25847
rect 22078 25783 22140 25847
rect 22204 25783 22260 25847
rect 22324 25783 22370 25847
rect 21970 22175 22370 25783
rect 21970 22111 22014 22175
rect 22078 22111 22140 22175
rect 22204 22111 22260 22175
rect 22324 22111 22370 22175
rect 21970 22057 22370 22111
rect 21970 21993 22014 22057
rect 22078 21993 22140 22057
rect 22204 21993 22260 22057
rect 22324 21993 22370 22057
rect 21970 18068 22370 21993
rect 21970 18004 22014 18068
rect 22078 18004 22140 18068
rect 22204 18004 22260 18068
rect 22324 18004 22370 18068
rect 21970 17950 22370 18004
rect 21970 17886 22014 17950
rect 22078 17886 22140 17950
rect 22204 17886 22260 17950
rect 22324 17886 22370 17950
rect 21970 14250 22370 17886
rect 21970 14186 22014 14250
rect 22078 14186 22140 14250
rect 22204 14186 22260 14250
rect 22324 14186 22370 14250
rect 21970 14132 22370 14186
rect 21970 14068 22014 14132
rect 22078 14068 22140 14132
rect 22204 14068 22260 14132
rect 22324 14068 22370 14132
rect 21970 10286 22370 14068
rect 21970 10222 22014 10286
rect 22078 10222 22140 10286
rect 22204 10222 22260 10286
rect 22324 10222 22370 10286
rect 21970 10168 22370 10222
rect 21970 10104 22014 10168
rect 22078 10104 22140 10168
rect 22204 10104 22260 10168
rect 22324 10104 22370 10168
rect 21970 6274 22370 10104
rect 21970 6210 22014 6274
rect 22078 6210 22140 6274
rect 22204 6210 22260 6274
rect 22324 6210 22370 6274
rect 21970 6156 22370 6210
rect 21970 6092 22014 6156
rect 22078 6092 22140 6156
rect 22204 6092 22260 6156
rect 22324 6092 22370 6156
rect 21970 2274 22370 6092
rect 21970 2210 22014 2274
rect 22078 2210 22140 2274
rect 22204 2210 22260 2274
rect 22324 2210 22370 2274
rect 21970 2156 22370 2210
rect 21970 2092 22014 2156
rect 22078 2092 22140 2156
rect 22204 2092 22260 2156
rect 22324 2092 22370 2156
rect 21970 0 22370 2092
use adc_noise_decoup_cell1  adc_noise_decoup_cell1_0
array 0 2 4000 0 0 0
timestamp 1515178157
transform 1 0 8527 0 1 32532
box 0 0 4000 4000
use adc_noise_decoup_cell1  adc_noise_decoup_cell1_1
array 0 4 4000 0 7 4000
timestamp 1515178157
transform 1 0 946 0 1 0
box 0 0 4000 4000
use adc_noise_decoup_cell1  adc_noise_decoup_cell1_3
array 0 4 4000 0 7 4000
timestamp 1515178157
transform 1 0 946 0 1 44000
box 0 0 4000 4000
use nfet_01v8_w500_l500_nf2  nfet_01v8_w500_l500_nf2_0
timestamp 1515178157
transform 1 0 2655 0 1 39031
box -213 -76 213 76
use nfet_01v8_w500_l500_nf2  nfet_01v8_w500_l500_nf2_1
timestamp 1515178157
transform 1 0 2210 0 1 39031
box -213 -76 213 76
use nfet_01v8_w500_l500_nf2  nfet_01v8_w500_l500_nf2_2
timestamp 1515178157
transform 1 0 2612 0 1 36975
box -213 -76 213 76
use nfet_01v8_w500_l500_nf2  nfet_01v8_w500_l500_nf2_3
timestamp 1515178157
transform 1 0 2132 0 1 36975
box -213 -76 213 76
use nfet_01v8_w500_l500_nf2  nfet_01v8_w500_l500_nf2_4
timestamp 1515178157
transform 1 0 1779 0 -1 39031
box -213 -76 213 76
use pfet_01v8_w500_l500_nf2  pfet_01v8_w500_l500_nf2_0
timestamp 1515178157
transform 1 0 2655 0 1 38693
box -224 -36 223 138
use pfet_01v8_w500_l500_nf2  pfet_01v8_w500_l500_nf2_1
timestamp 1515178157
transform 1 0 2210 0 1 38692
box -224 -36 223 138
use pfet_01v8_w500_l500_nf2  pfet_01v8_w500_l500_nf2_2
timestamp 1515178157
transform 1 0 2612 0 1 37213
box -224 -36 223 138
use pfet_01v8_w500_l500_nf2  pfet_01v8_w500_l500_nf2_3
timestamp 1515178157
transform 1 0 2132 0 1 37213
box -224 -36 223 138
use pfet_01v8_w500_l500_nf2  pfet_01v8_w500_l500_nf2_4
timestamp 1515178157
transform 1 0 1779 0 -1 38794
box -224 -36 223 138
use sky130_fd_sc_hd__buf_4  sky130_fd_sc_hd__buf_4_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform -1 0 4169 0 -1 39091
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  sky130_fd_sc_hd__buf_4_1
timestamp 1694700623
transform -1 0 3617 0 -1 39091
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  sky130_fd_sc_hd__buf_4_2
timestamp 1694700623
transform -1 0 4169 0 1 36915
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  sky130_fd_sc_hd__buf_4_3
timestamp 1694700623
transform -1 0 3617 0 1 36915
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s6s_1  sky130_fd_sc_hd__dlymetal6s6s_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 1961 0 1 38003
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s6s_1  sky130_fd_sc_hd__dlymetal6s6s_1_1
timestamp 1694700623
transform 1 0 1961 0 -1 38003
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s6s_1  sky130_fd_sc_hd__dlymetal6s6s_1_2
timestamp 1694700623
transform 1 0 2881 0 1 38003
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s6s_1  sky130_fd_sc_hd__dlymetal6s6s_1_3
timestamp 1694700623
transform 1 0 3801 0 1 38003
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s6s_1  sky130_fd_sc_hd__dlymetal6s6s_1_4
timestamp 1694700623
transform 1 0 2881 0 -1 38003
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s6s_1  sky130_fd_sc_hd__dlymetal6s6s_1_5
timestamp 1694700623
transform 1 0 3801 0 -1 38003
box -38 -48 958 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform -1 0 4721 0 -1 39091
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_1
timestamp 1694700623
transform -1 0 4721 0 1 36915
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_2
timestamp 1694700623
transform -1 0 4445 0 -1 39091
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_3
timestamp 1694700623
transform -1 0 4445 0 1 36915
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_4
timestamp 1694700623
transform 1 0 1409 0 -1 38003
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  sky130_fd_sc_hd__nand2_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform -1 0 1961 0 1 38003
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  sky130_fd_sc_hd__nand2_1_1
timestamp 1694700623
transform 1 0 1685 0 -1 38003
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 1593 0 1 38003
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_1
timestamp 1694700623
transform -1 0 3065 0 -1 39091
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_2
timestamp 1694700623
transform -1 0 3065 0 1 36915
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_3
timestamp 1694700623
transform 1 0 1317 0 -1 38003
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_4
timestamp 1694700623
transform 1 0 1501 0 1 36915
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_5
timestamp 1694700623
transform 1 0 1388 0 -1 39092
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_6
timestamp 1694700623
transform 1 0 4721 0 1 38003
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_7
timestamp 1694700623
transform 1 0 4721 0 -1 38003
box -38 -48 130 592
<< labels >>
flabel locali s 1339 38217 1373 38269 0 FreeSans 1000 0 0 0 clk
port 0 nsew
flabel metal1 s 2919 37023 2956 37058 0 FreeSans 400 180 0 0 phi2
port 3 nsew
flabel metal1 s 2900 38829 2937 38876 0 FreeSans 400 180 0 0 phi1_n
port 5 nsew
flabel metal1 s 2899 38946 2935 38981 0 FreeSans 400 180 0 0 phi1
port 7 nsew
flabel metal1 s 2867 37131 2904 37178 0 FreeSans 400 180 0 0 phi2_n
port 9 nsew
rlabel metal2 s 22306 36596 22370 36986 4 vcm
port 10 nsew
flabel metal4 s 0 0 400 76000 0 FreeSans 2000 90 0 0 VDD
port 11 nsew
flabel metal4 s 21502 0 21902 76000 0 FreeSans 2000 90 0 0 VDD
port 11 nsew
flabel metal4 s 463 0 863 76000 0 FreeSans 2000 90 0 0 VSS
port 12 nsew
flabel metal4 s 21028 0 21428 76000 0 FreeSans 2000 90 0 0 VSS
port 12 nsew
flabel metal4 s 2306 39775 2467 40000 0 FreeSans 600 90 0 0 mimtop1
port 15 nsew
flabel metal4 s 2493 32001 2737 32321 0 FreeSans 600 90 0 0 mimtop2
port 17 nsew
flabel metal4 s 4189 39754 4348 40000 0 FreeSans 600 90 0 0 mimbot1
port 19 nsew
<< properties >>
string GDS_END 2086350
string GDS_FILE adc_top.gds.gz
string GDS_START 1755836
<< end >>
