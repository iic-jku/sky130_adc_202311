magic
tech sky130A
magscale 1 2
timestamp 1699054381
<< metal3 >>
rect -30 100 30 157
rect -30 -157 30 -100
<< rmetal3 >>
rect -30 -100 30 100
<< properties >>
string gencell sky130_fd_pr__res_generic_m3
string library sky130
string parameters w 0.3 l 1.0 m 1 nx 1 wmin 0.30 lmin 0.30 rho 0.047 val 156.666m dummy 0 dw 0.0 term 0.0 roverlap 0
<< end >>
