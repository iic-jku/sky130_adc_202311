magic
tech sky130A
magscale 1 2
timestamp 1698999411
<< nwell >>
rect -8 69 506 390
<< pwell >>
rect 98 -154 400 -16
rect 36 -240 462 -154
<< nmos >>
rect 186 -126 216 -42
rect 282 -126 312 -42
<< pmos >>
rect 90 106 120 266
rect 186 106 216 266
rect 282 106 312 266
rect 378 106 408 266
<< ndiff >>
rect 124 -67 186 -42
rect 124 -101 136 -67
rect 170 -101 186 -67
rect 124 -126 186 -101
rect 216 -67 282 -42
rect 216 -101 232 -67
rect 266 -101 282 -67
rect 216 -126 282 -101
rect 312 -67 374 -42
rect 312 -101 328 -67
rect 362 -101 374 -67
rect 312 -126 374 -101
<< pdiff >>
rect 28 237 90 266
rect 28 203 40 237
rect 74 203 90 237
rect 28 169 90 203
rect 28 135 40 169
rect 74 135 90 169
rect 28 106 90 135
rect 120 237 186 266
rect 120 203 136 237
rect 170 203 186 237
rect 120 169 186 203
rect 120 135 136 169
rect 170 135 186 169
rect 120 106 186 135
rect 216 237 282 266
rect 216 203 232 237
rect 266 203 282 237
rect 216 169 282 203
rect 216 135 232 169
rect 266 135 282 169
rect 216 106 282 135
rect 312 237 378 266
rect 312 203 328 237
rect 362 203 378 237
rect 312 169 378 203
rect 312 135 328 169
rect 362 135 378 169
rect 312 106 378 135
rect 408 237 470 266
rect 408 203 424 237
rect 458 203 470 237
rect 408 169 470 203
rect 408 135 424 169
rect 458 135 470 169
rect 408 106 470 135
<< ndiffc >>
rect 136 -101 170 -67
rect 232 -101 266 -67
rect 328 -101 362 -67
<< pdiffc >>
rect 40 203 74 237
rect 40 135 74 169
rect 136 203 170 237
rect 136 135 170 169
rect 232 203 266 237
rect 232 135 266 169
rect 328 203 362 237
rect 328 135 362 169
rect 424 203 458 237
rect 424 135 458 169
<< psubdiff >>
rect 62 -214 96 -180
rect 130 -214 164 -180
rect 198 -214 232 -180
rect 266 -214 300 -180
rect 334 -214 368 -180
rect 402 -214 436 -180
<< nsubdiff >>
rect 40 320 96 354
rect 130 320 164 354
rect 198 320 232 354
rect 266 320 300 354
rect 334 320 368 354
rect 402 320 458 354
<< psubdiffcont >>
rect 96 -214 130 -180
rect 164 -214 198 -180
rect 232 -214 266 -180
rect 300 -214 334 -180
rect 368 -214 402 -180
<< nsubdiffcont >>
rect 96 320 130 354
rect 164 320 198 354
rect 232 320 266 354
rect 300 320 334 354
rect 368 320 402 354
<< poly >>
rect 90 266 120 293
rect 186 266 216 292
rect 282 266 312 293
rect 378 266 408 292
rect 90 60 120 106
rect 186 66 216 106
rect 52 44 120 60
rect 52 10 70 44
rect 104 10 120 44
rect 52 0 120 10
rect 162 56 222 66
rect 282 60 312 106
rect 378 66 408 106
rect 162 22 178 56
rect 212 22 222 56
rect 162 6 222 22
rect 276 45 336 60
rect 276 11 286 45
rect 320 11 336 45
rect 186 -42 216 6
rect 276 1 336 11
rect 378 56 446 66
rect 378 22 396 56
rect 430 22 446 56
rect 378 6 446 22
rect 282 -42 312 1
rect 186 -152 216 -126
rect 282 -152 312 -126
<< polycont >>
rect 70 10 104 44
rect 178 22 212 56
rect 286 11 320 45
rect 396 22 430 56
<< locali >>
rect 40 320 96 354
rect 130 320 164 354
rect 198 320 232 354
rect 266 320 300 354
rect 334 320 368 354
rect 402 320 458 354
rect 40 237 74 320
rect 40 169 74 203
rect 40 102 74 135
rect 136 237 170 270
rect 136 169 170 203
rect 136 102 170 135
rect 232 237 266 270
rect 232 189 266 203
rect 232 102 266 135
rect 328 237 362 270
rect 328 169 362 203
rect 328 102 362 135
rect 424 237 458 320
rect 424 169 458 203
rect 424 102 458 135
rect 52 44 120 60
rect 52 10 70 44
rect 104 10 120 44
rect 52 0 120 10
rect 162 56 230 66
rect 162 22 178 56
rect 212 22 230 56
rect 162 6 230 22
rect 268 45 336 60
rect 268 10 286 45
rect 320 10 336 45
rect 268 1 336 10
rect 378 56 446 66
rect 378 22 396 56
rect 430 22 446 56
rect 378 6 446 22
rect 136 -67 170 -38
rect 136 -180 170 -101
rect 232 -67 266 -38
rect 232 -130 266 -122
rect 328 -67 362 -38
rect 328 -180 362 -101
rect 62 -214 96 -180
rect 130 -214 164 -180
rect 198 -214 232 -180
rect 266 -214 300 -180
rect 334 -214 368 -180
rect 402 -214 436 -180
<< viali >>
rect 232 169 266 189
rect 232 155 266 169
rect 70 10 104 44
rect 178 22 212 56
rect 286 11 320 44
rect 286 10 320 11
rect 396 22 430 56
rect 232 -101 266 -88
rect 232 -122 266 -101
<< metal1 >>
rect 223 198 275 204
rect 223 140 275 146
rect 22 84 476 112
rect 168 56 220 84
rect 386 56 438 84
rect 61 44 113 56
rect 61 10 70 44
rect 104 10 113 44
rect 168 22 178 56
rect 212 22 220 56
rect 168 10 220 22
rect 276 44 336 56
rect 276 10 286 44
rect 320 10 336 44
rect 386 22 396 56
rect 430 22 438 56
rect 386 10 438 22
rect 61 -19 113 10
rect 276 -19 336 10
rect 22 -47 476 -19
rect 223 -86 275 -76
rect 223 -147 275 -138
<< via1 >>
rect 223 189 275 198
rect 223 155 232 189
rect 232 155 266 189
rect 266 155 275 189
rect 223 146 275 155
rect 223 -88 275 -86
rect 223 -122 232 -88
rect 232 -122 266 -88
rect 266 -122 275 -88
rect 223 -138 275 -122
<< metal2 >>
rect 221 198 277 209
rect 221 146 223 198
rect 275 146 277 198
rect 221 135 277 146
rect 223 -86 275 135
rect 22 -138 223 -119
rect 275 -138 476 -119
rect 22 -147 476 -138
<< labels >>
flabel metal1 s 22 84 476 112 0 FreeSans 200 0 0 0 a
port 1 nsew
flabel metal1 s 22 -47 476 -19 0 FreeSans 200 0 0 0 b
port 2 nsew
flabel locali s 62 -214 436 -180 0 FreeSans 200 0 0 0 VSS
port 3 nsew
flabel locali s 40 320 458 354 0 FreeSans 200 0 0 0 VDD
port 4 nsew
flabel metal2 s 22 -147 476 -119 0 FreeSans 200 0 0 0 q
port 5 nsew
<< end >>
