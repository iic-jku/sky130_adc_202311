magic
tech sky130A
magscale 1 2
timestamp 1698131850
use pa_nfet_w30_nf4  pa_nfet_w30_nf4_0
timestamp 1698131850
transform 1 0 2430 0 1 -8
box -54 -85 2428 1821
use pa_nfet_w30_nf4  pa_nfet_w30_nf4_1
timestamp 1698131850
transform 1 0 54 0 1 -8
box -54 -85 2428 1821
<< end >>
