magic
tech sky130A
magscale 1 2
timestamp 1699972208
<< locali >>
rect 8025 8637 9130 8657
rect 8025 7677 8045 8637
rect 8533 7677 9130 8637
rect 8025 7657 9130 7677
rect 8025 779 9130 799
rect 8025 -181 8045 779
rect 8533 -181 9130 779
rect 8025 -201 9130 -181
rect 8025 -7079 9130 -7059
rect 8025 -8039 8045 -7079
rect 8533 -8039 9130 -7079
rect 8025 -8059 9130 -8039
rect 8025 -11693 9130 -11673
rect 8025 -12653 8045 -11693
rect 8533 -12653 9130 -11693
rect 8025 -12673 9130 -12653
rect 8025 -14685 9130 -14665
rect 8025 -15645 8045 -14685
rect 8533 -15645 9130 -14685
rect 8025 -15665 9130 -15645
rect 8025 -17677 9205 -17657
rect 8025 -18637 8045 -17677
rect 8533 -18637 9205 -17677
rect 8025 -18657 9205 -18637
rect -298 -21732 2 -21500
rect -298 -22072 -268 -21732
rect -28 -22072 2 -21732
rect -298 -22250 2 -22072
rect 20706 -21732 21006 -21500
rect 20706 -22072 20736 -21732
rect 20976 -22072 21006 -21732
rect 20706 -22250 21006 -22072
rect 4880 -25376 5180 -25144
rect 4880 -25716 4910 -25376
rect 5150 -25716 5180 -25376
rect 4880 -25894 5180 -25716
rect 15532 -25376 15832 -25144
rect 15532 -25716 15562 -25376
rect 15802 -25716 15832 -25376
rect 15532 -25894 15832 -25716
rect 7466 -29020 7766 -28788
rect 7466 -29360 7496 -29020
rect 7736 -29360 7766 -29020
rect 7466 -29538 7766 -29360
rect 12942 -29020 13242 -28788
rect 12942 -29360 12972 -29020
rect 13212 -29360 13242 -29020
rect 12942 -29538 13242 -29360
rect 8025 -32452 9210 -32432
rect 8025 -33162 8045 -32452
rect 8533 -32664 9210 -32452
rect 8533 -33004 8790 -32664
rect 9030 -33004 9210 -32664
rect 8533 -33162 9210 -33004
rect 8025 -33182 9210 -33162
rect 11648 -32664 11948 -32432
rect 11648 -33004 11678 -32664
rect 11918 -33004 11948 -32664
rect 11648 -33182 11948 -33004
rect 8025 -47211 9617 -47091
rect 8025 -47971 8045 -47211
rect 8533 -47932 9359 -47211
rect 9429 -47932 9617 -47211
rect 8533 -47971 9617 -47932
rect 8025 -48091 9617 -47971
rect 8025 -49390 8055 -49104
rect 8523 -49390 8553 -49104
rect 8025 -49420 8553 -49390
rect 8025 -50103 9617 -50083
rect 8025 -51063 8045 -50103
rect 8533 -50195 9617 -50103
rect 8533 -50971 9359 -50195
rect 9429 -50971 9617 -50195
rect 8533 -51063 9617 -50971
rect 8025 -51083 9617 -51063
rect 8025 -53095 9617 -53075
rect 8025 -54055 8045 -53095
rect 8533 -53187 9617 -53095
rect 8533 -53963 9359 -53187
rect 9429 -53963 9617 -53187
rect 8533 -54055 9617 -53963
rect 8025 -54075 9617 -54055
rect 8025 -57709 9441 -57689
rect 8025 -58669 8045 -57709
rect 8533 -57801 9441 -57709
rect 8533 -58577 9359 -57801
rect 9429 -58577 9441 -57801
rect 8533 -58669 9441 -58577
rect 8025 -58689 9441 -58669
rect 8025 -65567 9441 -65547
rect 8025 -66527 8045 -65567
rect 8533 -65659 9441 -65567
rect 8533 -66435 9359 -65659
rect 9429 -66435 9441 -65659
rect 8533 -66527 9441 -66435
rect 8025 -66547 9441 -66527
rect 8025 -73425 9441 -73405
rect 8025 -74385 8045 -73425
rect 8533 -73517 9441 -73425
rect 8533 -74293 9359 -73517
rect 9429 -74293 9441 -73517
rect 8533 -74385 9441 -74293
rect 8025 -74405 9441 -74385
rect 48854 -79210 49254 -79170
rect 48854 -79658 48894 -79210
rect 49214 -79658 49254 -79210
rect 48854 -79698 49254 -79658
<< viali >>
rect 8045 7677 8533 8637
rect 9359 7769 9429 8545
rect 8045 -181 8533 779
rect 9359 -89 9429 687
rect 8045 -8039 8533 -7079
rect 9359 -7947 9429 -7171
rect 8045 -12653 8533 -11693
rect 9359 -12561 9429 -11785
rect 8045 -15645 8533 -14685
rect 9359 -15553 9429 -14777
rect 8045 -18637 8533 -17677
rect 9358 -18545 9428 -17769
rect -268 -22072 -28 -21732
rect 20736 -22072 20976 -21732
rect 4910 -25716 5150 -25376
rect 15562 -25716 15802 -25376
rect 7496 -29360 7736 -29020
rect 12972 -29360 13212 -29020
rect 8045 -33162 8533 -32452
rect 8790 -33004 9030 -32664
rect 11678 -33004 11918 -32664
rect 8045 -47971 8533 -47211
rect 9359 -47932 9429 -47211
rect 8055 -49390 8523 -49050
rect 8045 -51063 8533 -50103
rect 9359 -50971 9429 -50195
rect 8045 -54055 8533 -53095
rect 9359 -53963 9429 -53187
rect 8045 -58669 8533 -57709
rect 9359 -58577 9429 -57801
rect 8045 -66527 8533 -65567
rect 9359 -66435 9429 -65659
rect 8045 -74385 8533 -73425
rect 9359 -74293 9429 -73517
rect 48894 -79658 49214 -79210
<< metal1 >>
rect 10104 11126 10604 11156
rect 10104 10886 10134 11126
rect 10574 10886 10604 11126
rect 10104 10856 10604 10886
rect 8025 8637 8553 8657
rect 8025 7677 8045 8637
rect 8533 8557 8553 8637
rect 8533 8545 9441 8557
rect 8533 7769 9359 8545
rect 9429 7769 9441 8545
rect 8533 7757 9441 7769
rect 8533 7677 8553 7757
rect 8025 7657 8553 7677
rect 10284 7314 10382 7626
rect 8025 779 8553 799
rect 8025 -181 8045 779
rect 8533 699 8553 779
rect 8533 687 9441 699
rect 8533 -89 9359 687
rect 9429 -89 9441 687
rect 8533 -101 9441 -89
rect 8533 -181 8553 -101
rect 8025 -201 8553 -181
rect 10284 -544 10382 -232
rect 8025 -7079 8553 -7059
rect 8025 -8039 8045 -7079
rect 8533 -7159 8553 -7079
rect 8533 -7171 9441 -7159
rect 8533 -7947 9359 -7171
rect 9429 -7947 9441 -7171
rect 8533 -7959 9441 -7947
rect 8533 -8039 8553 -7959
rect 8025 -8059 8553 -8039
rect 10284 -8402 10382 -8090
rect 8025 -11693 8553 -11673
rect 8025 -12653 8045 -11693
rect 8533 -11773 8553 -11693
rect 8533 -11785 9441 -11773
rect 8533 -12561 9359 -11785
rect 9429 -12561 9441 -11785
rect 8533 -12573 9441 -12561
rect 8533 -12653 8553 -12573
rect 8025 -12673 8553 -12653
rect 10284 -13016 10382 -12704
rect 8025 -14685 8553 -14665
rect 8025 -15645 8045 -14685
rect 8533 -14765 8553 -14685
rect 8533 -14777 9441 -14765
rect 8533 -15553 9359 -14777
rect 9429 -15553 9441 -14777
rect 8533 -15565 9441 -15553
rect 8533 -15645 8553 -15565
rect 8025 -15665 8553 -15645
rect 10284 -16008 10382 -15696
rect 8025 -17677 8553 -17657
rect 8025 -18637 8045 -17677
rect 8533 -17757 8553 -17677
rect 8533 -17769 9441 -17757
rect 8533 -18545 9358 -17769
rect 9428 -18545 9441 -17769
rect 8533 -18557 9441 -18545
rect 8533 -18637 8553 -18557
rect 8025 -18657 8553 -18637
rect 10284 -19000 10382 -18688
rect -298 -21732 2 -21702
rect -298 -22072 -268 -21732
rect -28 -22072 2 -21732
rect -298 -22102 2 -22072
rect 20706 -21732 21006 -21702
rect 20706 -22072 20736 -21732
rect 20976 -22072 21006 -21732
rect 20706 -22102 21006 -22072
rect 4880 -25376 5180 -25346
rect 4880 -25716 4910 -25376
rect 5150 -25716 5180 -25376
rect 4880 -25746 5180 -25716
rect 15532 -25376 15832 -25346
rect 15532 -25716 15562 -25376
rect 15802 -25716 15832 -25376
rect 15532 -25746 15832 -25716
rect 7466 -29020 7766 -28990
rect 7466 -29360 7496 -29020
rect 7736 -29360 7766 -29020
rect 7466 -29390 7766 -29360
rect 12942 -29020 13242 -28990
rect 12942 -29360 12972 -29020
rect 13212 -29360 13242 -29020
rect 12942 -29390 13242 -29360
rect 8025 -32452 8553 -32432
rect 8025 -33162 8045 -32452
rect 8533 -33162 8553 -32452
rect 8760 -32664 9060 -32634
rect 8760 -33004 8790 -32664
rect 9030 -33004 9060 -32664
rect 8760 -33034 9060 -33004
rect 11648 -32664 11948 -32634
rect 11648 -33004 11678 -32664
rect 11918 -33004 11948 -32664
rect 11648 -33034 11948 -33004
rect 8025 -33182 8553 -33162
rect 6337 -34866 8764 -34834
rect 6337 -34930 8037 -34866
rect 8025 -34938 8037 -34930
rect 8541 -34930 8764 -34866
rect 11944 -34930 14292 -34834
rect 8541 -34938 8553 -34930
rect 8025 -34950 8553 -34938
rect 18654 -35144 19043 -35114
rect 18654 -35378 18684 -35144
rect 6416 -35474 8922 -35378
rect 11944 -35474 14450 -35378
rect 17472 -35444 18684 -35378
rect 19013 -35444 19043 -35144
rect 17472 -35474 19043 -35444
rect 4790 -35528 4862 -35522
rect 4790 -35612 4796 -35528
rect 4856 -35612 4862 -35528
rect 4790 -36622 4862 -35612
rect 10318 -35528 10390 -35522
rect 10318 -35612 10324 -35528
rect 10384 -35612 10390 -35528
rect 10318 -36622 10390 -35612
rect 15846 -35528 15918 -35522
rect 15846 -35612 15852 -35528
rect 15912 -35612 15918 -35528
rect 15846 -36622 15918 -35612
rect 6220 -37433 9080 -37337
rect 11185 -37433 14519 -37337
rect 6189 -37893 8991 -37881
rect 6189 -38400 8037 -37893
rect 8541 -38316 8991 -37893
rect 11755 -38316 14519 -37881
rect 8541 -38400 9049 -38316
rect 6189 -38412 9049 -38400
rect 11717 -38412 14519 -38316
rect 3425 -39114 19043 -38860
rect 3425 -39244 18684 -39114
rect 18654 -39414 18684 -39244
rect 19013 -39414 19043 -39114
rect 18654 -39444 19043 -39414
rect 10326 -47060 10424 -46748
rect 8025 -47211 9441 -47191
rect 8025 -47971 8045 -47211
rect 8533 -47932 9359 -47211
rect 9429 -47932 9441 -47211
rect 8533 -47971 9441 -47932
rect 8025 -47991 9441 -47971
rect 8025 -49050 8553 -49020
rect 8025 -49390 8055 -49050
rect 8523 -49390 8553 -49050
rect 8025 -49450 8553 -49390
rect 10326 -50052 10424 -49740
rect 8025 -50103 8553 -50083
rect 8025 -51063 8045 -50103
rect 8533 -50183 8553 -50103
rect 8533 -50195 9441 -50183
rect 8533 -50971 9359 -50195
rect 9429 -50971 9441 -50195
rect 8533 -50983 9441 -50971
rect 8533 -51063 8553 -50983
rect 8025 -51083 8553 -51063
rect 10326 -53044 10424 -52732
rect 8025 -53095 8553 -53075
rect 8025 -54055 8045 -53095
rect 8533 -53175 8553 -53095
rect 8533 -53187 9441 -53175
rect 8533 -53963 9359 -53187
rect 9429 -53963 9441 -53187
rect 8533 -53975 9441 -53963
rect 8533 -54055 8553 -53975
rect 8025 -54075 8553 -54055
rect 10326 -57658 10424 -57346
rect 8025 -57709 8553 -57689
rect 8025 -58669 8045 -57709
rect 8533 -57789 8553 -57709
rect 8533 -57801 9441 -57789
rect 8533 -58577 9359 -57801
rect 9429 -58577 9441 -57801
rect 19361 -58006 19905 -57960
rect 8533 -58589 9441 -58577
rect 8533 -58669 8553 -58589
rect 8025 -58689 8553 -58669
rect 19361 -62224 19905 -62178
rect 19361 -64398 19905 -64352
rect 10326 -65516 10424 -65204
rect 8025 -65567 8553 -65547
rect 19361 -65550 19905 -65504
rect 8025 -66527 8045 -65567
rect 8533 -65647 8553 -65567
rect 8533 -65659 9441 -65647
rect 8533 -66435 9359 -65659
rect 9429 -66435 9441 -65659
rect 8533 -66447 9441 -66435
rect 8533 -66527 8553 -66447
rect 8025 -66547 8553 -66527
rect 19361 -66572 19905 -66526
rect 19361 -67594 19905 -67548
rect 10326 -73374 10424 -73062
rect 8025 -73425 8553 -73405
rect 8025 -74385 8045 -73425
rect 8533 -73505 8553 -73425
rect 8533 -73517 9441 -73505
rect 8533 -74293 9359 -73517
rect 9429 -74293 9441 -73517
rect 8533 -74305 9441 -74293
rect 8533 -74385 8553 -74305
rect 8025 -74405 8553 -74385
rect 9557 -79200 11157 -79170
rect 9557 -79668 9587 -79200
rect 11127 -79668 11157 -79200
rect 9557 -79698 11157 -79668
rect 48854 -79210 49254 -79170
rect 48854 -79658 48894 -79210
rect 49214 -79658 49254 -79210
rect 48854 -79698 49254 -79658
<< via1 >>
rect 10134 10886 10574 11126
rect 8045 7777 8533 8537
rect 9359 7769 9429 8545
rect 8045 -81 8533 679
rect 9359 -89 9429 687
rect 8045 -7939 8533 -7179
rect 9359 -7947 9429 -7171
rect 8045 -12553 8533 -11793
rect 9359 -12561 9429 -11785
rect 8045 -15545 8533 -14785
rect 9359 -15553 9429 -14777
rect 8045 -18537 8533 -17777
rect 9358 -18545 9428 -17769
rect -268 -22072 -28 -21732
rect 20736 -22072 20976 -21732
rect 4910 -25716 5150 -25376
rect 15562 -25716 15802 -25376
rect 7496 -29360 7736 -29020
rect 12972 -29360 13212 -29020
rect 8790 -33004 9030 -32664
rect 11678 -33004 11918 -32664
rect 8037 -34938 8541 -34866
rect 18684 -35444 19013 -35144
rect 4796 -35612 4856 -35528
rect 10324 -35612 10384 -35528
rect 15852 -35612 15912 -35528
rect 8037 -38400 8541 -37893
rect 18684 -39414 19013 -39114
rect 8045 -47971 8533 -47211
rect 9359 -47932 9429 -47211
rect 8045 -50963 8533 -50203
rect 9359 -50971 9429 -50195
rect 8045 -53955 8533 -53195
rect 9359 -53963 9429 -53187
rect 8045 -58569 8533 -57809
rect 9359 -58577 9429 -57801
rect 8045 -66427 8533 -65667
rect 9359 -66435 9429 -65659
rect 8045 -74285 8533 -73525
rect 9359 -74293 9429 -73517
rect 9587 -79668 11127 -79200
rect 48894 -79658 49214 -79210
<< metal2 >>
rect 8025 9874 8553 11156
rect 10104 11126 10604 11156
rect 10104 10886 10134 11126
rect 10574 10886 10604 11126
rect 10104 10856 10604 10886
rect 8025 9534 8055 9874
rect 8523 9534 8553 9874
rect 8025 8557 8553 9534
rect 8025 8545 9441 8557
rect 8025 8537 9359 8545
rect 8025 7777 8045 8537
rect 8533 7777 9359 8537
rect 8025 7769 9359 7777
rect 9429 7769 9441 8545
rect 8025 7757 9441 7769
rect 8025 2128 8553 7757
rect 8025 1788 8055 2128
rect 8523 1788 8553 2128
rect 8025 699 8553 1788
rect 8025 687 9441 699
rect 8025 679 9359 687
rect 8025 -81 8045 679
rect 8533 -81 9359 679
rect 8025 -89 9359 -81
rect 9429 -89 9441 687
rect 8025 -101 9441 -89
rect 8025 -5730 8553 -101
rect 8025 -6070 8055 -5730
rect 8523 -6070 8553 -5730
rect 8025 -7159 8553 -6070
rect 8025 -7171 9441 -7159
rect 8025 -7179 9359 -7171
rect 8025 -7939 8045 -7179
rect 8533 -7939 9359 -7179
rect 8025 -7947 9359 -7939
rect 9429 -7947 9441 -7171
rect 8025 -7959 9441 -7947
rect 8025 -10344 8553 -7959
rect 8025 -10684 8055 -10344
rect 8523 -10684 8553 -10344
rect 8025 -11773 8553 -10684
rect 8025 -11785 9441 -11773
rect 8025 -11793 9359 -11785
rect 8025 -12553 8045 -11793
rect 8533 -12553 9359 -11793
rect 8025 -12561 9359 -12553
rect 9429 -12561 9441 -11785
rect 8025 -12573 9441 -12561
rect 8025 -13336 8553 -12573
rect 8025 -13676 8055 -13336
rect 8523 -13676 8553 -13336
rect 8025 -14765 8553 -13676
rect 8025 -14777 9441 -14765
rect 8025 -14785 9359 -14777
rect 8025 -15545 8045 -14785
rect 8533 -15545 9359 -14785
rect 8025 -15553 9359 -15545
rect 9429 -15553 9441 -14777
rect 8025 -15565 9441 -15553
rect 8025 -16328 8553 -15565
rect 8025 -16668 8055 -16328
rect 8523 -16668 8553 -16328
rect 8025 -17757 8553 -16668
rect 8025 -17769 9441 -17757
rect 8025 -17777 9358 -17769
rect 8025 -18537 8045 -17777
rect 8533 -18537 9358 -17777
rect 8025 -18545 9358 -18537
rect 9428 -18545 9441 -17769
rect 8025 -18557 9441 -18545
rect 8025 -19320 8553 -18557
rect 8025 -19660 8055 -19320
rect 8523 -19660 8553 -19320
rect 8025 -19690 8553 -19660
rect -298 -21732 21006 -21702
rect -298 -22072 -268 -21732
rect -28 -22072 8055 -21732
rect 8523 -22072 20736 -21732
rect 20976 -22072 21006 -21732
rect -298 -22102 21006 -22072
rect 4880 -25376 15832 -25346
rect 4880 -25716 4910 -25376
rect 5150 -25716 8055 -25376
rect 8523 -25716 15562 -25376
rect 15802 -25716 15832 -25376
rect 4880 -25746 15832 -25716
rect 5026 -26392 5180 -26296
rect 15532 -26306 15682 -26296
rect 15672 -26382 15682 -26306
rect 15532 -26392 15682 -26382
rect 5026 -26450 5180 -26440
rect 5026 -26526 5036 -26450
rect 5026 -26536 5180 -26526
rect 15532 -26536 15682 -26440
rect 7466 -29020 13242 -28990
rect 7466 -29360 7496 -29020
rect 7736 -29360 8055 -29020
rect 8523 -29360 12972 -29020
rect 13212 -29360 13242 -29020
rect 7466 -29390 13242 -29360
rect 2520 -30870 2529 -30774
rect 2625 -30870 12402 -30774
rect 12498 -30870 12507 -30774
rect 12718 -32034 12814 -32025
rect 8025 -32664 11948 -32634
rect 8025 -33004 8055 -32664
rect 8523 -33004 8790 -32664
rect 9030 -33004 11678 -32664
rect 11918 -33004 11948 -32664
rect 8025 -33034 11948 -33004
rect 1089 -33157 1098 -33061
rect 1194 -33157 7057 -33061
rect 452 -34103 461 -34007
rect 557 -34103 566 -34007
rect 461 -36550 557 -34103
rect 4787 -35528 4865 -35522
rect 4787 -35612 4796 -35528
rect 4856 -35612 4865 -35528
rect 4787 -35618 4865 -35612
rect 6961 -36550 7057 -33157
rect 8025 -34866 8553 -34854
rect 8025 -34938 8037 -34866
rect 8541 -34938 8553 -34866
rect 8025 -35224 8055 -34938
rect 8523 -35224 8553 -34938
rect 7387 -36550 7473 -36546
rect 425 -36646 6227 -36550
rect 6960 -36555 7478 -36550
rect 6960 -36641 7387 -36555
rect 7473 -36641 7478 -36555
rect 6960 -36646 7478 -36641
rect 7387 -36650 7473 -36646
rect 3425 -36790 6227 -36694
rect 3425 -36934 6227 -36838
rect 3425 -36992 6227 -36982
rect 3425 -37068 5509 -36992
rect 6217 -37068 6227 -36992
rect 3425 -37078 6227 -37068
rect 8025 -37893 8553 -35224
rect 10315 -35528 10393 -35522
rect 10315 -35612 10324 -35528
rect 10384 -35612 10393 -35528
rect 10315 -35618 10393 -35612
rect 12718 -36550 12814 -32130
rect 18654 -35144 19043 -35114
rect 18654 -35444 18684 -35144
rect 19013 -35444 19043 -35144
rect 18654 -35474 19043 -35444
rect 15843 -35528 15921 -35522
rect 15843 -35612 15852 -35528
rect 15912 -35612 15921 -35528
rect 15843 -35618 15921 -35612
rect 8767 -36646 8776 -36550
rect 8872 -36646 11755 -36550
rect 12718 -36646 17283 -36550
rect 8953 -36790 11755 -36694
rect 14481 -36790 17283 -36694
rect 8953 -36934 11755 -36838
rect 14481 -36934 17283 -36838
rect 8953 -36992 11755 -36982
rect 8953 -37068 11037 -36992
rect 11745 -37068 11755 -36992
rect 8953 -37078 11755 -37068
rect 14481 -36992 17283 -36982
rect 14481 -37068 16565 -36992
rect 17273 -37068 17283 -36992
rect 14481 -37078 17283 -37068
rect 8025 -38400 8037 -37893
rect 8541 -38400 8553 -37893
rect 8025 -39096 8553 -38400
rect 8025 -39436 8055 -39096
rect 8523 -39436 8553 -39096
rect 8025 -39466 8553 -39436
rect 18654 -39114 19043 -39084
rect 18654 -39414 18684 -39114
rect 19013 -39414 19043 -39114
rect 18654 -39444 19043 -39414
rect 9754 -40930 10154 -40900
rect 9754 -41170 9784 -40930
rect 10124 -41170 10154 -40930
rect 9754 -41200 10154 -41170
rect 8025 -42088 8553 -42058
rect 8025 -42370 8055 -42088
rect 7523 -42428 8055 -42370
rect 8523 -42370 8553 -42088
rect 8523 -42428 13548 -42370
rect 7523 -42466 13548 -42428
rect 8025 -42901 8553 -42466
rect 8025 -47191 8553 -46901
rect 8025 -47211 9441 -47191
rect 8025 -47971 8045 -47211
rect 8533 -47932 9359 -47211
rect 9429 -47932 9441 -47211
rect 8533 -47971 8553 -47932
rect 8025 -47972 8553 -47971
rect 19542 -48852 19614 -47598
rect 20134 -48918 20206 -47598
rect 8025 -49080 8553 -49050
rect 8025 -49362 8055 -49080
rect 7449 -49420 8055 -49362
rect 8523 -49362 8553 -49080
rect 8523 -49420 13455 -49362
rect 7449 -49458 13455 -49420
rect 8025 -50183 8553 -49458
rect 8025 -50195 9441 -50183
rect 8025 -50203 9359 -50195
rect 8025 -50963 8045 -50203
rect 8533 -50963 9359 -50203
rect 8025 -50971 9359 -50963
rect 9429 -50971 9441 -50195
rect 8025 -50983 9441 -50971
rect 8025 -52072 8553 -50983
rect 8025 -52412 8055 -52072
rect 8523 -52412 8553 -52072
rect 8025 -53175 8553 -52412
rect 8025 -53187 9441 -53175
rect 8025 -53195 9359 -53187
rect 8025 -53955 8045 -53195
rect 8533 -53955 9359 -53195
rect 8025 -53963 9359 -53955
rect 9429 -53963 9441 -53187
rect 8025 -53975 9441 -53963
rect 8025 -55064 8553 -53975
rect 8025 -55404 8055 -55064
rect 8523 -55404 8553 -55064
rect 8025 -57789 8553 -55404
rect 8025 -57801 9441 -57789
rect 8025 -57809 9359 -57801
rect 8025 -58569 8045 -57809
rect 8533 -58569 9359 -57809
rect 8025 -58577 9359 -58569
rect 9429 -58577 9441 -57801
rect 8025 -58589 9441 -58577
rect 8025 -59678 8553 -58589
rect 8025 -60018 8055 -59678
rect 8523 -60018 8553 -59678
rect 8025 -65647 8553 -60018
rect 8025 -65659 9441 -65647
rect 8025 -65667 9359 -65659
rect 8025 -66427 8045 -65667
rect 8533 -66427 9359 -65667
rect 8025 -66435 9359 -66427
rect 9429 -66435 9441 -65659
rect 8025 -66447 9441 -66435
rect 8025 -67536 8553 -66447
rect 8025 -67876 8055 -67536
rect 8523 -67876 8553 -67536
rect 8025 -73505 8553 -67876
rect 8025 -73517 9441 -73505
rect 8025 -73525 9359 -73517
rect 8025 -74285 8045 -73525
rect 8533 -74285 9359 -73525
rect 8025 -74293 9359 -74285
rect 9429 -74293 9441 -73517
rect 8025 -74305 9441 -74293
rect 8025 -75394 8553 -74305
rect 8025 -75734 8055 -75394
rect 8523 -75734 8553 -75394
rect 8025 -75764 8553 -75734
rect 48854 -78482 49254 -78442
rect 48854 -78930 48894 -78482
rect 49214 -78930 49254 -78482
rect 48854 -78970 49254 -78930
rect 9557 -79200 11157 -79170
rect 9557 -79668 9587 -79200
rect 11127 -79668 11157 -79200
rect 9557 -79698 11157 -79668
rect 48854 -79210 49254 -79170
rect 48854 -79658 48894 -79210
rect 49214 -79658 49254 -79210
rect 48854 -79698 49254 -79658
<< via2 >>
rect 10134 10886 10574 11126
rect 8055 9534 8523 9874
rect 8055 1788 8523 2128
rect 8055 -6070 8523 -5730
rect 8055 -10684 8523 -10344
rect 8055 -13676 8523 -13336
rect 8055 -16668 8523 -16328
rect 8055 -19660 8523 -19320
rect 8055 -22072 8523 -21732
rect 16892 -22738 17272 -22662
rect 3436 -22882 3816 -22806
rect 8055 -25716 8523 -25376
rect 15292 -26382 15672 -26306
rect 5036 -26526 5416 -26450
rect 8055 -29360 8523 -29020
rect 12552 -30026 12932 -29950
rect 7776 -30170 8156 -30094
rect 2529 -30870 2625 -30774
rect 12402 -30870 12498 -30774
rect 12718 -32130 12814 -32034
rect 8055 -33004 8523 -32664
rect 1098 -33157 1194 -33061
rect 461 -34103 557 -34007
rect 4796 -35612 4856 -35528
rect 11258 -33670 11638 -33594
rect 9070 -33814 9450 -33738
rect 8055 -34938 8523 -34884
rect 8055 -35224 8523 -34938
rect 7387 -36641 7473 -36555
rect 5509 -37068 6217 -36992
rect 10324 -35612 10384 -35528
rect 18684 -35444 19013 -35144
rect 15852 -35612 15912 -35528
rect 8776 -36646 8872 -36550
rect 11037 -37068 11745 -36992
rect 16565 -37068 17273 -36992
rect 8055 -39436 8523 -39096
rect 18684 -39414 19013 -39114
rect 10964 -39982 11344 -39810
rect 9364 -40270 9744 -40098
rect 9784 -41170 10124 -40930
rect 8055 -42428 8523 -42088
rect 10564 -44182 10944 -44010
rect 8055 -49420 8523 -49080
rect 8055 -52412 8523 -52072
rect 8055 -55404 8523 -55064
rect 8055 -60018 8523 -59678
rect 8055 -67876 8523 -67536
rect 8055 -75734 8523 -75394
rect 48894 -78930 49214 -78482
rect 9587 -79668 11127 -79200
rect 48894 -79658 49214 -79210
<< metal3 >>
rect -76647 330811 -74139 331063
rect -76647 326320 -75618 330811
rect -74320 326320 -74139 330811
rect -76647 326022 -74139 326320
rect -76012 278877 -73504 279074
rect -76012 274271 -75580 278877
rect -73782 274271 -73504 278877
rect -76012 274033 -73504 274271
rect -76304 226863 -73804 227026
rect -76304 222257 -75711 226863
rect -73913 222257 -73804 226863
rect -76304 222026 -73804 222257
rect 10104 11126 10604 11156
rect 10104 10886 10134 11126
rect 10574 10886 10604 11126
rect 10104 10856 10604 10886
rect 8025 9874 8553 9904
rect 8025 9534 8055 9874
rect 8523 9534 8553 9874
rect 8025 9504 8553 9534
rect 8025 2128 8553 2158
rect 8025 1788 8055 2128
rect 8523 1788 8553 2128
rect 8025 1758 8553 1788
rect 8025 -5730 8553 -5700
rect 8025 -6070 8055 -5730
rect 8523 -6070 8553 -5730
rect 8025 -6100 8553 -6070
rect 8025 -10344 8553 -10314
rect 8025 -10684 8055 -10344
rect 8523 -10684 8553 -10344
rect 8025 -10714 8553 -10684
rect 8025 -13336 8553 -13306
rect 8025 -13676 8055 -13336
rect 8523 -13676 8553 -13336
rect 8025 -13706 8553 -13676
rect 8025 -16328 8553 -16298
rect 8025 -16668 8055 -16328
rect 8523 -16668 8553 -16328
rect 8025 -16698 8553 -16668
rect 8025 -19320 8553 -19290
rect 8025 -19660 8055 -19320
rect 8523 -19660 8553 -19320
rect 8025 -19690 8553 -19660
rect 8025 -21732 8553 -21702
rect 8025 -22072 8055 -21732
rect 8523 -22072 8553 -21732
rect 8025 -22102 8553 -22072
rect 3426 -22538 3826 -22508
rect 3426 -22806 3456 -22538
rect 3796 -22806 3826 -22538
rect 3426 -22882 3436 -22806
rect 3816 -22882 3826 -22806
rect 3426 -22892 3826 -22882
rect 16882 -22538 17282 -22508
rect 16882 -22662 16912 -22538
rect 17252 -22662 17282 -22538
rect 16882 -22738 16892 -22662
rect 17272 -22738 17282 -22662
rect 16882 -22862 16912 -22738
rect 17252 -22862 17282 -22738
rect 16882 -22892 17282 -22862
rect 8025 -25376 8553 -25346
rect 8025 -25716 8055 -25376
rect 8523 -25716 8553 -25376
rect 8025 -25746 8553 -25716
rect 5026 -26182 5426 -26152
rect 5026 -26450 5056 -26182
rect 5396 -26450 5426 -26182
rect 5026 -26526 5036 -26450
rect 5416 -26526 5426 -26450
rect 5026 -26536 5426 -26526
rect 15282 -26182 15682 -26152
rect 15282 -26306 15312 -26182
rect 15652 -26306 15682 -26182
rect 15282 -26382 15292 -26306
rect 15672 -26382 15682 -26306
rect 15282 -26506 15312 -26382
rect 15652 -26506 15682 -26382
rect 15282 -26536 15682 -26506
rect 8025 -29020 8553 -28990
rect 8025 -29360 8055 -29020
rect 8523 -29360 8553 -29020
rect 8025 -29390 8553 -29360
rect 7766 -29826 8166 -29796
rect 455 -30067 461 -29971
rect 557 -30067 563 -29971
rect 461 -34002 557 -30067
rect 7766 -30094 7796 -29826
rect 8136 -30094 8166 -29826
rect 7766 -30170 7776 -30094
rect 8156 -30170 8166 -30094
rect 7766 -30180 8166 -30170
rect 12542 -29826 12942 -29796
rect 12542 -29950 12572 -29826
rect 12912 -29950 12942 -29826
rect 12542 -30026 12552 -29950
rect 12932 -30026 12942 -29950
rect 12542 -30150 12572 -30026
rect 12912 -30150 12942 -30026
rect 12542 -30180 12942 -30150
rect 1092 -30828 1098 -30732
rect 1194 -30828 1200 -30732
rect 1098 -33056 1194 -30828
rect 2518 -30865 2524 -30769
rect 2630 -30865 2636 -30769
rect 12397 -30774 12503 -30769
rect 2524 -30870 2529 -30865
rect 2625 -30870 2630 -30865
rect 2524 -30875 2630 -30870
rect 12397 -30870 12402 -30774
rect 12498 -30870 12814 -30774
rect 12397 -30875 12503 -30870
rect 12718 -32029 12814 -30870
rect 12713 -32034 12819 -32029
rect 12713 -32130 12718 -32034
rect 12814 -32130 12819 -32034
rect 12713 -32135 12819 -32130
rect 8025 -32664 8553 -32634
rect 8025 -33004 8055 -32664
rect 8523 -33004 8553 -32664
rect 8025 -33034 8553 -33004
rect 1093 -33061 1199 -33056
rect 1093 -33157 1098 -33061
rect 1194 -33157 1199 -33061
rect 1093 -33162 1199 -33157
rect 9060 -33470 9460 -33440
rect 9060 -33738 9090 -33470
rect 9430 -33738 9460 -33470
rect 9060 -33814 9070 -33738
rect 9450 -33814 9460 -33738
rect 9060 -33824 9460 -33814
rect 11248 -33470 11648 -33440
rect 11248 -33594 11278 -33470
rect 11618 -33594 11648 -33470
rect 11248 -33670 11258 -33594
rect 11638 -33670 11648 -33594
rect 11248 -33794 11278 -33670
rect 11618 -33794 11648 -33670
rect 11248 -33824 11648 -33794
rect 456 -34007 562 -34002
rect 456 -34103 461 -34007
rect 557 -34103 562 -34007
rect 456 -34108 562 -34103
rect 8764 -34210 11944 -34114
rect 8764 -34402 11944 -34306
rect 8764 -34594 11944 -34498
rect 8764 -34786 11944 -34690
rect 8025 -34884 8553 -34854
rect 8025 -35224 8055 -34884
rect 8523 -35224 8553 -34884
rect 8025 -35254 8553 -35224
rect 18654 -35144 19043 -35114
rect 18654 -35444 18684 -35144
rect 19013 -35444 19043 -35144
rect 18654 -35474 19043 -35444
rect 8771 -36550 8877 -36545
rect 7382 -36555 8776 -36550
rect 7382 -36641 7387 -36555
rect 7473 -36641 8776 -36555
rect 7382 -36646 8776 -36641
rect 8872 -36646 8877 -36550
rect 8771 -36651 8877 -36646
rect 5499 -36706 6227 -36694
rect 5499 -36970 5511 -36706
rect 6215 -36970 6227 -36706
rect 5499 -36992 6227 -36970
rect 5499 -37068 5509 -36992
rect 6217 -37068 6227 -36992
rect 5499 -37078 6227 -37068
rect 11027 -36992 11755 -36982
rect 11027 -37068 11037 -36992
rect 11745 -37068 11755 -36992
rect 11027 -37090 11755 -37068
rect 11027 -37354 11039 -37090
rect 11743 -37354 11755 -37090
rect 11027 -37366 11755 -37354
rect 16555 -36992 17283 -36982
rect 16555 -37068 16565 -36992
rect 17273 -37068 17283 -36992
rect 16555 -37090 17283 -37068
rect 16555 -37354 16567 -37090
rect 17271 -37354 17283 -37090
rect 16555 -37366 17283 -37354
rect 8025 -39096 8553 -39066
rect 8025 -39436 8055 -39096
rect 8523 -39436 8553 -39096
rect 18654 -39114 19043 -39084
rect 8025 -39466 8553 -39436
rect 9354 -39296 9754 -39266
rect 9354 -39536 9384 -39296
rect 9724 -39536 9754 -39296
rect 9354 -40098 9754 -39536
rect 9354 -40270 9364 -40098
rect 9744 -40270 9754 -40098
rect 9354 -40288 9754 -40270
rect 10954 -39296 11354 -39266
rect 10954 -39536 10984 -39296
rect 11324 -39536 11354 -39296
rect 18654 -39414 18684 -39114
rect 19013 -39414 19043 -39114
rect 18654 -39444 19043 -39414
rect 10954 -39810 11354 -39536
rect 10954 -39982 10964 -39810
rect 11344 -39982 11354 -39810
rect 10954 -40288 11354 -39982
rect 9754 -40930 10154 -40900
rect 9754 -41170 9784 -40930
rect 10124 -41170 10154 -40930
rect 8025 -42088 8553 -42058
rect 8025 -42428 8055 -42088
rect 8523 -42428 8553 -42088
rect 8025 -42458 8553 -42428
rect 9754 -44192 10154 -41170
rect 10554 -40930 10954 -40900
rect 10554 -41170 10584 -40930
rect 10924 -41170 10954 -40930
rect 10554 -44010 10954 -41170
rect 10554 -44182 10564 -44010
rect 10944 -44182 10954 -44010
rect 10554 -44192 10954 -44182
rect 8025 -49080 8553 -49050
rect 8025 -49420 8055 -49080
rect 8523 -49420 8553 -49080
rect 8025 -49450 8553 -49420
rect 8025 -52072 8553 -52042
rect 8025 -52412 8055 -52072
rect 8523 -52412 8553 -52072
rect 8025 -52442 8553 -52412
rect 8025 -55064 8553 -55034
rect 8025 -55404 8055 -55064
rect 8523 -55404 8553 -55064
rect 8025 -55434 8553 -55404
rect 8025 -59678 8553 -59648
rect 8025 -60018 8055 -59678
rect 8523 -60018 8553 -59678
rect 8025 -60048 8553 -60018
rect 8025 -67536 8553 -67506
rect 8025 -67876 8055 -67536
rect 8523 -67876 8553 -67536
rect 8025 -67906 8553 -67876
rect 18960 -69887 20784 -69838
rect 18856 -70962 20843 -69887
rect 18856 -72072 18982 -70962
rect 20728 -72072 20843 -70962
rect 18856 -72200 20843 -72072
rect 8025 -75394 8553 -75364
rect 8025 -75734 8055 -75394
rect 8523 -75734 8553 -75394
rect 8025 -75764 8553 -75734
rect 18856 -76276 20843 -76270
rect -7912 -76382 -5927 -76378
rect -7912 -76384 18856 -76382
rect -5927 -78263 18856 -76384
rect -5927 -78369 20843 -78263
rect -7912 -78375 -5927 -78369
rect 48854 -78482 49254 -78442
rect 48854 -78930 48894 -78482
rect 49214 -78930 49254 -78482
rect 48854 -78970 49254 -78930
rect 9557 -79200 11157 -79170
rect 9557 -79668 9587 -79200
rect 11127 -79668 11157 -79200
rect 9557 -79698 11157 -79668
rect 48854 -79210 49254 -79170
rect 48854 -79658 48894 -79210
rect 49214 -79658 49254 -79210
rect 48854 -79698 49254 -79658
rect -40129 -163739 -32599 -162711
rect -40129 -164544 -39416 -163739
rect -78304 -167004 -39416 -164544
rect -40129 -174544 -39416 -167004
rect -78304 -177004 -39416 -174544
rect -40129 -180752 -39416 -177004
rect -33277 -180752 -32599 -163739
rect -40129 -182076 -32599 -180752
rect 71128 -211254 71134 -206454
rect 75934 -211254 75940 -206454
rect 81128 -211254 81134 -206454
rect 85934 -211254 85940 -206454
rect -76304 -219640 -59804 -219374
rect -76304 -223736 -63767 -219640
rect -60342 -223736 -59804 -219640
rect -76304 -224374 -59804 -223736
rect 71134 -228320 75934 -211254
rect 81134 -228320 85934 -211254
<< via3 >>
rect -75618 326320 -74320 330811
rect -75580 274271 -73782 278877
rect -75711 222257 -73913 226863
rect 10134 10886 10574 11126
rect 8055 9534 8523 9874
rect 8055 1788 8523 2128
rect 8055 -6070 8523 -5730
rect 8055 -10684 8523 -10344
rect 8055 -13676 8523 -13336
rect 8055 -16668 8523 -16328
rect 8055 -19660 8523 -19320
rect 8055 -22072 8523 -21732
rect 3456 -22806 3796 -22538
rect 3456 -22862 3796 -22806
rect 16912 -22662 17252 -22538
rect 16912 -22738 17252 -22662
rect 16912 -22862 17252 -22738
rect 8055 -25716 8523 -25376
rect 5056 -26450 5396 -26182
rect 5056 -26506 5396 -26450
rect 15312 -26306 15652 -26182
rect 15312 -26382 15652 -26306
rect 15312 -26506 15652 -26382
rect 8055 -29360 8523 -29020
rect 461 -30067 557 -29971
rect 7796 -30094 8136 -29826
rect 7796 -30150 8136 -30094
rect 12572 -29950 12912 -29826
rect 12572 -30026 12912 -29950
rect 12572 -30150 12912 -30026
rect 1098 -30828 1194 -30732
rect 2524 -30774 2630 -30769
rect 2524 -30865 2529 -30774
rect 2529 -30865 2625 -30774
rect 2625 -30865 2630 -30774
rect 8055 -33004 8523 -32664
rect 9090 -33738 9430 -33470
rect 9090 -33794 9430 -33738
rect 11278 -33594 11618 -33470
rect 11278 -33670 11618 -33594
rect 11278 -33794 11618 -33670
rect 5838 -34198 6214 -34126
rect 14494 -34198 14870 -34126
rect 5838 -34390 6214 -34318
rect 14494 -34390 14870 -34318
rect 5838 -34582 6214 -34510
rect 14494 -34582 14870 -34510
rect 5838 -34774 6214 -34702
rect 14494 -34774 14870 -34702
rect 8055 -35224 8523 -34884
rect 18684 -35444 19013 -35144
rect 5836 -35800 6216 -35724
rect 11364 -35800 11744 -35724
rect 14492 -35800 14872 -35724
rect 5036 -35992 5416 -35916
rect 8964 -35992 9344 -35916
rect 15292 -35992 15672 -35916
rect 4236 -36184 4616 -36108
rect 9764 -36184 10144 -36108
rect 16092 -36184 16472 -36108
rect 3436 -36376 3816 -36300
rect 10564 -36376 10944 -36300
rect 16892 -36376 17272 -36300
rect 5511 -36970 6215 -36706
rect 11039 -37354 11743 -37090
rect 16567 -37354 17271 -37090
rect 8055 -39436 8523 -39096
rect 9384 -39536 9724 -39296
rect 10984 -39536 11324 -39296
rect 18684 -39414 19013 -39114
rect 9784 -41170 10124 -40930
rect 8055 -42428 8523 -42088
rect 10584 -41170 10924 -40930
rect 8055 -49420 8523 -49080
rect 8055 -52412 8523 -52072
rect 8055 -55404 8523 -55064
rect 18982 -72072 20728 -70962
rect 8055 -75734 8523 -75394
rect -7912 -78369 -5927 -76384
rect 18856 -78263 20843 -76276
rect 48894 -78930 49214 -78482
rect 9587 -79668 11127 -79200
rect 48894 -79658 49214 -79210
rect -39416 -180752 -33277 -163739
rect 71134 -211254 75934 -206454
rect 81134 -211254 85934 -206454
rect -63767 -223736 -60342 -219640
<< metal4 >>
rect -76647 330811 -74139 331063
rect -76647 326320 -75618 330811
rect -74320 326320 -74139 330811
rect -76647 326022 -74139 326320
rect -76012 278877 -73504 279074
rect -76012 274271 -75580 278877
rect -73782 274271 -73504 278877
rect -76012 274033 -73504 274271
rect -76304 226863 -73804 227026
rect -76304 222257 -75711 226863
rect -73913 222257 -73804 226863
rect -76304 222026 -73804 222257
rect 8025 11126 12610 11156
rect 8025 10886 8055 11126
rect 8523 10886 10134 11126
rect 10574 10886 12610 11126
rect 8025 10856 12610 10886
rect 8025 10626 12610 10656
rect 8025 10386 9884 10626
rect 10824 10386 12112 10626
rect 12580 10386 12610 10626
rect 8025 10356 12610 10386
rect 8025 9874 8553 9904
rect 8025 9534 8055 9874
rect 8523 9534 8553 9874
rect 8025 9504 8553 9534
rect 8025 2128 8553 2158
rect 8025 1788 8055 2128
rect 8523 1788 8553 2128
rect 8025 1758 8553 1788
rect 8025 -5730 8553 -5700
rect 8025 -6070 8055 -5730
rect 8523 -6070 8553 -5730
rect 8025 -6100 8553 -6070
rect 8025 -10344 8553 -10314
rect 8025 -10684 8055 -10344
rect 8523 -10684 8553 -10344
rect 8025 -10714 8553 -10684
rect 8025 -13336 8553 -13306
rect 8025 -13676 8055 -13336
rect 8523 -13676 8553 -13336
rect 8025 -13706 8553 -13676
rect 8025 -16328 8553 -16298
rect 8025 -16668 8055 -16328
rect 8523 -16668 8553 -16328
rect 8025 -16698 8553 -16668
rect 8025 -19320 8553 -19290
rect 8025 -19660 8055 -19320
rect 8523 -19660 8553 -19320
rect 8025 -19690 8553 -19660
rect 8025 -21732 8553 -21702
rect 8025 -22072 8055 -21732
rect 8523 -22072 8553 -21732
rect 8025 -22102 8553 -22072
rect 3426 -22538 3826 -22508
rect 3426 -22862 3456 -22538
rect 3796 -22862 3826 -22538
rect 3426 -22892 3826 -22862
rect 16882 -22538 17282 -22508
rect 16882 -22862 16912 -22538
rect 17252 -22862 17282 -22538
rect 16882 -22892 17282 -22862
rect 8025 -25376 8553 -25346
rect 8025 -25716 8055 -25376
rect 8523 -25716 8553 -25376
rect 8025 -25746 8553 -25716
rect 4226 -26182 5426 -26152
rect 4226 -26506 4256 -26182
rect 4596 -26506 5056 -26182
rect 5396 -26506 5426 -26182
rect 4226 -26536 5426 -26506
rect 15282 -26182 16482 -26152
rect 15282 -26506 15312 -26182
rect 15652 -26506 16112 -26182
rect 16452 -26506 16482 -26182
rect 15282 -26536 16482 -26506
rect 8025 -29020 8553 -28990
rect 8025 -29360 8055 -29020
rect 8523 -29360 8553 -29020
rect 8025 -29390 8553 -29360
rect 5026 -29826 8166 -29796
rect 5026 -30150 5056 -29826
rect 5396 -30150 7796 -29826
rect 8136 -30150 8166 -29826
rect 5026 -30180 8166 -30150
rect 12542 -29826 15682 -29796
rect 12542 -30150 12572 -29826
rect 12912 -30150 15312 -29826
rect 15652 -30150 15682 -29826
rect 12542 -30180 15682 -30150
rect 8025 -32664 8553 -32634
rect 8025 -33004 8055 -32664
rect 8523 -33004 8553 -32664
rect 8025 -33034 8553 -33004
rect 5826 -33470 9460 -33440
rect 5826 -33794 5856 -33470
rect 6196 -33794 9090 -33470
rect 9430 -33794 9460 -33470
rect 5826 -33824 9460 -33794
rect 11248 -33470 14882 -33440
rect 11248 -33794 11278 -33470
rect 11618 -33794 14512 -33470
rect 14852 -33794 14882 -33470
rect 11248 -33824 14882 -33794
rect 3236 -34126 17472 -34114
rect 3236 -34198 5838 -34126
rect 6214 -34198 14494 -34126
rect 14870 -34198 17472 -34126
rect 3236 -34210 17472 -34198
rect 3236 -34318 17472 -34306
rect 3236 -34390 5838 -34318
rect 6214 -34390 14494 -34318
rect 14870 -34390 17472 -34318
rect 3236 -34402 17472 -34390
rect 3236 -34510 17472 -34498
rect 3236 -34582 5838 -34510
rect 6214 -34582 14494 -34510
rect 14870 -34582 17472 -34510
rect 3236 -34594 17472 -34582
rect 3236 -34702 17472 -34690
rect 3236 -34774 5838 -34702
rect 6214 -34774 14494 -34702
rect 14870 -34774 17472 -34702
rect 3236 -34786 17472 -34774
rect 8025 -34884 8553 -34854
rect 8025 -35224 8055 -34884
rect 8523 -35224 8553 -34884
rect 8025 -35254 8553 -35224
rect 18654 -35144 19043 -35114
rect 5826 -35456 6226 -35426
rect 5026 -35648 5426 -35618
rect 4226 -35840 4626 -35810
rect 3426 -36032 3826 -36002
rect 3426 -36300 3456 -36032
rect 3796 -36300 3826 -36032
rect 4226 -36108 4256 -35840
rect 4596 -36108 4626 -35840
rect 5026 -35916 5056 -35648
rect 5396 -35916 5426 -35648
rect 5826 -35724 5856 -35456
rect 6196 -35724 6226 -35456
rect 11354 -35456 11754 -35426
rect 5826 -35800 5836 -35724
rect 6216 -35800 6226 -35724
rect 5826 -35810 6226 -35800
rect 8954 -35648 9354 -35618
rect 5026 -35992 5036 -35916
rect 5416 -35992 5426 -35916
rect 5026 -36002 5426 -35992
rect 8954 -35916 8984 -35648
rect 9324 -35916 9354 -35648
rect 11354 -35724 11384 -35456
rect 11724 -35724 11754 -35456
rect 11354 -35800 11364 -35724
rect 11744 -35800 11754 -35724
rect 11354 -35810 11754 -35800
rect 14482 -35456 14882 -35426
rect 14482 -35724 14512 -35456
rect 14852 -35724 14882 -35456
rect 18654 -35444 18684 -35144
rect 19013 -35444 19043 -35144
rect 18654 -35474 19043 -35444
rect 14482 -35800 14492 -35724
rect 14872 -35800 14882 -35724
rect 14482 -35810 14882 -35800
rect 15282 -35648 15682 -35618
rect 8954 -35992 8964 -35916
rect 9344 -35992 9354 -35916
rect 8954 -36002 9354 -35992
rect 9754 -35840 10154 -35810
rect 4226 -36184 4236 -36108
rect 4616 -36184 4626 -36108
rect 4226 -36194 4626 -36184
rect 9754 -36108 9784 -35840
rect 10124 -36108 10154 -35840
rect 15282 -35916 15312 -35648
rect 15652 -35916 15682 -35648
rect 15282 -35992 15292 -35916
rect 15672 -35992 15682 -35916
rect 15282 -36002 15682 -35992
rect 16082 -35840 16482 -35810
rect 9754 -36184 9764 -36108
rect 10144 -36184 10154 -36108
rect 9754 -36194 10154 -36184
rect 10554 -36032 10954 -36002
rect 3426 -36376 3436 -36300
rect 3816 -36376 3826 -36300
rect 3426 -36386 3826 -36376
rect 10554 -36300 10584 -36032
rect 10924 -36300 10954 -36032
rect 16082 -36108 16112 -35840
rect 16452 -36108 16482 -35840
rect 16082 -36184 16092 -36108
rect 16472 -36184 16482 -36108
rect 16082 -36194 16482 -36184
rect 16882 -36032 17282 -36002
rect 10554 -36376 10564 -36300
rect 10944 -36376 10954 -36300
rect 10554 -36386 10954 -36376
rect 16882 -36300 16912 -36032
rect 17252 -36300 17282 -36032
rect 16882 -36376 16892 -36300
rect 17272 -36376 17282 -36300
rect 16882 -36386 17282 -36376
rect -2021 -36706 22729 -36694
rect -2021 -36970 5511 -36706
rect 6215 -36718 22729 -36706
rect 6215 -36958 21436 -36718
rect 21788 -36958 22729 -36718
rect 6215 -36970 22729 -36958
rect -2021 -36982 22729 -36970
rect -2021 -37090 22729 -37078
rect -2021 -37354 11039 -37090
rect 11743 -37354 16567 -37090
rect 17271 -37102 22729 -37090
rect 17271 -37342 17958 -37102
rect 18310 -37342 22729 -37102
rect 17271 -37354 22729 -37342
rect -2021 -37366 22729 -37354
rect 8025 -39096 8553 -39066
rect 8025 -39436 8055 -39096
rect 8523 -39436 8553 -39096
rect 18654 -39114 19043 -39084
rect 8025 -39466 8553 -39436
rect 8954 -39296 9754 -39266
rect 8954 -39536 8984 -39296
rect 9324 -39536 9384 -39296
rect 9724 -39536 9754 -39296
rect 8954 -39566 9754 -39536
rect 10954 -39296 11754 -39266
rect 10954 -39536 10984 -39296
rect 11324 -39536 11384 -39296
rect 11724 -39536 11754 -39296
rect 18654 -39414 18684 -39114
rect 19013 -39414 19043 -39114
rect 18654 -39444 19043 -39414
rect 10954 -39566 11754 -39536
rect 9754 -40930 10154 -40900
rect 9754 -41170 9784 -40930
rect 10124 -41170 10154 -40930
rect 9754 -41200 10154 -41170
rect 10554 -40930 10954 -40900
rect 10554 -41170 10584 -40930
rect 10924 -41170 10954 -40930
rect 10554 -41200 10954 -41170
rect 8025 -42088 8553 -42058
rect 8025 -42428 8055 -42088
rect 8523 -42428 8553 -42088
rect 8025 -42458 8553 -42428
rect 18654 -46853 20913 -46823
rect 18654 -47273 18684 -46853
rect 19013 -47273 20463 -46853
rect 20883 -47273 20913 -46853
rect 18654 -47303 20913 -47273
rect 17934 -47628 18334 -47598
rect 8025 -49080 8553 -49050
rect -1006 -49274 -526 -49244
rect -1006 -50214 -976 -49274
rect -556 -50214 -526 -49274
rect -1006 -50244 -526 -50214
rect 2198 -49274 2678 -49244
rect 2198 -50214 2228 -49274
rect 2648 -50214 2678 -49274
rect 8025 -49420 8055 -49080
rect 8523 -49420 8553 -49080
rect 8025 -49450 8553 -49420
rect 2198 -50244 2678 -50214
rect 17934 -50022 17964 -47628
rect 18304 -50022 18334 -47628
rect 17934 -50244 18334 -50022
rect 21412 -47628 21812 -47598
rect 21412 -50022 21442 -47628
rect 21782 -50022 21812 -47628
rect 21412 -50244 21812 -50022
rect 8025 -52072 8553 -52042
rect 8025 -52412 8055 -52072
rect 8523 -52412 8553 -52072
rect 8025 -52442 8553 -52412
rect 8025 -55064 8553 -55034
rect 8025 -55404 8055 -55064
rect 8523 -55404 8553 -55064
rect 8025 -55434 8553 -55404
rect 8025 -59678 8553 -59648
rect 8025 -60018 8055 -59678
rect 8523 -60018 8553 -59678
rect 8025 -60048 8553 -60018
rect 8025 -67536 8553 -67506
rect 8025 -67876 8055 -67536
rect 8523 -67876 8553 -67536
rect 8025 -67906 8553 -67876
rect 18856 -70962 20844 -70864
rect 18856 -72072 18982 -70962
rect 20728 -72072 20844 -70962
rect 18856 -72200 20844 -72072
rect -1006 -75394 21714 -75364
rect -1006 -75734 -976 -75394
rect -556 -75734 2228 -75394
rect 2648 -75734 8055 -75394
rect 8523 -75734 18060 -75394
rect 18480 -75734 21714 -75394
rect -1006 -75764 21714 -75734
rect -7913 -76384 -5926 -76383
rect -7913 -78369 -7912 -76384
rect -5927 -78369 -5926 -76384
rect 18855 -78263 18856 -78262
rect 20843 -78263 20844 -78262
rect 18855 -78264 20844 -78263
rect -7913 -124560 -5926 -78369
rect 6626 -78472 49254 -78442
rect 6626 -78940 9884 -78472
rect 10824 -78940 12112 -78472
rect 12580 -78482 49254 -78472
rect 12580 -78493 48894 -78482
rect 12580 -78884 27900 -78493
rect 35299 -78884 48894 -78493
rect 12580 -78930 48894 -78884
rect 49214 -78930 49254 -78482
rect 12580 -78940 49254 -78930
rect 6626 -78970 49254 -78940
rect 6626 -79200 49254 -79170
rect 6626 -79668 8055 -79200
rect 8523 -79668 9587 -79200
rect 11127 -79210 49254 -79200
rect 11127 -79230 48894 -79210
rect 11127 -79621 37890 -79230
rect 45289 -79621 48894 -79230
rect 11127 -79658 48894 -79621
rect 49214 -79658 49254 -79210
rect 11127 -79668 49254 -79658
rect 6626 -79698 49254 -79668
rect -40129 -163739 -32599 -162711
rect -40129 -180752 -39416 -163739
rect -33277 -180752 -32599 -163739
rect -40129 -182076 -32599 -180752
rect -63991 -219640 -60155 -219417
rect -63991 -223736 -63767 -219640
rect -60342 -223736 -60155 -219640
rect -63991 -224071 -60155 -223736
<< via4 >>
rect -75618 326320 -74320 330811
rect -75580 274271 -73782 278877
rect -75711 222257 -73913 226863
rect 8055 10886 8523 11126
rect 9884 10386 10824 10626
rect 12112 10386 12580 10626
rect 8055 9534 8523 9874
rect 8055 1788 8523 2128
rect 8055 -6070 8523 -5730
rect 8055 -10684 8523 -10344
rect 8055 -13676 8523 -13336
rect 8055 -16668 8523 -16328
rect 8055 -19660 8523 -19320
rect 8055 -22072 8523 -21732
rect 3456 -22862 3796 -22538
rect 16912 -22862 17252 -22538
rect 8055 -25716 8523 -25376
rect 4256 -26506 4596 -26182
rect 16112 -26506 16452 -26182
rect 8055 -29360 8523 -29020
rect 349 -29971 669 -29859
rect 349 -30067 461 -29971
rect 461 -30067 557 -29971
rect 557 -30067 669 -29971
rect 349 -30179 669 -30067
rect 5056 -30150 5396 -29826
rect 15312 -30150 15652 -29826
rect 986 -30732 1306 -30620
rect 986 -30828 1098 -30732
rect 1098 -30828 1194 -30732
rect 1194 -30828 1306 -30732
rect 986 -30940 1306 -30828
rect 2417 -30769 2737 -30657
rect 2417 -30865 2524 -30769
rect 2524 -30865 2630 -30769
rect 2630 -30865 2737 -30769
rect 2417 -30977 2737 -30865
rect 8055 -33004 8523 -32664
rect 5856 -33794 6196 -33470
rect 14512 -33794 14852 -33470
rect 8055 -35224 8523 -34884
rect 3456 -36300 3796 -36032
rect 4256 -36108 4596 -35840
rect 5056 -35916 5396 -35648
rect 5856 -35724 6196 -35456
rect 5856 -35780 6196 -35724
rect 5056 -35972 5396 -35916
rect 8984 -35916 9324 -35648
rect 11384 -35724 11724 -35456
rect 11384 -35780 11724 -35724
rect 14512 -35724 14852 -35456
rect 18684 -35444 19013 -35144
rect 14512 -35780 14852 -35724
rect 8984 -35972 9324 -35916
rect 4256 -36164 4596 -36108
rect 9784 -36108 10124 -35840
rect 15312 -35916 15652 -35648
rect 15312 -35972 15652 -35916
rect 9784 -36164 10124 -36108
rect 3456 -36356 3796 -36300
rect 10584 -36300 10924 -36032
rect 16112 -36108 16452 -35840
rect 16112 -36164 16452 -36108
rect 10584 -36356 10924 -36300
rect 16912 -36300 17252 -36032
rect 16912 -36356 17252 -36300
rect 21436 -36958 21788 -36718
rect 17958 -37342 18310 -37102
rect 8055 -39436 8523 -39096
rect 8984 -39536 9324 -39296
rect 11384 -39536 11724 -39296
rect 18684 -39414 19013 -39114
rect 9784 -41170 10124 -40930
rect 10584 -41170 10924 -40930
rect 8055 -42428 8523 -42088
rect 18684 -47273 19013 -46853
rect 20463 -47273 20883 -46853
rect -976 -50214 -556 -49274
rect 2228 -50214 2648 -49274
rect 8055 -49420 8523 -49080
rect 17964 -50022 18304 -47628
rect 21442 -50022 21782 -47628
rect 8055 -52412 8523 -52072
rect 8055 -55404 8523 -55064
rect 8055 -60018 8523 -59678
rect 8055 -67876 8523 -67536
rect 18982 -72072 20728 -70962
rect -976 -75734 -556 -75394
rect 2228 -75734 2648 -75394
rect 8055 -75734 8523 -75394
rect 18060 -75734 18480 -75394
rect 18855 -76276 20844 -76275
rect 18855 -78262 18856 -76276
rect 18856 -78262 20843 -76276
rect 20843 -78262 20844 -76276
rect 9884 -78940 10824 -78472
rect 12112 -78940 12580 -78472
rect 27900 -78884 35299 -78493
rect 8055 -79668 8523 -79200
rect 37890 -79621 45289 -79230
rect -7913 -125347 -5926 -124560
rect -39416 -180752 -33277 -163739
rect 71133 -206454 75935 -206453
rect 71133 -211254 71134 -206454
rect 71134 -211254 75934 -206454
rect 75934 -211254 75935 -206454
rect 71133 -211255 75935 -211254
rect 81133 -206454 85935 -206453
rect 81133 -211254 81134 -206454
rect 81134 -211254 85934 -206454
rect 85934 -211254 85935 -206454
rect 81133 -211255 85935 -211254
rect -63767 -223736 -60342 -219640
<< metal5 >>
rect -76647 330811 -74139 331063
rect -76647 326320 -75618 330811
rect -74320 328634 -74139 330811
rect -74320 328314 -54182 328634
rect -74320 326320 -74139 328314
rect -76647 326022 -74139 326320
rect -76012 278877 -73504 279074
rect -76012 274271 -75580 278877
rect -73782 276691 -73504 278877
rect -73782 276354 -55909 276691
rect -73782 274271 -73504 276354
rect -76012 274033 -73504 274271
rect -76304 226863 -73804 227026
rect -76304 222257 -75711 226863
rect -73913 225775 -73804 226863
rect -73913 225455 -57660 225775
rect -73913 222257 -73804 225455
rect -76304 222026 -73804 222257
rect -57980 -4564 -57660 225455
rect -56246 -3227 -55909 276354
rect -54502 -1563 -54182 328314
rect 8025 11126 8553 11156
rect 8025 10886 8055 11126
rect 8523 10886 8553 11126
rect 8025 9874 8553 10886
rect 9854 10626 10854 10856
rect 9854 10386 9884 10626
rect 10824 10386 10854 10626
rect 9854 10356 10854 10386
rect 12082 10626 12610 11156
rect 12082 10386 12112 10626
rect 12580 10386 12610 10626
rect 8025 9534 8055 9874
rect 8523 9534 8553 9874
rect 8025 2128 8553 9534
rect 8025 1788 8055 2128
rect 8523 1788 8553 2128
rect -54502 -1883 2737 -1563
rect -56246 -3564 1651 -3227
rect -57980 -4884 669 -4564
rect 349 -29835 669 -4884
rect 325 -29859 693 -29835
rect 325 -30179 349 -29859
rect 669 -30179 693 -29859
rect 325 -30203 693 -30179
rect 1314 -30596 1651 -3564
rect 962 -30620 1651 -30596
rect 962 -30940 986 -30620
rect 1306 -30940 1651 -30620
rect 2417 -30633 2737 -1883
rect 8025 -5730 8553 1788
rect 8025 -6070 8055 -5730
rect 8523 -6070 8553 -5730
rect 8025 -10344 8553 -6070
rect 8025 -10684 8055 -10344
rect 8523 -10684 8553 -10344
rect 8025 -13336 8553 -10684
rect 8025 -13676 8055 -13336
rect 8523 -13676 8553 -13336
rect 8025 -16328 8553 -13676
rect 8025 -16668 8055 -16328
rect 8523 -16668 8553 -16328
rect 8025 -19320 8553 -16668
rect 8025 -19660 8055 -19320
rect 8523 -19660 8553 -19320
rect 8025 -21732 8553 -19660
rect 8025 -22072 8055 -21732
rect 8523 -22072 8553 -21732
rect 3426 -22538 3826 -22508
rect 3426 -22862 3456 -22538
rect 3796 -22862 3826 -22538
rect 962 -30949 1651 -30940
rect 2393 -30657 2761 -30633
rect 962 -30964 1330 -30949
rect 2393 -30977 2417 -30657
rect 2737 -30977 2761 -30657
rect 2393 -31001 2761 -30977
rect 3426 -36032 3826 -22862
rect 3426 -36356 3456 -36032
rect 3796 -36356 3826 -36032
rect 3426 -36426 3826 -36356
rect 4226 -26182 4626 -22508
rect 4226 -26506 4256 -26182
rect 4596 -26506 4626 -26182
rect 4226 -35840 4626 -26506
rect 4226 -36164 4256 -35840
rect 4596 -36164 4626 -35840
rect 4226 -36426 4626 -36164
rect 5026 -29826 5426 -22508
rect 5026 -30150 5056 -29826
rect 5396 -30150 5426 -29826
rect 5026 -35648 5426 -30150
rect 5026 -35972 5056 -35648
rect 5396 -35972 5426 -35648
rect 5026 -36426 5426 -35972
rect 5826 -33470 6226 -22508
rect 5826 -33794 5856 -33470
rect 6196 -33794 6226 -33470
rect 5826 -35456 6226 -33794
rect 5826 -35780 5856 -35456
rect 6196 -35780 6226 -35456
rect 5826 -36426 6226 -35780
rect 8025 -25376 8553 -22072
rect 8025 -25716 8055 -25376
rect 8523 -25716 8553 -25376
rect 8025 -29020 8553 -25716
rect 8025 -29360 8055 -29020
rect 8523 -29360 8553 -29020
rect 8025 -32664 8553 -29360
rect 8025 -33004 8055 -32664
rect 8523 -33004 8553 -32664
rect 8025 -34884 8553 -33004
rect 8025 -35224 8055 -34884
rect 8523 -35224 8553 -34884
rect 8025 -39096 8553 -35224
rect 8025 -39436 8055 -39096
rect 8523 -39436 8553 -39096
rect 8025 -42088 8553 -39436
rect 8954 -35648 9354 -34035
rect 8954 -35972 8984 -35648
rect 9324 -35972 9354 -35648
rect 8954 -39296 9354 -35972
rect 8954 -39536 8984 -39296
rect 9324 -39536 9354 -39296
rect 8954 -41200 9354 -39536
rect 9754 -35840 10154 -34035
rect 9754 -36164 9784 -35840
rect 10124 -36164 10154 -35840
rect 9754 -40930 10154 -36164
rect 9754 -41170 9784 -40930
rect 10124 -41170 10154 -40930
rect 9754 -41200 10154 -41170
rect 10554 -36032 10954 -34035
rect 10554 -36356 10584 -36032
rect 10924 -36356 10954 -36032
rect 10554 -40930 10954 -36356
rect 10554 -41170 10584 -40930
rect 10924 -41170 10954 -40930
rect 10554 -41200 10954 -41170
rect 11354 -35456 11754 -34035
rect 11354 -35780 11384 -35456
rect 11724 -35780 11754 -35456
rect 11354 -39296 11754 -35780
rect 11354 -39536 11384 -39296
rect 11724 -39536 11754 -39296
rect 11354 -41200 11754 -39536
rect 8025 -42428 8055 -42088
rect 8523 -42428 8553 -42088
rect 8025 -49080 8553 -42428
rect -1006 -49274 -526 -49244
rect -1006 -50214 -976 -49274
rect -556 -50214 -526 -49274
rect -1006 -50510 -526 -50214
rect 2198 -49274 2678 -49244
rect 2198 -50214 2228 -49274
rect 2648 -50214 2678 -49274
rect 2198 -50510 2678 -50214
rect 8025 -49420 8055 -49080
rect 8523 -49420 8553 -49080
rect 8025 -52072 8553 -49420
rect 8025 -52412 8055 -52072
rect 8523 -52412 8553 -52072
rect 8025 -55064 8553 -52412
rect 8025 -55404 8055 -55064
rect 8523 -55404 8553 -55064
rect -1006 -75394 -526 -70006
rect -1006 -75734 -976 -75394
rect -556 -75734 -526 -75394
rect -1006 -75764 -526 -75734
rect 2198 -75394 2678 -56572
rect 2198 -75734 2228 -75394
rect 2648 -75734 2678 -75394
rect 2198 -75764 2678 -75734
rect 8025 -59678 8553 -55404
rect 8025 -60018 8055 -59678
rect 8523 -60018 8553 -59678
rect 8025 -67536 8553 -60018
rect 8025 -67876 8055 -67536
rect 8523 -67876 8553 -67536
rect 8025 -75394 8553 -67876
rect 8025 -75734 8055 -75394
rect 8523 -75734 8553 -75394
rect 8025 -79200 8553 -75734
rect 8025 -79668 8055 -79200
rect 8523 -79668 8553 -79200
rect 8025 -79698 8553 -79668
rect 9854 -78472 10854 -78442
rect 9854 -78940 9884 -78472
rect 10824 -78940 10854 -78472
rect 9854 -79698 10854 -78940
rect 12082 -78472 12610 10386
rect 14482 -33470 14882 -22508
rect 14482 -33794 14512 -33470
rect 14852 -33794 14882 -33470
rect 14482 -35456 14882 -33794
rect 14482 -35780 14512 -35456
rect 14852 -35780 14882 -35456
rect 14482 -36426 14882 -35780
rect 15282 -29826 15682 -22508
rect 15282 -30150 15312 -29826
rect 15652 -30150 15682 -29826
rect 15282 -35648 15682 -30150
rect 15282 -35972 15312 -35648
rect 15652 -35972 15682 -35648
rect 15282 -36426 15682 -35972
rect 16082 -26182 16482 -22508
rect 16082 -26506 16112 -26182
rect 16452 -26506 16482 -26182
rect 16082 -35840 16482 -26506
rect 16082 -36164 16112 -35840
rect 16452 -36164 16482 -35840
rect 16082 -36426 16482 -36164
rect 16882 -22538 17282 -22508
rect 16882 -22862 16912 -22538
rect 17252 -22862 17282 -22538
rect 16882 -36032 17282 -22862
rect 16882 -36356 16912 -36032
rect 17252 -36356 17282 -36032
rect 16882 -36426 17282 -36356
rect 18654 -35144 19043 -33440
rect 18654 -35444 18684 -35144
rect 19013 -35444 19043 -35144
rect 17934 -37102 18334 -36694
rect 17934 -37342 17958 -37102
rect 18310 -37342 18334 -37102
rect 17934 -47628 18334 -37342
rect 18654 -39114 19043 -35444
rect 18654 -39414 18684 -39114
rect 19013 -39414 19043 -39114
rect 18654 -46853 19043 -39414
rect 21412 -36718 21812 -36694
rect 21412 -36958 21436 -36718
rect 21788 -36958 21812 -36718
rect 18654 -47273 18684 -46853
rect 19013 -47273 19043 -46853
rect 20433 -46853 20913 -46823
rect 20433 -47273 20463 -46853
rect 20883 -47273 20913 -46853
rect 18654 -47303 19043 -47273
rect 17934 -50022 17964 -47628
rect 18304 -50022 18334 -47628
rect 17934 -50052 18334 -50022
rect 21412 -47628 21812 -36958
rect 21412 -50022 21442 -47628
rect 21782 -50022 21812 -47628
rect 21412 -50052 21812 -50022
rect 18030 -75394 18510 -70006
rect 18030 -75734 18060 -75394
rect 18480 -75734 18510 -75394
rect 18030 -75764 18510 -75734
rect 18856 -70962 20843 -70867
rect 18856 -72072 18982 -70962
rect 20728 -72072 20843 -70962
rect 18856 -76251 20843 -72072
rect 21234 -75764 21714 -56572
rect 18831 -76275 20868 -76251
rect 18831 -78262 18855 -76275
rect 20844 -78262 20868 -76275
rect 18831 -78286 20868 -78262
rect 12082 -78940 12112 -78472
rect 12580 -78940 12610 -78472
rect 12082 -79698 12610 -78940
rect 27822 -78493 35352 -77265
rect 27822 -78884 27900 -78493
rect 35299 -78884 35352 -78493
rect -13104 -90973 -11014 -89973
rect -13104 -102827 -11014 -101827
rect -64045 -124560 -5513 -124452
rect -64045 -125347 -7913 -124560
rect -5926 -125347 -5513 -124560
rect -64045 -128455 -5513 -125347
rect -64045 -219640 -60042 -128455
rect 27822 -133596 35352 -78884
rect -57969 -141119 35352 -133596
rect -57969 -206166 -50446 -141119
rect 27822 -141131 35352 -141119
rect 37822 -79230 45352 -78884
rect 37822 -79621 37890 -79230
rect 45289 -79621 45352 -79230
rect 37822 -145968 45352 -79621
rect -40055 -153498 45352 -145968
rect -40055 -162711 -32525 -153498
rect -40129 -163739 -32525 -162711
rect -40129 -180752 -39416 -163739
rect -33277 -180752 -32525 -163739
rect -40129 -182039 -32525 -180752
rect -40129 -182076 -32599 -182039
rect -57969 -206453 86125 -206166
rect -57969 -211255 71133 -206453
rect 75935 -211255 81133 -206453
rect 85935 -211255 86125 -206453
rect -57969 -213689 86125 -211255
rect -64045 -223736 -63767 -219640
rect -60342 -223736 -60042 -219640
rect -64045 -224129 -60042 -223736
use capbank  capbank_0
timestamp 1698052002
transform -1 0 12625 0 -1 -55628
box -4432 -9038 8974 20462
use capbank  capbank_1
timestamp 1698052002
transform -1 0 12625 0 1 -10120
box -4432 -9038 8974 20462
use gc  gc_0
timestamp 1699972208
transform 1 0 14824 0 -1 -34882
box -532 -847 2650 1544
use gc  gc_2
timestamp 1699972208
transform -1 0 5884 0 -1 -34882
box -532 -847 2650 1544
use gc  gc_4
timestamp 1699972208
transform -1 0 11412 0 -1 -34882
box -532 -847 2650 1544
use mux21  mux21_0
timestamp 1699972208
transform 1 0 14523 0 1 -38290
box -42 -666 2760 1744
use mux21  mux21_2
timestamp 1699972208
transform 1 0 3467 0 1 -38290
box -42 -666 2760 1744
use mux21  mux21_3
timestamp 1699972208
transform 1 0 8995 0 1 -38290
box -42 -666 2760 1744
use osc_total  osc_total_1
timestamp 1699263546
transform 1 0 4 0 1 -27894
box -2821 -7596 22925 58950
use pa_total  pa_total_0
timestamp 1699369155
transform 1 0 -4393 0 1 -67194
box -72403 -55994 31999 32036
use startup  startup_0
timestamp 1699972208
transform -1 0 2640 0 -1 -47596
box -179 -352 3825 23026
use startup  startup_2
timestamp 1699972208
transform 1 0 18068 0 -1 -47596
box -179 -352 3825 23026
use uwb_noise_decoup_cell1  uwb_noise_decoup_cell1_0
timestamp 1663849571
transform 1 0 53254 0 1 -44190
box 0 0 4000 4000
use uwb_noise_decoup_cell1  uwb_noise_decoup_cell1_1
timestamp 1663849571
transform 1 0 33254 0 1 -96190
box 0 0 4000 4000
use uwb_noise_decoup_cell1  uwb_noise_decoup_cell1_2
timestamp 1663849571
transform 1 0 53254 0 1 -76190
box 0 0 4000 4000
use uwb_noise_decoup_cell1  uwb_noise_decoup_cell1_3
timestamp 1663849571
transform 1 0 53254 0 1 -72190
box 0 0 4000 4000
use uwb_noise_decoup_cell1  uwb_noise_decoup_cell1_4
timestamp 1663849571
transform 1 0 53254 0 1 -68190
box 0 0 4000 4000
use uwb_noise_decoup_cell1  uwb_noise_decoup_cell1_5
timestamp 1663849571
transform 1 0 53254 0 1 -64190
box 0 0 4000 4000
use uwb_noise_decoup_cell1  uwb_noise_decoup_cell1_6
timestamp 1663849571
transform 1 0 53254 0 1 -60190
box 0 0 4000 4000
use uwb_noise_decoup_cell1  uwb_noise_decoup_cell1_7
timestamp 1663849571
transform 1 0 53254 0 1 -56190
box 0 0 4000 4000
use uwb_noise_decoup_cell1  uwb_noise_decoup_cell1_8
timestamp 1663849571
transform 1 0 53254 0 1 -52190
box 0 0 4000 4000
use uwb_noise_decoup_cell1  uwb_noise_decoup_cell1_9
timestamp 1663849571
transform 1 0 53254 0 1 -48190
box 0 0 4000 4000
use uwb_noise_decoup_cell1  uwb_noise_decoup_cell1_10
timestamp 1663849571
transform 1 0 53254 0 1 -28190
box 0 0 4000 4000
use uwb_noise_decoup_cell1  uwb_noise_decoup_cell1_11
timestamp 1663849571
transform 1 0 49254 0 1 -32190
box 0 0 4000 4000
use uwb_noise_decoup_cell1  uwb_noise_decoup_cell1_12
timestamp 1663849571
transform 1 0 53254 0 1 -36190
box 0 0 4000 4000
use uwb_noise_decoup_cell1  uwb_noise_decoup_cell1_13
timestamp 1663849571
transform 1 0 53254 0 1 -32190
box 0 0 4000 4000
use uwb_noise_decoup_cell1  uwb_noise_decoup_cell1_14
timestamp 1663849571
transform 1 0 53254 0 1 -16190
box 0 0 4000 4000
use uwb_noise_decoup_cell1  uwb_noise_decoup_cell1_15
timestamp 1663849571
transform 1 0 53254 0 1 -24190
box 0 0 4000 4000
use uwb_noise_decoup_cell1  uwb_noise_decoup_cell1_16
timestamp 1663849571
transform 1 0 53254 0 1 -20190
box 0 0 4000 4000
use uwb_noise_decoup_cell1  uwb_noise_decoup_cell1_17
timestamp 1663849571
transform 1 0 53254 0 1 -190
box 0 0 4000 4000
use uwb_noise_decoup_cell1  uwb_noise_decoup_cell1_18
timestamp 1663849571
transform 1 0 53254 0 1 -12190
box 0 0 4000 4000
use uwb_noise_decoup_cell1  uwb_noise_decoup_cell1_19
timestamp 1663849571
transform 1 0 53254 0 1 -8190
box 0 0 4000 4000
use uwb_noise_decoup_cell1  uwb_noise_decoup_cell1_20
timestamp 1663849571
transform 1 0 53254 0 1 -4190
box 0 0 4000 4000
use uwb_noise_decoup_cell1  uwb_noise_decoup_cell1_22
timestamp 1663849571
transform 1 0 53254 0 1 3810
box 0 0 4000 4000
use uwb_noise_decoup_cell1  uwb_noise_decoup_cell1_23
timestamp 1663849571
transform 1 0 53254 0 1 7810
box 0 0 4000 4000
use uwb_noise_decoup_cell1  uwb_noise_decoup_cell1_29
timestamp 1663849571
transform 1 0 53254 0 1 -80190
box 0 0 4000 4000
use uwb_noise_decoup_cell1  uwb_noise_decoup_cell1_30
timestamp 1663849571
transform 1 0 53254 0 1 -84190
box 0 0 4000 4000
use uwb_noise_decoup_cell1  uwb_noise_decoup_cell1_31
timestamp 1663849571
transform 1 0 33254 0 1 -92190
box 0 0 4000 4000
use uwb_noise_decoup_cell1  uwb_noise_decoup_cell1_32
timestamp 1663849571
transform 1 0 53254 0 1 -92190
box 0 0 4000 4000
use uwb_noise_decoup_cell1  uwb_noise_decoup_cell1_33
timestamp 1663849571
transform 1 0 33254 0 1 -112190
box 0 0 4000 4000
use uwb_noise_decoup_cell1  uwb_noise_decoup_cell1_34
timestamp 1663849571
transform 1 0 37254 0 1 -96190
box 0 0 4000 4000
use uwb_noise_decoup_cell1  uwb_noise_decoup_cell1_35
timestamp 1663849571
transform 1 0 41254 0 1 -96190
box 0 0 4000 4000
use uwb_noise_decoup_cell1  uwb_noise_decoup_cell1_36
timestamp 1663849571
transform 1 0 45254 0 1 -96190
box 0 0 4000 4000
use uwb_noise_decoup_cell1  uwb_noise_decoup_cell1_37
timestamp 1663849571
transform 1 0 53254 0 1 -88190
box 0 0 4000 4000
use uwb_noise_decoup_cell1  uwb_noise_decoup_cell1_38
timestamp 1663849571
transform 1 0 33254 0 1 -88190
box 0 0 4000 4000
use uwb_noise_decoup_cell1  uwb_noise_decoup_cell1_39
timestamp 1663849571
transform 1 0 45254 0 1 -92190
box 0 0 4000 4000
use uwb_noise_decoup_cell1  uwb_noise_decoup_cell1_40
timestamp 1663849571
transform 1 0 41254 0 1 -92190
box 0 0 4000 4000
use uwb_noise_decoup_cell1  uwb_noise_decoup_cell1_41
timestamp 1663849571
transform 1 0 37254 0 1 -92190
box 0 0 4000 4000
use uwb_noise_decoup_cell1  uwb_noise_decoup_cell1_42
timestamp 1663849571
transform 1 0 45254 0 1 -88190
box 0 0 4000 4000
use uwb_noise_decoup_cell1  uwb_noise_decoup_cell1_43
timestamp 1663849571
transform 1 0 41254 0 1 -88190
box 0 0 4000 4000
use uwb_noise_decoup_cell1  uwb_noise_decoup_cell1_44
timestamp 1663849571
transform 1 0 37254 0 1 -88190
box 0 0 4000 4000
use uwb_noise_decoup_cell1  uwb_noise_decoup_cell1_45
timestamp 1663849571
transform 1 0 61254 0 1 -112190
box 0 0 4000 4000
use uwb_noise_decoup_cell1  uwb_noise_decoup_cell1_46
timestamp 1663849571
transform 1 0 45254 0 1 -112190
box 0 0 4000 4000
use uwb_noise_decoup_cell1  uwb_noise_decoup_cell1_47
timestamp 1663849571
transform 1 0 41254 0 1 -112190
box 0 0 4000 4000
use uwb_noise_decoup_cell1  uwb_noise_decoup_cell1_48
timestamp 1663849571
transform 1 0 37254 0 1 -112190
box 0 0 4000 4000
use uwb_noise_decoup_cell1  uwb_noise_decoup_cell1_49
timestamp 1663849571
transform 1 0 53254 0 1 -96190
box 0 0 4000 4000
use uwb_noise_decoup_cell1  uwb_noise_decoup_cell1_50
timestamp 1663849571
transform 1 0 53254 0 1 -100190
box 0 0 4000 4000
use uwb_noise_decoup_cell1  uwb_noise_decoup_cell1_51
timestamp 1663849571
transform 1 0 45254 0 1 -100190
box 0 0 4000 4000
use uwb_noise_decoup_cell1  uwb_noise_decoup_cell1_52
timestamp 1663849571
transform 1 0 41254 0 1 -100190
box 0 0 4000 4000
use uwb_noise_decoup_cell1  uwb_noise_decoup_cell1_53
timestamp 1663849571
transform 1 0 37254 0 1 -100190
box 0 0 4000 4000
use uwb_noise_decoup_cell1  uwb_noise_decoup_cell1_54
timestamp 1663849571
transform 1 0 33254 0 1 -100190
box 0 0 4000 4000
use uwb_noise_decoup_cell1  uwb_noise_decoup_cell1_55
timestamp 1663849571
transform 1 0 33254 0 1 -104190
box 0 0 4000 4000
use uwb_noise_decoup_cell1  uwb_noise_decoup_cell1_56
timestamp 1663849571
transform 1 0 37254 0 1 -104190
box 0 0 4000 4000
use uwb_noise_decoup_cell1  uwb_noise_decoup_cell1_57
timestamp 1663849571
transform 1 0 41254 0 1 -104190
box 0 0 4000 4000
use uwb_noise_decoup_cell1  uwb_noise_decoup_cell1_58
timestamp 1663849571
transform 1 0 45254 0 1 -104190
box 0 0 4000 4000
use uwb_noise_decoup_cell1  uwb_noise_decoup_cell1_59
timestamp 1663849571
transform 1 0 53254 0 1 -104190
box 0 0 4000 4000
use uwb_noise_decoup_cell1  uwb_noise_decoup_cell1_60
timestamp 1663849571
transform 1 0 33254 0 1 -108190
box 0 0 4000 4000
use uwb_noise_decoup_cell1  uwb_noise_decoup_cell1_61
timestamp 1663849571
transform 1 0 37254 0 1 -108190
box 0 0 4000 4000
use uwb_noise_decoup_cell1  uwb_noise_decoup_cell1_62
timestamp 1663849571
transform 1 0 41254 0 1 -108190
box 0 0 4000 4000
use uwb_noise_decoup_cell1  uwb_noise_decoup_cell1_63
timestamp 1663849571
transform 1 0 45254 0 1 -108190
box 0 0 4000 4000
use uwb_noise_decoup_cell1  uwb_noise_decoup_cell1_64
timestamp 1663849571
transform 1 0 61254 0 1 -108190
box 0 0 4000 4000
use uwb_noise_decoup_cell1  uwb_noise_decoup_cell1_65
timestamp 1663849571
transform 1 0 53254 0 1 15810
box 0 0 4000 4000
use uwb_noise_decoup_cell1  uwb_noise_decoup_cell1_66
timestamp 1663849571
transform 1 0 53254 0 1 11810
box 0 0 4000 4000
use uwb_noise_decoup_cell1  uwb_noise_decoup_cell1_67
timestamp 1663849571
transform 1 0 53254 0 1 23810
box 0 0 4000 4000
use uwb_noise_decoup_cell1  uwb_noise_decoup_cell1_68
timestamp 1663849571
transform 1 0 53254 0 1 19810
box 0 0 4000 4000
use uwb_noise_decoup_cell1  uwb_noise_decoup_cell1_69
timestamp 1663849571
transform 1 0 53254 0 1 31810
box 0 0 4000 4000
use uwb_noise_decoup_cell1  uwb_noise_decoup_cell1_70
timestamp 1663849571
transform 1 0 53254 0 1 27810
box 0 0 4000 4000
use uwb_noise_decoup_cell1  uwb_noise_decoup_cell1_71
timestamp 1663849571
transform 1 0 45254 0 1 11810
box 0 0 4000 4000
use uwb_noise_decoup_cell1  uwb_noise_decoup_cell1_72
timestamp 1663849571
transform 1 0 45254 0 1 15810
box 0 0 4000 4000
use uwb_noise_decoup_cell1  uwb_noise_decoup_cell1_73
timestamp 1663849571
transform 1 0 45254 0 1 19810
box 0 0 4000 4000
use uwb_noise_decoup_cell1  uwb_noise_decoup_cell1_74
timestamp 1663849571
transform 1 0 45254 0 1 23810
box 0 0 4000 4000
use uwb_noise_decoup_cell1  uwb_noise_decoup_cell1_75
timestamp 1663849571
transform 1 0 45254 0 1 27810
box 0 0 4000 4000
use uwb_noise_decoup_cell1  uwb_noise_decoup_cell1_76
timestamp 1663849571
transform 1 0 45254 0 1 31810
box 0 0 4000 4000
use uwb_noise_decoup_cell1  uwb_noise_decoup_cell1_77
timestamp 1663849571
transform 1 0 41254 0 1 11810
box 0 0 4000 4000
use uwb_noise_decoup_cell1  uwb_noise_decoup_cell1_78
timestamp 1663849571
transform 1 0 41254 0 1 15810
box 0 0 4000 4000
use uwb_noise_decoup_cell1  uwb_noise_decoup_cell1_79
timestamp 1663849571
transform 1 0 41254 0 1 19810
box 0 0 4000 4000
use uwb_noise_decoup_cell1  uwb_noise_decoup_cell1_80
timestamp 1663849571
transform 1 0 41254 0 1 23810
box 0 0 4000 4000
use uwb_noise_decoup_cell1  uwb_noise_decoup_cell1_81
timestamp 1663849571
transform 1 0 41254 0 1 27810
box 0 0 4000 4000
use uwb_noise_decoup_cell1  uwb_noise_decoup_cell1_82
timestamp 1663849571
transform 1 0 41254 0 1 31810
box 0 0 4000 4000
use uwb_noise_decoup_cell1  uwb_noise_decoup_cell1_83
timestamp 1663849571
transform 1 0 37254 0 1 15810
box 0 0 4000 4000
use uwb_noise_decoup_cell1  uwb_noise_decoup_cell1_84
timestamp 1663849571
transform 1 0 37254 0 1 11810
box 0 0 4000 4000
use uwb_noise_decoup_cell1  uwb_noise_decoup_cell1_85
timestamp 1663849571
transform 1 0 37254 0 1 19810
box 0 0 4000 4000
use uwb_noise_decoup_cell1  uwb_noise_decoup_cell1_86
timestamp 1663849571
transform 1 0 37254 0 1 23810
box 0 0 4000 4000
use uwb_noise_decoup_cell1  uwb_noise_decoup_cell1_87
timestamp 1663849571
transform 1 0 37254 0 1 27810
box 0 0 4000 4000
use uwb_noise_decoup_cell1  uwb_noise_decoup_cell1_88
timestamp 1663849571
transform 1 0 37254 0 1 31810
box 0 0 4000 4000
use uwb_noise_decoup_cell1  uwb_noise_decoup_cell1_89
timestamp 1663849571
transform 1 0 33254 0 1 23810
box 0 0 4000 4000
use uwb_noise_decoup_cell1  uwb_noise_decoup_cell1_90
timestamp 1663849571
transform 1 0 33254 0 1 19810
box 0 0 4000 4000
use uwb_noise_decoup_cell1  uwb_noise_decoup_cell1_91
timestamp 1663849571
transform 1 0 33254 0 1 11810
box 0 0 4000 4000
use uwb_noise_decoup_cell1  uwb_noise_decoup_cell1_92
timestamp 1663849571
transform 1 0 33254 0 1 15810
box 0 0 4000 4000
use uwb_noise_decoup_cell1  uwb_noise_decoup_cell1_93
timestamp 1663849571
transform 1 0 33254 0 1 27810
box 0 0 4000 4000
use uwb_noise_decoup_cell1  uwb_noise_decoup_cell1_94
timestamp 1663849571
transform 1 0 33254 0 1 31810
box 0 0 4000 4000
use uwb_noise_decoup_cell1  uwb_noise_decoup_cell1_101
timestamp 1663849571
transform 1 0 49254 0 1 -112190
box 0 0 4000 4000
use uwb_noise_decoup_cell1  uwb_noise_decoup_cell1_102
timestamp 1663849571
transform 1 0 49254 0 1 -108190
box 0 0 4000 4000
use uwb_noise_decoup_cell1  uwb_noise_decoup_cell1_103
timestamp 1663849571
transform 1 0 49254 0 1 -104190
box 0 0 4000 4000
use uwb_noise_decoup_cell1  uwb_noise_decoup_cell1_104
timestamp 1663849571
transform 1 0 49254 0 1 -100190
box 0 0 4000 4000
use uwb_noise_decoup_cell1  uwb_noise_decoup_cell1_105
timestamp 1663849571
transform 1 0 49254 0 1 -96190
box 0 0 4000 4000
use uwb_noise_decoup_cell1  uwb_noise_decoup_cell1_106
timestamp 1663849571
transform 1 0 49254 0 1 -92190
box 0 0 4000 4000
use uwb_noise_decoup_cell1  uwb_noise_decoup_cell1_107
timestamp 1663849571
transform 1 0 49254 0 1 -88190
box 0 0 4000 4000
use uwb_noise_decoup_cell1  uwb_noise_decoup_cell1_108
timestamp 1663849571
transform 1 0 49254 0 1 -84190
box 0 0 4000 4000
use uwb_noise_decoup_cell1  uwb_noise_decoup_cell1_109
timestamp 1663849571
transform 1 0 49254 0 1 -80190
box 0 0 4000 4000
use uwb_noise_decoup_cell1  uwb_noise_decoup_cell1_110
timestamp 1663849571
transform 1 0 49254 0 1 -76190
box 0 0 4000 4000
use uwb_noise_decoup_cell1  uwb_noise_decoup_cell1_111
timestamp 1663849571
transform 1 0 49254 0 1 -72190
box 0 0 4000 4000
use uwb_noise_decoup_cell1  uwb_noise_decoup_cell1_112
timestamp 1663849571
transform 1 0 49254 0 1 -68190
box 0 0 4000 4000
use uwb_noise_decoup_cell1  uwb_noise_decoup_cell1_113
timestamp 1663849571
transform 1 0 49254 0 1 -64190
box 0 0 4000 4000
use uwb_noise_decoup_cell1  uwb_noise_decoup_cell1_114
timestamp 1663849571
transform 1 0 49254 0 1 -60190
box 0 0 4000 4000
use uwb_noise_decoup_cell1  uwb_noise_decoup_cell1_115
timestamp 1663849571
transform 1 0 49254 0 1 -56190
box 0 0 4000 4000
use uwb_noise_decoup_cell1  uwb_noise_decoup_cell1_116
timestamp 1663849571
transform 1 0 49254 0 1 -52190
box 0 0 4000 4000
use uwb_noise_decoup_cell1  uwb_noise_decoup_cell1_117
timestamp 1663849571
transform 1 0 49254 0 1 -48190
box 0 0 4000 4000
use uwb_noise_decoup_cell1  uwb_noise_decoup_cell1_118
timestamp 1663849571
transform 1 0 49254 0 1 -44190
box 0 0 4000 4000
use uwb_noise_decoup_cell1  uwb_noise_decoup_cell1_119
timestamp 1663849571
transform 1 0 49254 0 1 -36190
box 0 0 4000 4000
use uwb_noise_decoup_cell1  uwb_noise_decoup_cell1_120
timestamp 1663849571
transform 1 0 53254 0 1 -40190
box 0 0 4000 4000
use uwb_noise_decoup_cell1  uwb_noise_decoup_cell1_121
timestamp 1663849571
transform 1 0 61254 0 1 -36190
box 0 0 4000 4000
use uwb_noise_decoup_cell1  uwb_noise_decoup_cell1_122
timestamp 1663849571
transform 1 0 49254 0 1 -28190
box 0 0 4000 4000
use uwb_noise_decoup_cell1  uwb_noise_decoup_cell1_123
timestamp 1663849571
transform 1 0 49254 0 1 -20190
box 0 0 4000 4000
use uwb_noise_decoup_cell1  uwb_noise_decoup_cell1_124
timestamp 1663849571
transform 1 0 49254 0 1 -24190
box 0 0 4000 4000
use uwb_noise_decoup_cell1  uwb_noise_decoup_cell1_125
timestamp 1663849571
transform 1 0 49254 0 1 -16190
box 0 0 4000 4000
use uwb_noise_decoup_cell1  uwb_noise_decoup_cell1_126
timestamp 1663849571
transform 1 0 49254 0 1 -8190
box 0 0 4000 4000
use uwb_noise_decoup_cell1  uwb_noise_decoup_cell1_127
timestamp 1663849571
transform 1 0 49254 0 1 -12190
box 0 0 4000 4000
use uwb_noise_decoup_cell1  uwb_noise_decoup_cell1_128
timestamp 1663849571
transform 1 0 49254 0 1 -190
box 0 0 4000 4000
use uwb_noise_decoup_cell1  uwb_noise_decoup_cell1_129
timestamp 1663849571
transform 1 0 49254 0 1 -4190
box 0 0 4000 4000
use uwb_noise_decoup_cell1  uwb_noise_decoup_cell1_130
timestamp 1663849571
transform 1 0 49254 0 1 11810
box 0 0 4000 4000
use uwb_noise_decoup_cell1  uwb_noise_decoup_cell1_131
timestamp 1663849571
transform 1 0 49254 0 1 7810
box 0 0 4000 4000
use uwb_noise_decoup_cell1  uwb_noise_decoup_cell1_132
timestamp 1663849571
transform 1 0 49254 0 1 3810
box 0 0 4000 4000
use uwb_noise_decoup_cell1  uwb_noise_decoup_cell1_133
timestamp 1663849571
transform 1 0 49254 0 1 15810
box 0 0 4000 4000
use uwb_noise_decoup_cell1  uwb_noise_decoup_cell1_134
timestamp 1663849571
transform 1 0 49254 0 1 19810
box 0 0 4000 4000
use uwb_noise_decoup_cell1  uwb_noise_decoup_cell1_135
timestamp 1663849571
transform 1 0 49254 0 1 27810
box 0 0 4000 4000
use uwb_noise_decoup_cell1  uwb_noise_decoup_cell1_136
timestamp 1663849571
transform 1 0 49254 0 1 31810
box 0 0 4000 4000
use uwb_noise_decoup_cell1  uwb_noise_decoup_cell1_137
timestamp 1663849571
transform 1 0 49254 0 1 23810
box 0 0 4000 4000
use uwb_noise_decoup_cell1  uwb_noise_decoup_cell1_138
timestamp 1663849571
transform 1 0 53254 0 1 -108190
box 0 0 4000 4000
use uwb_noise_decoup_cell1  uwb_noise_decoup_cell1_139
timestamp 1663849571
transform 1 0 53254 0 1 -112190
box 0 0 4000 4000
use uwb_noise_decoup_cell1  uwb_noise_decoup_cell1_140
timestamp 1663849571
transform 1 0 61254 0 1 -100190
box 0 0 4000 4000
use uwb_noise_decoup_cell1  uwb_noise_decoup_cell1_141
timestamp 1663849571
transform 1 0 61254 0 1 -104190
box 0 0 4000 4000
use uwb_noise_decoup_cell1  uwb_noise_decoup_cell1_142
timestamp 1663849571
transform 1 0 61254 0 1 -92190
box 0 0 4000 4000
use uwb_noise_decoup_cell1  uwb_noise_decoup_cell1_143
timestamp 1663849571
transform 1 0 61254 0 1 -96190
box 0 0 4000 4000
use uwb_noise_decoup_cell1  uwb_noise_decoup_cell1_144
timestamp 1663849571
transform 1 0 61254 0 1 -80190
box 0 0 4000 4000
use uwb_noise_decoup_cell1  uwb_noise_decoup_cell1_145
timestamp 1663849571
transform 1 0 61254 0 1 -84190
box 0 0 4000 4000
use uwb_noise_decoup_cell1  uwb_noise_decoup_cell1_146
timestamp 1663849571
transform 1 0 61254 0 1 -88190
box 0 0 4000 4000
use uwb_noise_decoup_cell1  uwb_noise_decoup_cell1_147
timestamp 1663849571
transform 1 0 61254 0 1 -72190
box 0 0 4000 4000
use uwb_noise_decoup_cell1  uwb_noise_decoup_cell1_148
timestamp 1663849571
transform 1 0 61254 0 1 -76190
box 0 0 4000 4000
use uwb_noise_decoup_cell1  uwb_noise_decoup_cell1_149
timestamp 1663849571
transform 1 0 61254 0 1 -60190
box 0 0 4000 4000
use uwb_noise_decoup_cell1  uwb_noise_decoup_cell1_150
timestamp 1663849571
transform 1 0 61254 0 1 -64190
box 0 0 4000 4000
use uwb_noise_decoup_cell1  uwb_noise_decoup_cell1_151
timestamp 1663849571
transform 1 0 61254 0 1 -68190
box 0 0 4000 4000
use uwb_noise_decoup_cell1  uwb_noise_decoup_cell1_152
timestamp 1663849571
transform 1 0 61254 0 1 -52190
box 0 0 4000 4000
use uwb_noise_decoup_cell1  uwb_noise_decoup_cell1_153
timestamp 1663849571
transform 1 0 61254 0 1 -56190
box 0 0 4000 4000
use uwb_noise_decoup_cell1  uwb_noise_decoup_cell1_154
timestamp 1663849571
transform 1 0 57254 0 1 -36190
box 0 0 4000 4000
use uwb_noise_decoup_cell1  uwb_noise_decoup_cell1_155
timestamp 1663849571
transform 1 0 61254 0 1 -44190
box 0 0 4000 4000
use uwb_noise_decoup_cell1  uwb_noise_decoup_cell1_156
timestamp 1663849571
transform 1 0 61254 0 1 -48190
box 0 0 4000 4000
use uwb_noise_decoup_cell1  uwb_noise_decoup_cell1_157
timestamp 1663849571
transform 1 0 61254 0 1 -32190
box 0 0 4000 4000
use uwb_noise_decoup_cell1  uwb_noise_decoup_cell1_158
timestamp 1663849571
transform 1 0 49254 0 1 -40190
box 0 0 4000 4000
use uwb_noise_decoup_cell1  uwb_noise_decoup_cell1_159
timestamp 1663849571
transform 1 0 61254 0 1 -28190
box 0 0 4000 4000
use uwb_noise_decoup_cell1  uwb_noise_decoup_cell1_160
timestamp 1663849571
transform 1 0 61254 0 1 -20190
box 0 0 4000 4000
use uwb_noise_decoup_cell1  uwb_noise_decoup_cell1_161
timestamp 1663849571
transform 1 0 61254 0 1 -24190
box 0 0 4000 4000
use uwb_noise_decoup_cell1  uwb_noise_decoup_cell1_162
timestamp 1663849571
transform 1 0 61254 0 1 -8190
box 0 0 4000 4000
use uwb_noise_decoup_cell1  uwb_noise_decoup_cell1_163
timestamp 1663849571
transform 1 0 61254 0 1 -12190
box 0 0 4000 4000
use uwb_noise_decoup_cell1  uwb_noise_decoup_cell1_164
timestamp 1663849571
transform 1 0 61254 0 1 -16190
box 0 0 4000 4000
use uwb_noise_decoup_cell1  uwb_noise_decoup_cell1_165
timestamp 1663849571
transform 1 0 61254 0 1 -190
box 0 0 4000 4000
use uwb_noise_decoup_cell1  uwb_noise_decoup_cell1_166
timestamp 1663849571
transform 1 0 61254 0 1 -4190
box 0 0 4000 4000
use uwb_noise_decoup_cell1  uwb_noise_decoup_cell1_167
timestamp 1663849571
transform 1 0 61254 0 1 11810
box 0 0 4000 4000
use uwb_noise_decoup_cell1  uwb_noise_decoup_cell1_168
timestamp 1663849571
transform 1 0 61254 0 1 7810
box 0 0 4000 4000
use uwb_noise_decoup_cell1  uwb_noise_decoup_cell1_169
timestamp 1663849571
transform 1 0 61254 0 1 3810
box 0 0 4000 4000
use uwb_noise_decoup_cell1  uwb_noise_decoup_cell1_170
timestamp 1663849571
transform 1 0 61254 0 1 19810
box 0 0 4000 4000
use uwb_noise_decoup_cell1  uwb_noise_decoup_cell1_171
timestamp 1663849571
transform 1 0 61254 0 1 15810
box 0 0 4000 4000
use uwb_noise_decoup_cell1  uwb_noise_decoup_cell1_172
timestamp 1663849571
transform 1 0 61254 0 1 31810
box 0 0 4000 4000
use uwb_noise_decoup_cell1  uwb_noise_decoup_cell1_173
timestamp 1663849571
transform 1 0 61254 0 1 27810
box 0 0 4000 4000
use uwb_noise_decoup_cell1  uwb_noise_decoup_cell1_174
timestamp 1663849571
transform 1 0 61254 0 1 23810
box 0 0 4000 4000
use uwb_noise_decoup_cell1  uwb_noise_decoup_cell1_175
timestamp 1663849571
transform 1 0 57254 0 1 -112190
box 0 0 4000 4000
use uwb_noise_decoup_cell1  uwb_noise_decoup_cell1_176
timestamp 1663849571
transform 1 0 57254 0 1 -108190
box 0 0 4000 4000
use uwb_noise_decoup_cell1  uwb_noise_decoup_cell1_177
timestamp 1663849571
transform 1 0 57254 0 1 -100190
box 0 0 4000 4000
use uwb_noise_decoup_cell1  uwb_noise_decoup_cell1_178
timestamp 1663849571
transform 1 0 57254 0 1 -104190
box 0 0 4000 4000
use uwb_noise_decoup_cell1  uwb_noise_decoup_cell1_179
timestamp 1663849571
transform 1 0 57254 0 1 -92190
box 0 0 4000 4000
use uwb_noise_decoup_cell1  uwb_noise_decoup_cell1_180
timestamp 1663849571
transform 1 0 57254 0 1 -96190
box 0 0 4000 4000
use uwb_noise_decoup_cell1  uwb_noise_decoup_cell1_181
timestamp 1663849571
transform 1 0 57254 0 1 -80190
box 0 0 4000 4000
use uwb_noise_decoup_cell1  uwb_noise_decoup_cell1_182
timestamp 1663849571
transform 1 0 57254 0 1 -84190
box 0 0 4000 4000
use uwb_noise_decoup_cell1  uwb_noise_decoup_cell1_183
timestamp 1663849571
transform 1 0 57254 0 1 -88190
box 0 0 4000 4000
use uwb_noise_decoup_cell1  uwb_noise_decoup_cell1_184
timestamp 1663849571
transform 1 0 57254 0 1 -72190
box 0 0 4000 4000
use uwb_noise_decoup_cell1  uwb_noise_decoup_cell1_185
timestamp 1663849571
transform 1 0 57254 0 1 -76190
box 0 0 4000 4000
use uwb_noise_decoup_cell1  uwb_noise_decoup_cell1_186
timestamp 1663849571
transform 1 0 57254 0 1 -60190
box 0 0 4000 4000
use uwb_noise_decoup_cell1  uwb_noise_decoup_cell1_187
timestamp 1663849571
transform 1 0 57254 0 1 -64190
box 0 0 4000 4000
use uwb_noise_decoup_cell1  uwb_noise_decoup_cell1_188
timestamp 1663849571
transform 1 0 57254 0 1 -68190
box 0 0 4000 4000
use uwb_noise_decoup_cell1  uwb_noise_decoup_cell1_189
timestamp 1663849571
transform 1 0 57254 0 1 -52190
box 0 0 4000 4000
use uwb_noise_decoup_cell1  uwb_noise_decoup_cell1_190
timestamp 1663849571
transform 1 0 57254 0 1 -56190
box 0 0 4000 4000
use uwb_noise_decoup_cell1  uwb_noise_decoup_cell1_191
timestamp 1663849571
transform 1 0 61254 0 1 -40190
box 0 0 4000 4000
use uwb_noise_decoup_cell1  uwb_noise_decoup_cell1_192
timestamp 1663849571
transform 1 0 57254 0 1 -44190
box 0 0 4000 4000
use uwb_noise_decoup_cell1  uwb_noise_decoup_cell1_193
timestamp 1663849571
transform 1 0 57254 0 1 -48190
box 0 0 4000 4000
use uwb_noise_decoup_cell1  uwb_noise_decoup_cell1_194
timestamp 1663849571
transform 1 0 57254 0 1 -32190
box 0 0 4000 4000
use uwb_noise_decoup_cell1  uwb_noise_decoup_cell1_195
timestamp 1663849571
transform 1 0 57254 0 1 -40190
box 0 0 4000 4000
use uwb_noise_decoup_cell1  uwb_noise_decoup_cell1_196
timestamp 1663849571
transform 1 0 57254 0 1 -28190
box 0 0 4000 4000
use uwb_noise_decoup_cell1  uwb_noise_decoup_cell1_197
timestamp 1663849571
transform 1 0 57254 0 1 -20190
box 0 0 4000 4000
use uwb_noise_decoup_cell1  uwb_noise_decoup_cell1_198
timestamp 1663849571
transform 1 0 57254 0 1 -24190
box 0 0 4000 4000
use uwb_noise_decoup_cell1  uwb_noise_decoup_cell1_199
timestamp 1663849571
transform 1 0 57254 0 1 -8190
box 0 0 4000 4000
use uwb_noise_decoup_cell1  uwb_noise_decoup_cell1_200
timestamp 1663849571
transform 1 0 57254 0 1 -12190
box 0 0 4000 4000
use uwb_noise_decoup_cell1  uwb_noise_decoup_cell1_201
timestamp 1663849571
transform 1 0 57254 0 1 -16190
box 0 0 4000 4000
use uwb_noise_decoup_cell1  uwb_noise_decoup_cell1_202
timestamp 1663849571
transform 1 0 57254 0 1 -190
box 0 0 4000 4000
use uwb_noise_decoup_cell1  uwb_noise_decoup_cell1_203
timestamp 1663849571
transform 1 0 57254 0 1 -4190
box 0 0 4000 4000
use uwb_noise_decoup_cell1  uwb_noise_decoup_cell1_204
timestamp 1663849571
transform 1 0 57254 0 1 11810
box 0 0 4000 4000
use uwb_noise_decoup_cell1  uwb_noise_decoup_cell1_205
timestamp 1663849571
transform 1 0 57254 0 1 7810
box 0 0 4000 4000
use uwb_noise_decoup_cell1  uwb_noise_decoup_cell1_206
timestamp 1663849571
transform 1 0 57254 0 1 3810
box 0 0 4000 4000
use uwb_noise_decoup_cell1  uwb_noise_decoup_cell1_207
timestamp 1663849571
transform 1 0 57254 0 1 19810
box 0 0 4000 4000
use uwb_noise_decoup_cell1  uwb_noise_decoup_cell1_208
timestamp 1663849571
transform 1 0 57254 0 1 15810
box 0 0 4000 4000
use uwb_noise_decoup_cell1  uwb_noise_decoup_cell1_209
timestamp 1663849571
transform 1 0 57254 0 1 31810
box 0 0 4000 4000
use uwb_noise_decoup_cell1  uwb_noise_decoup_cell1_210
timestamp 1663849571
transform 1 0 57254 0 1 27810
box 0 0 4000 4000
use uwb_noise_decoup_cell1  uwb_noise_decoup_cell1_211
timestamp 1663849571
transform 1 0 57254 0 1 23810
box 0 0 4000 4000
<< labels >>
flabel metal1 10284 7314 10382 7626 0 FreeSans 1600 0 0 0 osc_tune[5]
port 20 nsew
flabel metal1 10284 -544 10382 -232 0 FreeSans 1600 0 0 0 osc_tune[4]
port 21 nsew
flabel metal1 10284 -8402 10382 -8090 0 FreeSans 1600 0 0 0 osc_tune[3]
port 22 nsew
flabel metal1 10284 -13016 10382 -12704 0 FreeSans 1600 0 0 0 osc_tune[2]
port 23 nsew
flabel metal1 10284 -16008 10382 -15696 0 FreeSans 1600 0 0 0 osc_tune[1]
port 24 nsew
flabel metal1 10284 -19000 10382 -18688 0 FreeSans 1600 0 0 0 osc_tune[0]
port 25 nsew
flabel metal3 8764 -34210 11944 -34114 0 FreeSans 1600 0 0 0 pa_gain[3]
port 26 nsew
flabel metal3 8764 -34402 11944 -34306 0 FreeSans 1600 0 0 0 pa_gain[2]
port 27 nsew
flabel metal3 8764 -34594 11944 -34498 0 FreeSans 1600 0 0 0 pa_gain[1]
port 28 nsew
flabel metal3 8764 -34786 11944 -34690 0 FreeSans 1600 0 0 0 pa_gain[0]
port 29 nsew
flabel metal4 14870 -34210 17472 -34114 0 FreeSans 1600 0 0 0 osc_gain[3]
port 30 nsew
flabel metal4 14870 -34402 17472 -34306 0 FreeSans 1600 0 0 0 osc_gain[2]
port 31 nsew
flabel metal4 14870 -34594 17472 -34498 0 FreeSans 1600 0 0 0 osc_gain[1]
port 32 nsew
flabel metal4 14870 -34786 17472 -34690 0 FreeSans 1600 0 0 0 osc_gain[0]
port 33 nsew
flabel metal2 8953 -36934 11755 -36838 0 FreeSans 1600 0 0 0 pa_trig1_en
port 35 nsew
flabel metal2 8953 -36790 11755 -36694 0 FreeSans 1600 0 0 0 pa_trig1_test_en
port 36 nsew
flabel metal2 14481 -36790 17283 -36694 0 FreeSans 1600 0 0 0 osc_trig1_test_en
port 39 nsew
flabel metal2 14481 -36934 17283 -36838 0 FreeSans 1600 0 0 0 osc_trig1_en
port 38 nsew
flabel metal2 14481 -36646 17283 -36550 0 FreeSans 1600 0 0 0 osc_trig1_test
port 40 nsew
flabel metal2 3425 -36646 6227 -36550 0 FreeSans 1600 0 0 0 osc_trig2_test
port 41 nsew
flabel metal2 3425 -36790 6227 -36694 0 FreeSans 1600 0 0 0 osc_trig2_test_en
port 42 nsew
flabel metal2 3425 -36934 6227 -36838 0 FreeSans 1600 0 0 0 osc_trig2_en
port 43 nsew
flabel metal5 18654 -35144 19043 -33440 0 FreeSans 1600 0 0 0 vdd1v8
port 44 nsew
flabel metal4 8523 -79698 9587 -79170 0 FreeSans 1600 0 0 0 vss
port 0 nsew
flabel metal4 10824 -78970 12112 -78442 0 FreeSans 1600 0 0 0 vdd1v0
port 2 nsew
flabel metal1 10326 -73374 10424 -73062 0 FreeSans 1600 0 0 0 pa_tune[5]
port 14 nsew
flabel metal1 10326 -65516 10424 -65204 0 FreeSans 1600 0 0 0 pa_tune[4]
port 15 nsew
flabel metal1 10326 -57658 10424 -57346 0 FreeSans 1600 0 0 0 pa_tune[3]
port 16 nsew
flabel metal1 10326 -53044 10424 -52732 0 FreeSans 1600 0 0 0 pa_tune[2]
port 17 nsew
flabel metal1 10326 -50052 10424 -49740 0 FreeSans 1600 0 0 0 pa_tune[1]
port 18 nsew
flabel metal2 19542 -48852 19614 -47598 0 FreeSans 1600 90 0 0 trigger_line[0]
port 13 nsew
flabel metal2 20134 -48918 20206 -47598 0 FreeSans 1600 90 0 0 trigger_line[1]
port 12 nsew
flabel metal3 18960 -69934 20784 -69838 0 FreeSans 1600 0 0 0 in_uwb
port 3 nsew
flabel metal1 19361 -58006 19905 -57960 0 FreeSans 1600 0 0 0 delayline[5]
port 6 nsew
flabel metal1 19361 -62224 19905 -62178 0 FreeSans 1600 0 0 0 delayline[4]
port 7 nsew
flabel metal1 19361 -65550 19905 -65504 0 FreeSans 1600 0 0 0 delayline[2]
port 9 nsew
flabel metal1 19361 -64398 19905 -64352 0 FreeSans 1600 0 0 0 delayline[3]
port 8 nsew
flabel metal1 19361 -66572 19905 -66526 0 FreeSans 1600 0 0 0 delayline[1]
port 10 nsew
flabel metal1 19361 -67594 19905 -67548 0 FreeSans 1600 0 0 0 delayline[0]
port 11 nsew
flabel metal5 -13104 -102827 -11014 -101827 0 FreeSans 1600 0 0 0 outp_uwb
port 46 nsew
flabel metal5 -13104 -90973 -11014 -89973 0 FreeSans 1600 0 0 0 outn_uwb
port 45 nsew
flabel metal1 10326 -47060 10424 -46748 0 FreeSans 1600 0 0 0 pa_tune[0]
port 19 nsew
flabel metal2 8953 -36646 11755 -36550 0 FreeSans 1600 0 0 0 pa_trig1_test
port 37 nsew
<< end >>
